library ieee;
use ieee.std_logic_1164.all;

entity top is
port(
    dest_x: in std_logic_vector(29 downto 0);
    dest_y: in std_logic_vector(29 downto 0);
    outport: out std_logic_vector(29 downto 0));
	end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256: std_logic;

begin

w0 <= not dest_x(9) and not dest_x(10);
w1 <= dest_x(9) and dest_x(10);
w2 <= not w0 and not w1;
w3 <= dest_x(11) and not w0;
w4 <= not dest_x(11) and w0;
w5 <= not w3 and not w4;
w6 <= not dest_x(12) and not w3;
w7 <= dest_x(12) and w3;
w8 <= not w6 and not w7;
w9 <= not dest_x(13) and w6;
w10 <= dest_x(13) and not w6;
w11 <= not w9 and not w10;
w12 <= dest_x(14) and not w9;
w13 <= not dest_x(14) and w9;
w14 <= not w12 and not w13;
w15 <= dest_x(15) and not w12;
w16 <= not dest_x(15) and w12;
w17 <= not w15 and not w16;
w18 <= dest_x(15) and w12;
w19 <= not dest_x(16) and not w18;
w20 <= dest_x(16) and w18;
w21 <= not w19 and not w20;
w22 <= dest_x(17) and not w19;
w23 <= not dest_x(17) and w19;
w24 <= not w22 and not w23;
w25 <= not dest_x(18) and not w22;
w26 <= dest_x(18) and w22;
w27 <= not w25 and not w26;
w28 <= dest_x(19) and not w25;
w29 <= not dest_x(19) and w25;
w30 <= not w28 and not w29;
w31 <= dest_x(20) and not w28;
w32 <= not dest_x(20) and w28;
w33 <= not w31 and not w32;
w34 <= dest_x(20) and w28;
w35 <= not dest_x(21) and not w34;
w36 <= dest_x(21) and w34;
w37 <= not w35 and not w36;
w38 <= not dest_x(22) and w35;
w39 <= dest_x(22) and not w35;
w40 <= not w38 and not w39;
w41 <= dest_x(23) and not w38;
w42 <= not dest_x(23) and w38;
w43 <= not w41 and not w42;
w44 <= dest_x(24) and not w41;
w45 <= not dest_x(24) and w41;
w46 <= not w44 and not w45;
w47 <= dest_x(24) and w41;
w48 <= dest_x(25) and not w47;
w49 <= not dest_x(25) and w47;
w50 <= not w48 and not w49;
w51 <= dest_x(25) and w47;
w52 <= not dest_x(26) and not w51;
w53 <= dest_x(26) and w51;
w54 <= not w52 and not w53;
w55 <= dest_x(27) and not w52;
w56 <= not dest_x(27) and w52;
w57 <= not w55 and not w56;
w58 <= dest_x(28) and not w55;
w59 <= not dest_x(28) and w55;
w60 <= not w58 and not w59;
w61 <= dest_x(28) and w55;
w62 <= not dest_x(29) and w61;
w63 <= dest_x(29) and not w61;
w64 <= not w62 and not w63;
w65 <= not dest_x(9) and not w64;
w66 <= not w60 and w65;
w67 <= w57 and w66;
w68 <= not w54 and w67;
w69 <= not w50 and w68;
w70 <= not w46 and w69;
w71 <= w43 and w70;
w72 <= not w40 and w71;
w73 <= not w37 and w72;
w74 <= not w33 and w73;
w75 <= w30 and w74;
w76 <= not w27 and w75;
w77 <= w24 and w76;
w78 <= not w21 and w77;
w79 <= not w17 and w78;
w80 <= w14 and w79;
w81 <= not w11 and w80;
w82 <= not w8 and w81;
w83 <= w5 and w82;
w84 <= not w2 and w83;
w85 <= dest_x(8) and w84;
w86 <= dest_x(7) and w85;
w87 <= dest_x(6) and w86;
w88 <= dest_x(5) and w87;
w89 <= dest_x(4) and w88;
w90 <= dest_x(3) and w89;
w91 <= dest_x(2) and w90;
w92 <= dest_x(1) and w91;
w93 <= dest_x(0) and w92;
w94 <= dest_x(29) and w61;
w95 <= not w93 and not w94;
w96 <= not dest_x(1) and not dest_x(2);
w97 <= not dest_x(3) and w96;
w98 <= not dest_x(4) and w97;
w99 <= not dest_x(5) and w98;
w100 <= not dest_x(6) and w99;
w101 <= not dest_x(7) and w100;
w102 <= not dest_x(8) and w101;
w103 <= w2 and w102;
w104 <= not w5 and w103;
w105 <= w8 and w104;
w106 <= w11 and w105;
w107 <= not w14 and w106;
w108 <= w17 and w107;
w109 <= w21 and w108;
w110 <= not w24 and w109;
w111 <= w27 and w110;
w112 <= not w30 and w111;
w113 <= w33 and w112;
w114 <= w37 and w113;
w115 <= w40 and w114;
w116 <= not w43 and w115;
w117 <= w46 and w116;
w118 <= w50 and w117;
w119 <= w54 and w118;
w120 <= not w57 and w119;
w121 <= w60 and w120;
w122 <= dest_x(9) and w121;
w123 <= w94 and not w122;
w124 <= not w95 and not w123;
w125 <= not dest_y(9) and not dest_y(10);
w126 <= dest_y(11) and not w125;
w127 <= not dest_y(12) and not w126;
w128 <= not dest_y(13) and w127;
w129 <= dest_y(14) and not w128;
w130 <= dest_y(15) and w129;
w131 <= not dest_y(16) and not w130;
w132 <= dest_y(17) and not w131;
w133 <= not dest_y(18) and not w132;
w134 <= dest_y(19) and not w133;
w135 <= dest_y(20) and w134;
w136 <= not dest_y(21) and not w135;
w137 <= not dest_y(22) and w136;
w138 <= dest_y(23) and not w137;
w139 <= dest_y(24) and w138;
w140 <= dest_y(25) and w139;
w141 <= not dest_y(26) and not w140;
w142 <= dest_y(27) and not w141;
w143 <= dest_y(28) and w142;
w144 <= dest_y(29) and w143;
w145 <= dest_x(0) and not w144;
w146 <= not dest_x(0) and not dest_y(0);
w147 <= w144 and not w146;
w148 <= dest_y(9) and dest_y(10);
w149 <= not w125 and not w148;
w150 <= not dest_y(11) and w125;
w151 <= not w126 and not w150;
w152 <= dest_y(12) and w126;
w153 <= not w127 and not w152;
w154 <= dest_y(13) and not w127;
w155 <= not w128 and not w154;
w156 <= not dest_y(14) and w128;
w157 <= not w129 and not w156;
w158 <= dest_y(15) and not w129;
w159 <= not dest_y(15) and w129;
w160 <= not w158 and not w159;
w161 <= dest_y(16) and w130;
w162 <= not w131 and not w161;
w163 <= not dest_y(17) and w131;
w164 <= not w132 and not w163;
w165 <= dest_y(18) and w132;
w166 <= not w133 and not w165;
w167 <= not dest_y(19) and w133;
w168 <= not w134 and not w167;
w169 <= dest_y(20) and not w134;
w170 <= not dest_y(20) and w134;
w171 <= not w169 and not w170;
w172 <= dest_y(21) and w135;
w173 <= not w136 and not w172;
w174 <= dest_y(22) and not w136;
w175 <= not w137 and not w174;
w176 <= not dest_y(23) and w137;
w177 <= not w138 and not w176;
w178 <= dest_y(24) and not w138;
w179 <= not dest_y(24) and w138;
w180 <= not w178 and not w179;
w181 <= dest_y(25) and not w139;
w182 <= not dest_y(25) and w139;
w183 <= not w181 and not w182;
w184 <= dest_y(26) and w140;
w185 <= not w141 and not w184;
w186 <= not dest_y(27) and w141;
w187 <= not w142 and not w186;
w188 <= dest_y(28) and not w142;
w189 <= not dest_y(28) and w142;
w190 <= not w188 and not w189;
w191 <= dest_y(0) and not dest_y(9);
w192 <= dest_y(29) and w191;
w193 <= not w190 and w192;
w194 <= w187 and w193;
w195 <= not w185 and w194;
w196 <= not w183 and w195;
w197 <= not w180 and w196;
w198 <= w177 and w197;
w199 <= not w175 and w198;
w200 <= not w173 and w199;
w201 <= not w171 and w200;
w202 <= w168 and w201;
w203 <= not w166 and w202;
w204 <= w164 and w203;
w205 <= not w162 and w204;
w206 <= not w160 and w205;
w207 <= w157 and w206;
w208 <= not w155 and w207;
w209 <= not w153 and w208;
w210 <= w151 and w209;
w211 <= not w149 and w210;
w212 <= dest_y(8) and w211;
w213 <= dest_y(7) and w212;
w214 <= dest_y(6) and w213;
w215 <= dest_y(5) and w214;
w216 <= dest_y(4) and w215;
w217 <= dest_y(3) and w216;
w218 <= dest_y(2) and w217;
w219 <= dest_y(1) and w218;
w220 <= not dest_y(1) and not dest_y(2);
w221 <= not dest_y(3) and w220;
w222 <= not dest_y(4) and w221;
w223 <= not dest_y(5) and w222;
w224 <= not dest_y(6) and w223;
w225 <= not dest_y(7) and w224;
w226 <= not dest_y(8) and w225;
w227 <= w149 and w226;
w228 <= not w151 and w227;
w229 <= w153 and w228;
w230 <= w155 and w229;
w231 <= not w157 and w230;
w232 <= w160 and w231;
w233 <= w162 and w232;
w234 <= not w164 and w233;
w235 <= w166 and w234;
w236 <= not w168 and w235;
w237 <= w171 and w236;
w238 <= w173 and w237;
w239 <= w175 and w238;
w240 <= not w177 and w239;
w241 <= w180 and w240;
w242 <= w183 and w241;
w243 <= w185 and w242;
w244 <= not w187 and w243;
w245 <= w190 and w244;
w246 <= dest_y(9) and w245;
w247 <= w144 and not w246;
w248 <= not w219 and not w247;
w249 <= not w147 and w248;
w250 <= not w95 and not w249;
w251 <= not w145 and w250;
w252 <= not w123 and not w251;
w253 <= dest_x(0) and w144;
w254 <= dest_y(0) and w253;
w255 <= not w247 and not w254;
w256 <= w124 and not w255;
one <= '1';
outport(0) <= not w124;-- level 52
outport(1) <= w252;-- level 54
outport(2) <= w256;-- level 53
outport(3) <= not one;-- level 0
outport(4) <= not one;-- level 0
outport(5) <= not one;-- level 0
outport(6) <= not one;-- level 0
outport(7) <= not one;-- level 0
outport(8) <= not one;-- level 0
outport(9) <= not one;-- level 0
outport(10) <= not one;-- level 0
outport(11) <= not one;-- level 0
outport(12) <= not one;-- level 0
outport(13) <= not one;-- level 0
outport(14) <= not one;-- level 0
outport(15) <= not one;-- level 0
outport(16) <= not one;-- level 0
outport(17) <= not one;-- level 0
outport(18) <= not one;-- level 0
outport(19) <= not one;-- level 0
outport(20) <= not one;-- level 0
outport(21) <= not one;-- level 0
outport(22) <= not one;-- level 0
outport(23) <= not one;-- level 0
outport(24) <= not one;-- level 0
outport(25) <= not one;-- level 0
outport(26) <= not one;-- level 0
outport(27) <= not one;-- level 0
outport(28) <= not one;-- level 0
outport(29) <= not one;-- level 0
end Behavioral;
