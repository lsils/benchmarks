module mem_ctrl ( 
    pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008,
    pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017,
    pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026,
    pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035,
    pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044,
    pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053,
    pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
    pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
    pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080,
    pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089,
    pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098,
    pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107,
    pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116,
    pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125,
    pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
    pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
    pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152,
    pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161,
    pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170,
    pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179,
    pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188,
    pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197,
    pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
    pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
    pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224,
    pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233,
    pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242,
    pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251,
    pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260,
    pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269,
    pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
    pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
    pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296,
    pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305,
    pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314,
    pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323,
    pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332,
    pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341,
    pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
    pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
    pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368,
    pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377,
    pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386,
    pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395,
    pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404,
    pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413,
    pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
    pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
    pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440,
    pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449,
    pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458,
    pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467,
    pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476,
    pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485,
    pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
    pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
    pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512,
    pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521,
    pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530,
    pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539,
    pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548,
    pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557,
    pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
    pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
    pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584,
    pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593,
    pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602,
    pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611,
    pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620,
    pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629,
    pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
    pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
    pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656,
    pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665,
    pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674,
    pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683,
    pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692,
    pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701,
    pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
    pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
    pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728,
    pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737,
    pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746,
    pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755,
    pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764,
    pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773,
    pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
    pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
    pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800,
    pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809,
    pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818,
    pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827,
    pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836,
    pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845,
    pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
    pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
    pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872,
    pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881,
    pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890,
    pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899,
    pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908,
    pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917,
    pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
    pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
    pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944,
    pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953,
    pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962,
    pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971,
    pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980,
    pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989,
    pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
    pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230  );
  input  pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
    pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016,
    pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025,
    pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034,
    pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043,
    pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052,
    pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061,
    pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
    pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
    pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088,
    pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097,
    pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106,
    pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115,
    pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124,
    pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133,
    pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
    pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
    pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160,
    pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169,
    pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178,
    pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187,
    pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196,
    pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205,
    pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
    pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
    pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232,
    pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241,
    pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250,
    pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259,
    pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268,
    pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277,
    pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
    pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
    pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304,
    pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313,
    pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322,
    pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331,
    pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340,
    pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349,
    pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
    pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
    pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376,
    pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385,
    pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394,
    pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403,
    pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412,
    pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421,
    pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
    pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
    pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448,
    pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457,
    pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466,
    pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475,
    pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484,
    pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493,
    pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
    pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
    pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520,
    pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529,
    pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538,
    pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547,
    pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556,
    pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565,
    pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
    pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
    pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592,
    pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601,
    pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610,
    pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619,
    pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628,
    pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637,
    pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
    pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
    pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664,
    pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673,
    pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682,
    pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691,
    pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700,
    pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709,
    pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
    pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
    pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736,
    pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745,
    pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754,
    pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763,
    pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772,
    pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781,
    pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
    pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
    pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808,
    pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817,
    pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826,
    pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835,
    pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844,
    pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853,
    pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
    pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
    pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880,
    pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889,
    pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898,
    pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907,
    pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916,
    pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925,
    pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
    pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
    pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952,
    pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961,
    pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970,
    pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979,
    pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988,
    pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997,
    pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
    n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
    n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
    n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
    n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
    n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
    n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
    n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
    n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
    n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
    n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
    n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
    n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
    n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
    n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
    n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
    n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
    n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
    n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
    n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
    n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
    n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
    n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
    n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
    n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
    n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
    n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
    n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
    n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
    n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
    n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
    n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
    n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
    n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
    n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
    n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
    n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
    n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
    n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
    n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
    n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
    n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
    n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
    n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
    n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
    n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
    n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
    n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
    n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
    n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
    n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
    n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
    n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
    n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
    n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
    n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
    n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
    n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
    n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
    n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
    n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
    n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
    n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
    n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
    n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
    n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
    n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
    n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
    n3307, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
    n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
    n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
    n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
    n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
    n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
    n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
    n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
    n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
    n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
    n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
    n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
    n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
    n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
    n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
    n3538, n3539, n3540, n3541, n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
    n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
    n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
    n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
    n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
    n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
    n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
    n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
    n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
    n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
    n3709, n3710, n3711, n3712, n3714, n3715, n3716, n3717, n3718, n3719,
    n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
    n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
    n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
    n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
    n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
    n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
    n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
    n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
    n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
    n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
    n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
    n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
    n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
    n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
    n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3942, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
    n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
    n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
    n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
    n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
    n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
    n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
    n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
    n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
    n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
    n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
    n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
    n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
    n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
    n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
    n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
    n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
    n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4171,
    n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
    n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
    n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
    n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
    n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
    n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
    n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
    n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
    n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
    n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
    n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
    n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
    n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
    n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
    n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
    n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
    n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
    n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
    n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
    n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
    n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
    n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
    n4392, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
    n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
    n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
    n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
    n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
    n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
    n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
    n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
    n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
    n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
    n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
    n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
    n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
    n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
    n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
    n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
    n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
    n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
    n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
    n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
    n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
    n4613, n4614, n4615, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
    n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
    n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
    n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
    n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
    n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
    n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
    n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
    n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
    n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
    n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
    n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
    n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
    n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
    n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
    n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
    n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
    n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
    n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
    n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
    n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
    n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
    n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
    n4844, n4845, n4846, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
    n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
    n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
    n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
    n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
    n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
    n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
    n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
    n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
    n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
    n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
    n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
    n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
    n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
    n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
    n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
    n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
    n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
    n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
    n5065, n5066, n5067, n5068, n5069, n5071, n5072, n5073, n5074, n5075,
    n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
    n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
    n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
    n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
    n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
    n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
    n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
    n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
    n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
    n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
    n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
    n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
    n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
    n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
    n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
    n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
    n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
    n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
    n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
    n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
    n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5294, n5295, n5296,
    n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
    n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
    n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
    n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
    n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
    n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
    n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
    n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
    n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
    n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
    n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
    n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
    n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
    n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
    n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
    n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
    n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
    n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
    n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
    n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
    n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
    n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
    n5527, n5528, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
    n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
    n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
    n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
    n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
    n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
    n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
    n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
    n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
    n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
    n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
    n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
    n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
    n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
    n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
    n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
    n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
    n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
    n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
    n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
    n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
    n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
    n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
    n5758, n5759, n5760, n5761, n5762, n5763, n5765, n5766, n5767, n5768,
    n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
    n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
    n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
    n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
    n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
    n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
    n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
    n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
    n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
    n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
    n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
    n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
    n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
    n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
    n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
    n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
    n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
    n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
    n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
    n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
    n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
    n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
    n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
    n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
    n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
    n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
    n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
    n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
    n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
    n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
    n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
    n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
    n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
    n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
    n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
    n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
    n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
    n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
    n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
    n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
    n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
    n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
    n6190, n6191, n6192, n6193, n6194, n6195, n6197, n6198, n6199, n6200,
    n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
    n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
    n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
    n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
    n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
    n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
    n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
    n6271, n6272, n6273, n6275, n6276, n6277, n6279, n6280, n6281, n6282,
    n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
    n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
    n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
    n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
    n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
    n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
    n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
    n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
    n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
    n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
    n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
    n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
    n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
    n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
    n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
    n6434, n6435, n6436, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
    n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
    n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
    n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
    n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
    n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
    n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
    n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
    n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
    n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
    n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
    n6565, n6566, n6567, n6568, n6569, n6570, n6572, n6573, n6574, n6575,
    n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
    n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
    n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
    n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
    n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
    n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
    n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
    n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
    n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6695, n6696,
    n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
    n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
    n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
    n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
    n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
    n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
    n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
    n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
    n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
    n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
    n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
    n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6825, n6826, n6827,
    n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
    n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
    n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
    n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
    n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
    n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
    n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
    n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
    n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
    n6918, n6919, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
    n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
    n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
    n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
    n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
    n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
    n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
    n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
    n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
    n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7017, n7018, n7019,
    n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
    n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
    n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
    n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
    n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
    n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
    n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
    n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
    n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
    n7110, n7111, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
    n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
    n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
    n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
    n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
    n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
    n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
    n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
    n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
    n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7209, n7210, n7211,
    n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
    n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
    n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
    n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
    n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
    n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
    n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
    n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
    n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7301, n7302,
    n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
    n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
    n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
    n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
    n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7353,
    n7354, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
    n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
    n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
    n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
    n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
    n7406, n7407, n7408, n7409, n7411, n7413, n7415, n7417, n7418, n7419,
    n7420, n7421, n7422, n7423, n7424, n7425, n7427, n7428, n7429, n7430,
    n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
    n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
    n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
    n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
    n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
    n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
    n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
    n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
    n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
    n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
    n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
    n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
    n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
    n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
    n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
    n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
    n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
    n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
    n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
    n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
    n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
    n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
    n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
    n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
    n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
    n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
    n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
    n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
    n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
    n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
    n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
    n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
    n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
    n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
    n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
    n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
    n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
    n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
    n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
    n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
    n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
    n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
    n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
    n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
    n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
    n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
    n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
    n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
    n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
    n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
    n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
    n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
    n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
    n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
    n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
    n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
    n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
    n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
    n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
    n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
    n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
    n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
    n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
    n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
    n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
    n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
    n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
    n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
    n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
    n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
    n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
    n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
    n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
    n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
    n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
    n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
    n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
    n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
    n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
    n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
    n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
    n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
    n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
    n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
    n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
    n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
    n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
    n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
    n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
    n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
    n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
    n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
    n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
    n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
    n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
    n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
    n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
    n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
    n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
    n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
    n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
    n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
    n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
    n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
    n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
    n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
    n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
    n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
    n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
    n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
    n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
    n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
    n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
    n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
    n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
    n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
    n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
    n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
    n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
    n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
    n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
    n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
    n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
    n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
    n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
    n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
    n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
    n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
    n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
    n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
    n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
    n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
    n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
    n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
    n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
    n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
    n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
    n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
    n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
    n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
    n8871, n8872, n8873, n8874, n8875, n8876, n8878, n8879, n8880, n8881,
    n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
    n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
    n8902, n8903, n8904, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
    n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
    n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
    n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
    n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
    n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
    n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
    n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
    n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
    n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
    n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
    n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
    n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
    n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
    n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
    n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
    n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
    n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
    n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
    n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
    n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
    n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
    n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
    n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
    n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
    n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
    n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
    n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
    n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
    n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
    n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
    n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
    n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
    n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
    n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
    n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
    n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
    n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
    n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
    n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
    n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
    n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
    n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
    n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
    n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
    n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
    n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
    n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
    n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
    n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
    n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
    n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
    n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
    n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
    n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
    n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
    n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
    n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
    n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
    n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
    n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
    n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
    n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
    n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
    n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
    n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
    n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
    n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
    n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
    n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
    n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
    n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
    n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
    n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
    n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
    n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
    n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
    n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
    n9684, n9685, n9686, n9687, n9688, n9689, n9691, n9692, n9693, n9694,
    n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
    n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
    n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
    n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
    n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
    n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
    n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
    n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
    n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
    n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
    n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
    n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
    n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
    n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
    n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
    n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
    n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
    n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
    n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
    n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
    n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
    n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
    n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
    n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
    n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
    n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
    n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
    n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
    n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
    n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
    n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
    n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
    n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
    n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
    n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
    n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
    n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10067,
    n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
    n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
    n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
    n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
    n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
    n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
    n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
    n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
    n10140, n10141, n10142, n10143, n10144, n10145, n10147, n10148, n10149,
    n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
    n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
    n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
    n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
    n10196, n10197, n10198, n10200, n10201, n10202, n10203, n10204, n10205,
    n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
    n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
    n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
    n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
    n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
    n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
    n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
    n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
    n10278, n10279, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
    n10288, n10289, n10290, n10291, n10292, n10293, n10295, n10296, n10297,
    n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
    n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
    n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
    n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
    n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
    n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
    n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
    n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
    n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
    n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
    n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
    n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
    n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
    n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
    n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
    n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
    n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
    n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
    n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
    n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
    n10478, n10479, n10480, n10481, n10482, n10484, n10485, n10486, n10487,
    n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
    n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
    n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
    n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
    n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
    n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
    n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
    n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
    n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
    n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
    n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
    n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
    n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
    n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
    n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
    n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
    n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
    n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
    n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
    n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
    n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
    n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
    n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
    n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
    n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
    n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
    n10722, n10723, n10724, n10725, n10726, n10727, n10729, n10730, n10731,
    n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
    n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
    n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
    n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
    n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
    n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
    n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
    n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
    n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
    n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
    n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
    n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
    n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
    n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
    n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
    n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
    n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
    n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
    n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
    n10903, n10904, n10905, n10907, n10908, n10909, n10910, n10911, n10912,
    n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
    n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
    n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
    n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
    n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
    n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
    n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
    n10976, n10977, n10978, n10979, n10980, n10982, n10983, n10984, n10986,
    n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
    n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
    n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
    n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
    n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
    n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
    n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11051,
    n11052, n11053, n11054, n11055, n11057, n11058, n11059, n11060, n11061,
    n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
    n11071, n11072, n11073, n11074, n11076, n11077, n11078, n11079, n11080,
    n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
    n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
    n11099, n11100, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
    n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
    n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
    n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
    n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
    n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
    n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
    n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
    n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
    n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
    n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
    n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
    n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
    n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
    n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
    n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
    n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
    n11254, n11255, n11256, n11257, n11258, n11259, n11261, n11262, n11263,
    n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11273,
    n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
    n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
    n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
    n11302, n11303, n11304, n11305, n11307, n11308, n11309, n11310, n11311,
    n11312, n11313, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
    n11322, n11323, n11325, n11326, n11328, n11329, n11330, n11331, n11332,
    n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11343,
    n11344, n11345, n11346, n11348, n11349, n11350, n11351, n11353, n11354,
    n11355, n11356, n11357, n11359, n11360, n11361, n11362, n11363, n11364,
    n11365, n11366, n11367, n11369, n11370, n11371, n11373, n11374, n11375,
    n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
    n11385, n11386, n11387, n11388, n11390, n11391, n11392, n11393, n11395,
    n11396, n11397, n11398, n11399, n11400, n11401, n11403, n11404, n11405,
    n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
    n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
    n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
    n11434, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
    n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
    n11453, n11454, n11455, n11456, n11458, n11459, n11460, n11461, n11462,
    n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
    n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
    n11482, n11483, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
    n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11500, n11501,
    n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11510, n11511,
    n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
    n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
    n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
    n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
    n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
    n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
    n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
    n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
    n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
    n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
    n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
    n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
    n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
    n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
    n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
    n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
    n11656, n11657, n11658, n11659, n11660, n11661, n11663, n11664, n11665,
    n11666, n11667, n11668, n11669, n11670, n11671, n11673, n11675, n11676,
    n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
    n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
    n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
    n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
    n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
    n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
    n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
    n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
    n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
    n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
    n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
    n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
    n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
    n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
    n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
    n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
    n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
    n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
    n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
    n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
    n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
    n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
    n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
    n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
    n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
    n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
    n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
    n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
    n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
    n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
    n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
    n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
    n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
    n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
    n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
    n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
    n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
    n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
    n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
    n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
    n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
    n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
    n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
    n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
    n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
    n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
    n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
    n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
    n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
    n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
    n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
    n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
    n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
    n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
    n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
    n12172, n12173, n12174, n12175, n12176, n12178, n12179, n12180, n12181,
    n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
    n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
    n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
    n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
    n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
    n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
    n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
    n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
    n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
    n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
    n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
    n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
    n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
    n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
    n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
    n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
    n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
    n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
    n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
    n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
    n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
    n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
    n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
    n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
    n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
    n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
    n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
    n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
    n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
    n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
    n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
    n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
    n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
    n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
    n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
    n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
    n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
    n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
    n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
    n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
    n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
    n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
    n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
    n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
    n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
    n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
    n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
    n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
    n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
    n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
    n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
    n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
    n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
    n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
    n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
    n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
    n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
    n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
    n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
    n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
    n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
    n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
    n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
    n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
    n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
    n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
    n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
    n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
    n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
    n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
    n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
    n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
    n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
    n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
    n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
    n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
    n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
    n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
    n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
    n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
    n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
    n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
    n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
    n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
    n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
    n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
    n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
    n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
    n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
    n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
    n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
    n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
    n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
    n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
    n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
    n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13047, n13048,
    n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
    n13058, n13059, n13061, n13062, n13063, n13064, n13065, n13067, n13068,
    n13069, n13070, n13072, n13073, n13074, n13076, n13077, n13078, n13080,
    n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
    n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
    n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
    n13110, n13111, n13112, n13113, n13115, n13116, n13117, n13118, n13119,
    n13120, n13121, n13122, n13123, n13124, n13125, n13127, n13128, n13129,
    n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13139,
    n13140, n13141, n13142, n13143, n13144, n13146, n13147, n13148, n13149,
    n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
    n13159, n13160, n13161, n13162, n13164, n13165, n13166, n13167, n13168,
    n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
    n13178, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
    n13188, n13189, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
    n13198, n13199, n13201, n13202, n13203, n13204, n13206, n13207, n13208,
    n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
    n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
    n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
    n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
    n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
    n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
    n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
    n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
    n13281, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
    n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13300,
    n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
    n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
    n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
    n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
    n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
    n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
    n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
    n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
    n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13381, n13383,
    n13384, n13385, n13386, n13387, n13388, n13389, n13391, n13392, n13393,
    n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
    n13403, n13404, n13405, n13406, n13407, n13409, n13410, n13411, n13412,
    n13413, n13414, n13415, n13416, n13417, n13419, n13421, n13422, n13423,
    n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
    n13433, n13434, n13435, n13436, n13437, n13439, n13441, n13442, n13443,
    n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13452, n13453,
    n13454, n13455, n13456, n13459, n13460, n13461, n13462, n13463, n13464,
    n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
    n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
    n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
    n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
    n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
    n13510, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
    n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
    n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
    n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
    n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13555, n13556,
    n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
    n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
    n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
    n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
    n13593, n13594, n13595, n13597, n13598, n13599, n13600, n13601, n13602,
    n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
    n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
    n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
    n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
    n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13648,
    n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
    n13658, n13659, n13660, n13661, n13662, n13664, n13665, n13666, n13667,
    n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
    n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
    n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
    n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
    n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
    n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
    n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
    n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
    n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
    n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
    n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
    n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
    n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
    n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
    n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
    n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
    n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
    n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
    n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
    n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
    n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
    n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
    n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
    n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
    n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
    n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
    n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
    n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
    n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
    n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
    n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
    n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
    n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
    n13965, n13966, n13967, n13969, n13970, n13971, n13972, n13973, n13974,
    n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
    n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
    n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
    n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
    n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
    n14020, n14021, n14022, n14024, n14025, n14026, n14027, n14028, n14029,
    n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
    n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
    n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
    n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
    n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
    n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
    n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
    n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
    n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
    n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
    n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
    n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
    n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
    n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
    n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
    n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
    n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
    n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
    n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
    n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
    n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
    n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
    n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
    n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
    n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
    n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
    n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
    n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
    n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
    n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
    n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
    n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
    n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
    n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
    n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
    n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
    n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
    n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
    n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
    n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
    n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
    n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
    n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
    n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
    n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
    n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
    n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
    n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
    n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
    n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
    n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
    n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
    n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
    n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
    n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
    n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
    n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
    n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
    n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
    n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
    n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
    n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
    n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
    n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
    n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
    n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
    n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
    n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
    n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
    n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
    n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
    n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
    n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
    n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
    n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
    n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
    n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
    n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
    n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
    n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
    n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
    n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
    n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
    n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
    n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
    n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
    n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
    n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
    n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
    n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
    n14841, n14842, n14843, n14844, n14845, n14847, n14848, n14849, n14850,
    n14851, n14852, n14853, n14855, n14856, n14857, n14858, n14859, n14860,
    n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
    n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
    n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
    n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
    n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
    n14906, n14907, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
    n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
    n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
    n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
    n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
    n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
    n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
    n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
    n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
    n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
    n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
    n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
    n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
    n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
    n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
    n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
    n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
    n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
    n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
    n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
    n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
    n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
    n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
    n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
    n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
    n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
    n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
    n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
    n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
    n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
    n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
    n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
    n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
    n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
    n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
    n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
    n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
    n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
    n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
    n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
    n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
    n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
    n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
    n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
    n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
    n15312, n15313, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
    n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
    n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
    n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
    n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
    n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
    n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
    n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
    n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
    n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
    n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
    n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
    n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
    n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
    n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
    n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
    n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
    n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
    n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
    n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
    n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
    n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
    n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
    n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
    n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
    n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
    n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
    n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
    n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
    n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
    n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
    n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
    n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
    n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15618, n15619,
    n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
    n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
    n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
    n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
    n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
    n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
    n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
    n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
    n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
    n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
    n15710, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
    n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
    n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15737, n15738,
    n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
    n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
    n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
    n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
    n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
    n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
    n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
    n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
    n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
    n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
    n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
    n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
    n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
    n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
    n15865, n15866, n15867, n15868, n15869, n15870, n15872, n15873, n15874,
    n15875, n15876, n15877, n15878, n15880, n15881, n15882, n15883, n15884,
    n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
    n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
    n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
    n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
    n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
    n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
    n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
    n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
    n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
    n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
    n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
    n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
    n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
    n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
    n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
    n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
    n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
    n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
    n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
    n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
    n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
    n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
    n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
    n16092, n16093, n16094, n16096, n16097, n16098, n16099, n16100, n16101,
    n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
    n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
    n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
    n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
    n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
    n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
    n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
    n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
    n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
    n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
    n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
    n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
    n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
    n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
    n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
    n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
    n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
    n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
    n16265, n16266, n16267, n16268, n16269, n16271, n16272, n16273, n16274,
    n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
    n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
    n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
    n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
    n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
    n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
    n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
    n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
    n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
    n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
    n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
    n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
    n16383, n16384, n16385, n16386, n16387, n16388, n16390, n16391, n16392,
    n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
    n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
    n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
    n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
    n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
    n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
    n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
    n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
    n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
    n16474, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
    n16484, n16485, n16486, n16487, n16489, n16490, n16491, n16492, n16493,
    n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
    n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
    n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
    n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
    n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
    n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
    n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
    n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
    n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16574, n16575,
    n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
    n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
    n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
    n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
    n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
    n16621, n16622, n16623, n16624, n16625, n16626, n16628, n16629, n16630,
    n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
    n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
    n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
    n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
    n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
    n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
    n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
    n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
    n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
    n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
    n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
    n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
    n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
    n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
    n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
    n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
    n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
    n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
    n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
    n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
    n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
    n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
    n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
    n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
    n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
    n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
    n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
    n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
    n16883, n16884, n16885, n16886, n16887, n16889, n16890, n16891, n16892,
    n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
    n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
    n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
    n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
    n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
    n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
    n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
    n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
    n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
    n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
    n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
    n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
    n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
    n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
    n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
    n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
    n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
    n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
    n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
    n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
    n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
    n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
    n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
    n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
    n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
    n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
    n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
    n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
    n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
    n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
    n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
    n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
    n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
    n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
    n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
    n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
    n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
    n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
    n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
    n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
    n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
    n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
    n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
    n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
    n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
    n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
    n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
    n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
    n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
    n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
    n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
    n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
    n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
    n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
    n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
    n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
    n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
    n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
    n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
    n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
    n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
    n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
    n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
    n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
    n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
    n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
    n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
    n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
    n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
    n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
    n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
    n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
    n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
    n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
    n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
    n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
    n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
    n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
    n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
    n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
    n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
    n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
    n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
    n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
    n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
    n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
    n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
    n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
    n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
    n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
    n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
    n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
    n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
    n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
    n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
    n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
    n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
    n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
    n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
    n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
    n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
    n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
    n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
    n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
    n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
    n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
    n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
    n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
    n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
    n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
    n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
    n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
    n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
    n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
    n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
    n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
    n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
    n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
    n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
    n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
    n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
    n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
    n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
    n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
    n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
    n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
    n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
    n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
    n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
    n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
    n18063, n18064, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
    n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
    n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
    n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
    n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
    n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
    n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
    n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
    n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
    n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
    n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
    n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
    n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
    n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
    n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
    n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
    n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
    n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
    n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
    n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
    n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
    n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
    n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
    n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
    n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
    n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
    n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
    n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
    n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
    n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
    n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
    n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
    n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
    n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
    n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
    n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
    n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
    n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
    n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
    n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
    n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
    n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
    n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
    n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
    n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
    n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
    n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
    n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
    n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
    n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
    n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
    n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
    n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
    n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
    n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
    n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
    n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
    n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
    n18586, n18587, n18588, n18589, n18591, n18592, n18593, n18594, n18595,
    n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
    n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
    n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
    n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
    n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
    n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
    n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
    n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
    n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
    n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
    n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
    n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
    n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
    n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
    n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
    n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
    n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
    n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
    n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
    n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
    n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
    n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
    n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
    n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
    n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
    n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
    n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
    n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
    n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
    n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
    n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
    n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
    n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
    n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
    n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
    n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
    n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
    n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
    n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
    n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
    n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
    n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
    n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
    n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
    n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
    n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
    n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
    n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
    n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
    n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
    n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
    n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
    n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
    n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
    n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
    n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
    n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
    n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
    n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
    n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
    n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
    n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
    n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
    n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
    n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
    n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
    n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
    n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
    n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
    n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
    n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
    n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
    n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
    n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
    n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
    n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
    n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
    n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
    n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
    n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
    n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
    n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
    n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
    n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
    n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
    n19361, n19362, n19363, n19364, n19366, n19367, n19368, n19369, n19370,
    n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
    n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
    n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
    n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
    n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
    n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
    n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
    n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
    n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
    n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
    n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
    n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
    n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
    n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
    n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
    n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
    n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
    n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
    n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
    n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
    n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
    n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
    n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
    n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
    n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
    n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
    n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
    n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
    n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
    n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
    n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
    n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
    n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
    n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
    n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
    n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
    n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
    n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
    n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
    n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
    n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
    n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
    n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
    n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
    n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
    n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
    n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
    n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
    n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
    n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
    n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
    n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
    n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
    n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
    n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
    n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
    n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
    n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19892, n19893,
    n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
    n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
    n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
    n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
    n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
    n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
    n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
    n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
    n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
    n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
    n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
    n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
    n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
    n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
    n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
    n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
    n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
    n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
    n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
    n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
    n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
    n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
    n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
    n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
    n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
    n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
    n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
    n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
    n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
    n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
    n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
    n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
    n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
    n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
    n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
    n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
    n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
    n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
    n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
    n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
    n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
    n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
    n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
    n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
    n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
    n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
    n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
    n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
    n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
    n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
    n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
    n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
    n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
    n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
    n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
    n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
    n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
    n20407, n20408, n20409, n20411, n20412, n20413, n20414, n20415, n20416,
    n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
    n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
    n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
    n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
    n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
    n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
    n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
    n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
    n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
    n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
    n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
    n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
    n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
    n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
    n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
    n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
    n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
    n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
    n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
    n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
    n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
    n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
    n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
    n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
    n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
    n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
    n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
    n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
    n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
    n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
    n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
    n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
    n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
    n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
    n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
    n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
    n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
    n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
    n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
    n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
    n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
    n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
    n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
    n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
    n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
    n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
    n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
    n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
    n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
    n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
    n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
    n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
    n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
    n20894, n20895, n20896, n20897, n20899, n20900, n20901, n20902, n20903,
    n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
    n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
    n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
    n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
    n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
    n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
    n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
    n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
    n20976, n20977, n20978, n20980, n20981, n20982, n20983, n20984, n20985,
    n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
    n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
    n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
    n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
    n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
    n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
    n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,
    n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
    n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
    n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
    n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
    n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
    n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
    n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
    n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120,
    n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21129, n21130,
    n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
    n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
    n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
    n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
    n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
    n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184,
    n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21193, n21194,
    n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
    n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
    n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
    n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
    n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
    n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248,
    n21249, n21250, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
    n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
    n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
    n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
    n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294,
    n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303,
    n21304, n21305, n21306, n21308, n21309, n21310, n21311, n21312, n21313,
    n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
    n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
    n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
    n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
    n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
    n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367,
    n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376,
    n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21386,
    n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
    n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404,
    n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413,
    n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422,
    n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431,
    n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,
    n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
    n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
    n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
    n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476,
    n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485,
    n21486, n21487, n21489, n21490, n21491, n21492, n21493, n21494, n21495,
    n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504,
    n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
    n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522,
    n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
    n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540,
    n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549,
    n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558,
    n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567,
    n21568, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
    n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
    n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
    n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
    n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613,
    n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21622, n21623,
    n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632,
    n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
    n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650,
    n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
    n21660, n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669,
    n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678,
    n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687,
    n21688, n21689, n21690, n21692, n21693, n21694, n21695, n21696, n21697,
    n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706,
    n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
    n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724,
    n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733,
    n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742,
    n21743, n21744, n21745, n21746, n21747, n21749, n21750, n21751, n21752,
    n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
    n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770,
    n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
    n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788,
    n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797,
    n21798, n21799, n21800, n21801, n21802, n21803, n21805, n21806, n21807,
    n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816,
    n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
    n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834,
    n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
    n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852,
    n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21861, n21862,
    n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
    n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880,
    n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
    n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898,
    n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
    n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
    n21917, n21918, n21920, n21921, n21922, n21923, n21924, n21925, n21926,
    n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
    n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944,
    n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
    n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962,
    n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971,
    n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980,
    n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989,
    n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998,
    n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
    n22008, n22009, n22010, n22011, n22012, n22013, n22015, n22016, n22017,
    n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026,
    n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035,
    n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044,
    n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053,
    n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062,
    n22063, n22064, n22065, n22066, n22067, n22068, n22070, n22071, n22072,
    n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
    n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090,
    n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
    n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108,
    n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117,
    n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126,
    n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136,
    n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
    n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154,
    n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
    n22164, n22165, n22166, n22168, n22169, n22170, n22171, n22172, n22173,
    n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182,
    n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191,
    n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200,
    n22201, n22202, n22203, n22204, n22205, n22206, n22208, n22209, n22210,
    n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
    n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228,
    n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237,
    n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246,
    n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255,
    n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264,
    n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
    n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282,
    n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291,
    n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300,
    n22301, n22302, n22303, n22305, n22306, n22307, n22308, n22309, n22310,
    n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319,
    n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328,
    n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
    n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346,
    n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356,
    n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365,
    n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374,
    n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383,
    n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392,
    n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
    n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410,
    n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419,
    n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22429,
    n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438,
    n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447,
    n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456,
    n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
    n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474,
    n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483,
    n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492,
    n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501,
    n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22510, n22511,
    n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520,
    n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
    n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538,
    n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547,
    n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556,
    n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565,
    n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574,
    n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583,
    n22584, n22585, n22586, n22587, n22588, n22590, n22591, n22592, n22593,
    n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602,
    n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611,
    n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620,
    n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629,
    n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638,
    n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647,
    n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656,
    n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
    n22666, n22667, n22668, n22669, n22671, n22672, n22673, n22674, n22675,
    n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684,
    n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693,
    n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702,
    n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711,
    n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720,
    n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
    n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738,
    n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747,
    n22748, n22749, n22750, n22752, n22753, n22754, n22755, n22756, n22757,
    n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766,
    n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775,
    n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784,
    n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
    n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802,
    n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811,
    n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820,
    n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829,
    n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838,
    n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847,
    n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856,
    n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
    n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874,
    n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883,
    n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892,
    n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901,
    n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910,
    n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919,
    n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928,
    n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
    n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946,
    n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955,
    n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964,
    n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973,
    n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982,
    n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991,
    n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000,
    n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
    n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018,
    n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027,
    n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036,
    n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045,
    n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054,
    n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063,
    n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072,
    n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
    n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090,
    n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099,
    n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108,
    n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117,
    n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126,
    n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135,
    n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144,
    n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
    n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162,
    n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171,
    n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180,
    n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189,
    n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198,
    n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207,
    n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216,
    n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
    n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235,
    n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244,
    n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253,
    n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262,
    n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271,
    n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280,
    n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
    n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298,
    n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307,
    n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316,
    n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325,
    n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334,
    n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343,
    n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352,
    n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
    n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370,
    n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379,
    n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388,
    n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397,
    n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406,
    n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415,
    n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424,
    n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
    n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442,
    n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451,
    n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460,
    n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469,
    n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478,
    n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487,
    n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496,
    n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
    n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514,
    n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
    n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532,
    n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541,
    n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550,
    n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559,
    n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568,
    n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
    n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586,
    n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595,
    n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604,
    n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613,
    n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622,
    n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631,
    n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640,
    n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
    n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658,
    n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667,
    n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676,
    n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685,
    n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694,
    n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703,
    n23704, n23705, n23706, n23707, n23708, n23709, n23711, n23712, n23713,
    n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722,
    n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731,
    n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740,
    n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749,
    n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758,
    n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767,
    n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776,
    n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
    n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794,
    n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803,
    n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812,
    n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821,
    n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830,
    n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839,
    n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848,
    n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
    n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866,
    n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
    n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884,
    n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893,
    n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902,
    n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911,
    n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920,
    n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
    n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938,
    n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
    n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956,
    n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965,
    n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974,
    n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983,
    n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992,
    n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
    n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010,
    n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019,
    n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028,
    n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037,
    n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046,
    n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055,
    n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064,
    n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
    n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082,
    n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091,
    n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100,
    n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109,
    n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118,
    n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127,
    n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136,
    n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
    n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154,
    n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163,
    n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172,
    n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181,
    n24182, n24183, n24184, n24185, n24186, n24187, n24189, n24190, n24191,
    n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200,
    n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
    n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218,
    n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227,
    n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236,
    n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245,
    n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254,
    n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263,
    n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272,
    n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
    n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290,
    n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
    n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308,
    n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317,
    n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326,
    n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335,
    n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344,
    n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
    n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362,
    n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
    n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380,
    n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389,
    n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398,
    n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407,
    n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416,
    n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
    n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434,
    n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
    n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452,
    n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461,
    n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470,
    n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479,
    n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488,
    n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
    n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506,
    n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515,
    n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524,
    n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533,
    n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542,
    n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551,
    n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560,
    n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
    n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578,
    n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587,
    n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596,
    n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605,
    n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614,
    n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623,
    n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632,
    n24633, n24634, n24635, n24636, n24637, n24639, n24640, n24641, n24642,
    n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651,
    n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660,
    n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669,
    n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678,
    n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687,
    n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696,
    n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
    n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714,
    n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723,
    n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732,
    n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741,
    n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750,
    n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759,
    n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768,
    n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
    n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786,
    n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795,
    n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804,
    n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813,
    n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822,
    n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831,
    n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840,
    n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
    n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858,
    n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867,
    n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876,
    n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885,
    n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894,
    n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903,
    n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912,
    n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
    n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930,
    n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939,
    n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948,
    n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957,
    n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966,
    n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975,
    n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984,
    n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
    n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002,
    n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011,
    n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020,
    n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029,
    n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038,
    n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047,
    n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056,
    n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
    n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074,
    n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083,
    n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092,
    n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101,
    n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110,
    n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119,
    n25120, n25121, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
    n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138,
    n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147,
    n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156,
    n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165,
    n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174,
    n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183,
    n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192,
    n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
    n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210,
    n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219,
    n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228,
    n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237,
    n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246,
    n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255,
    n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264,
    n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
    n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
    n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291,
    n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300,
    n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309,
    n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318,
    n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327,
    n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336,
    n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
    n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354,
    n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
    n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372,
    n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381,
    n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390,
    n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399,
    n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408,
    n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
    n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426,
    n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435,
    n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444,
    n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453,
    n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462,
    n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471,
    n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480,
    n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
    n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498,
    n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
    n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516,
    n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525,
    n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534,
    n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543,
    n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552,
    n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
    n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570,
    n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
    n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588,
    n25589, n25590, n25591, n25592, n25594, n25595, n25596, n25597, n25598,
    n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607,
    n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616,
    n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
    n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634,
    n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643,
    n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652,
    n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661,
    n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670,
    n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679,
    n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688,
    n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
    n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706,
    n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715,
    n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724,
    n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732, n25733,
    n25734, n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742,
    n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751,
    n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760,
    n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
    n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778,
    n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787,
    n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796,
    n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805,
    n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814,
    n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823,
    n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832,
    n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
    n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850,
    n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859,
    n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868,
    n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877,
    n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886,
    n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895,
    n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904,
    n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
    n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922,
    n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
    n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940,
    n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949,
    n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958,
    n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967,
    n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976,
    n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
    n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994,
    n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003,
    n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012,
    n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021,
    n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030,
    n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039,
    n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048,
    n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
    n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066,
    n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26076,
    n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085,
    n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094,
    n26095, n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103,
    n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112,
    n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
    n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130,
    n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139,
    n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148,
    n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157,
    n26158, n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166,
    n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175,
    n26176, n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184,
    n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
    n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202,
    n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211,
    n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220,
    n26221, n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229,
    n26230, n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238,
    n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247,
    n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256,
    n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
    n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274,
    n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283,
    n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292,
    n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301,
    n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310,
    n26311, n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319,
    n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328,
    n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
    n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346,
    n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355,
    n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364,
    n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373,
    n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26382,
    n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391,
    n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400,
    n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
    n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418,
    n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427,
    n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436,
    n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445,
    n26446, n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454,
    n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463,
    n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472,
    n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
    n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490,
    n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499,
    n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508,
    n26509, n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517,
    n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526,
    n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535,
    n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544,
    n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26553, n26554,
    n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563,
    n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572,
    n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581,
    n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590,
    n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599,
    n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608,
    n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
    n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626,
    n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635,
    n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644,
    n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653,
    n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661, n26662,
    n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671,
    n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680,
    n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
    n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698,
    n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707,
    n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716,
    n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725,
    n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734,
    n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743,
    n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752,
    n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
    n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770,
    n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779,
    n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788,
    n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797,
    n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806,
    n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815,
    n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824,
    n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
    n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
    n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851,
    n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860,
    n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869,
    n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878,
    n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887,
    n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896,
    n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
    n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914,
    n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923,
    n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932,
    n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941,
    n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950,
    n26951, n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959,
    n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968,
    n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
    n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986,
    n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995,
    n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004,
    n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013,
    n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022,
    n27023, n27024, n27025, n27026, n27027, n27028, n27030, n27031, n27032,
    n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
    n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050,
    n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059,
    n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068,
    n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077,
    n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086,
    n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095,
    n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104,
    n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
    n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122,
    n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131,
    n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140,
    n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149,
    n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27158,
    n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167,
    n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176,
    n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
    n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194,
    n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203,
    n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212,
    n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221,
    n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230,
    n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239,
    n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248,
    n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
    n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266,
    n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275,
    n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284,
    n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293,
    n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302,
    n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311,
    n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320,
    n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
    n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338,
    n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347,
    n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356,
    n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365,
    n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374,
    n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383,
    n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392,
    n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
    n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410,
    n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419,
    n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428,
    n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437,
    n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446,
    n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455,
    n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464,
    n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
    n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482,
    n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491,
    n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27501,
    n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510,
    n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519,
    n27520, n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528,
    n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
    n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546,
    n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555,
    n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564,
    n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573,
    n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582,
    n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591,
    n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600,
    n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
    n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618,
    n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627,
    n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636,
    n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645,
    n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654,
    n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663,
    n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672,
    n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
    n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690,
    n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699,
    n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708,
    n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717,
    n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726,
    n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734, n27735,
    n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743, n27744,
    n27745, n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
    n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762,
    n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771,
    n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780,
    n27781, n27782, n27783, n27784, n27785, n27786, n27787, n27788, n27789,
    n27790, n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798,
    n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806, n27807,
    n27808, n27809, n27810, n27811, n27812, n27813, n27814, n27815, n27816,
    n27817, n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
    n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834,
    n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843,
    n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852,
    n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860, n27861,
    n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870,
    n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879,
    n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887, n27888,
    n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
    n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906,
    n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915,
    n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924,
    n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933,
    n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942,
    n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950, n27951,
    n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959, n27960,
    n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
    n27970, n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979,
    n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988,
    n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997,
    n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006,
    n28007, n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015,
    n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024,
    n28025, n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
    n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042,
    n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051,
    n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060,
    n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069,
    n28070, n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078,
    n28079, n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087,
    n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095, n28096,
    n28097, n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
    n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114,
    n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123,
    n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132,
    n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141,
    n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149, n28150,
    n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159,
    n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167, n28168,
    n28169, n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
    n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186,
    n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195,
    n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204,
    n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213,
    n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222,
    n28223, n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231,
    n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239, n28240,
    n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
    n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258,
    n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267,
    n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276,
    n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285,
    n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294,
    n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303,
    n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312,
    n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
    n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330,
    n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339,
    n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348,
    n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357,
    n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366,
    n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375,
    n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384,
    n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
    n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402,
    n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411,
    n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420,
    n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429,
    n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438,
    n28439, n28440, n28441, n28443, n28444, n28445, n28446, n28447, n28448,
    n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
    n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466,
    n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475,
    n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484,
    n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493,
    n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28502,
    n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511,
    n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519, n28520,
    n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
    n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538,
    n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547,
    n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556,
    n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565,
    n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574,
    n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583,
    n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592,
    n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
    n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610,
    n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619,
    n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628,
    n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637,
    n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646,
    n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655,
    n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664,
    n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
    n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682,
    n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691,
    n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700,
    n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709,
    n28710, n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718,
    n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727,
    n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736,
    n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
    n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754,
    n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763,
    n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772,
    n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780, n28781,
    n28782, n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790,
    n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799,
    n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808,
    n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
    n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826,
    n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835,
    n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844,
    n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852, n28853,
    n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862,
    n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871,
    n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880,
    n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
    n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898,
    n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907,
    n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916,
    n28917, n28918, n28920, n28921, n28922, n28923, n28924, n28925, n28926,
    n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935,
    n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944,
    n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
    n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962,
    n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971,
    n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980,
    n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989,
    n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998,
    n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007,
    n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016,
    n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
    n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034,
    n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043,
    n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052,
    n29053, n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061,
    n29062, n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070,
    n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079,
    n29080, n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088,
    n29089, n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
    n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106,
    n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115,
    n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124,
    n29125, n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133,
    n29134, n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142,
    n29143, n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151,
    n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160,
    n29161, n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
    n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178,
    n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187,
    n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196,
    n29197, n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205,
    n29206, n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214,
    n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223,
    n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232,
    n29233, n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
    n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250,
    n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259,
    n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267, n29268,
    n29269, n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29277,
    n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286,
    n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295,
    n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304,
    n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
    n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322,
    n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331,
    n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340,
    n29341, n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349,
    n29350, n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358,
    n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367,
    n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376,
    n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
    n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29395,
    n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404,
    n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413,
    n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422,
    n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431,
    n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440,
    n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
    n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458,
    n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467,
    n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476,
    n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485,
    n29486, n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494,
    n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503,
    n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512,
    n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
    n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530,
    n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539,
    n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548,
    n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557,
    n29558, n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566,
    n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575,
    n29576, n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584,
    n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
    n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602,
    n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611,
    n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620,
    n29621, n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629,
    n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638,
    n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647,
    n29648, n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656,
    n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
    n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674,
    n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683,
    n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692,
    n29693, n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701,
    n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710,
    n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719,
    n29720, n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728,
    n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
    n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746,
    n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755,
    n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763, n29764,
    n29765, n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773,
    n29774, n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782,
    n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791,
    n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800,
    n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
    n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818,
    n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827,
    n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836,
    n29837, n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845,
    n29846, n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854,
    n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863,
    n29864, n29865, n29866, n29867, n29868, n29870, n29871, n29872, n29873,
    n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881, n29882,
    n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891,
    n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899, n29900,
    n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908, n29909,
    n29910, n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918,
    n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926, n29927,
    n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29936,
    n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
    n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954,
    n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963,
    n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971, n29972,
    n29973, n29974, n29975, n29976, n29977, n29978, n29979, n29980, n29981,
    n29982, n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990,
    n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999,
    n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008,
    n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
    n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026,
    n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035,
    n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043, n30044,
    n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052, n30053,
    n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062,
    n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070, n30071,
    n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080,
    n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
    n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098,
    n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107,
    n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115, n30116,
    n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124, n30125,
    n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134,
    n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142, n30143,
    n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151, n30152,
    n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
    n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170,
    n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179,
    n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187, n30188,
    n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196, n30197,
    n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206,
    n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214, n30215,
    n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223, n30224,
    n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
    n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241, n30242,
    n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251,
    n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259, n30260,
    n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268, n30269,
    n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278,
    n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286, n30287,
    n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296,
    n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
    n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313, n30314,
    n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323,
    n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331, n30332,
    n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340, n30341,
    n30342, n30343, n30345, n30346, n30347, n30348, n30349, n30350, n30351,
    n30352, n30353, n30354, n30355, n30356, n30357, n30358, n30359, n30360,
    n30361, n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
    n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377, n30378,
    n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387,
    n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395, n30396,
    n30397, n30398, n30399, n30400, n30401, n30402, n30403, n30404, n30405,
    n30406, n30407, n30408, n30409, n30410, n30411, n30412, n30413, n30414,
    n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422, n30423,
    n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431, n30432,
    n30433, n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
    n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449, n30450,
    n30451, n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459,
    n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467, n30468,
    n30469, n30470, n30471, n30472, n30473, n30474, n30475, n30476, n30477,
    n30478, n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486,
    n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494, n30495,
    n30496, n30497, n30498, n30499, n30500, n30501, n30502, n30503, n30504,
    n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
    n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521, n30522,
    n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531,
    n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539, n30540,
    n30541, n30542, n30543, n30544, n30545, n30546, n30547, n30548, n30549,
    n30550, n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558,
    n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567,
    n30568, n30569, n30570, n30571, n30572, n30573, n30574, n30575, n30576,
    n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
    n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593, n30594,
    n30595, n30596, n30597, n30598, n30599, n30600, n30601, n30602, n30603,
    n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611, n30612,
    n30613, n30614, n30615, n30616, n30617, n30618, n30619, n30620, n30621,
    n30622, n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630,
    n30631, n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639,
    n30640, n30641, n30642, n30643, n30644, n30645, n30646, n30647, n30648,
    n30649, n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
    n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665, n30666,
    n30667, n30668, n30669, n30670, n30671, n30672, n30673, n30674, n30675,
    n30676, n30677, n30678, n30679, n30680, n30681, n30682, n30683, n30684,
    n30685, n30686, n30687, n30688, n30689, n30690, n30691, n30692, n30693,
    n30694, n30695, n30696, n30697, n30698, n30699, n30700, n30701, n30702,
    n30703, n30704, n30705, n30706, n30707, n30708, n30709, n30710, n30711,
    n30712, n30713, n30714, n30715, n30716, n30717, n30718, n30719, n30720,
    n30721, n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
    n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737, n30738,
    n30739, n30740, n30741, n30742, n30743, n30744, n30745, n30746, n30747,
    n30748, n30749, n30750, n30751, n30752, n30753, n30754, n30755, n30756,
    n30757, n30758, n30759, n30760, n30761, n30762, n30763, n30764, n30765,
    n30766, n30767, n30768, n30769, n30770, n30771, n30772, n30773, n30774,
    n30775, n30776, n30777, n30778, n30779, n30780, n30781, n30782, n30783,
    n30784, n30785, n30786, n30787, n30788, n30789, n30790, n30791, n30792,
    n30793, n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
    n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809, n30810,
    n30811, n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819,
    n30820, n30821, n30822, n30824, n30825, n30826, n30827, n30828, n30829,
    n30830, n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838,
    n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847,
    n30848, n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856,
    n30857, n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
    n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874,
    n30875, n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883,
    n30884, n30885, n30886, n30887, n30888, n30889, n30890, n30891, n30892,
    n30893, n30894, n30895, n30896, n30897, n30898, n30899, n30900, n30901,
    n30902, n30903, n30904, n30905, n30906, n30907, n30908, n30909, n30910,
    n30911, n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919,
    n30920, n30921, n30922, n30923, n30924, n30925, n30926, n30927, n30928,
    n30929, n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
    n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945, n30946,
    n30947, n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955,
    n30956, n30957, n30958, n30959, n30960, n30961, n30962, n30963, n30964,
    n30965, n30966, n30967, n30968, n30969, n30970, n30971, n30972, n30973,
    n30974, n30975, n30976, n30977, n30978, n30979, n30980, n30981, n30982,
    n30983, n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991,
    n30992, n30993, n30994, n30995, n30996, n30997, n30998, n30999, n31000,
    n31001, n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
    n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017, n31018,
    n31019, n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027,
    n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035, n31036,
    n31037, n31038, n31039, n31040, n31041, n31042, n31043, n31044, n31045,
    n31046, n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054,
    n31055, n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063,
    n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072,
    n31073, n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
    n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089, n31090,
    n31091, n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099,
    n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107, n31108,
    n31109, n31110, n31111, n31112, n31113, n31114, n31115, n31116, n31117,
    n31118, n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126,
    n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135,
    n31136, n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144,
    n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
    n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162,
    n31163, n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171,
    n31172, n31173, n31174, n31175, n31176, n31177, n31178, n31179, n31180,
    n31181, n31182, n31183, n31184, n31185, n31186, n31187, n31188, n31189,
    n31190, n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198,
    n31199, n31200, n31201, n31202, n31203, n31204, n31205, n31206, n31207,
    n31208, n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216,
    n31217, n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
    n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233, n31234,
    n31235, n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243,
    n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251, n31252,
    n31253, n31254, n31255, n31256, n31257, n31258, n31259, n31260, n31261,
    n31262, n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270,
    n31271, n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279,
    n31280, n31281, n31282, n31283, n31284, n31285, n31286, n31287, n31288,
    n31289, n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
    n31298, n31299, n31301, n31302, n31303, n31304, n31305, n31306, n31307,
    n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315, n31316,
    n31317, n31318, n31319, n31320, n31321, n31322, n31323, n31324, n31325,
    n31326, n31327, n31328, n31329, n31330, n31331, n31332, n31333, n31334,
    n31335, n31336, n31337, n31338, n31339, n31340, n31341, n31342, n31343,
    n31344, n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352,
    n31353, n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
    n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370,
    n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378, n31379,
    n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387, n31388,
    n31389, n31390, n31391, n31392, n31393, n31394, n31395, n31396, n31397,
    n31398, n31399, n31400, n31401, n31402, n31403, n31404, n31405, n31406,
    n31407, n31408, n31409, n31410, n31411, n31412, n31413, n31414, n31415,
    n31416, n31417, n31418, n31419, n31420, n31421, n31422, n31423, n31424,
    n31425, n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
    n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441, n31442,
    n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450, n31451,
    n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459, n31460,
    n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468, n31469,
    n31470, n31471, n31472, n31473, n31474, n31475, n31476, n31477, n31478,
    n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486, n31487,
    n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495, n31496,
    n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
    n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514,
    n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523,
    n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531, n31532,
    n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31540, n31541,
    n31542, n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550,
    n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558, n31559,
    n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567, n31568,
    n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
    n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585, n31586,
    n31587, n31588, n31589, n31590, n31591, n31592, n31593, n31594, n31595,
    n31596, n31597, n31598, n31599, n31600, n31601, n31602, n31603, n31604,
    n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612, n31613,
    n31614, n31615, n31616, n31617, n31618, n31619, n31620, n31621, n31622,
    n31623, n31624, n31625, n31626, n31627, n31628, n31629, n31630, n31631,
    n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639, n31640,
    n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
    n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657, n31658,
    n31659, n31660, n31661, n31662, n31663, n31664, n31665, n31666, n31667,
    n31668, n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676,
    n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684, n31685,
    n31686, n31687, n31688, n31689, n31690, n31691, n31692, n31693, n31694,
    n31695, n31696, n31697, n31698, n31699, n31700, n31701, n31702, n31703,
    n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711, n31712,
    n31713, n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
    n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729, n31730,
    n31731, n31732, n31733, n31734, n31735, n31736, n31737, n31738, n31739,
    n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747, n31748,
    n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756, n31757,
    n31758, n31759, n31760, n31761, n31762, n31763, n31764, n31765, n31766,
    n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774, n31775,
    n31776, n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
    n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793, n31794,
    n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802, n31803,
    n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811, n31812,
    n31813, n31814, n31815, n31816, n31817, n31818, n31819, n31820, n31821,
    n31822, n31823, n31824, n31825, n31826, n31827, n31828, n31829, n31830,
    n31831, n31832, n31833, n31834, n31835, n31836, n31837, n31838, n31839,
    n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847, n31848,
    n31849, n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
    n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865, n31866,
    n31867, n31868, n31869, n31870, n31871, n31872, n31873, n31874, n31875,
    n31876, n31877, n31878, n31879, n31880, n31881, n31882, n31883, n31884,
    n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892, n31893,
    n31894, n31895, n31896, n31897, n31898, n31899, n31900, n31901, n31902,
    n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910, n31911,
    n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919, n31920,
    n31921, n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
    n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937, n31938,
    n31939, n31940, n31941, n31942, n31943, n31944, n31945, n31946, n31947,
    n31948, n31949, n31950, n31951, n31952, n31953, n31954, n31955, n31956,
    n31957, n31958, n31959, n31960, n31961, n31962, n31963, n31964, n31965,
    n31966, n31967, n31968, n31969, n31970, n31971, n31972, n31973, n31974,
    n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982, n31983,
    n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991, n31992,
    n31993, n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
    n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009, n32010,
    n32011, n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019,
    n32020, n32021, n32022, n32023, n32024, n32025, n32026, n32027, n32028,
    n32029, n32030, n32031, n32032, n32033, n32034, n32035, n32036, n32037,
    n32038, n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046,
    n32047, n32048, n32049, n32050, n32051, n32052, n32053, n32054, n32055,
    n32056, n32057, n32058, n32059, n32060, n32061, n32062, n32063, n32064,
    n32065, n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
    n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081, n32082,
    n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090, n32091,
    n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099, n32100,
    n32101, n32102, n32103, n32104, n32105, n32106, n32107, n32108, n32109,
    n32110, n32111, n32112, n32113, n32114, n32115, n32116, n32117, n32118,
    n32119, n32120, n32121, n32122, n32123, n32124, n32125, n32126, n32127,
    n32128, n32129, n32130, n32131, n32132, n32133, n32134, n32135, n32136,
    n32137, n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
    n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154,
    n32155, n32156, n32157, n32158, n32159, n32160, n32161, n32162, n32163,
    n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32171, n32172,
    n32173, n32174, n32175, n32176, n32177, n32178, n32179, n32180, n32181,
    n32182, n32183, n32184, n32185, n32186, n32187, n32188, n32189, n32190,
    n32191, n32192, n32193, n32194, n32195, n32196, n32197, n32198, n32199,
    n32200, n32201, n32202, n32203, n32204, n32205, n32206, n32207, n32208,
    n32209, n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
    n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225, n32226,
    n32227, n32228, n32229, n32230, n32231, n32232, n32233, n32234, n32235,
    n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243, n32244,
    n32245, n32246, n32247, n32248, n32249, n32250, n32251, n32252, n32253,
    n32255, n32256, n32257, n32258, n32259, n32260, n32261, n32262, n32263,
    n32264, n32265, n32266, n32267, n32268, n32269, n32270, n32271, n32272,
    n32273, n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
    n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289, n32290,
    n32291, n32292, n32293, n32294, n32295, n32296, n32297, n32298, n32299,
    n32300, n32301, n32302, n32303, n32304, n32305, n32306, n32307, n32308,
    n32309, n32310, n32311, n32312, n32313, n32314, n32315, n32316, n32317,
    n32318, n32319, n32320, n32321, n32322, n32323, n32324, n32325, n32326,
    n32327, n32328, n32329, n32330, n32331, n32332, n32333, n32334, n32335,
    n32336, n32337, n32338, n32339, n32340, n32341, n32342, n32343, n32344,
    n32345, n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
    n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362,
    n32363, n32364, n32365, n32366, n32367, n32368, n32369, n32370, n32371,
    n32372, n32373, n32374, n32375, n32376, n32377, n32378, n32379, n32380,
    n32381, n32382, n32383, n32384, n32385, n32386, n32387, n32388, n32389,
    n32390, n32391, n32392, n32393, n32394, n32395, n32396, n32397, n32398,
    n32399, n32400, n32401, n32402, n32403, n32404, n32405, n32406, n32407,
    n32408, n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416,
    n32417, n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
    n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433, n32434,
    n32435, n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443,
    n32444, n32445, n32446, n32447, n32448, n32449, n32450, n32451, n32452,
    n32453, n32454, n32455, n32456, n32457, n32458, n32459, n32460, n32461,
    n32462, n32463, n32464, n32465, n32466, n32467, n32468, n32469, n32470,
    n32471, n32472, n32473, n32474, n32475, n32476, n32477, n32478, n32479,
    n32480, n32481, n32482, n32483, n32484, n32485, n32486, n32487, n32488,
    n32489, n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
    n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505, n32506,
    n32507, n32508, n32509, n32510, n32511, n32512, n32513, n32514, n32515,
    n32516, n32517, n32518, n32519, n32520, n32521, n32522, n32523, n32524,
    n32525, n32526, n32527, n32528, n32529, n32530, n32531, n32532, n32533,
    n32534, n32535, n32536, n32537, n32538, n32539, n32540, n32541, n32542,
    n32543, n32544, n32545, n32546, n32547, n32548, n32549, n32550, n32551,
    n32552, n32553, n32554, n32555, n32556, n32557, n32558, n32559, n32560,
    n32561, n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
    n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577, n32578,
    n32579, n32580, n32581, n32582, n32583, n32584, n32585, n32586, n32587,
    n32588, n32589, n32590, n32591, n32592, n32593, n32594, n32595, n32596,
    n32597, n32598, n32599, n32600, n32601, n32602, n32603, n32604, n32605,
    n32606, n32607, n32608, n32609, n32610, n32611, n32612, n32613, n32614,
    n32615, n32616, n32617, n32618, n32619, n32620, n32621, n32622, n32623,
    n32624, n32625, n32626, n32627, n32628, n32629, n32630, n32631, n32632,
    n32633, n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
    n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649, n32650,
    n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32658, n32659,
    n32660, n32661, n32662, n32663, n32664, n32665, n32666, n32667, n32668,
    n32669, n32670, n32671, n32672, n32673, n32674, n32675, n32676, n32677,
    n32678, n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686,
    n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694, n32695,
    n32696, n32697, n32698, n32699, n32700, n32701, n32702, n32703, n32704,
    n32705, n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
    n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722,
    n32723, n32724, n32725, n32727, n32728, n32729, n32730, n32731, n32732,
    n32733, n32734, n32735, n32736, n32737, n32738, n32739, n32740, n32741,
    n32742, n32743, n32744, n32745, n32746, n32747, n32748, n32749, n32750,
    n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758, n32759,
    n32760, n32761, n32762, n32763, n32764, n32765, n32766, n32767, n32768,
    n32769, n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
    n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785, n32786,
    n32787, n32788, n32789, n32790, n32791, n32792, n32793, n32794, n32795,
    n32796, n32797, n32798, n32799, n32800, n32801, n32802, n32803, n32804,
    n32805, n32806, n32807, n32808, n32809, n32810, n32811, n32812, n32813,
    n32814, n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822,
    n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830, n32831,
    n32832, n32833, n32834, n32835, n32836, n32837, n32838, n32839, n32840,
    n32841, n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
    n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857, n32858,
    n32859, n32860, n32861, n32862, n32863, n32864, n32865, n32866, n32867,
    n32868, n32869, n32870, n32871, n32872, n32873, n32874, n32875, n32876,
    n32877, n32878, n32879, n32880, n32881, n32882, n32883, n32884, n32885,
    n32886, n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894,
    n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902, n32903,
    n32904, n32905, n32906, n32907, n32908, n32909, n32910, n32911, n32912,
    n32913, n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
    n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930,
    n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938, n32939,
    n32940, n32941, n32942, n32943, n32944, n32945, n32946, n32947, n32948,
    n32949, n32950, n32951, n32952, n32953, n32954, n32955, n32956, n32957,
    n32958, n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966,
    n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974, n32975,
    n32976, n32977, n32978, n32979, n32980, n32981, n32982, n32983, n32984,
    n32985, n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
    n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001, n33002,
    n33003, n33004, n33005, n33006, n33007, n33008, n33009, n33010, n33011,
    n33012, n33013, n33014, n33015, n33016, n33017, n33018, n33019, n33020,
    n33021, n33022, n33023, n33024, n33025, n33026, n33027, n33028, n33029,
    n33030, n33031, n33032, n33033, n33034, n33035, n33036, n33037, n33038,
    n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046, n33047,
    n33048, n33049, n33050, n33051, n33052, n33053, n33054, n33055, n33056,
    n33057, n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
    n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073, n33074,
    n33075, n33076, n33077, n33078, n33079, n33080, n33081, n33082, n33083,
    n33084, n33085, n33086, n33087, n33088, n33089, n33090, n33091, n33092,
    n33093, n33094, n33095, n33096, n33097, n33098, n33099, n33100, n33101,
    n33102, n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110,
    n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118, n33119,
    n33120, n33121, n33122, n33123, n33124, n33125, n33126, n33127, n33128,
    n33129, n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
    n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145, n33146,
    n33147, n33148, n33149, n33150, n33151, n33152, n33153, n33154, n33155,
    n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163, n33164,
    n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172, n33173,
    n33174, n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182,
    n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190, n33191,
    n33192, n33193, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
    n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209, n33210,
    n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219,
    n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228,
    n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236, n33237,
    n33238, n33239, n33240, n33241, n33242, n33243, n33245, n33246, n33247,
    n33248, n33249, n33250, n33251, n33252, n33253, n33254, n33255, n33256,
    n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
    n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274,
    n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283,
    n33284, n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292,
    n33293, n33294, n33295, n33296, n33297, n33298, n33299, n33300, n33301,
    n33302, n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310,
    n33311, n33312, n33314, n33315, n33316, n33317, n33318, n33319, n33320,
    n33321, n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
    n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337, n33338,
    n33339, n33340, n33341, n33342, n33343, n33344, n33345, n33346, n33347,
    n33348, n33349, n33350, n33351, n33352, n33353, n33354, n33355, n33356,
    n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364, n33365,
    n33366, n33367, n33368, n33369, n33370, n33371, n33372, n33373, n33375,
    n33376, n33377, n33378, n33379, n33380, n33381, n33382, n33383, n33384,
    n33385, n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
    n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401, n33402,
    n33403, n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411,
    n33412, n33413, n33414, n33415, n33416, n33417, n33418, n33419, n33420,
    n33421, n33422, n33423, n33424, n33425, n33426, n33427, n33428, n33429,
    n33430, n33431, n33432, n33433, n33434, n33435, n33436, n33437, n33438,
    n33439, n33440, n33441, n33442, n33443, n33444, n33445, n33446, n33447,
    n33448, n33449, n33450, n33451, n33452, n33453, n33454, n33455, n33456,
    n33457, n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
    n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473, n33474,
    n33475, n33476, n33477, n33478, n33479, n33480, n33481, n33482, n33483,
    n33484, n33485, n33486, n33487, n33488, n33489, n33490, n33491, n33492,
    n33493, n33494, n33495, n33496, n33497, n33498, n33499, n33500, n33501,
    n33502, n33503, n33504, n33505, n33506, n33507, n33508, n33509, n33510,
    n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33518, n33519,
    n33520, n33521, n33522, n33523, n33524, n33525, n33526, n33527, n33528,
    n33529, n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
    n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545, n33546,
    n33547, n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555,
    n33556, n33557, n33558, n33559, n33560, n33561, n33562, n33563, n33564,
    n33565, n33566, n33567, n33568, n33569, n33570, n33571, n33572, n33573,
    n33574, n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582,
    n33583, n33584, n33585, n33586, n33587, n33588, n33589, n33590, n33591,
    n33592, n33593, n33594, n33595, n33596, n33597, n33598, n33599, n33600,
    n33601, n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
    n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617, n33618,
    n33619, n33620, n33621, n33622, n33623, n33624, n33625, n33626, n33627,
    n33628, n33629, n33630, n33631, n33632, n33633, n33634, n33635, n33636,
    n33637, n33638, n33639, n33640, n33641, n33642, n33643, n33644, n33645,
    n33646, n33647, n33648, n33649, n33650, n33651, n33652, n33653, n33654,
    n33655, n33656, n33657, n33658, n33659, n33660, n33661, n33662, n33663,
    n33664, n33665, n33666, n33667, n33668, n33669, n33670, n33671, n33672,
    n33673, n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
    n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689, n33690,
    n33691, n33692, n33693, n33694, n33695, n33696, n33697, n33698, n33699,
    n33700, n33701, n33702, n33703, n33704, n33705, n33706, n33707, n33708,
    n33709, n33710, n33711, n33712, n33713, n33714, n33715, n33716, n33717,
    n33718, n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726,
    n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734, n33735,
    n33736, n33737, n33738, n33739, n33740, n33741, n33742, n33743, n33744,
    n33745, n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
    n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761, n33762,
    n33763, n33764, n33765, n33766, n33767, n33768, n33769, n33770, n33771,
    n33772, n33773, n33774, n33775, n33776, n33777, n33778, n33779, n33780,
    n33781, n33782, n33783, n33784, n33785, n33786, n33787, n33788, n33789,
    n33790, n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798,
    n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806, n33807,
    n33808, n33809, n33810, n33811, n33812, n33813, n33814, n33815, n33816,
    n33817, n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
    n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833, n33834,
    n33835, n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843,
    n33844, n33845, n33846, n33847, n33848, n33849, n33850, n33851, n33852,
    n33853, n33854, n33855, n33856, n33857, n33858, n33859, n33860, n33861,
    n33862, n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870,
    n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878, n33879,
    n33880, n33881, n33882, n33883, n33884, n33885, n33886, n33887, n33888,
    n33889, n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
    n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905, n33906,
    n33907, n33908, n33909, n33910, n33911, n33912, n33913, n33914, n33915,
    n33916, n33917, n33918, n33919, n33920, n33921, n33922, n33923, n33924,
    n33925, n33926, n33927, n33928, n33929, n33930, n33931, n33932, n33933,
    n33934, n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942,
    n33943, n33944, n33945, n33946, n33947, n33948, n33949, n33950, n33951,
    n33952, n33953, n33954, n33955, n33956, n33957, n33958, n33959, n33960,
    n33961, n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
    n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977, n33978,
    n33979, n33980, n33981, n33982, n33983, n33984, n33985, n33986, n33987,
    n33988, n33989, n33990, n33991, n33992, n33993, n33994, n33995, n33996,
    n33997, n33998, n33999, n34000, n34001, n34002, n34003, n34004, n34005,
    n34006, n34007, n34008, n34009, n34011, n34012, n34013, n34014, n34015,
    n34016, n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024,
    n34025, n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
    n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042,
    n34043, n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051,
    n34052, n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060,
    n34061, n34062, n34063, n34064, n34065, n34066, n34067, n34068, n34069,
    n34070, n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078,
    n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086, n34087,
    n34088, n34089, n34090, n34091, n34092, n34093, n34094, n34095, n34096,
    n34097, n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
    n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113, n34114,
    n34115, n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123,
    n34124, n34125, n34126, n34127, n34128, n34129, n34130, n34131, n34132,
    n34133, n34134, n34135, n34136, n34137, n34138, n34139, n34140, n34141,
    n34142, n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150,
    n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158, n34159,
    n34160, n34161, n34162, n34163, n34164, n34165, n34166, n34167, n34168,
    n34169, n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
    n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185, n34186,
    n34187, n34188, n34189, n34190, n34191, n34192, n34193, n34194, n34195,
    n34196, n34197, n34198, n34199, n34200, n34201, n34202, n34203, n34204,
    n34205, n34206, n34207, n34208, n34209, n34210, n34211, n34212, n34213,
    n34214, n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222,
    n34223, n34224, n34225, n34226, n34227, n34228, n34229, n34230, n34231,
    n34232, n34233, n34234, n34235, n34236, n34237, n34238, n34239, n34240,
    n34241, n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
    n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257, n34258,
    n34259, n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267,
    n34268, n34269, n34270, n34271, n34272, n34273, n34274, n34275, n34276,
    n34277, n34278, n34279, n34280, n34281, n34282, n34283, n34284, n34285,
    n34286, n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294,
    n34295, n34296, n34297, n34298, n34299, n34300, n34302, n34303, n34304,
    n34305, n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
    n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321, n34322,
    n34323, n34324, n34325, n34326, n34327, n34328, n34329, n34330, n34331,
    n34332, n34333, n34334, n34335, n34336, n34337, n34338, n34339, n34340,
    n34341, n34342, n34343, n34344, n34345, n34346, n34347, n34348, n34349,
    n34350, n34351, n34352, n34353, n34354, n34355, n34356, n34357, n34358,
    n34359, n34360, n34361, n34362, n34363, n34364, n34365, n34366, n34367,
    n34368, n34369, n34370, n34371, n34372, n34373, n34374, n34375, n34376,
    n34377, n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
    n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393, n34394,
    n34395, n34396, n34397, n34398, n34399, n34400, n34401, n34402, n34403,
    n34404, n34405, n34406, n34407, n34408, n34409, n34410, n34411, n34412,
    n34413, n34414, n34415, n34416, n34417, n34418, n34419, n34420, n34421,
    n34422, n34423, n34424, n34425, n34426, n34427, n34428, n34429, n34430,
    n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438, n34439,
    n34440, n34441, n34442, n34443, n34444, n34445, n34446, n34447, n34448,
    n34449, n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
    n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465, n34466,
    n34467, n34468, n34469, n34470, n34471, n34472, n34473, n34474, n34475,
    n34476, n34477, n34478, n34479, n34480, n34481, n34482, n34483, n34484,
    n34485, n34486, n34487, n34488, n34489, n34490, n34491, n34492, n34493,
    n34494, n34495, n34496, n34497, n34498, n34499, n34500, n34501, n34502,
    n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510, n34511,
    n34512, n34513, n34514, n34515, n34516, n34517, n34518, n34519, n34520,
    n34521, n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
    n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537, n34538,
    n34539, n34540, n34541, n34542, n34543, n34544, n34545, n34546, n34547,
    n34548, n34549, n34550, n34551, n34552, n34553, n34554, n34555, n34556,
    n34557, n34558, n34559, n34560, n34561, n34562, n34563, n34564, n34565,
    n34566, n34567, n34568, n34569, n34570, n34571, n34572, n34573, n34574,
    n34575, n34576, n34577, n34578, n34579, n34580, n34581, n34583, n34584,
    n34585, n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
    n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601, n34602,
    n34603, n34604, n34605, n34606, n34607, n34608, n34609, n34610, n34611,
    n34612, n34613, n34614, n34615, n34616, n34617, n34618, n34619, n34620,
    n34621, n34622, n34623, n34624, n34625, n34626, n34627, n34628, n34629,
    n34630, n34631, n34632, n34633, n34634, n34635, n34636, n34637, n34638,
    n34639, n34640, n34641, n34642, n34643, n34644, n34645, n34646, n34647,
    n34648, n34649, n34650, n34651, n34652, n34653, n34654, n34655, n34656,
    n34657, n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
    n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673, n34674,
    n34675, n34676, n34677, n34678, n34679, n34680, n34681, n34682, n34683,
    n34684, n34685, n34686, n34687, n34688, n34689, n34690, n34691, n34692,
    n34693, n34694, n34695, n34696, n34697, n34698, n34699, n34700, n34701,
    n34702, n34703, n34704, n34705, n34706, n34707, n34708, n34709, n34710,
    n34711, n34712, n34713, n34714, n34715, n34716, n34717, n34718, n34719,
    n34720, n34721, n34722, n34723, n34724, n34725, n34726, n34727, n34728,
    n34729, n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
    n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745, n34746,
    n34747, n34748, n34749, n34750, n34751, n34752, n34753, n34754, n34755,
    n34756, n34757, n34758, n34759, n34760, n34761, n34762, n34763, n34764,
    n34765, n34766, n34767, n34768, n34769, n34770, n34771, n34772, n34773,
    n34774, n34775, n34776, n34778, n34779, n34780, n34781, n34782, n34783,
    n34784, n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34794,
    n34795, n34796, n34797, n34798, n34799, n34800, n34801, n34802, n34803,
    n34804, n34805, n34806, n34807, n34808, n34809, n34810, n34811, n34812,
    n34813, n34814, n34815, n34816, n34817, n34818, n34819, n34820, n34821,
    n34822, n34823, n34824, n34825, n34826, n34827, n34828, n34829, n34830,
    n34831, n34832, n34833, n34834, n34835, n34836, n34837, n34838, n34839,
    n34840, n34841, n34842, n34843, n34844, n34845, n34846, n34847, n34848,
    n34849, n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
    n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865, n34866,
    n34867, n34868, n34869, n34870, n34871, n34872, n34873, n34874, n34875,
    n34876, n34877, n34878, n34879, n34880, n34881, n34882, n34883, n34884,
    n34885, n34886, n34887, n34888, n34889, n34890, n34891, n34892, n34893,
    n34894, n34895, n34896, n34897, n34898, n34899, n34900, n34901, n34903,
    n34904, n34905, n34906, n34907, n34908, n34910, n34911, n34912, n34913,
    n34914, n34915, n34916, n34918, n34919, n34920, n34921, n34922, n34923,
    n34924, n34925, n34926, n34927, n34928, n34929, n34930, n34931, n34932,
    n34933, n34934, n34935, n34936, n34937, n34938, n34939, n34940, n34941,
    n34942, n34943, n34944, n34945, n34946, n34947, n34948, n34949, n34950,
    n34951, n34952, n34953, n34954, n34955, n34956, n34957, n34958, n34959,
    n34960, n34961, n34962, n34963, n34964, n34965, n34966, n34967, n34968,
    n34969, n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
    n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985, n34986,
    n34987, n34988, n34989, n34990, n34991, n34992, n34993, n34994, n34995,
    n34996, n34997, n34998, n34999, n35000, n35001, n35002, n35003, n35004,
    n35005, n35006, n35007, n35008, n35009, n35010, n35011, n35012, n35013,
    n35014, n35015, n35016, n35017, n35018, n35019, n35020, n35021, n35022,
    n35023, n35024, n35025, n35026, n35027, n35028, n35029, n35030, n35031,
    n35032, n35033, n35034, n35035, n35036, n35037, n35038, n35039, n35040,
    n35041, n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
    n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057, n35058,
    n35059, n35060, n35061, n35062, n35063, n35064, n35065, n35066, n35067,
    n35068, n35069, n35070, n35071, n35072, n35073, n35074, n35075, n35076,
    n35077, n35078, n35079, n35080, n35081, n35082, n35083, n35084, n35085,
    n35086, n35087, n35088, n35089, n35090, n35091, n35092, n35093, n35094,
    n35095, n35096, n35097, n35098, n35099, n35100, n35101, n35102, n35103,
    n35104, n35105, n35106, n35107, n35108, n35109, n35110, n35111, n35112,
    n35113, n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
    n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129, n35130,
    n35131, n35132, n35133, n35134, n35135, n35136, n35137, n35138, n35139,
    n35140, n35141, n35142, n35143, n35144, n35145, n35146, n35147, n35148,
    n35149, n35150, n35151, n35152, n35153, n35154, n35155, n35156, n35157,
    n35158, n35159, n35160, n35161, n35162, n35163, n35164, n35165, n35166,
    n35167, n35168, n35169, n35170, n35171, n35172, n35173, n35174, n35175,
    n35176, n35177, n35178, n35179, n35180, n35181, n35182, n35183, n35184,
    n35185, n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
    n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201, n35202,
    n35203, n35204, n35205, n35206, n35207, n35208, n35209, n35210, n35211,
    n35212, n35213, n35214, n35215, n35216, n35217, n35218, n35219, n35220,
    n35221, n35222, n35223, n35224, n35225, n35226, n35227, n35228, n35229,
    n35230, n35231, n35232, n35233, n35234, n35235, n35236, n35237, n35238,
    n35239, n35240, n35241, n35242, n35243, n35244, n35245, n35246, n35247,
    n35248, n35249, n35250, n35251, n35252, n35253, n35254, n35255, n35256,
    n35257, n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
    n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273, n35274,
    n35275, n35276, n35277, n35278, n35279, n35280, n35281, n35282, n35283,
    n35284, n35285, n35286, n35287, n35288, n35289, n35290, n35291, n35292,
    n35293, n35294, n35295, n35296, n35297, n35298, n35299, n35300, n35301,
    n35302, n35303, n35304, n35305, n35306, n35307, n35308, n35309, n35310,
    n35311, n35312, n35313, n35314, n35315, n35316, n35317, n35318, n35319,
    n35320, n35321, n35322, n35323, n35324, n35325, n35326, n35327, n35328,
    n35329, n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
    n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345, n35346,
    n35347, n35348, n35349, n35350, n35351, n35352, n35353, n35354, n35355,
    n35356, n35357, n35358, n35359, n35360, n35361, n35362, n35363, n35364,
    n35365, n35366, n35367, n35368, n35369, n35370, n35371, n35372, n35373,
    n35374, n35375, n35376, n35377, n35378, n35379, n35380, n35381, n35382,
    n35383, n35384, n35385, n35386, n35387, n35388, n35389, n35390, n35391,
    n35392, n35393, n35394, n35395, n35396, n35397, n35398, n35399, n35400,
    n35401, n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35410,
    n35411, n35412, n35413, n35414, n35415, n35416, n35417, n35418, n35419,
    n35420, n35421, n35422, n35423, n35424, n35425, n35426, n35427, n35428,
    n35429, n35430, n35431, n35432, n35433, n35434, n35435, n35436, n35437,
    n35438, n35439, n35440, n35441, n35442, n35443, n35444, n35445, n35446,
    n35447, n35448, n35449, n35450, n35451, n35452, n35453, n35454, n35455,
    n35456, n35457, n35458, n35459, n35460, n35461, n35462, n35463, n35464,
    n35465, n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
    n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481, n35482,
    n35483, n35485, n35486, n35487, n35488, n35489, n35490, n35491, n35492,
    n35493, n35494, n35495, n35496, n35497, n35498, n35499, n35500, n35501,
    n35502, n35503, n35504, n35505, n35506, n35507, n35508, n35509, n35510,
    n35511, n35512, n35513, n35514, n35515, n35516, n35517, n35518, n35519,
    n35520, n35521, n35522, n35523, n35524, n35525, n35526, n35527, n35528,
    n35529, n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
    n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545, n35546,
    n35547, n35548, n35549, n35550, n35551, n35552, n35553, n35554, n35555,
    n35556, n35557, n35558, n35559, n35560, n35561, n35562, n35563, n35564,
    n35565, n35566, n35567, n35568, n35569, n35570, n35571, n35572, n35573,
    n35574, n35575, n35576, n35577, n35578, n35579, n35580, n35581, n35582,
    n35583, n35584, n35585, n35586, n35587, n35588, n35589, n35590, n35591,
    n35592, n35593, n35594, n35595, n35596, n35597, n35598, n35599, n35600,
    n35601, n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
    n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617, n35618,
    n35619, n35620, n35621, n35622, n35623, n35624, n35625, n35626, n35627,
    n35628, n35629, n35630, n35631, n35632, n35633, n35634, n35635, n35636,
    n35637, n35638, n35639, n35640, n35641, n35642, n35643, n35645, n35646,
    n35647, n35648, n35649, n35650, n35651, n35652, n35653, n35654, n35655,
    n35656, n35657, n35658, n35659, n35660, n35661, n35662, n35663, n35664,
    n35665, n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
    n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681, n35682,
    n35683, n35684, n35685, n35686, n35687, n35688, n35689, n35690, n35691,
    n35692, n35693, n35694, n35695, n35696, n35697, n35698, n35699, n35700,
    n35701, n35702, n35703, n35704, n35705, n35706, n35707, n35708, n35709,
    n35710, n35711, n35712, n35713, n35714, n35715, n35716, n35717, n35718,
    n35719, n35720, n35721, n35722, n35723, n35724, n35725, n35726, n35727,
    n35728, n35729, n35730, n35731, n35732, n35733, n35734, n35735, n35736,
    n35737, n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
    n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753, n35754,
    n35755, n35756, n35757, n35758, n35759, n35760, n35761, n35762, n35763,
    n35764, n35765, n35766, n35767, n35768, n35769, n35771, n35772, n35773,
    n35774, n35775, n35776, n35777, n35778, n35779, n35780, n35781, n35782,
    n35783, n35784, n35785, n35786, n35787, n35788, n35789, n35790, n35791,
    n35792, n35793, n35794, n35795, n35796, n35798, n35799, n35800, n35801,
    n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809, n35810,
    n35811, n35812, n35813, n35814, n35815, n35816, n35817, n35819, n35820,
    n35821, n35822, n35823, n35824, n35825, n35826, n35827, n35828, n35829,
    n35830, n35831, n35832, n35833, n35834, n35835, n35836, n35837, n35838,
    n35840, n35841, n35842, n35843, n35844, n35845, n35846, n35847, n35848,
    n35849, n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
    n35858, n35859, n35861, n35862, n35863, n35864, n35865, n35866, n35867,
    n35868, n35869, n35870, n35871, n35872, n35873, n35874, n35875, n35876,
    n35877, n35878, n35879, n35880, n35881, n35882, n35883, n35884, n35885,
    n35886, n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894,
    n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903,
    n35904, n35905, n35906, n35907, n35908, n35909, n35910, n35911, n35912,
    n35913, n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
    n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929, n35930,
    n35931, n35932, n35933, n35934, n35935, n35936, n35937, n35938, n35939,
    n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947, n35948,
    n35949, n35950, n35951, n35952, n35953, n35954, n35955, n35956, n35957,
    n35958, n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966,
    n35967, n35968, n35969, n35970, n35971, n35972, n35973, n35974, n35975,
    n35977, n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
    n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993, n35994,
    n35995, n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003,
    n36004, n36005, n36006, n36007, n36008, n36009, n36010, n36011, n36012,
    n36013, n36014, n36015, n36016, n36017, n36018, n36019, n36020, n36021,
    n36022, n36023, n36024, n36025, n36026, n36027, n36028, n36029, n36030,
    n36031, n36032, n36033, n36034, n36035, n36036, n36037, n36038, n36039,
    n36040, n36041, n36042, n36043, n36044, n36045, n36046, n36047, n36048,
    n36049, n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
    n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065, n36066,
    n36067, n36068, n36069, n36070, n36071, n36072, n36073, n36074, n36075,
    n36076, n36077, n36078, n36079, n36080, n36081, n36082, n36083, n36084,
    n36085, n36086, n36088, n36089, n36090, n36091, n36092, n36093, n36094,
    n36095, n36096, n36097, n36098, n36099, n36100, n36101, n36102, n36103,
    n36104, n36105, n36107, n36108, n36109, n36110, n36111, n36112, n36114,
    n36115, n36116, n36117, n36118, n36119, n36120, n36121, n36122, n36123,
    n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36131, n36132,
    n36133, n36135, n36136, n36137, n36138, n36139, n36140, n36142, n36143,
    n36144, n36145, n36146, n36147, n36148, n36149, n36150, n36151, n36152,
    n36153, n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
    n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169, n36170,
    n36171, n36172, n36173, n36174, n36175, n36176, n36177, n36178, n36179,
    n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187, n36188,
    n36189, n36190, n36191, n36192, n36193, n36194, n36195, n36196, n36197,
    n36198, n36199, n36200, n36201, n36202, n36203, n36204, n36205, n36206,
    n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214, n36215,
    n36216, n36217, n36218, n36219, n36220, n36221, n36222, n36223, n36224,
    n36225, n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
    n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241, n36242,
    n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36251, n36252,
    n36253, n36254, n36255, n36256, n36257, n36258, n36259, n36260, n36261,
    n36262, n36263, n36264, n36265, n36266, n36267, n36268, n36269, n36270,
    n36271, n36272, n36273, n36274, n36275, n36276, n36277, n36278, n36279,
    n36280, n36281, n36282, n36283, n36284, n36285, n36286, n36287, n36288,
    n36289, n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
    n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305, n36306,
    n36307, n36308, n36309, n36310, n36311, n36312, n36313, n36314, n36315,
    n36316, n36317, n36318, n36319, n36320, n36321, n36322, n36323, n36324,
    n36325, n36326, n36327, n36328, n36329, n36330, n36331, n36332, n36333,
    n36334, n36335, n36336, n36337, n36338, n36339, n36340, n36341, n36342,
    n36343, n36344, n36345, n36346, n36347, n36348, n36349, n36350, n36351,
    n36352, n36353, n36354, n36355, n36356, n36357, n36358, n36359, n36360,
    n36361, n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
    n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377, n36378,
    n36379, n36380, n36381, n36382, n36383, n36384, n36385, n36386, n36387,
    n36388, n36389, n36390, n36391, n36392, n36393, n36394, n36395, n36396,
    n36397, n36398, n36399, n36400, n36401, n36402, n36403, n36404, n36405,
    n36406, n36407, n36408, n36409, n36410, n36411, n36412, n36413, n36414,
    n36415, n36416, n36417, n36418, n36419, n36420, n36421, n36422, n36423,
    n36424, n36425, n36426, n36427, n36428, n36429, n36430, n36431, n36432,
    n36433, n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
    n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450,
    n36451, n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459,
    n36460, n36461, n36462, n36463, n36464, n36465, n36466, n36467, n36468,
    n36469, n36470, n36471, n36472, n36473, n36474, n36475, n36476, n36477,
    n36478, n36479, n36480, n36481, n36482, n36483, n36484, n36485, n36486,
    n36487, n36488, n36489, n36490, n36491, n36492, n36493, n36494, n36495,
    n36496, n36497, n36498, n36499, n36500, n36501, n36502, n36503, n36504,
    n36505, n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
    n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521, n36522,
    n36523, n36524, n36525, n36526, n36527, n36528, n36529, n36530, n36531,
    n36532, n36533, n36534, n36535, n36536, n36537, n36538, n36539, n36540,
    n36541, n36542, n36543, n36544, n36545, n36546, n36547, n36548, n36549,
    n36550, n36551, n36552, n36553, n36554, n36555, n36556, n36557, n36558,
    n36559, n36560, n36561, n36562, n36563, n36564, n36565, n36566, n36567,
    n36568, n36569, n36570, n36571, n36572, n36573, n36574, n36575, n36576,
    n36577, n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
    n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594,
    n36595, n36596, n36597, n36598, n36599, n36600, n36601, n36602, n36603,
    n36604, n36605, n36606, n36607, n36608, n36609, n36610, n36611, n36612,
    n36613, n36614, n36615, n36616, n36617, n36618, n36619, n36620, n36621,
    n36622, n36623, n36624, n36625, n36626, n36627, n36628, n36629, n36630,
    n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638, n36639,
    n36640, n36641, n36642, n36643, n36644, n36645, n36646, n36647, n36648,
    n36649, n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
    n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665, n36666,
    n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675,
    n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683, n36684,
    n36685, n36686, n36687, n36688, n36689, n36690, n36691, n36692, n36693,
    n36694, n36695, n36696, n36697, n36698, n36699, n36700, n36701, n36702,
    n36703, n36704, n36705, n36706, n36707, n36708, n36709, n36710, n36711,
    n36712, n36713, n36714, n36715, n36716, n36717, n36718, n36719, n36720,
    n36721, n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
    n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738,
    n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746, n36747,
    n36748, n36749, n36750, n36751, n36752, n36753, n36754, n36755, n36756,
    n36757, n36758, n36759, n36760, n36761, n36762, n36763, n36764, n36765,
    n36766, n36767, n36768, n36769, n36770, n36771, n36772, n36773, n36774,
    n36775, n36776, n36777, n36778, n36779, n36780, n36781, n36782, n36783,
    n36784, n36785, n36786, n36787, n36788, n36789, n36790, n36791, n36792,
    n36793, n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801,
    n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809, n36810,
    n36811, n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819,
    n36820, n36821, n36822, n36823, n36824, n36825, n36826, n36827, n36828,
    n36829, n36830, n36831, n36832, n36833, n36834, n36835, n36836, n36837,
    n36838, n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846,
    n36847, n36848, n36849, n36850, n36851, n36852, n36853, n36854, n36855,
    n36856, n36857, n36858, n36859, n36860, n36861, n36862, n36863, n36864,
    n36865, n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873,
    n36874, n36875, n36877, n36878, n36879, n36880, n36881, n36882, n36883,
    n36884, n36885, n36886, n36887, n36888, n36889, n36890, n36891, n36892,
    n36893, n36894, n36895, n36896, n36897, n36898, n36899, n36900, n36901,
    n36902, n36903, n36904, n36905, n36906, n36907, n36908, n36909, n36910,
    n36911, n36912, n36913, n36914, n36915, n36916, n36917, n36918, n36919,
    n36920, n36921, n36922, n36923, n36924, n36925, n36926, n36927, n36928,
    n36929, n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
    n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945, n36946,
    n36947, n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955,
    n36956, n36957, n36958, n36959, n36960, n36961, n36962, n36963, n36964,
    n36965, n36966, n36967, n36968, n36969, n36970, n36971, n36972, n36973,
    n36974, n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982,
    n36983, n36984, n36985, n36986, n36987, n36988, n36989, n36990, n36991,
    n36992, n36993, n36994, n36995, n36996, n36997, n36998, n36999, n37000,
    n37001, n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
    n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017, n37018,
    n37019, n37020, n37021, n37022, n37023, n37024, n37025, n37026, n37027,
    n37028, n37029, n37030, n37031, n37032, n37033, n37034, n37035, n37036,
    n37037, n37038, n37039, n37040, n37041, n37042, n37043, n37044, n37045,
    n37046, n37047, n37048, n37049, n37050, n37051, n37052, n37053, n37054,
    n37055, n37056, n37057, n37058, n37059, n37060, n37061, n37062, n37063,
    n37064, n37065, n37066, n37067, n37068, n37069, n37070, n37071, n37072,
    n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
    n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37090,
    n37091, n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099,
    n37100, n37101, n37102, n37103, n37104, n37105, n37106, n37107, n37108,
    n37109, n37110, n37111, n37112, n37113, n37114, n37115, n37116, n37117,
    n37118, n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126,
    n37127, n37128, n37129, n37130, n37131, n37132, n37133, n37134, n37135,
    n37136, n37137, n37138, n37139, n37140, n37141, n37142, n37143, n37144,
    n37145, n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
    n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37162,
    n37163, n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171,
    n37172, n37173, n37174, n37175, n37176, n37177, n37178, n37179, n37180,
    n37181, n37182, n37183, n37184, n37185, n37186, n37187, n37188, n37189,
    n37190, n37191, n37192, n37193, n37194, n37195, n37196, n37197, n37198,
    n37199, n37200, n37201, n37202, n37203, n37204, n37205, n37206, n37207,
    n37208, n37209, n37210, n37211, n37212, n37213, n37214, n37215, n37216,
    n37217, n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
    n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234,
    n37235, n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243,
    n37244, n37245, n37246, n37247, n37248, n37249, n37250, n37251, n37252,
    n37253, n37254, n37255, n37256, n37257, n37258, n37259, n37260, n37261,
    n37262, n37263, n37264, n37265, n37266, n37267, n37268, n37269, n37270,
    n37271, n37272, n37273, n37274, n37275, n37276, n37277, n37278, n37279,
    n37280, n37281, n37282, n37283, n37284, n37285, n37286, n37287, n37288,
    n37289, n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
    n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305, n37306,
    n37307, n37308, n37309, n37310, n37311, n37312, n37313, n37314, n37315,
    n37316, n37317, n37318, n37319, n37320, n37321, n37322, n37323, n37324,
    n37325, n37326, n37327, n37328, n37329, n37330, n37331, n37332, n37333,
    n37334, n37335, n37336, n37337, n37338, n37339, n37340, n37341, n37342,
    n37343, n37344, n37345, n37346, n37347, n37348, n37349, n37350, n37351,
    n37352, n37353, n37354, n37355, n37356, n37357, n37358, n37359, n37360,
    n37361, n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
    n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377, n37378,
    n37379, n37380, n37381, n37382, n37383, n37384, n37385, n37386, n37387,
    n37388, n37389, n37390, n37391, n37392, n37393, n37394, n37395, n37396,
    n37397, n37398, n37399, n37400, n37401, n37402, n37403, n37404, n37405,
    n37406, n37407, n37408, n37409, n37410, n37411, n37412, n37413, n37414,
    n37415, n37416, n37417, n37418, n37419, n37420, n37421, n37422, n37423,
    n37424, n37425, n37426, n37427, n37428, n37429, n37430, n37431, n37432,
    n37433, n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
    n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449, n37450,
    n37451, n37452, n37453, n37454, n37455, n37456, n37457, n37459, n37460,
    n37461, n37462, n37463, n37464, n37465, n37466, n37467, n37468, n37469,
    n37470, n37471, n37472, n37473, n37474, n37475, n37476, n37477, n37478,
    n37479, n37480, n37481, n37482, n37483, n37484, n37485, n37486, n37487,
    n37488, n37489, n37490, n37491, n37492, n37493, n37494, n37495, n37496,
    n37497, n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505,
    n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513, n37514,
    n37515, n37516, n37517, n37518, n37519, n37520, n37521, n37522, n37523,
    n37524, n37525, n37526, n37527, n37528, n37529, n37530, n37531, n37532,
    n37533, n37534, n37535, n37536, n37537, n37538, n37539, n37540, n37541,
    n37542, n37543, n37544, n37545, n37546, n37547, n37548, n37549, n37550,
    n37551, n37552, n37553, n37554, n37555, n37556, n37557, n37558, n37559,
    n37560, n37561, n37562, n37563, n37564, n37565, n37566, n37567, n37568,
    n37569, n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577,
    n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585, n37586,
    n37587, n37588, n37589, n37590, n37591, n37592, n37593, n37594, n37595,
    n37596, n37597, n37598, n37599, n37600, n37601, n37602, n37603, n37604,
    n37605, n37606, n37607, n37608, n37609, n37610, n37611, n37612, n37613,
    n37614, n37615, n37616, n37617, n37618, n37619, n37620, n37621, n37622,
    n37623, n37624, n37625, n37626, n37627, n37628, n37629, n37630, n37631,
    n37632, n37633, n37634, n37635, n37636, n37637, n37638, n37639, n37640,
    n37641, n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649,
    n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657, n37658,
    n37659, n37660, n37661, n37662, n37663, n37664, n37665, n37666, n37667,
    n37668, n37669, n37670, n37671, n37672, n37673, n37674, n37675, n37676,
    n37677, n37678, n37679, n37680, n37681, n37682, n37683, n37684, n37685,
    n37686, n37687, n37688, n37689, n37690, n37691, n37692, n37693, n37694,
    n37695, n37696, n37697, n37698, n37699, n37700, n37701, n37702, n37703,
    n37704, n37705, n37706, n37707, n37708, n37709, n37710, n37711, n37712,
    n37713, n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
    n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729, n37730,
    n37731, n37732, n37733, n37734, n37735, n37736, n37737, n37738, n37739,
    n37740, n37741, n37742, n37743, n37744, n37745, n37746, n37747, n37748,
    n37749, n37750, n37751, n37752, n37753, n37754, n37755, n37756, n37757,
    n37758, n37759, n37760, n37761, n37762, n37763, n37764, n37765, n37766,
    n37767, n37768, n37769, n37770, n37771, n37772, n37773, n37774, n37775,
    n37776, n37777, n37778, n37779, n37780, n37781, n37782, n37783, n37784,
    n37785, n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793,
    n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801, n37802,
    n37803, n37804, n37805, n37806, n37807, n37808, n37809, n37810, n37811,
    n37812, n37813, n37814, n37815, n37816, n37817, n37818, n37819, n37820,
    n37821, n37822, n37823, n37824, n37825, n37826, n37827, n37828, n37829,
    n37830, n37831, n37832, n37833, n37834, n37835, n37836, n37837, n37838,
    n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846, n37847,
    n37848, n37849, n37850, n37851, n37852, n37853, n37854, n37855, n37856,
    n37857, n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865,
    n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873, n37874,
    n37875, n37876, n37877, n37878, n37879, n37880, n37881, n37882, n37883,
    n37884, n37885, n37886, n37887, n37888, n37889, n37890, n37891, n37892,
    n37893, n37894, n37895, n37896, n37897, n37898, n37899, n37900, n37901,
    n37902, n37903, n37904, n37905, n37906, n37907, n37908, n37909, n37910,
    n37911, n37912, n37913, n37914, n37915, n37916, n37917, n37918, n37919,
    n37920, n37921, n37922, n37923, n37924, n37925, n37926, n37927, n37928,
    n37929, n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937,
    n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945, n37946,
    n37947, n37948, n37949, n37950, n37951, n37952, n37953, n37954, n37955,
    n37956, n37957, n37958, n37959, n37960, n37961, n37962, n37963, n37964,
    n37965, n37966, n37967, n37968, n37969, n37970, n37971, n37972, n37973,
    n37974, n37975, n37976, n37977, n37978, n37979, n37980, n37981, n37982,
    n37983, n37984, n37985, n37986, n37987, n37988, n37989, n37990, n37991,
    n37992, n37993, n37994, n37995, n37996, n37997, n37998, n37999, n38000,
    n38001, n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009,
    n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017, n38018,
    n38019, n38020, n38021, n38022, n38023, n38024, n38025, n38026, n38027,
    n38028, n38029, n38030, n38031, n38032, n38033, n38034, n38035, n38036,
    n38037, n38038, n38039, n38040, n38041, n38042, n38043, n38044, n38045,
    n38046, n38048, n38049, n38050, n38051, n38052, n38053, n38054, n38055,
    n38056, n38057, n38058, n38059, n38060, n38061, n38062, n38063, n38064,
    n38065, n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073,
    n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081, n38082,
    n38083, n38084, n38085, n38086, n38087, n38088, n38089, n38090, n38091,
    n38092, n38093, n38094, n38095, n38096, n38097, n38098, n38099, n38100,
    n38101, n38102, n38103, n38104, n38105, n38106, n38107, n38108, n38109,
    n38110, n38111, n38112, n38113, n38114, n38115, n38116, n38117, n38118,
    n38119, n38120, n38121, n38122, n38123, n38124, n38125, n38126, n38127,
    n38128, n38129, n38130, n38131, n38132, n38133, n38134, n38135, n38136,
    n38137, n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145,
    n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153, n38154,
    n38155, n38156, n38157, n38158, n38159, n38160, n38161, n38162, n38163,
    n38164, n38165, n38166, n38167, n38168, n38169, n38170, n38171, n38173,
    n38174, n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182,
    n38183, n38184, n38185, n38186, n38187, n38188, n38189, n38190, n38191,
    n38192, n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38200,
    n38201, n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209,
    n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217, n38218,
    n38219, n38220, n38221, n38222, n38223, n38224, n38226, n38227, n38228,
    n38229, n38230, n38231, n38232, n38233, n38234, n38235, n38236, n38237,
    n38238, n38239, n38240, n38241, n38242, n38243, n38244, n38245, n38246,
    n38247, n38248, n38249, n38250, n38251, n38252, n38253, n38254, n38255,
    n38257, n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265,
    n38266, n38267, n38269, n38270, n38271, n38272, n38273, n38274, n38275,
    n38276, n38277, n38278, n38279, n38280, n38281, n38282, n38283, n38284,
    n38285, n38286, n38287, n38288, n38289, n38290, n38291, n38292, n38293,
    n38294, n38295, n38296, n38297, n38298, n38299, n38300, n38301, n38302,
    n38303, n38304, n38305, n38306, n38307, n38308, n38309, n38310, n38311,
    n38312, n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320,
    n38321, n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329,
    n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338,
    n38339, n38340, n38341, n38342, n38343, n38344, n38345, n38346, n38347,
    n38348, n38349, n38350, n38352, n38353, n38354, n38355, n38356, n38357,
    n38358, n38359, n38360, n38361, n38362, n38363, n38364, n38365, n38366,
    n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374, n38375,
    n38376, n38377, n38378, n38379, n38380, n38381, n38382, n38383, n38384,
    n38385, n38386, n38387, n38389, n38390, n38391, n38392, n38393, n38394,
    n38395, n38396, n38397, n38398, n38399, n38400, n38401, n38402, n38403,
    n38404, n38405, n38406, n38407, n38408, n38409, n38410, n38412, n38413,
    n38414, n38415, n38416, n38417, n38418, n38419, n38420, n38421, n38422,
    n38423, n38424, n38425, n38426, n38427, n38428, n38429, n38430, n38431,
    n38432, n38433, n38434, n38435, n38436, n38437, n38438, n38439, n38440,
    n38441, n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449,
    n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457, n38458,
    n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466, n38467,
    n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475, n38476,
    n38477, n38478, n38479, n38480, n38481, n38482, n38483, n38484, n38485,
    n38486, n38487, n38488, n38489, n38490, n38491, n38492, n38493, n38494,
    n38495, n38496, n38497, n38498, n38499, n38500, n38501, n38502, n38503,
    n38504, n38505, n38506, n38507, n38508, n38509, n38510, n38511, n38512,
    n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
    n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529, n38530,
    n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538, n38539,
    n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547, n38548,
    n38549, n38550, n38551, n38552, n38553, n38554, n38555, n38556, n38557,
    n38558, n38559, n38560, n38561, n38562, n38563, n38564, n38565, n38566,
    n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574, n38575,
    n38576, n38577, n38578, n38579, n38580, n38581, n38582, n38583, n38584,
    n38585, n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593,
    n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601, n38602,
    n38603, n38604, n38605, n38606, n38607, n38608, n38609, n38610, n38611,
    n38612, n38613, n38614, n38615, n38616, n38617, n38618, n38619, n38620,
    n38621, n38622, n38623, n38624, n38625, n38626, n38627, n38628, n38629,
    n38630, n38631, n38632, n38633, n38634, n38635, n38636, n38637, n38638,
    n38639, n38640, n38641, n38642, n38643, n38644, n38645, n38646, n38647,
    n38648, n38649, n38650, n38651, n38652, n38653, n38654, n38655, n38656,
    n38657, n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665,
    n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673, n38674,
    n38675, n38676, n38677, n38678, n38679, n38680, n38681, n38682, n38683,
    n38684, n38685, n38686, n38687, n38688, n38689, n38690, n38691, n38692,
    n38693, n38694, n38695, n38696, n38697, n38698, n38699, n38700, n38701,
    n38702, n38703, n38704, n38705, n38706, n38707, n38708, n38709, n38710,
    n38711, n38712, n38713, n38714, n38715, n38716, n38717, n38718, n38719,
    n38720, n38721, n38722, n38723, n38724, n38725, n38726, n38727, n38728,
    n38729, n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737,
    n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745, n38746,
    n38747, n38748, n38749, n38750, n38751, n38752, n38753, n38754, n38755,
    n38756, n38757, n38758, n38759, n38760, n38761, n38762, n38763, n38764,
    n38765, n38766, n38767, n38768, n38769, n38770, n38771, n38772, n38773,
    n38774, n38775, n38776, n38777, n38778, n38779, n38780, n38781, n38782,
    n38783, n38784, n38785, n38786, n38787, n38788, n38789, n38790, n38791,
    n38792, n38793, n38794, n38795, n38796, n38797, n38798, n38799, n38800,
    n38801, n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809,
    n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817, n38818,
    n38819, n38820, n38821, n38822, n38824, n38825, n38826, n38827, n38828,
    n38829, n38830, n38831, n38832, n38833, n38834, n38835, n38836, n38837,
    n38838, n38839, n38840, n38841, n38842, n38843, n38844, n38845, n38846,
    n38847, n38848, n38849, n38850, n38851, n38852, n38853, n38854, n38855,
    n38856, n38857, n38858, n38859, n38860, n38861, n38862, n38863, n38864,
    n38865, n38866, n38867, n38868, n38869, n38870, n38871, n38872, n38873,
    n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881, n38882,
    n38883, n38884, n38885, n38886, n38887, n38888, n38889, n38890, n38891,
    n38892, n38893, n38894, n38895, n38896, n38897, n38898, n38899, n38900,
    n38901, n38902, n38903, n38904, n38905, n38906, n38907, n38908, n38909,
    n38910, n38911, n38912, n38913, n38914, n38915, n38916, n38917, n38918,
    n38919, n38920, n38921, n38922, n38923, n38924, n38925, n38926, n38927,
    n38928, n38929, n38930, n38931, n38932, n38933, n38934, n38935, n38936,
    n38937, n38938, n38939, n38940, n38941, n38942, n38943, n38944, n38945,
    n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953, n38954,
    n38955, n38956, n38957, n38958, n38959, n38960, n38961, n38962, n38963,
    n38964, n38965, n38966, n38967, n38968, n38969, n38970, n38971, n38972,
    n38973, n38974, n38975, n38976, n38977, n38978, n38979, n38980, n38981,
    n38982, n38983, n38984, n38985, n38986, n38987, n38988, n38989, n38990,
    n38991, n38992, n38993, n38994, n38995, n38996, n38997, n38998, n38999,
    n39000, n39001, n39002, n39003, n39004, n39005, n39006, n39007, n39008,
    n39009, n39010, n39011, n39012, n39013, n39014, n39015, n39016, n39017,
    n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025, n39026,
    n39027, n39028, n39029, n39030, n39031, n39032, n39033, n39034, n39035,
    n39036, n39037, n39038, n39039, n39040, n39041, n39042, n39043, n39044,
    n39045, n39046, n39047, n39048, n39049, n39050, n39051, n39052, n39053,
    n39054, n39055, n39056, n39057, n39058, n39059, n39060, n39061, n39062,
    n39063, n39064, n39065, n39066, n39067, n39068, n39069, n39070, n39071,
    n39072, n39073, n39074, n39075, n39076, n39077, n39078, n39079, n39080,
    n39081, n39082, n39083, n39084, n39085, n39086, n39087, n39088, n39089,
    n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097, n39098,
    n39099, n39100, n39101, n39102, n39103, n39104, n39105, n39106, n39107,
    n39108, n39109, n39110, n39111, n39112, n39113, n39114, n39115, n39116,
    n39117, n39118, n39119, n39120, n39121, n39122, n39123, n39124, n39125,
    n39126, n39127, n39128, n39129, n39130, n39131, n39132, n39133, n39134,
    n39135, n39136, n39137, n39138, n39139, n39140, n39141, n39142, n39143,
    n39144, n39145, n39146, n39147, n39148, n39149, n39150, n39151, n39152,
    n39153, n39154, n39155, n39156, n39158, n39159, n39160, n39161, n39162,
    n39163, n39164, n39165, n39166, n39167, n39168, n39169, n39170, n39171,
    n39172, n39173, n39174, n39175, n39176, n39177, n39178, n39179, n39180,
    n39181, n39182, n39183, n39184, n39185, n39186, n39187, n39188, n39189,
    n39190, n39191, n39192, n39193, n39194, n39195, n39196, n39197, n39198,
    n39199, n39200, n39201, n39202, n39203, n39204, n39205, n39206, n39207,
    n39208, n39209, n39210, n39211, n39212, n39213, n39214, n39215, n39216,
    n39217, n39218, n39219, n39220, n39221, n39222, n39223, n39224, n39225,
    n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233, n39234,
    n39235, n39236, n39237, n39238, n39239, n39240, n39241, n39242, n39243,
    n39244, n39245, n39246, n39247, n39248, n39249, n39250, n39251, n39252,
    n39253, n39254, n39255, n39256, n39257, n39258, n39259, n39260, n39261,
    n39262, n39263, n39264, n39265, n39266, n39267, n39268, n39269, n39270,
    n39271, n39272, n39273, n39274, n39275, n39276, n39277, n39278, n39279,
    n39280, n39281, n39282, n39283, n39284, n39285, n39286, n39287, n39288,
    n39289, n39290, n39291, n39292, n39293, n39294, n39295, n39296, n39297,
    n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305, n39306,
    n39307, n39308, n39309, n39310, n39311, n39312, n39313, n39314, n39315,
    n39316, n39317, n39318, n39319, n39320, n39321, n39322, n39323, n39324,
    n39325, n39326, n39327, n39328, n39329, n39330, n39331, n39332, n39333,
    n39334, n39335, n39336, n39337, n39338, n39339, n39340, n39341, n39342,
    n39343, n39344, n39345, n39346, n39347, n39348, n39349, n39350, n39351,
    n39352, n39353, n39354, n39356, n39357, n39358, n39359, n39360, n39361,
    n39362, n39363, n39364, n39365, n39366, n39367, n39369, n39370, n39371,
    n39372, n39373, n39374, n39375, n39376, n39377, n39378, n39379, n39380,
    n39381, n39382, n39383, n39384, n39385, n39386, n39387, n39388, n39389,
    n39390, n39391, n39392, n39393, n39394, n39395, n39396, n39397, n39398,
    n39399, n39400, n39401, n39402, n39403, n39404, n39405, n39406, n39407,
    n39408, n39409, n39410, n39411, n39412, n39413, n39414, n39415, n39416,
    n39417, n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425,
    n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433, n39434,
    n39435, n39436, n39437, n39438, n39439, n39440, n39441, n39442, n39443,
    n39444, n39445, n39446, n39447, n39448, n39449, n39450, n39451, n39452,
    n39453, n39454, n39455, n39456, n39457, n39458, n39459, n39460, n39461,
    n39462, n39463, n39464, n39465, n39466, n39467, n39468, n39469, n39470,
    n39471, n39472, n39473, n39474, n39475, n39476, n39477, n39478, n39479,
    n39480, n39481, n39482, n39483, n39484, n39485, n39486, n39487, n39488,
    n39489, n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497,
    n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505, n39506,
    n39507, n39508, n39509, n39510, n39511, n39512, n39513, n39514, n39515,
    n39516, n39517, n39518, n39519, n39520, n39521, n39522, n39523, n39524,
    n39525, n39526, n39527, n39528, n39529, n39530, n39531, n39532, n39533,
    n39534, n39535, n39536, n39537, n39538, n39539, n39540, n39541, n39542,
    n39543, n39544, n39545, n39546, n39547, n39548, n39549, n39550, n39551,
    n39552, n39553, n39554, n39555, n39556, n39557, n39558, n39559, n39560,
    n39561, n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569,
    n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577, n39578,
    n39579, n39580, n39581, n39582, n39583, n39584, n39585, n39586, n39587,
    n39588, n39589, n39590, n39591, n39592, n39593, n39594, n39595, n39596,
    n39597, n39598, n39599, n39600, n39601, n39602, n39603, n39604, n39605,
    n39606, n39607, n39608, n39609, n39610, n39611, n39612, n39613, n39614,
    n39615, n39616, n39617, n39618, n39619, n39620, n39621, n39622, n39623,
    n39624, n39625, n39626, n39627, n39628, n39629, n39631, n39632, n39633,
    n39634, n39635, n39636, n39637, n39638, n39639, n39640, n39641, n39642,
    n39643, n39644, n39645, n39646, n39647, n39648, n39649, n39650, n39651,
    n39652, n39653, n39654, n39655, n39656, n39657, n39658, n39659, n39660,
    n39661, n39662, n39663, n39664, n39665, n39666, n39667, n39668, n39669,
    n39670, n39671, n39672, n39673, n39674, n39675, n39676, n39677, n39678,
    n39679, n39680, n39681, n39682, n39683, n39684, n39685, n39686, n39687,
    n39688, n39689, n39690, n39691, n39692, n39693, n39694, n39695, n39696,
    n39697, n39698, n39699, n39700, n39701, n39702, n39703, n39704, n39705,
    n39706, n39707, n39708, n39709, n39710, n39711, n39712, n39713, n39714,
    n39715, n39716, n39717, n39718, n39719, n39720, n39721, n39722, n39723,
    n39724, n39725, n39726, n39727, n39728, n39729, n39730, n39731, n39732,
    n39733, n39734, n39735, n39736, n39737, n39738, n39739, n39740, n39741,
    n39742, n39743, n39744, n39745, n39746, n39747, n39748, n39749, n39750,
    n39751, n39752, n39753, n39754, n39755, n39756, n39757, n39758, n39759,
    n39760, n39761, n39762, n39763, n39764, n39765, n39766, n39767, n39768,
    n39769, n39770, n39771, n39772, n39773, n39774, n39775, n39776, n39777,
    n39778, n39779, n39780, n39781, n39782, n39783, n39784, n39785, n39786,
    n39787, n39788, n39789, n39790, n39791, n39792, n39793, n39794, n39795,
    n39796, n39797, n39798, n39799, n39800, n39801, n39802, n39803, n39804,
    n39805, n39806, n39807, n39808, n39809, n39810, n39811, n39812, n39813,
    n39814, n39815, n39816, n39817, n39818, n39819, n39820, n39821, n39822,
    n39823, n39824, n39825, n39826, n39827, n39828, n39829, n39830, n39831,
    n39832, n39833, n39834, n39835, n39836, n39837, n39838, n39839, n39840,
    n39841, n39842, n39843, n39844, n39845, n39846, n39847, n39848, n39849,
    n39850, n39851, n39852, n39853, n39854, n39855, n39856, n39857, n39858,
    n39859, n39860, n39861, n39862, n39863, n39864, n39865, n39866, n39867,
    n39868, n39869, n39870, n39871, n39872, n39873, n39874, n39875, n39876,
    n39877, n39878, n39879, n39880, n39881, n39882, n39883, n39884, n39885,
    n39886, n39887, n39888, n39889, n39890, n39891, n39892, n39893, n39894,
    n39895, n39896, n39897, n39898, n39899, n39900, n39901, n39902, n39903,
    n39904, n39905, n39906, n39907, n39908, n39909, n39910, n39911, n39912,
    n39913, n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921,
    n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929, n39930,
    n39931, n39932, n39933, n39934, n39935, n39936, n39937, n39938, n39939,
    n39940, n39941, n39942, n39943, n39944, n39945, n39946, n39947, n39948,
    n39949, n39950, n39951, n39952, n39953, n39954, n39955, n39956, n39957,
    n39958, n39959, n39960, n39961, n39962, n39963, n39964, n39965, n39966,
    n39967, n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976,
    n39977, n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985,
    n39986, n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994,
    n39995, n39996, n39997, n39998, n39999, n40000, n40001, n40002, n40003,
    n40004, n40005, n40006, n40007, n40008, n40009, n40010, n40011, n40012,
    n40013, n40014, n40015, n40016, n40017, n40018, n40019, n40020, n40021,
    n40022, n40023, n40024, n40025, n40026, n40027, n40028, n40029, n40030,
    n40031, n40032, n40033, n40034, n40035, n40036, n40037, n40038, n40039,
    n40040, n40041, n40042, n40043, n40044, n40045, n40046, n40047, n40048,
    n40049, n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057,
    n40058, n40060, n40061, n40062, n40063, n40064, n40065, n40066, n40067,
    n40068, n40069, n40070, n40071, n40072, n40073, n40074, n40075, n40076,
    n40077, n40078, n40079, n40080, n40081, n40082, n40083, n40084, n40085,
    n40086, n40087, n40088, n40089, n40090, n40091, n40092, n40093, n40094,
    n40095, n40096, n40097, n40098, n40099, n40100, n40101, n40102, n40103,
    n40104, n40105, n40106, n40107, n40108, n40109, n40110, n40111, n40112,
    n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121,
    n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129, n40130,
    n40131, n40132, n40133, n40134, n40135, n40136, n40137, n40138, n40139,
    n40140, n40141, n40142, n40143, n40144, n40145, n40146, n40147, n40148,
    n40149, n40150, n40151, n40152, n40153, n40154, n40155, n40156, n40157,
    n40158, n40159, n40160, n40161, n40162, n40163, n40164, n40165, n40166,
    n40167, n40168, n40169, n40170, n40171, n40172, n40173, n40174, n40175,
    n40176, n40177, n40178, n40179, n40180, n40181, n40182, n40183, n40184,
    n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193,
    n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201, n40202,
    n40203, n40204, n40205, n40206, n40207, n40208, n40209, n40210, n40211,
    n40212, n40213, n40214, n40215, n40216, n40217, n40218, n40219, n40220,
    n40221, n40222, n40223, n40224, n40225, n40226, n40227, n40228, n40229,
    n40230, n40231, n40232, n40233, n40234, n40235, n40236, n40237, n40238,
    n40239, n40240, n40241, n40242, n40243, n40244, n40245, n40246, n40247,
    n40248, n40249, n40250, n40251, n40252, n40253, n40254, n40255, n40256,
    n40257, n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265,
    n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273, n40274,
    n40275, n40276, n40277, n40278, n40279, n40280, n40281, n40282, n40283,
    n40284, n40285, n40286, n40287, n40288, n40289, n40290, n40291, n40292,
    n40293, n40294, n40295, n40296, n40297, n40298, n40299, n40300, n40301,
    n40302, n40303, n40304, n40305, n40306, n40307, n40308, n40309, n40310,
    n40311, n40312, n40313, n40314, n40315, n40316, n40317, n40318, n40319,
    n40320, n40321, n40322, n40323, n40324, n40325, n40326, n40327, n40328,
    n40329, n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337,
    n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345, n40346,
    n40347, n40348, n40349, n40350, n40351, n40352, n40353, n40354, n40355,
    n40356, n40357, n40358, n40359, n40360, n40361, n40362, n40363, n40364,
    n40365, n40366, n40367, n40368, n40369, n40370, n40371, n40372, n40373,
    n40374, n40375, n40376, n40377, n40378, n40379, n40380, n40381, n40382,
    n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390, n40391,
    n40392, n40393, n40394, n40395, n40396, n40397, n40398, n40399, n40400,
    n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409,
    n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417, n40418,
    n40419, n40420, n40421, n40422, n40423, n40424, n40425, n40426, n40427,
    n40428, n40429, n40430, n40431, n40432, n40433, n40434, n40435, n40436,
    n40437, n40438, n40439, n40440, n40441, n40442, n40443, n40444, n40445,
    n40446, n40447, n40448, n40449, n40450, n40451, n40452, n40453, n40454,
    n40455, n40456, n40457, n40458, n40459, n40460, n40461, n40462, n40463,
    n40464, n40465, n40466, n40467, n40468, n40469, n40470, n40471, n40472,
    n40473, n40474, n40475, n40476, n40477, n40478, n40479, n40481, n40482,
    n40483, n40484, n40485, n40486, n40487, n40488, n40489, n40490, n40491,
    n40492, n40493, n40494, n40495, n40496, n40497, n40498, n40499, n40500,
    n40501, n40502, n40503, n40504, n40505, n40506, n40507, n40508, n40509,
    n40510, n40511, n40512, n40513, n40514, n40515, n40516, n40517, n40518,
    n40519, n40520, n40521, n40522, n40523, n40524, n40525, n40526, n40527,
    n40528, n40529, n40530, n40531, n40532, n40533, n40534, n40535, n40536,
    n40537, n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40545,
    n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553, n40554,
    n40555, n40556, n40557, n40558, n40559, n40560, n40561, n40562, n40563,
    n40564, n40565, n40566, n40567, n40568, n40569, n40570, n40571, n40572,
    n40573, n40574, n40575, n40576, n40577, n40578, n40579, n40580, n40581,
    n40582, n40583, n40584, n40585, n40586, n40587, n40588, n40589, n40590,
    n40591, n40592, n40593, n40594, n40595, n40596, n40597, n40598, n40599,
    n40600, n40601, n40602, n40603, n40604, n40605, n40606, n40607, n40608,
    n40609, n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617,
    n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625, n40626,
    n40627, n40628, n40629, n40630, n40631, n40632, n40633, n40634, n40635,
    n40636, n40637, n40638, n40639, n40640, n40641, n40642, n40643, n40644,
    n40645, n40646, n40647, n40648, n40649, n40650, n40651, n40652, n40653,
    n40654, n40655, n40656, n40657, n40658, n40659, n40660, n40661, n40662,
    n40663, n40664, n40665, n40666, n40667, n40668, n40669, n40670, n40671,
    n40672, n40673, n40674, n40675, n40676, n40677, n40678, n40679, n40680,
    n40681, n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689,
    n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698,
    n40699, n40700, n40701, n40702, n40703, n40704, n40705, n40706, n40707,
    n40708, n40709, n40710, n40711, n40712, n40713, n40714, n40715, n40716,
    n40717, n40718, n40719, n40720, n40721, n40722, n40723, n40724, n40725,
    n40726, n40727, n40728, n40729, n40730, n40731, n40732, n40733, n40734,
    n40735, n40736, n40737, n40738, n40739, n40740, n40741, n40742, n40743,
    n40744, n40745, n40746, n40747, n40748, n40749, n40750, n40751, n40752,
    n40753, n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761,
    n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40770, n40771,
    n40772, n40773, n40774, n40775, n40776, n40777, n40778, n40779, n40780,
    n40781, n40782, n40783, n40784, n40785, n40786, n40787, n40788, n40789,
    n40790, n40791, n40792, n40793, n40794, n40795, n40796, n40797, n40798,
    n40799, n40800, n40801, n40802, n40803, n40804, n40805, n40806, n40807,
    n40808, n40809, n40810, n40811, n40812, n40813, n40814, n40815, n40816,
    n40817, n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825,
    n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833, n40834,
    n40835, n40836, n40837, n40838, n40839, n40840, n40841, n40842, n40843,
    n40844, n40845, n40846, n40847, n40848, n40849, n40850, n40851, n40852,
    n40853, n40854, n40855, n40856, n40857, n40859, n40860, n40861, n40862,
    n40863, n40864, n40865, n40866, n40867, n40868, n40869, n40870, n40871,
    n40872, n40873, n40874, n40875, n40876, n40877, n40878, n40879, n40880,
    n40881, n40882, n40883, n40884, n40885, n40886, n40887, n40888, n40889,
    n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897, n40898,
    n40899, n40900, n40901, n40902, n40903, n40904, n40905, n40906, n40907,
    n40908, n40909, n40910, n40911, n40912, n40913, n40914, n40915, n40916,
    n40917, n40918, n40919, n40920, n40921, n40922, n40923, n40924, n40925,
    n40926, n40927, n40928, n40929, n40930, n40931, n40932, n40933, n40934,
    n40935, n40936, n40937, n40938, n40939, n40940, n40941, n40942, n40943,
    n40944, n40945, n40946, n40947, n40948, n40949, n40950, n40951, n40952,
    n40953, n40954, n40955, n40956, n40957, n40958, n40959, n40960, n40961,
    n40962, n40963, n40964, n40965, n40966, n40967, n40968, n40969, n40970,
    n40971, n40972, n40973, n40974, n40975, n40976, n40977, n40978, n40979,
    n40980, n40981, n40982, n40983, n40984, n40985, n40986, n40987, n40988,
    n40989, n40990, n40991, n40992, n40993, n40994, n40995, n40996, n40997,
    n40998, n40999, n41000, n41001, n41002, n41003, n41004, n41005, n41006,
    n41007, n41008, n41009, n41010, n41011, n41012, n41013, n41014, n41015,
    n41016, n41017, n41018, n41019, n41020, n41021, n41022, n41023, n41024,
    n41025, n41026, n41027, n41028, n41029, n41030, n41031, n41032, n41033,
    n41034, n41035, n41036, n41037, n41038, n41039, n41040, n41041, n41042,
    n41043, n41044, n41045, n41046, n41047, n41048, n41049, n41050, n41051,
    n41052, n41053, n41054, n41055, n41056, n41057, n41058, n41059, n41060,
    n41061, n41062, n41063, n41064, n41065, n41066, n41067, n41068, n41069,
    n41070, n41071, n41072, n41073, n41074, n41075, n41076, n41077, n41078,
    n41079, n41080, n41081, n41082, n41083, n41084, n41085, n41086, n41087,
    n41088, n41089, n41090, n41091, n41092, n41093, n41094, n41095, n41096,
    n41097, n41098, n41099, n41100, n41101, n41102, n41103, n41104, n41105,
    n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113, n41114,
    n41115, n41116, n41117, n41118, n41119, n41120, n41121, n41122, n41123,
    n41124, n41125, n41126, n41127, n41128, n41129, n41130, n41131, n41132,
    n41133, n41134, n41135, n41136, n41137, n41138, n41139, n41140, n41141,
    n41142, n41143, n41144, n41145, n41146, n41147, n41148, n41149, n41150,
    n41151, n41152, n41153, n41154, n41155, n41156, n41157, n41158, n41159,
    n41160, n41161, n41162, n41163, n41164, n41165, n41166, n41167, n41168,
    n41170, n41171, n41172, n41173, n41174, n41175, n41176, n41177, n41178,
    n41179, n41180, n41181, n41182, n41183, n41184, n41185, n41186, n41187,
    n41188, n41189, n41190, n41191, n41192, n41193, n41194, n41195, n41196,
    n41197, n41198, n41199, n41200, n41201, n41202, n41203, n41204, n41205,
    n41206, n41207, n41208, n41209, n41210, n41211, n41212, n41213, n41214,
    n41215, n41216, n41217, n41218, n41219, n41220, n41221, n41223, n41224,
    n41225, n41226, n41227, n41228, n41229, n41230, n41231, n41232, n41233,
    n41234, n41235, n41236, n41237, n41238, n41239, n41240, n41241, n41242,
    n41243, n41244, n41245, n41246, n41247, n41248, n41249, n41250, n41251,
    n41252, n41253, n41254, n41255, n41256, n41257, n41258, n41259, n41260,
    n41261, n41262, n41263, n41264, n41265, n41266, n41267, n41268, n41269,
    n41270, n41271, n41272, n41273, n41274, n41275, n41276, n41277, n41278,
    n41279, n41280, n41281, n41282, n41283, n41284, n41285, n41286, n41287,
    n41288, n41289, n41290, n41291, n41292, n41293, n41294, n41295, n41296,
    n41297, n41298, n41299, n41300, n41301, n41302, n41303, n41304, n41305,
    n41306, n41307, n41308, n41309, n41310, n41311, n41312, n41313, n41314,
    n41315, n41316, n41317, n41318, n41319, n41320, n41321, n41322, n41323,
    n41324, n41325, n41326, n41327, n41328, n41329, n41330, n41331, n41332,
    n41333, n41334, n41335, n41336, n41337, n41338, n41339, n41340, n41341,
    n41342, n41343, n41344, n41345, n41346, n41347, n41348, n41349, n41350,
    n41351, n41352, n41353, n41354, n41355, n41356, n41357, n41358, n41359,
    n41360, n41361, n41362, n41363, n41364, n41365, n41366, n41367, n41368,
    n41369, n41370, n41371, n41372, n41373, n41374, n41375, n41376, n41377,
    n41378, n41379, n41380, n41381, n41382, n41383, n41384, n41385, n41386,
    n41387, n41388, n41389, n41390, n41391, n41392, n41393, n41394, n41395,
    n41396, n41397, n41398, n41399, n41400, n41401, n41402, n41403, n41404,
    n41405, n41406, n41407, n41408, n41409, n41410, n41411, n41412, n41413,
    n41414, n41415, n41416, n41417, n41418, n41419, n41420, n41421, n41422,
    n41423, n41424, n41425, n41426, n41427, n41428, n41429, n41430, n41431,
    n41432, n41433, n41434, n41435, n41436, n41437, n41438, n41439, n41440,
    n41441, n41442, n41443, n41444, n41445, n41446, n41447, n41448, n41449,
    n41450, n41451, n41452, n41453, n41454, n41455, n41456, n41457, n41458,
    n41459, n41460, n41461, n41462, n41463, n41464, n41465, n41466, n41467,
    n41468, n41470, n41471, n41472, n41473, n41474, n41475, n41476, n41477,
    n41478, n41479, n41480, n41481, n41482, n41483, n41484, n41485, n41486,
    n41487, n41488, n41489, n41490, n41491, n41492, n41493, n41494, n41495,
    n41496, n41497, n41498, n41499, n41500, n41501, n41502, n41503, n41504,
    n41505, n41506, n41507, n41508, n41509, n41510, n41511, n41512, n41513,
    n41514, n41515, n41516, n41517, n41518, n41519, n41520, n41521, n41522,
    n41523, n41524, n41525, n41526, n41527, n41528, n41529, n41530, n41531,
    n41532, n41533, n41534, n41535, n41536, n41537, n41538, n41539, n41540,
    n41541, n41542, n41543, n41544, n41545, n41546, n41547, n41548, n41549,
    n41550, n41551, n41552, n41553, n41554, n41555, n41556, n41557, n41558,
    n41559, n41560, n41561, n41562, n41563, n41564, n41565, n41566, n41567,
    n41568, n41569, n41570, n41571, n41572, n41573, n41574, n41575, n41576,
    n41577, n41578, n41579, n41580, n41581, n41582, n41583, n41584, n41585,
    n41586, n41587, n41588, n41589, n41590, n41591, n41592, n41593, n41594,
    n41595, n41596, n41597, n41598, n41599, n41600, n41601, n41602, n41603,
    n41604, n41605, n41606, n41607, n41608, n41609, n41610, n41611, n41612,
    n41613, n41614, n41615, n41616, n41617, n41618, n41619, n41620, n41621,
    n41622, n41623, n41624, n41625, n41626, n41627, n41628, n41629, n41630,
    n41631, n41632, n41633, n41634, n41635, n41636, n41637, n41638, n41639,
    n41640, n41641, n41642, n41643, n41644, n41645, n41646, n41647, n41648,
    n41649, n41650, n41651, n41652, n41653, n41654, n41655, n41656, n41657,
    n41658, n41659, n41660, n41661, n41662, n41663, n41664, n41665, n41666,
    n41667, n41668, n41669, n41670, n41671, n41672, n41673, n41674, n41675,
    n41676, n41677, n41678, n41679, n41680, n41681, n41682, n41683, n41684,
    n41685, n41686, n41687, n41688, n41689, n41690, n41691, n41692, n41693,
    n41694, n41695, n41696, n41697, n41698, n41699, n41700, n41701, n41702,
    n41703, n41704, n41705, n41706, n41707, n41708, n41709, n41710, n41711,
    n41712, n41713, n41714, n41715, n41716, n41717, n41718, n41719, n41720,
    n41721, n41722, n41723, n41724, n41725, n41726, n41727, n41728, n41729,
    n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737, n41738,
    n41739, n41740, n41741, n41742, n41744, n41745, n41746, n41747, n41748,
    n41749, n41750, n41751, n41752, n41753, n41754, n41755, n41756, n41757,
    n41758, n41759, n41760, n41761, n41762, n41763, n41764, n41765, n41766,
    n41767, n41768, n41769, n41770, n41771, n41772, n41773, n41774, n41775,
    n41776, n41777, n41778, n41779, n41780, n41781, n41782, n41783, n41784,
    n41785, n41786, n41787, n41788, n41789, n41790, n41791, n41792, n41793,
    n41794, n41795, n41796, n41797, n41798, n41799, n41800, n41801, n41802,
    n41803, n41804, n41805, n41806, n41807, n41808, n41809, n41810, n41811,
    n41812, n41813, n41814, n41815, n41816, n41817, n41818, n41819, n41820,
    n41821, n41822, n41823, n41824, n41825, n41826, n41827, n41828, n41829,
    n41830, n41831, n41832, n41833, n41834, n41835, n41836, n41837, n41838,
    n41839, n41840, n41841, n41842, n41843, n41844, n41845, n41846, n41847,
    n41848, n41849, n41850, n41851, n41852, n41853, n41854, n41855, n41856,
    n41857, n41858, n41859, n41860, n41861, n41862, n41863, n41864, n41865,
    n41866, n41867, n41868, n41869, n41870, n41871, n41872, n41873, n41874,
    n41875, n41876, n41877, n41878, n41879, n41880, n41881, n41882, n41883,
    n41884, n41885, n41886, n41887, n41888, n41889, n41890, n41891, n41892,
    n41893, n41894, n41895, n41896, n41897, n41898, n41899, n41900, n41901,
    n41902, n41903, n41904, n41905, n41906, n41907, n41908, n41909, n41910,
    n41911, n41912, n41913, n41914, n41915, n41916, n41917, n41918, n41919,
    n41920, n41921, n41922, n41923, n41924, n41925, n41926, n41927, n41928,
    n41929, n41930, n41931, n41932, n41933, n41934, n41935, n41936, n41937,
    n41938, n41939, n41940, n41941, n41942, n41943, n41944, n41945, n41946,
    n41947, n41948, n41949, n41950, n41951, n41952, n41953, n41954, n41955,
    n41956, n41957, n41958, n41959, n41960, n41961, n41962, n41963, n41964,
    n41965, n41966, n41967, n41968, n41969, n41970, n41971, n41972, n41974,
    n41975, n41976, n41977, n41978, n41979, n41980, n41981, n41982, n41983,
    n41984, n41985, n41986, n41987, n41988, n41989, n41990, n41991, n41992,
    n41993, n41994, n41995, n41996, n41997, n41998, n41999, n42000, n42001,
    n42002, n42003, n42004, n42005, n42006, n42007, n42008, n42009, n42010,
    n42011, n42012, n42013, n42014, n42015, n42016, n42017, n42018, n42019,
    n42020, n42021, n42022, n42023, n42024, n42025, n42026, n42027, n42028,
    n42029, n42030, n42031, n42032, n42033, n42034, n42035, n42036, n42037,
    n42038, n42039, n42040, n42041, n42042, n42043, n42044, n42045, n42046,
    n42047, n42048, n42049, n42050, n42051, n42052, n42053, n42054, n42055,
    n42056, n42057, n42058, n42059, n42060, n42061, n42062, n42063, n42064,
    n42065, n42066, n42067, n42068, n42069, n42070, n42071, n42072, n42073,
    n42074, n42075, n42076, n42077, n42078, n42079, n42080, n42081, n42082,
    n42083, n42084, n42085, n42086, n42087, n42088, n42089, n42090, n42091,
    n42092, n42093, n42094, n42095, n42096, n42097, n42098, n42099, n42100,
    n42101, n42102, n42103, n42104, n42105, n42106, n42107, n42108, n42109,
    n42110, n42111, n42112, n42113, n42114, n42115, n42116, n42117, n42118,
    n42119, n42120, n42121, n42122, n42123, n42124, n42125, n42126, n42127,
    n42128, n42129, n42130, n42131, n42132, n42133, n42134, n42135, n42137,
    n42138, n42139, n42140, n42141, n42142, n42143, n42144, n42145, n42146,
    n42147, n42148, n42149, n42150, n42151, n42152, n42153, n42154, n42155,
    n42156, n42157, n42158, n42159, n42160, n42161, n42162, n42163, n42164,
    n42165, n42166, n42167, n42168, n42169, n42170, n42171, n42172, n42173,
    n42174, n42175, n42176, n42177, n42178, n42179, n42180, n42181, n42182,
    n42183, n42184, n42185, n42186, n42187, n42188, n42189, n42190, n42191,
    n42192, n42193, n42194, n42195, n42196, n42197, n42198, n42199, n42200,
    n42201, n42202, n42203, n42204, n42205, n42206, n42207, n42208, n42209,
    n42210, n42211, n42212, n42213, n42214, n42215, n42216, n42217, n42218,
    n42219, n42220, n42221, n42222, n42223, n42224, n42225, n42226, n42227,
    n42228, n42229, n42230, n42231, n42232, n42233, n42234, n42235, n42236,
    n42237, n42238, n42239, n42240, n42241, n42242, n42243, n42244, n42245,
    n42246, n42247, n42248, n42249, n42250, n42251, n42252, n42253, n42254,
    n42255, n42256, n42257, n42258, n42259, n42260, n42261, n42262, n42263,
    n42264, n42265, n42266, n42267, n42268, n42269, n42270, n42271, n42272,
    n42273, n42274, n42275, n42276, n42277, n42278, n42279, n42280, n42281,
    n42282, n42283, n42284, n42285, n42286, n42287, n42288, n42289, n42290,
    n42291, n42292, n42293, n42294, n42295, n42296, n42297, n42298, n42299,
    n42300, n42301, n42302, n42303, n42304, n42305, n42306, n42307, n42308,
    n42309, n42310, n42311, n42312, n42313, n42314, n42315, n42316, n42317,
    n42318, n42319, n42320, n42321, n42322, n42323, n42325, n42326, n42327,
    n42328, n42329, n42330, n42331, n42333, n42334, n42335, n42336, n42337,
    n42338, n42339, n42340, n42341, n42343, n42344, n42345, n42346, n42347,
    n42348, n42349, n42350, n42351, n42352, n42353, n42354, n42355, n42356,
    n42357, n42358, n42359, n42360, n42361, n42362, n42363, n42364, n42365,
    n42366, n42367, n42368, n42369, n42370, n42371, n42372, n42373, n42374,
    n42375, n42376, n42377, n42378, n42379, n42380, n42381, n42382, n42383,
    n42385, n42386, n42387, n42388, n42389, n42390, n42391, n42392, n42393,
    n42394, n42395, n42396, n42397, n42398, n42399, n42400, n42401, n42402,
    n42403, n42404, n42405, n42406, n42407, n42408, n42409, n42410, n42411,
    n42412, n42413, n42414, n42415, n42416, n42417, n42418, n42419, n42420,
    n42421, n42422, n42423, n42424, n42425, n42426, n42427, n42428, n42429,
    n42430, n42431, n42432, n42433, n42434, n42435, n42436, n42437, n42438,
    n42439, n42440, n42441, n42442, n42443, n42444, n42445, n42446, n42447,
    n42448, n42449, n42450, n42451, n42452, n42453, n42454, n42455, n42456,
    n42457, n42458, n42459, n42460, n42461, n42462, n42463, n42464, n42465,
    n42466, n42467, n42468, n42469, n42470, n42471, n42472, n42473, n42474,
    n42475, n42476, n42477, n42478, n42479, n42480, n42481, n42482, n42483,
    n42484, n42485, n42486, n42487, n42488, n42489, n42490, n42491, n42492,
    n42493, n42494, n42495, n42496, n42497, n42498, n42499, n42500, n42501,
    n42502, n42503, n42504, n42505, n42506, n42507, n42508, n42509, n42510,
    n42511, n42512, n42513, n42514, n42515, n42516, n42517, n42518, n42519,
    n42520, n42521, n42522, n42523, n42524, n42525, n42526, n42527, n42528,
    n42529, n42530, n42531, n42532, n42533, n42534, n42535, n42536, n42537,
    n42538, n42539, n42540, n42541, n42542, n42543, n42544, n42545, n42546,
    n42547, n42548, n42549, n42550, n42551, n42552, n42553, n42554, n42555,
    n42556, n42557, n42558, n42559, n42560, n42561, n42562, n42563, n42564,
    n42565, n42566, n42567, n42568, n42569, n42570, n42571, n42572, n42573,
    n42574, n42575, n42576, n42577, n42578, n42579, n42580, n42581, n42582,
    n42583, n42584, n42585, n42586, n42587, n42588, n42589, n42590, n42591,
    n42592, n42593, n42594, n42595, n42596, n42597, n42598, n42599, n42600,
    n42601, n42602, n42603, n42604, n42605, n42606, n42607, n42608, n42609,
    n42610, n42611, n42612, n42613, n42614, n42615, n42616, n42617, n42618,
    n42619, n42621, n42622, n42623, n42624, n42625, n42626, n42627, n42628,
    n42629, n42630, n42631, n42632, n42633, n42634, n42635, n42636, n42637,
    n42638, n42639, n42640, n42641, n42642, n42643, n42644, n42645, n42646,
    n42647, n42648, n42649, n42650, n42651, n42652, n42653, n42654, n42655,
    n42656, n42657, n42658, n42659, n42660, n42661, n42662, n42663, n42664,
    n42665, n42666, n42667, n42668, n42669, n42670, n42671, n42672, n42673,
    n42674, n42675, n42676, n42677, n42678, n42679, n42680, n42681, n42682,
    n42683, n42684, n42685, n42686, n42687, n42688, n42689, n42690, n42691,
    n42692, n42693, n42694, n42695, n42696, n42697, n42698, n42699, n42700,
    n42701, n42702, n42703, n42704, n42705, n42706, n42707, n42708, n42709,
    n42710, n42711, n42712, n42713, n42714, n42715, n42716, n42717, n42718,
    n42719, n42720, n42721, n42722, n42723, n42724, n42725, n42726, n42727,
    n42728, n42729, n42730, n42731, n42732, n42733, n42734, n42735, n42736,
    n42737, n42738, n42739, n42740, n42741, n42742, n42743, n42744, n42745,
    n42746, n42747, n42748, n42749, n42750, n42751, n42752, n42753, n42754,
    n42755, n42756, n42757, n42758, n42759, n42760, n42761, n42762, n42763,
    n42764, n42765, n42766, n42767, n42768, n42769, n42770, n42771, n42772,
    n42773, n42774, n42775, n42776, n42777, n42778, n42779, n42780, n42781,
    n42782, n42783, n42784, n42785, n42786, n42787, n42788, n42789, n42790,
    n42791, n42792, n42793, n42794, n42795, n42796, n42797, n42798, n42799,
    n42800, n42801, n42802, n42803, n42804, n42805, n42806, n42807, n42808,
    n42809, n42810, n42811, n42812, n42813, n42814, n42815, n42816, n42817,
    n42818, n42819, n42820, n42821, n42822, n42823, n42824, n42825, n42826,
    n42827, n42828, n42829, n42830, n42831, n42832, n42833, n42834, n42835,
    n42836, n42837, n42838, n42839, n42840, n42841, n42842, n42843, n42844,
    n42845, n42847, n42848, n42849, n42850, n42851, n42853, n42854, n42855,
    n42856, n42857, n42859, n42860, n42861, n42862, n42863, n42865, n42866,
    n42867, n42868, n42869, n42871, n42872, n42873, n42874, n42875, n42877,
    n42878, n42879, n42880, n42881, n42882, n42884, n42885, n42886, n42887,
    n42888, n42889, n42891, n42892, n42893, n42894, n42895, n42896, n42897,
    n42898, n42899, n42900, n42901, n42902, n42903, n42904, n42905, n42906,
    n42907, n42908, n42909, n42910, n42911, n42912, n42913, n42914, n42915,
    n42916, n42917, n42918, n42919, n42920, n42921, n42922, n42923, n42925,
    n42926, n42927, n42928, n42929, n42930, n42931, n42932, n42933, n42934,
    n42935, n42936, n42937, n42938, n42939, n42940, n42941, n42942, n42943,
    n42944, n42945, n42946, n42947, n42948, n42949, n42950, n42951, n42952,
    n42953, n42954, n42955, n42956, n42957, n42958, n42959, n42960, n42961,
    n42962, n42963, n42964, n42965, n42966, n42967, n42968, n42969, n42970,
    n42971, n42972, n42973, n42974, n42975, n42976, n42977, n42978, n42979,
    n42980, n42981, n42982, n42983, n42984, n42985, n42986, n42987, n42988,
    n42989, n42990, n42991, n42992, n42993, n42994, n42995, n42996, n42997,
    n42998, n42999, n43000, n43001, n43002, n43003, n43004, n43005, n43006,
    n43007, n43008, n43009, n43010, n43011, n43012, n43013, n43014, n43015,
    n43016, n43017, n43018, n43019, n43020, n43021, n43022, n43023, n43024,
    n43025, n43026, n43027, n43028, n43029, n43030, n43031, n43032, n43033,
    n43034, n43035, n43036, n43037, n43038, n43039, n43040, n43041, n43042,
    n43043, n43044, n43045, n43046, n43047, n43048, n43049, n43050, n43051,
    n43052, n43053, n43054, n43055, n43056, n43057, n43058, n43059, n43060,
    n43061, n43062, n43063, n43064, n43065, n43066, n43067, n43068, n43069,
    n43070, n43071, n43072, n43073, n43074, n43075, n43076, n43077, n43078,
    n43079, n43080, n43081, n43082, n43083, n43084, n43085, n43086, n43087,
    n43088, n43089, n43090, n43091, n43092, n43093, n43094, n43095, n43096,
    n43097, n43098, n43099, n43100, n43101, n43102, n43103, n43104, n43105,
    n43106, n43107, n43108, n43109, n43110, n43111, n43112, n43113, n43114,
    n43115, n43116, n43117, n43118, n43119, n43120, n43121, n43122, n43123,
    n43124, n43125, n43126, n43127, n43128, n43129, n43130, n43131, n43132,
    n43133, n43135, n43136, n43137, n43138, n43139, n43140, n43141, n43142,
    n43143, n43144, n43145, n43146, n43147, n43148, n43149, n43150, n43151,
    n43152, n43153, n43154, n43155, n43156, n43157, n43158, n43159, n43160,
    n43161, n43162, n43163, n43164, n43165, n43166, n43167, n43168, n43169,
    n43170, n43171, n43172, n43173, n43174, n43175, n43176, n43177, n43178,
    n43180, n43181, n43182, n43183, n43184, n43185, n43186, n43187, n43188,
    n43189, n43190, n43191, n43192, n43193, n43194, n43195, n43196, n43197,
    n43198, n43199, n43200, n43201, n43202, n43203, n43204, n43205, n43206,
    n43207, n43208, n43209, n43210, n43211, n43212, n43213, n43214, n43215,
    n43216, n43217, n43218, n43219, n43221, n43222, n43223, n43224, n43225,
    n43226, n43227, n43228, n43229, n43230, n43231, n43232, n43233, n43234,
    n43235, n43236, n43237, n43238, n43239, n43240, n43241, n43242, n43243,
    n43244, n43245, n43246, n43247, n43248, n43249, n43250, n43251, n43252,
    n43253, n43254, n43255, n43256, n43257, n43258, n43259, n43260, n43261,
    n43262, n43263, n43264, n43265, n43266, n43267, n43268, n43269, n43270,
    n43271, n43272, n43273, n43274, n43275, n43276, n43277, n43278, n43279,
    n43280, n43281, n43282, n43283, n43284, n43285, n43286, n43288, n43289,
    n43290, n43291, n43292, n43293, n43294, n43295, n43296, n43297, n43298,
    n43299, n43300, n43301, n43302, n43303, n43304, n43305, n43306, n43307,
    n43308, n43309, n43310, n43311, n43312, n43313, n43314, n43315, n43316,
    n43317, n43318, n43319, n43320, n43321, n43322, n43323, n43324, n43325,
    n43326, n43327, n43328, n43329, n43330, n43331, n43332, n43333, n43334,
    n43335, n43336, n43337, n43338, n43339, n43340, n43341, n43342, n43343,
    n43344, n43345, n43346, n43347, n43348, n43349, n43350, n43351, n43352,
    n43353, n43354, n43355, n43356, n43357, n43358, n43359, n43360, n43361,
    n43362, n43363, n43364, n43365, n43366, n43367, n43368, n43369, n43370,
    n43371, n43372, n43373, n43374, n43375, n43376, n43377, n43378, n43379,
    n43380, n43381, n43382, n43383, n43384, n43385, n43386, n43387, n43388,
    n43389, n43390, n43391, n43392, n43393, n43394, n43395, n43396, n43397,
    n43398, n43399, n43400, n43401, n43402, n43403, n43404, n43405, n43406,
    n43407, n43408, n43409, n43410, n43411, n43412, n43413, n43414, n43415,
    n43416, n43417, n43418, n43419, n43420, n43421, n43422, n43423, n43424,
    n43425, n43426, n43427, n43428, n43429, n43430, n43431, n43432, n43433,
    n43434, n43435, n43436, n43437, n43438, n43439, n43440, n43441, n43442,
    n43443, n43444, n43445, n43446, n43447, n43448, n43449, n43450, n43451,
    n43452, n43453, n43454, n43455, n43456, n43457, n43458, n43459, n43460,
    n43461, n43462, n43463, n43464, n43465, n43466, n43467, n43468, n43469,
    n43470, n43471, n43472, n43473, n43474, n43475, n43476, n43477, n43478,
    n43479, n43480, n43481, n43482, n43483, n43484, n43485, n43486, n43487,
    n43488, n43489, n43490, n43491, n43492, n43493, n43495, n43496, n43497,
    n43498, n43499, n43500, n43501, n43502, n43503, n43504, n43505, n43506,
    n43507, n43508, n43509, n43510, n43511, n43512, n43513, n43514, n43515,
    n43516, n43517, n43518, n43519, n43520, n43521, n43522, n43523, n43524,
    n43525, n43526, n43527, n43528, n43529, n43530, n43531, n43532, n43533,
    n43534, n43535, n43536, n43537, n43538, n43539, n43540, n43541, n43542,
    n43543, n43544, n43545, n43546, n43547, n43548, n43549, n43550, n43551,
    n43552, n43553, n43554, n43555, n43556, n43557, n43558, n43559, n43560,
    n43561, n43562, n43563, n43564, n43565, n43566, n43567, n43568, n43569,
    n43570, n43571, n43572, n43573, n43574, n43575, n43576, n43577, n43578,
    n43579, n43580, n43581, n43582, n43583, n43584, n43585, n43586, n43587,
    n43588, n43589, n43590, n43591, n43592, n43593, n43594, n43595, n43596,
    n43597, n43598, n43599, n43600, n43601, n43602, n43603, n43604, n43605,
    n43606, n43607, n43608, n43609, n43610, n43611, n43612, n43613, n43614,
    n43615, n43616, n43617, n43618, n43619, n43620, n43621, n43622, n43623,
    n43624, n43625, n43626, n43627, n43628, n43629, n43630, n43631, n43632,
    n43633, n43634, n43635, n43636, n43637, n43638, n43639, n43640, n43641,
    n43642, n43643, n43644, n43645, n43646, n43647, n43648, n43649, n43650,
    n43652, n43653, n43654, n43655, n43656, n43657, n43658, n43659, n43660,
    n43661, n43662, n43663, n43664, n43665, n43666, n43667, n43668, n43669,
    n43670, n43671, n43672, n43673, n43674, n43675, n43676, n43677, n43678,
    n43679, n43680, n43681, n43682, n43683, n43684, n43685, n43686, n43687,
    n43688, n43689, n43690, n43691, n43692, n43693, n43694, n43695, n43697,
    n43698, n43699, n43700, n43701, n43702, n43703, n43704, n43705, n43706,
    n43707, n43708, n43709, n43710, n43711, n43712, n43713, n43714, n43715,
    n43716, n43717, n43718, n43719, n43720, n43721, n43722, n43723, n43724,
    n43725, n43726, n43727, n43728, n43729, n43730, n43731, n43732, n43733,
    n43734, n43735, n43736, n43737, n43738, n43739, n43741, n43742, n43743,
    n43744, n43745, n43746, n43747, n43748, n43749, n43750, n43751, n43752,
    n43753, n43754, n43755, n43756, n43757, n43758, n43759, n43760, n43761,
    n43762, n43763, n43764, n43765, n43766, n43767, n43768, n43769, n43770,
    n43771, n43772, n43773, n43774, n43775, n43776, n43777, n43778, n43779,
    n43780, n43781, n43782, n43783, n43784, n43785, n43786, n43787, n43788,
    n43790, n43791, n43792, n43793, n43794, n43795, n43796, n43797, n43798,
    n43799, n43800, n43801, n43802, n43803, n43804, n43805, n43806, n43807,
    n43808, n43809, n43810, n43811, n43812, n43813, n43814, n43815, n43816,
    n43817, n43818, n43819, n43820, n43821, n43822, n43823, n43824, n43825,
    n43826, n43827, n43828, n43829, n43830, n43831, n43832, n43833, n43834,
    n43835, n43836, n43837, n43838, n43839, n43840, n43841, n43842, n43843,
    n43844, n43845, n43846, n43847, n43848, n43849, n43850, n43851, n43852,
    n43853, n43854, n43855, n43856, n43857, n43858, n43859, n43860, n43861,
    n43862, n43863, n43864, n43865, n43866, n43867, n43868, n43869, n43870,
    n43871, n43872, n43873, n43874, n43875, n43876, n43877, n43878, n43879,
    n43880, n43881, n43882, n43883, n43884, n43885, n43886, n43887, n43888,
    n43889, n43891, n43892, n43893, n43894, n43895, n43896, n43897, n43898,
    n43899, n43900, n43901, n43902, n43903, n43904, n43905, n43906, n43907,
    n43908, n43909, n43910, n43911, n43912, n43913, n43914, n43915, n43916,
    n43917, n43918, n43919, n43920, n43921, n43922, n43923, n43924, n43925,
    n43926, n43927, n43928, n43929, n43930, n43931, n43932, n43933, n43934,
    n43935, n43936, n43937, n43938, n43939, n43940, n43941, n43942, n43943,
    n43944, n43945, n43946, n43947, n43948, n43949, n43950, n43951, n43952,
    n43954, n43955, n43956, n43957, n43958, n43959, n43960, n43961, n43962,
    n43963, n43964, n43965, n43966, n43967, n43968, n43969, n43970, n43971,
    n43972, n43973, n43974, n43975, n43976, n43977, n43978, n43979, n43980,
    n43981, n43982, n43983, n43984, n43985, n43986, n43987, n43988, n43989,
    n43990, n43991, n43992, n43993, n43995, n43996, n43997, n43998, n43999,
    n44000, n44001, n44002, n44003, n44004, n44005, n44006, n44007, n44008,
    n44009, n44010, n44011, n44012, n44013, n44014, n44015, n44016, n44017,
    n44018, n44019, n44020, n44021, n44022, n44023, n44024, n44025, n44026,
    n44027, n44028, n44029, n44030, n44031, n44032, n44033, n44034, n44035,
    n44036, n44037, n44038, n44039, n44040, n44041, n44042, n44043, n44044,
    n44045, n44046, n44047, n44048, n44049, n44050, n44051, n44052, n44053,
    n44054, n44055, n44056, n44057, n44058, n44059, n44060, n44061, n44062,
    n44063, n44064, n44065, n44066, n44067, n44069, n44070, n44071, n44072,
    n44073, n44074, n44075, n44076, n44077, n44078, n44079, n44080, n44081,
    n44082, n44083, n44084, n44085, n44086, n44087, n44088, n44089, n44090,
    n44091, n44092, n44093, n44094, n44095, n44096, n44098, n44099, n44100,
    n44101, n44102, n44103, n44104, n44105, n44106, n44107, n44108, n44109,
    n44110, n44111, n44112, n44113, n44114, n44115, n44116, n44117, n44118,
    n44119, n44120, n44121, n44122, n44123, n44124, n44125, n44126, n44127,
    n44128, n44129, n44130, n44131, n44132, n44133, n44134, n44135, n44136,
    n44137, n44138, n44139, n44141, n44142, n44143, n44144, n44145, n44146,
    n44147, n44148, n44149, n44150, n44151, n44152, n44153, n44154, n44155,
    n44156, n44157, n44158, n44159, n44160, n44161, n44162, n44163, n44164,
    n44165, n44166, n44167, n44168, n44169, n44170, n44171, n44172, n44173,
    n44174, n44175, n44176, n44177, n44178, n44179, n44180, n44181, n44182,
    n44183, n44184, n44185, n44186, n44187, n44188, n44189, n44190, n44191,
    n44192, n44193, n44194, n44195, n44196, n44197, n44198, n44199, n44200,
    n44201, n44202, n44203, n44204, n44205, n44206, n44207, n44208, n44210,
    n44211, n44212, n44213, n44214, n44215, n44216, n44217, n44218, n44219,
    n44220, n44221, n44222, n44223, n44224, n44225, n44226, n44227, n44228,
    n44229, n44230, n44231, n44232, n44233, n44234, n44235, n44236, n44237,
    n44238, n44239, n44240, n44241, n44242, n44243, n44244, n44245, n44246,
    n44247, n44248, n44249, n44250, n44251, n44252, n44253, n44254, n44255,
    n44256, n44257, n44258, n44259, n44260, n44261, n44262, n44263, n44264,
    n44265, n44266, n44267, n44269, n44270, n44271, n44272, n44273, n44274,
    n44275, n44276, n44277, n44278, n44279, n44280, n44281, n44282, n44283,
    n44284, n44285, n44286, n44287, n44288, n44289, n44290, n44291, n44292,
    n44293, n44294, n44295, n44296, n44297, n44298, n44299, n44300, n44301,
    n44302, n44303, n44304, n44305, n44306, n44307, n44308, n44309, n44310,
    n44311, n44313, n44314, n44315, n44316, n44317, n44318, n44319, n44320,
    n44321, n44322, n44323, n44324, n44325, n44326, n44327, n44328, n44329,
    n44330, n44331, n44332, n44333, n44334, n44335, n44336, n44337, n44338,
    n44339, n44340, n44341, n44342, n44343, n44344, n44345, n44346, n44347,
    n44348, n44349, n44350, n44352, n44353, n44354, n44355, n44356, n44357,
    n44358, n44359, n44360, n44361, n44362, n44363, n44364, n44365, n44366,
    n44367, n44368, n44369, n44370, n44371, n44372, n44373, n44374, n44375,
    n44376, n44377, n44378, n44379, n44380, n44381, n44382, n44383, n44384,
    n44385, n44386, n44387, n44388, n44389, n44391, n44392, n44393, n44394,
    n44395, n44396, n44397, n44398, n44399, n44400, n44401, n44402, n44403,
    n44404, n44405, n44406, n44407, n44408, n44409, n44410, n44411, n44412,
    n44413, n44414, n44415, n44416, n44417, n44418, n44419, n44420, n44421,
    n44422, n44423, n44424, n44425, n44426, n44427, n44428, n44429, n44430,
    n44431, n44432, n44433, n44434, n44435, n44436, n44437, n44438, n44439,
    n44440, n44441, n44442, n44443, n44444, n44445, n44446, n44447, n44448,
    n44450, n44451, n44452, n44454, n44455, n44456, n44457, n44458, n44459,
    n44460, n44461, n44462, n44463, n44464, n44465, n44466, n44467, n44468,
    n44469, n44470, n44472, n44473, n44474, n44475, n44476, n44477, n44478,
    n44479, n44480, n44481, n44482, n44483, n44484, n44485, n44486, n44487,
    n44488, n44490, n44492, n44493, n44495, n44496, n44497, n44499, n44500,
    n44501, n44502, n44503, n44504, n44505, n44506, n44507, n44508, n44509,
    n44510, n44511, n44512, n44514, n44515, n44517, n44518, n44520, n44521,
    n44523, n44524, n44526, n44527, n44529, n44530, n44532, n44533, n44535,
    n44536, n44538, n44539, n44541, n44542, n44543, n44544, n44545, n44546,
    n44547, n44549, n44550, n44551, n44552, n44553, n44554, n44556, n44557,
    n44558, n44560, n44561, n44562, n44563, n44564, n44565, n44566, n44567,
    n44568, n44569, n44570, n44571, n44572, n44573, n44574, n44575, n44576,
    n44577, n44578, n44579, n44580, n44582, n44583, n44585, n44586, n44588,
    n44589, n44591, n44592, n44594, n44595, n44597, n44598, n44600, n44601,
    n44603, n44604, n44605, n44606, n44607, n44608, n44609, n44610, n44611,
    n44612, n44613, n44614, n44615, n44616, n44617, n44618, n44619, n44620,
    n44621, n44622, n44623, n44624, n44625, n44626, n44627, n44628, n44630,
    n44631, n44632, n44634, n44635, n44637, n44638, n44639, n44641, n44642,
    n44644, n44645, n44646, n44647, n44648, n44649, n44650, n44651, n44652,
    n44653, n44654, n44656, n44657, n44658, n44659, n44661, n44662, n44664,
    n44665, n44666, n44668, n44669, n44670, n44671, n44673, n44674, n44676,
    n44677, n44679, n44680, n44682, n44683, n44685, n44686, n44688, n44689,
    n44691, n44692, n44694, n44695, n44697, n44698, n44700, n44701, n44703,
    n44704, n44706, n44707, n44708, n44709, n44710, n44711, n44712, n44714,
    n44715, n44716, n44717, n44719, n44720, n44721, n44722, n44723, n44724,
    n44725, n44726, n44727, n44728, n44729, n44731, n44732, n44734, n44735,
    n44737, n44738, n44740, n44741, n44743, n44744, n44746, n44747, n44749,
    n44750, n44752, n44753, n44754, n44755, n44756, n44758, n44759, n44761,
    n44762, n44764, n44765, n44767, n44768, n44770, n44771, n44773, n44774,
    n44776, n44777, n44779, n44780, n44782, n44783, n44785, n44786, n44788,
    n44789, n44791, n44792, n44794, n44795, n44797, n44798, n44800, n44801,
    n44803, n44804, n44806, n44807, n44809, n44810, n44812, n44813, n44815,
    n44816, n44818, n44819, n44821, n44822, n44824, n44825, n44827, n44828,
    n44830, n44831, n44833, n44834, n44836, n44837, n44839, n44840, n44842,
    n44843, n44845, n44846, n44848, n44849, n44851, n44852, n44854, n44855,
    n44857, n44858, n44860, n44861, n44863, n44864, n44866, n44867, n44869,
    n44870, n44872, n44873, n44875, n44876, n44878, n44879, n44881, n44882,
    n44884, n44885, n44887, n44888, n44890, n44891, n44893, n44894, n44896,
    n44897, n44899, n44900, n44902, n44903, n44905, n44906, n44908, n44909,
    n44911, n44912, n44914, n44915, n44917, n44918, n44920, n44921, n44923,
    n44924, n44926, n44927, n44929, n44930, n44932, n44933, n44935, n44936,
    n44938, n44939, n44941, n44942, n44944, n44945, n44947, n44948, n44950,
    n44951, n44953, n44954, n44956, n44957, n44959, n44960, n44962, n44963,
    n44965, n44966, n44968, n44969, n44971, n44972, n44974, n44975, n44977,
    n44978, n44979, n44981, n44982, n44984, n44985, n44987, n44988, n44990,
    n44991, n44993, n44994, n44996, n44997, n44999, n45000, n45002, n45003,
    n45005, n45006, n45008, n45009, n45011, n45012, n45014, n45015, n45017,
    n45018, n45020, n45021, n45023, n45024, n45026, n45027, n45029, n45030,
    n45032, n45033, n45035, n45036, n45038, n45039, n45041, n45042, n45044,
    n45045, n45047, n45048, n45050, n45051, n45053, n45054, n45056, n45057,
    n45059, n45060, n45062, n45063, n45065, n45066, n45068, n45069, n45071,
    n45072, n45074, n45075, n45077, n45078, n45080, n45081, n45083, n45084,
    n45086, n45087, n45089, n45090, n45092, n45093, n45095, n45096, n45098,
    n45099, n45101, n45102, n45104, n45105, n45107, n45108, n45109, n45110,
    n45111, n45112, n45113, n45114, n45115, n45116, n45117, n45118, n45119,
    n45120, n45121, n45122, n45123, n45124, n45125, n45126, n45127, n45128,
    n45129, n45131, n45132, n45134, n45135, n45137, n45138, n45140, n45141,
    n45143, n45144, n45146, n45147, n45149, n45150, n45152, n45153, n45154,
    n45155, n45156, n45157, n45158, n45159, n45160, n45161, n45162, n45163,
    n45164, n45165, n45166, n45167, n45168, n45169, n45170, n45171, n45172,
    n45173, n45174, n45175, n45177, n45178, n45179, n45180, n45181, n45182,
    n45183, n45184, n45185, n45186, n45187, n45188, n45189, n45190, n45191,
    n45192, n45193, n45195, n45196, n45197, n45198, n45199, n45200, n45201,
    n45202, n45203, n45204, n45205, n45206, n45207, n45208, n45209, n45210,
    n45211, n45212, n45213, n45214, n45215, n45216, n45217, n45218, n45219,
    n45220, n45221, n45222, n45223, n45225, n45226, n45227, n45228, n45229,
    n45231, n45232, n45233, n45234, n45235, n45236, n45237, n45238, n45239,
    n45240, n45241, n45242, n45243, n45244, n45245, n45246, n45247, n45248,
    n45249, n45251, n45252, n45253, n45254, n45255, n45256, n45257, n45258,
    n45259, n45260, n45261, n45262, n45263, n45264, n45265, n45266, n45267,
    n45268, n45269, n45271, n45272, n45273, n45274, n45275, n45276, n45277,
    n45278, n45279, n45280, n45281, n45282, n45283, n45284, n45285, n45286,
    n45287, n45288, n45289, n45291, n45292, n45293, n45294, n45295, n45296,
    n45297, n45298, n45299, n45300, n45301, n45302, n45303, n45304, n45305,
    n45306, n45307, n45308, n45309, n45311, n45312, n45313, n45314, n45315,
    n45316, n45317, n45318, n45319, n45320, n45322, n45323, n45324, n45325,
    n45326, n45327, n45328, n45329, n45330, n45331, n45333, n45334, n45335,
    n45336, n45337, n45338, n45339, n45340, n45341, n45342, n45344, n45345,
    n45346, n45347, n45348, n45349, n45350, n45351, n45352, n45353, n45354,
    n45357, n45358, n45360, n45361, n45363, n45364, n45366, n45367, n45369,
    n45370, n45372, n45373, n45375, n45376, n45378, n45379, n45381, n45382,
    n45384, n45385, n45387, n45388, n45390, n45391, n45393, n45394, n45396,
    n45397, n45399, n45400, n45402, n45403, n45405, n45406, n45408, n45409,
    n45411, n45412, n45414, n45415, n45417, n45418, n45420, n45421, n45423,
    n45424, n45426, n45427, n45429, n45430, n45431, n45432, n45433, n45434,
    n45435, n45436, n45438, n45439, n45441, n45442, n45444, n45445, n45447,
    n45448, n45450, n45451, n45453, n45454, n45455, n45456, n45457, n45459,
    n45460, n45462, n45463, n45465, n45466, n45468, n45469, n45471, n45472,
    n45474, n45475, n45477, n45478, n45479, n45480, n45481, n45483, n45484,
    n45486, n45487, n45489, n45490, n45492, n45493, n45495, n45496, n45497,
    n45498, n45500, n45501, n45503, n45504, n45506, n45507, n45509, n45510,
    n45512, n45513, n45515, n45516, n45518, n45519, n45521, n45522, n45524,
    n45525, n45527, n45528, n45530, n45531, n45533, n45534, n45536, n45537,
    n45539, n45540, n45542, n45543, n45545, n45546, n45548, n45549, n45551,
    n45552, n45554, n45555, n45557, n45558, n45560, n45561, n45562, n45563,
    n45565, n45566, n45568, n45569, n45571, n45572, n45574, n45575, n45577,
    n45578, n45580, n45581, n45583, n45584, n45586, n45587, n45589, n45590,
    n45592, n45593, n45595, n45596, n45598, n45599, n45601, n45602, n45603,
    n45604, n45606, n45607, n45609, n45610, n45612, n45613, n45615, n45616,
    n45618, n45619, n45621, n45622, n45624, n45625, n45627, n45628, n45630,
    n45631, n45633, n45634, n45635, n45636, n45637, n45638, n45639, n45640,
    n45641, n45642, n45643, n45644, n45645, n45646, n45647, n45648, n45649,
    n45650, n45651, n45652, n45653, n45654, n45655, n45656, n45657, n45658,
    n45659, n45660, n45661, n45662, n45663, n45664, n45665, n45666, n45667,
    n45668, n45669, n45670, n45671, n45672, n45673, n45674, n45675, n45676,
    n45677, n45678, n45679, n45680, n45681, n45682, n45683, n45684, n45685,
    n45686, n45687, n45688, n45689, n45690, n45691, n45692, n45693, n45694,
    n45695, n45696, n45697, n45698, n45699, n45700, n45701, n45702, n45703,
    n45704, n45705, n45706, n45707, n45708, n45709, n45710, n45711, n45712,
    n45713, n45714, n45715, n45716, n45717, n45718, n45719, n45720, n45721,
    n45722, n45723, n45724, n45725, n45726, n45727, n45728, n45729, n45730,
    n45731, n45732, n45733, n45734, n45735, n45736, n45737, n45738, n45739,
    n45740, n45741, n45742, n45744, n45745, n45747, n45748, n45750, n45751,
    n45752, n45753, n45755, n45756, n45758, n45759, n45761, n45762, n45764,
    n45765, n45767, n45768, n45770, n45771, n45773, n45774, n45776, n45777,
    n45779, n45780, n45782, n45783, n45785, n45786, n45788, n45789, n45791,
    n45792, n45794, n45795, n45797, n45798, n45800, n45801, n45802, n45803,
    n45804, n45805, n45807, n45808, n45809, n45810, n45812, n45813, n45814,
    n45815, n45816, n45817, n45818, n45819, n45820, n45821, n45822, n45823,
    n45824, n45825, n45826, n45827, n45828, n45829, n45830, n45831, n45833,
    n45834, n45835, n45837, n45838, n45839, n45841, n45842, n45843, n45845,
    n45846, n45847, n45848, n45849, n45850, n45851, n45852, n45853, n45854,
    n45855, n45856, n45857, n45858, n45859, n45860, n45861, n45862, n45863,
    n45864, n45865, n45866, n45867, n45868, n45869, n45870, n45871, n45872,
    n45873, n45874, n45875, n45876, n45877, n45878, n45879, n45880, n45881,
    n45882, n45883, n45884, n45885, n45886, n45887, n45888, n45889, n45890,
    n45891, n45892, n45893, n45894, n45895, n45896, n45897, n45898, n45899,
    n45900, n45901, n45902, n45903, n45904, n45905, n45906, n45907, n45908,
    n45909, n45910, n45911, n45912, n45913, n45914, n45915, n45916, n45917,
    n45918, n45919, n45920, n45921, n45922, n45923, n45924, n45925, n45926,
    n45927, n45928, n45929, n45930, n45931, n45932, n45933, n45934, n45935,
    n45936, n45937, n45938, n45939, n45940, n45941, n45942, n45943, n45944,
    n45945, n45946, n45947, n45948, n45949, n45950, n45951, n45952, n45953,
    n45954, n45955, n45956, n45957, n45958, n45959, n45960, n45961, n45962,
    n45963, n45964, n45965, n45966, n45967, n45968, n45969, n45970, n45971,
    n45972, n45973, n45974, n45975, n45976, n45977, n45978, n45979, n45980,
    n45981, n45982, n45983, n45984, n45985, n45986, n45987, n45988, n45989,
    n45990, n45991, n45992, n45993, n45994, n45995, n45996, n45997, n45998,
    n45999, n46000, n46001, n46002, n46003, n46004, n46005, n46006, n46007,
    n46008, n46009, n46010, n46011, n46012, n46013, n46014, n46015, n46016,
    n46017, n46018, n46019, n46020, n46021, n46022, n46023, n46024, n46025,
    n46026, n46027, n46028, n46029, n46030, n46031, n46032, n46033, n46034,
    n46035, n46036, n46037, n46038, n46039, n46040, n46041, n46042, n46043,
    n46044, n46045, n46046, n46047, n46048, n46049, n46050, n46051, n46052,
    n46053, n46054, n46055, n46056, n46057, n46058, n46059, n46060, n46061,
    n46062, n46063, n46064, n46065, n46066, n46067, n46068, n46069, n46070,
    n46071, n46072, n46073, n46074, n46075, n46076, n46077, n46078, n46079,
    n46080, n46081, n46082, n46083, n46084, n46085, n46086, n46087, n46088,
    n46089, n46090, n46091, n46092, n46093, n46094, n46095, n46096, n46097,
    n46098, n46099, n46100, n46101, n46102, n46103, n46104, n46105, n46106,
    n46107, n46108, n46109, n46110, n46111, n46112, n46113, n46114, n46115,
    n46116, n46117, n46118, n46119, n46120, n46121, n46122, n46123, n46124,
    n46125, n46126, n46127, n46128, n46129, n46130, n46131, n46132, n46133,
    n46134, n46135, n46136, n46137, n46138, n46139, n46140, n46141, n46142,
    n46143, n46144, n46145, n46146, n46147, n46148, n46149, n46150, n46151,
    n46152, n46153, n46154, n46155, n46156, n46157, n46158, n46159, n46160,
    n46161, n46162, n46163, n46164, n46165, n46166, n46167, n46168, n46169,
    n46170, n46171, n46172, n46173, n46174, n46175, n46176, n46177, n46178,
    n46179, n46180, n46181, n46182, n46183, n46184, n46185, n46186, n46187,
    n46188, n46189, n46190, n46191, n46192, n46193, n46194, n46195, n46196,
    n46197, n46198, n46199, n46200, n46201, n46202, n46203, n46204, n46205,
    n46206, n46207, n46208, n46209, n46210, n46211, n46212, n46213, n46214,
    n46215, n46216, n46217, n46218, n46219, n46220, n46221, n46222, n46223,
    n46224, n46225, n46226, n46227, n46228, n46229, n46230, n46231, n46232,
    n46233, n46234, n46235, n46236, n46237, n46238, n46239, n46240, n46241,
    n46242, n46243, n46244, n46245, n46246, n46247, n46248, n46249, n46250,
    n46251, n46252, n46253, n46254, n46255, n46256, n46257, n46258, n46259,
    n46260, n46261, n46262, n46263, n46264, n46265, n46266, n46267, n46268,
    n46269, n46270, n46271, n46272, n46273, n46274, n46275, n46276, n46277,
    n46278, n46279, n46280, n46281, n46282, n46283, n46284, n46285, n46286,
    n46287, n46288, n46289, n46290, n46291, n46292, n46293, n46294, n46295,
    n46296, n46297, n46298, n46299, n46300, n46301, n46302, n46303, n46304,
    n46305, n46306, n46307, n46308, n46309, n46310, n46311, n46312, n46313,
    n46314, n46315, n46316, n46317, n46318, n46319, n46320, n46321, n46322,
    n46323, n46324, n46325, n46326, n46327, n46328, n46329, n46330, n46331,
    n46332, n46333, n46334, n46335, n46336, n46337, n46338, n46339, n46340,
    n46341, n46342, n46343, n46344, n46345, n46346, n46347, n46348, n46349,
    n46350, n46351, n46352, n46353, n46354, n46355, n46356, n46357, n46358,
    n46359, n46360, n46361, n46362, n46363, n46364, n46365, n46366, n46367,
    n46368, n46369, n46370, n46371, n46372, n46373, n46374, n46375, n46376,
    n46377, n46378, n46379, n46380, n46381, n46382, n46383, n46384, n46385,
    n46386, n46387, n46388, n46389, n46390, n46391, n46392, n46393, n46394,
    n46395, n46396, n46397, n46398, n46399, n46400, n46401, n46402, n46403,
    n46404, n46405, n46406, n46407, n46408, n46409, n46410, n46411, n46412,
    n46413, n46414, n46415, n46416, n46417, n46418, n46419, n46420, n46421,
    n46422, n46423, n46424, n46425, n46426, n46427, n46428, n46429, n46430,
    n46431, n46432, n46433, n46434, n46435, n46436, n46437, n46438, n46439,
    n46440, n46441, n46442, n46443, n46444, n46445, n46446, n46447, n46448,
    n46449, n46450, n46451, n46452, n46453, n46454, n46455, n46456, n46457,
    n46458, n46459, n46460, n46461, n46462, n46463, n46464, n46465, n46466,
    n46467, n46468, n46469, n46470, n46471, n46472, n46473, n46474, n46475,
    n46476, n46477, n46478, n46479, n46480, n46481, n46482, n46483, n46484,
    n46485, n46486, n46487, n46488, n46489, n46490, n46491, n46492, n46493,
    n46494, n46495, n46496, n46497, n46498, n46499, n46500, n46501, n46502,
    n46503, n46504, n46505, n46506, n46507, n46508, n46509, n46510, n46511,
    n46512, n46513, n46514, n46515, n46516, n46517, n46518, n46519, n46520,
    n46521, n46522, n46523, n46524, n46525, n46526, n46527, n46528, n46529,
    n46530, n46531, n46532, n46533, n46534, n46535, n46536, n46537, n46538,
    n46539, n46540, n46541, n46542, n46543, n46544, n46545, n46546, n46547,
    n46548, n46549, n46550, n46551, n46552, n46553, n46554, n46555, n46556,
    n46557, n46558, n46559, n46560, n46561, n46562, n46563, n46564, n46565,
    n46566, n46567, n46568, n46569, n46570, n46571, n46572, n46573, n46574,
    n46575, n46576, n46577, n46578, n46579, n46580, n46581, n46582, n46583,
    n46584, n46585, n46586, n46587, n46588, n46589, n46590, n46591, n46592,
    n46593, n46594, n46595, n46596, n46597, n46598, n46599, n46600, n46601,
    n46602, n46603, n46604, n46605, n46606, n46607, n46608, n46609, n46610,
    n46611, n46612, n46613, n46614, n46615, n46616, n46617, n46618, n46619,
    n46620, n46621, n46622, n46623, n46624, n46625, n46626, n46627, n46628,
    n46629, n46630, n46631, n46632, n46633, n46634, n46635, n46636, n46637,
    n46638, n46639, n46640, n46641, n46642, n46643, n46644, n46645, n46646,
    n46647, n46648, n46649, n46650, n46651, n46652, n46653, n46654, n46655,
    n46656, n46657, n46658, n46659, n46660, n46661, n46662, n46663, n46664,
    n46665, n46666, n46667, n46668, n46669, n46670, n46671, n46672, n46673,
    n46674, n46675, n46676, n46677, n46678, n46679, n46680, n46681, n46682,
    n46683, n46684, n46685, n46686, n46687, n46688, n46689, n46690, n46691,
    n46692, n46693, n46694, n46695, n46696, n46697, n46698, n46699, n46700,
    n46701, n46702, n46703, n46704, n46705, n46706, n46707, n46708, n46709,
    n46710, n46711, n46712, n46713, n46714, n46715, n46716, n46717, n46718,
    n46719, n46720, n46721, n46722, n46724, n46725, n46726, n46727, n46728,
    n46729, n46731, n46732, n46733, n46734, n46735, n46737, n46738, n46739,
    n46740, n46741, n46743, n46744, n46745, n46747, n46748, n46749, n46750,
    n46751, n46753, n46754, n46755, n46757, n46758, n46760, n46761, n46762,
    n46764, n46765, n46766, n46767, n46768, n46769, n46770, n46771, n46772,
    n46773, n46774, n46776, n46777, n46778, n46779, n46780, n46781, n46782,
    n46783, n46785, n46786, n46787, n46788, n46790, n46791, n46792, n46793,
    n46794, n46795, n46797, n46798, n46800, n46801, n46802, n46803, n46804,
    n46806, n46807, n46808, n46810, n46811, n46812, n46814, n46815, n46816,
    n46818, n46819, n46820, n46822, n46823, n46824, n46826, n46827, n46828,
    n46830, n46831, n46832, n46834, n46835, n46836, n46837, n46839, n46840,
    n46841, n46842, n46844, n46845, n46846, n46847, n46849, n46850, n46851,
    n46852, n46853, n46855, n46856, n46857, n46859, n46860, n46861, n46863,
    n46864, n46865, n46867, n46868, n46869, n46871, n46872, n46873, n46875,
    n46876, n46877, n46879, n46880, n46881, n46882, n46883, n46885, n46886,
    n46887, n46888, n46890, n46891, n46892, n46894, n46895, n46896, n46898,
    n46899, n46900, n46902, n46903, n46904, n46906, n46907, n46908, n46910,
    n46911, n46912, n46914, n46915, n46916, n46918, n46919, n46920, n46922,
    n46923, n46924, n46926, n46927, n46928, n46930, n46931, n46932, n46934,
    n46935, n46936, n46938, n46939, n46940, n46942, n46943, n46944, n46946,
    n46947, n46948, n46950, n46951, n46952, n46954, n46955, n46956, n46958,
    n46959, n46960, n46962, n46963, n46964, n46966, n46967, n46968, n46970,
    n46971, n46972, n46974, n46975, n46976, n46978, n46979, n46980, n46982,
    n46983, n46984, n46986, n46987, n46988, n46990, n46991, n46992, n46994,
    n46995, n46996, n46998, n46999, n47000, n47002, n47003, n47004, n47006,
    n47007, n47008, n47010, n47011, n47012, n47014, n47015, n47016, n47018,
    n47019, n47020, n47022, n47023, n47024, n47026, n47027, n47028, n47029,
    n47030, n47031, n47032, n47033, n47034, n47036, n47038, n47039, n47040,
    n47042, n47043, n47044, n47046, n47047, n47048, n47050, n47051, n47052,
    n47053, n47054, n47055, n47056, n47057, n47058, n47059, n47060, n47061,
    n47062, n47063, n47064, n47065, n47066, n47067, n47068, n47069, n47070,
    n47071, n47072, n47073, n47074, n47075, n47076, n47077, n47078, n47079,
    n47080, n47081, n47082, n47083, n47084, n47085, n47086, n47087, n47088,
    n47089, n47090, n47091, n47092, n47093, n47094, n47095, n47096, n47097,
    n47099, n47100, n47101, n47102, n47103, n47104, n47105, n47106, n47107,
    n47108, n47109, n47110, n47111, n47112, n47113, n47114, n47115, n47116,
    n47117, n47118, n47119, n47120, n47121, n47122, n47123, n47124, n47125,
    n47126, n47127, n47128, n47129, n47130, n47131, n47132, n47133, n47134,
    n47135, n47136, n47137, n47138, n47139, n47141, n47142, n47143, n47145,
    n47146, n47147, n47148, n47149, n47150, n47151, n47152, n47153, n47154,
    n47155, n47156, n47157, n47158, n47159, n47160, n47161, n47162, n47163,
    n47164, n47165, n47166, n47167, n47168, n47169, n47170, n47171, n47172,
    n47173, n47174, n47175, n47176, n47177, n47178, n47179, n47181, n47182,
    n47183, n47184, n47185, n47186, n47187, n47188, n47189, n47190, n47191,
    n47192, n47193, n47194, n47195, n47196, n47197, n47198, n47199, n47200,
    n47201, n47202, n47203, n47204, n47205, n47206, n47207, n47208, n47209,
    n47210, n47211, n47212, n47213, n47214, n47215, n47216, n47218, n47219,
    n47220, n47221, n47222, n47223, n47224, n47225, n47226, n47227, n47228,
    n47229, n47230, n47231, n47232, n47233, n47234, n47235, n47236, n47237,
    n47238, n47239, n47240, n47241, n47242, n47243, n47244, n47245, n47246,
    n47247, n47248, n47249, n47250, n47251, n47252, n47254, n47255, n47256,
    n47258, n47259, n47260, n47261, n47262, n47263, n47264, n47265, n47266,
    n47267, n47268, n47269, n47270, n47271, n47272, n47273, n47274, n47275,
    n47276, n47277, n47278, n47279, n47280, n47281, n47282, n47283, n47284,
    n47285, n47286, n47287, n47288, n47289, n47291, n47292, n47293, n47294,
    n47295, n47296, n47297, n47298, n47299, n47300, n47301, n47302, n47303,
    n47304, n47305, n47306, n47307, n47308, n47309, n47310, n47311, n47312,
    n47313, n47314, n47315, n47316, n47317, n47318, n47319, n47320, n47321,
    n47323, n47324, n47325, n47326, n47327, n47328, n47329, n47330, n47331,
    n47332, n47333, n47334, n47335, n47336, n47337, n47338, n47339, n47340,
    n47341, n47342, n47343, n47344, n47345, n47346, n47347, n47348, n47349,
    n47350, n47351, n47352, n47353, n47354, n47355, n47356, n47357, n47359,
    n47360, n47361, n47362, n47363, n47364, n47365, n47366, n47367, n47368,
    n47369, n47370, n47371, n47372, n47373, n47374, n47375, n47376, n47377,
    n47378, n47379, n47380, n47381, n47382, n47383, n47384, n47385, n47386,
    n47387, n47388, n47389, n47390, n47391, n47392, n47393, n47395, n47396,
    n47397, n47398, n47399, n47400, n47401, n47402, n47403, n47404, n47405,
    n47406, n47407, n47408, n47409, n47410, n47411, n47412, n47413, n47414,
    n47415, n47416, n47417, n47418, n47419, n47420, n47421, n47422, n47423,
    n47424, n47425, n47426, n47427, n47428, n47429, n47430, n47431, n47433,
    n47434, n47435, n47436, n47437, n47438, n47439, n47440, n47441, n47442,
    n47443, n47444, n47445, n47446, n47447, n47448, n47449, n47450, n47451,
    n47452, n47453, n47454, n47455, n47456, n47457, n47458, n47459, n47460,
    n47461, n47462, n47463, n47464, n47465, n47466, n47467, n47469, n47470,
    n47471, n47472, n47473, n47474, n47475, n47476, n47477, n47478, n47479,
    n47480, n47481, n47482, n47483, n47484, n47485, n47486, n47487, n47488,
    n47489, n47490, n47491, n47492, n47493, n47494, n47495, n47496, n47497,
    n47498, n47499, n47500, n47501, n47502, n47503, n47505, n47506, n47507,
    n47508, n47509, n47510, n47511, n47512, n47513, n47514, n47515, n47516,
    n47517, n47518, n47519, n47520, n47521, n47522, n47523, n47524, n47525,
    n47526, n47527, n47528, n47529, n47530, n47531, n47532, n47533, n47534,
    n47535, n47537, n47538, n47539, n47540, n47541, n47542, n47543, n47544,
    n47545, n47546, n47547, n47548, n47549, n47550, n47551, n47552, n47553,
    n47554, n47555, n47556, n47557, n47558, n47559, n47560, n47561, n47562,
    n47563, n47564, n47565, n47566, n47567, n47569, n47570, n47571, n47572,
    n47573, n47574, n47575, n47576, n47577, n47578, n47579, n47580, n47581,
    n47582, n47583, n47584, n47585, n47586, n47587, n47588, n47589, n47590,
    n47591, n47592, n47593, n47594, n47595, n47596, n47597, n47598, n47599,
    n47600, n47601, n47602, n47603, n47604, n47606, n47607, n47608, n47610,
    n47611, n47612, n47614, n47615, n47616, n47617, n47618, n47619, n47620,
    n47621, n47622, n47623, n47624, n47625, n47626, n47627, n47628, n47629,
    n47630, n47631, n47632, n47633, n47634, n47635, n47636, n47637, n47638,
    n47639, n47640, n47641, n47642, n47643, n47644, n47647, n47648, n47649,
    n47651, n47652, n47653, n47654, n47655, n47656, n47657, n47658, n47659,
    n47660, n47661, n47662, n47663, n47664, n47665, n47666, n47667, n47668,
    n47669, n47670, n47671, n47672, n47673, n47674, n47675, n47676, n47677,
    n47678, n47679, n47680, n47681, n47682, n47683, n47684, n47685, n47686,
    n47687, n47688, n47689, n47691, n47692, n47693, n47695, n47696, n47697,
    n47699, n47700, n47701, n47703, n47704, n47705, n47706, n47707, n47708,
    n47709, n47710, n47711, n47712, n47713, n47714, n47715, n47716, n47717,
    n47718, n47719, n47720, n47721, n47722, n47723, n47724, n47725, n47726,
    n47727, n47728, n47729, n47730, n47731, n47732, n47733, n47734, n47735,
    n47737, n47738, n47739, n47741, n47742, n47743, n47745, n47746, n47747,
    n47748, n47749, n47750, n47751, n47752, n47753, n47754, n47755, n47756,
    n47757, n47758, n47759, n47760, n47761, n47762, n47763, n47764, n47765,
    n47766, n47767, n47768, n47769, n47770, n47771, n47772, n47773, n47774,
    n47775, n47776, n47777, n47778, n47780, n47781, n47782, n47784, n47785,
    n47786, n47788, n47789, n47790, n47792, n47793, n47794, n47796, n47797,
    n47798, n47800, n47801, n47802, n47804, n47805, n47806, n47808, n47809,
    n47810, n47812, n47813, n47814, n47816, n47817, n47818, n47820, n47821,
    n47822, n47824, n47825, n47826, n47828, n47829, n47830, n47832, n47833,
    n47834, n47836, n47837, n47838, n47839, n47840, n47841, n47842, n47843,
    n47844, n47845, n47846, n47847, n47848, n47849, n47850, n47851, n47852,
    n47853, n47854, n47855, n47856, n47857, n47858, n47859, n47860, n47861,
    n47862, n47863, n47864, n47865, n47866, n47867, n47868, n47869, n47870,
    n47872, n47873, n47874, n47875, n47876, n47877, n47878, n47879, n47880,
    n47881, n47882, n47883, n47884, n47885, n47886, n47887, n47888, n47889,
    n47890, n47891, n47892, n47893, n47894, n47895, n47896, n47897, n47898,
    n47899, n47900, n47901, n47902, n47903, n47904, n47905, n47906, n47907,
    n47908, n47909, n47910, n47912, n47913, n47914, n47916, n47917, n47918,
    n47920, n47921, n47922, n47923, n47924, n47925, n47926, n47927, n47928,
    n47929, n47930, n47931, n47932, n47933, n47934, n47935, n47936, n47937,
    n47938, n47939, n47940, n47941, n47942, n47943, n47944, n47945, n47946,
    n47947, n47948, n47949, n47950, n47951, n47952, n47954, n47955, n47956,
    n47957, n47958, n47959, n47960, n47961, n47962, n47963, n47964, n47965,
    n47966, n47967, n47968, n47969, n47970, n47971, n47972, n47973, n47974,
    n47975, n47976, n47977, n47978, n47979, n47980, n47981, n47982, n47983,
    n47984, n47985, n47986, n47987, n47989, n47990, n47991, n47992, n47993,
    n47994, n47995, n47996, n47997, n47998, n47999, n48000, n48001, n48002,
    n48003, n48004, n48005, n48006, n48007, n48008, n48009, n48010, n48011,
    n48012, n48013, n48014, n48015, n48016, n48017, n48018, n48019, n48020,
    n48021, n48023, n48024, n48025, n48026, n48027, n48028, n48029, n48030,
    n48031, n48032, n48033, n48034, n48035, n48036, n48037, n48038, n48039,
    n48040, n48041, n48042, n48043, n48044, n48045, n48046, n48047, n48048,
    n48049, n48050, n48051, n48052, n48053, n48054, n48055, n48056, n48058,
    n48059, n48060, n48062, n48063, n48064, n48065, n48066, n48067, n48068,
    n48069, n48070, n48071, n48072, n48073, n48074, n48075, n48076, n48077,
    n48078, n48079, n48080, n48081, n48082, n48083, n48084, n48085, n48086,
    n48087, n48088, n48089, n48090, n48091, n48092, n48093, n48094, n48095,
    n48096, n48098, n48099, n48100, n48101, n48102, n48103, n48104, n48105,
    n48106, n48107, n48108, n48109, n48110, n48111, n48112, n48113, n48114,
    n48115, n48116, n48117, n48118, n48119, n48120, n48121, n48122, n48123,
    n48124, n48125, n48126, n48127, n48128, n48129, n48130, n48132, n48133,
    n48134, n48135, n48136, n48137, n48138, n48139, n48140, n48141, n48142,
    n48143, n48144, n48145, n48146, n48147, n48148, n48149, n48150, n48151,
    n48152, n48153, n48154, n48155, n48156, n48157, n48158, n48159, n48160,
    n48161, n48162, n48163, n48164, n48165, n48166, n48168, n48169, n48170,
    n48171, n48172, n48173, n48174, n48175, n48176, n48177, n48178, n48179,
    n48180, n48181, n48182, n48183, n48184, n48185, n48186, n48187, n48188,
    n48189, n48190, n48191, n48192, n48193, n48194, n48195, n48196, n48197,
    n48198, n48199, n48200, n48202, n48203, n48204, n48205, n48206, n48207,
    n48208, n48209, n48210, n48211, n48212, n48213, n48214, n48215, n48216,
    n48217, n48218, n48219, n48220, n48221, n48222, n48223, n48224, n48225,
    n48226, n48227, n48228, n48229, n48230, n48231, n48232, n48233, n48234,
    n48235, n48237, n48238, n48239, n48240, n48241, n48242, n48243, n48244,
    n48245, n48246, n48247, n48248, n48249, n48250, n48251, n48252, n48253,
    n48254, n48255, n48256, n48257, n48258, n48259, n48260, n48261, n48262,
    n48263, n48264, n48265, n48266, n48267, n48268, n48269, n48270, n48271,
    n48272, n48273, n48274, n48275, n48276, n48277, n48278, n48279, n48280,
    n48281, n48282, n48283, n48284, n48285, n48286, n48287, n48288, n48289,
    n48290, n48291, n48293, n48294, n48295, n48296, n48297, n48298, n48299,
    n48300, n48301, n48302, n48303, n48304, n48305, n48306, n48307, n48308,
    n48309, n48310, n48311, n48312, n48313, n48314, n48315, n48316, n48317,
    n48318, n48319, n48320, n48321, n48322, n48323, n48324, n48325, n48326,
    n48328, n48329, n48330, n48332, n48333, n48334, n48336, n48337, n48338,
    n48340, n48341, n48342, n48344, n48345, n48346, n48348, n48349, n48350,
    n48352, n48353, n48354, n48356, n48357, n48358, n48360, n48361, n48362,
    n48363, n48364, n48365, n48366, n48367, n48368, n48369, n48370, n48371,
    n48372, n48373, n48374, n48375, n48377, n48378, n48379, n48381, n48382,
    n48383, n48384, n48385, n48386, n48387, n48388, n48389, n48390, n48391,
    n48392, n48393, n48394, n48395, n48396, n48397, n48398, n48399, n48400,
    n48401, n48402, n48403, n48404, n48405, n48406, n48407, n48408, n48409,
    n48410, n48411, n48412, n48413, n48414, n48415, n48417, n48418, n48419,
    n48421, n48422, n48423, n48425, n48426, n48427, n48429, n48430, n48431,
    n48433, n48434, n48435, n48437, n48438, n48440, n48441, n48442, n48444,
    n48445, n48446, n48448, n48449, n48450, n48452, n48453, n48454, n48456,
    n48457, n48458, n48460, n48461, n48462, n48464, n48465, n48466, n48468,
    n48469, n48470, n48471, n48472, n48473, n48474, n48475, n48476, n48477,
    n48478, n48479, n48481, n48482, n48483, n48485, n48486, n48487, n48489,
    n48490, n48491, n48493, n48494, n48495, n48497, n48498, n48499, n48501,
    n48502, n48503, n48505, n48506, n48507, n48509, n48510, n48511, n48513,
    n48514, n48515, n48517, n48518, n48519, n48521, n48522, n48523, n48525,
    n48526, n48527, n48529, n48530, n48531, n48533, n48534, n48535, n48537,
    n48538, n48539, n48541, n48542, n48543, n48545, n48546, n48547, n48550,
    n48551, n48552, n48553, n48554, n48555, n48556, n48557, n48558, n48559,
    n48560, n48561, n48562, n48563, n48564, n48565, n48566, n48567, n48568,
    n48569, n48570, n48571, n48573, n48574, n48575, n48577, n48578, n48579,
    n48581, n48582, n48583, n48585, n48586, n48587, n48588, n48589, n48590,
    n48591, n48592, n48593, n48594, n48595, n48596, n48597, n48598, n48599,
    n48600, n48602, n48603, n48604, n48606, n48607, n48608, n48609, n48611,
    n48612, n48613, n48614, n48616, n48617, n48618, n48620, n48621, n48622,
    n48623, n48624, n48625, n48626, n48628, n48629, n48630, n48632, n48633,
    n48634, n48635, n48636, n48637, n48638, n48639, n48640, n48641, n48642,
    n48643, n48644, n48645, n48646, n48647, n48649, n48650, n48651, n48653,
    n48654, n48655, n48657, n48658, n48659, n48660, n48661, n48662, n48663,
    n48667, n48668, n48670, n48672, n48673, n48675, n48676, n48678, n48679,
    n48681, n48682, n48684, n48685, n48687, n48688, n48690, n48691, n48693,
    n48694, n48696, n48697, n48699, n48700, n48702, n48703, n48704, n48706,
    n48707, n48709, n48710, n48711, n48712, n48713, n48714, n48715, n48716,
    n48718, n48719, n48721, n48722, n48724, n48725, n48727, n48728, n48730,
    n48731, n48733, n48734, n48736, n48737, n48738, n48740, n48741, n48743,
    n48744, n48746, n48747, n48749, n48750, n48752, n48753, n48755, n48756,
    n48758, n48759, n48761, n48762, n48764, n48765, n48767, n48768, n48770,
    n48772, n48774, n48776, n48779, n48780, n48781, n48783, n48784, n48785,
    n48786, n48787, n48788, n48789, n48790, n48791, n48792, n48793, n48794,
    n48795, n48796, n48797, n48798, n48799, n48800, n48801, n48802, n48803,
    n48804, n48805, n48806, n48807, n48808, n48809, n48810, n48812, n48813,
    n48814, n48815, n48816, n48817, n48818, n48819, n48820, n48821, n48822,
    n48823, n48824, n48825, n48826, n48827, n48828, n48829, n48830, n48831,
    n48832, n48833, n48834, n48835, n48836, n48837, n48838, n48840, n48841,
    n48842, n48843, n48844, n48845, n48846, n48847, n48848, n48849, n48850,
    n48851, n48852, n48853, n48854, n48855, n48856, n48857, n48858, n48859,
    n48860, n48861, n48862, n48863, n48864, n48865, n48866, n48868, n48869,
    n48870, n48871, n48872, n48873, n48874, n48875, n48876, n48877, n48878,
    n48879, n48880, n48881, n48882, n48883, n48884, n48885, n48886, n48887,
    n48888, n48889, n48890, n48891, n48892, n48893, n48894, n48896, n48897,
    n48899, n48901, n48902, n48904, n48907, n48909, n48910, n48912, n48913,
    n48915, n48916, n48918, n48919, n48922, n48923, n48925, n48926, n48928,
    n48929, n48931, n48932, n48934, n48935, n48937, n48938, n48940, n48941,
    n48943, n48944, n48946, n48947, n48949, n48950, n48952, n48953, n48955,
    n48956, n48958, n48959, n48961, n48962, n48964, n48965, n48967, n48968,
    n48970, n48971, n48973, n48974, n48976, n48977, n48979, n48980, n48981,
    n48982, n48983, n48984, n48985, n48986, n48988, n48989, n48991, n48992,
    n48994, n48995, n48997, n48998, n49000, n49001, n49003, n49004, n49006,
    n49007, n49009, n49010, n49011, n49012, n49013, n49014, n49015, n49016,
    n49018, n49019, n49021, n49022, n49024, n49025, n49027, n49028, n49030,
    n49031, n49033, n49034, n49035, n49036, n49037, n49038, n49039, n49040,
    n49042, n49043, n49045, n49046, n49047, n49048, n49049, n49050, n49051,
    n49052, n49054, n49055, n49056, n49057, n49058, n49059, n49060, n49061,
    n49063, n49064, n49065, n49066, n49067, n49068, n49069, n49070, n49072,
    n49073, n49075, n49076, n49078, n49080, n49081, n49083, n49084, n49086,
    n49087, n49089, n49091, n49092, n49094, n49095, n49097, n49098, n49100,
    n49101, n49103, n49104, n49106, n49107, n49109, n49110, n49112, n49113,
    n49115, n49116, n49118, n49120, n49121, n49123, n49124, n49126, n49127,
    n49129, n49131, n49133, n49134, n49136, n49137, n49138, n49139, n49140,
    n49141, n49142, n49143, n49144, n49145, n49147, n49149, n49150, n49152,
    n49153, n49155, n49156, n49158, n49160, n49161, n49163, n49165, n49166,
    n49168, n49170, n49171, n49173, n49174, n49176, n49177, n49179, n49180,
    n49182, n49184, n49185, n49187, n49188, n49190, n49191, n49193, n49194,
    n49196, n49197, n49199, n49200, n49202, n49204, n49205, n49207, n49208,
    n49210, n49211, n49213, n49215, n49217, n49218, n49220, n49222, n49223,
    n49225, n49226, n49228, n49230, n49231, n49233, n49235, n49236, n49238,
    n49239, n49241, n49242, n49244, n49245, n49248, n49250, n49252, n49253,
    n49256;
  assign n2437 = ~pi0332 & ~pi1144;
  assign n2438 = pi0215 & ~n2437;
  assign n2439 = pi0265 & ~pi0332;
  assign n2440 = pi0216 & ~n2439;
  assign n2441 = pi0105 & pi0228;
  assign n2442 = pi0095 & ~pi0479;
  assign n2443 = pi0234 & n2442;
  assign n2444 = ~pi0332 & ~n2443;
  assign n2445 = n2441 & n2444;
  assign n2446 = pi0153 & ~pi0332;
  assign n2447 = ~n2441 & n2446;
  assign n2448 = ~pi0216 & ~n2447;
  assign n2449 = ~n2445 & n2448;
  assign n2450 = ~n2440 & ~n2449;
  assign n2451 = ~pi0221 & ~n2450;
  assign n2452 = ~pi0216 & pi0833;
  assign n2453 = pi1144 & ~n2452;
  assign n2454 = pi0929 & n2452;
  assign n2455 = ~pi0332 & ~n2453;
  assign n2456 = ~n2454 & n2455;
  assign n2457 = pi0221 & ~n2456;
  assign n2458 = ~n2451 & ~n2457;
  assign n2459 = ~pi0215 & ~n2458;
  assign n2460 = ~n2438 & ~n2459;
  assign n2461 = ~pi0058 & ~pi0090;
  assign n2462 = ~pi0088 & ~pi0098;
  assign n2463 = ~pi0077 & n2462;
  assign n2464 = ~pi0050 & n2463;
  assign n2465 = ~pi0102 & n2464;
  assign n2466 = ~pi0065 & ~pi0071;
  assign n2467 = ~pi0083 & ~pi0103;
  assign n2468 = ~pi0067 & ~pi0069;
  assign n2469 = ~pi0066 & ~pi0073;
  assign n2470 = ~pi0061 & ~pi0076;
  assign n2471 = ~pi0085 & ~pi0106;
  assign n2472 = n2470 & n2471;
  assign n2473 = ~pi0048 & n2472;
  assign n2474 = ~pi0089 & n2473;
  assign n2475 = ~pi0049 & n2474;
  assign n2476 = ~pi0104 & n2475;
  assign n2477 = ~pi0045 & n2476;
  assign n2478 = ~pi0068 & ~pi0084;
  assign n2479 = ~pi0082 & ~pi0111;
  assign n2480 = ~pi0036 & n2479;
  assign n2481 = n2478 & n2480;
  assign n2482 = n2477 & n2481;
  assign n2483 = n2469 & n2482;
  assign n2484 = n2468 & n2483;
  assign n2485 = n2467 & n2484;
  assign n2486 = n2466 & n2485;
  assign n2487 = ~pi0063 & ~pi0107;
  assign n2488 = n2486 & n2487;
  assign n2489 = ~pi0064 & n2488;
  assign n2490 = ~pi0081 & n2489;
  assign n2491 = n2465 & n2490;
  assign n2492 = ~pi0047 & ~pi0091;
  assign n2493 = ~pi0109 & ~pi0110;
  assign n2494 = ~pi0053 & ~pi0060;
  assign n2495 = ~pi0086 & n2494;
  assign n2496 = ~pi0097 & ~pi0108;
  assign n2497 = ~pi0094 & n2496;
  assign n2498 = ~pi0046 & n2495;
  assign n2499 = n2497 & n2498;
  assign n2500 = n2493 & n2499;
  assign n2501 = n2492 & n2500;
  assign n2502 = n2491 & n2501;
  assign n2503 = n2461 & n2502;
  assign n2504 = ~pi0035 & ~pi0093;
  assign n2505 = n2503 & n2504;
  assign n2506 = ~pi0072 & ~pi0096;
  assign n2507 = ~pi0051 & ~pi0070;
  assign n2508 = n2506 & n2507;
  assign n2509 = n2505 & n2508;
  assign n2510 = ~pi0032 & ~pi0040;
  assign n2511 = n2509 & n2510;
  assign n2512 = ~pi0095 & n2511;
  assign n2513 = ~n2442 & ~n2512;
  assign n2514 = pi0234 & ~n2513;
  assign n2515 = ~pi0070 & n2505;
  assign n2516 = ~pi0051 & ~pi0096;
  assign n2517 = ~pi0040 & ~pi0072;
  assign n2518 = ~pi0032 & ~pi0095;
  assign n2519 = n2517 & n2518;
  assign n2520 = n2516 & n2519;
  assign n2521 = n2515 & n2520;
  assign n2522 = ~pi0234 & n2521;
  assign n2523 = ~n2514 & ~n2522;
  assign n2524 = pi0137 & ~n2523;
  assign n2525 = n2444 & ~n2524;
  assign n2526 = ~pi0215 & ~pi0221;
  assign n2527 = n2448 & n2526;
  assign n2528 = ~n2525 & n2527;
  assign n2529 = ~pi0056 & ~pi0062;
  assign n2530 = ~pi0038 & ~pi0039;
  assign n2531 = ~pi0100 & n2530;
  assign n2532 = ~pi0054 & ~pi0074;
  assign n2533 = ~pi0075 & ~pi0087;
  assign n2534 = ~pi0092 & n2533;
  assign n2535 = n2532 & n2534;
  assign n2536 = ~pi0055 & n2535;
  assign n2537 = n2531 & n2536;
  assign n2538 = n2529 & n2537;
  assign n2539 = n2528 & n2538;
  assign n2540 = pi0059 & n2460;
  assign n2541 = ~n2539 & n2540;
  assign n2542 = n2460 & ~n2537;
  assign n2543 = ~pi0105 & ~n2446;
  assign n2544 = pi0105 & ~n2525;
  assign n2545 = ~n2543 & ~n2544;
  assign n2546 = pi0228 & ~n2545;
  assign n2547 = pi0137 & n2521;
  assign n2548 = n2446 & ~n2547;
  assign n2549 = ~pi0332 & n2512;
  assign n2550 = ~pi0137 & ~pi0153;
  assign n2551 = n2549 & n2550;
  assign n2552 = ~pi0228 & ~n2548;
  assign n2553 = ~n2551 & n2552;
  assign n2554 = ~n2546 & ~n2553;
  assign n2555 = ~pi0216 & ~n2554;
  assign n2556 = ~n2440 & ~n2555;
  assign n2557 = ~pi0221 & ~n2556;
  assign n2558 = ~n2457 & ~n2557;
  assign n2559 = ~pi0215 & ~n2558;
  assign n2560 = ~n2438 & ~n2559;
  assign n2561 = n2537 & n2560;
  assign n2562 = ~n2542 & ~n2561;
  assign n2563 = ~pi0056 & ~n2562;
  assign n2564 = pi0056 & n2460;
  assign n2565 = pi0062 & ~n2564;
  assign n2566 = ~n2563 & n2565;
  assign n2567 = pi0056 & ~n2562;
  assign n2568 = ~pi0087 & ~pi0100;
  assign n2569 = ~pi0075 & ~pi0092;
  assign n2570 = n2532 & n2569;
  assign n2571 = n2568 & n2570;
  assign n2572 = n2530 & n2571;
  assign n2573 = n2460 & ~n2572;
  assign n2574 = pi0228 & ~n2543;
  assign n2575 = ~pi0332 & n2523;
  assign n2576 = pi0105 & ~n2575;
  assign n2577 = n2574 & ~n2576;
  assign n2578 = ~pi0228 & n2446;
  assign n2579 = ~n2521 & n2578;
  assign n2580 = ~pi0216 & ~n2579;
  assign n2581 = ~n2577 & n2580;
  assign n2582 = ~n2440 & ~n2581;
  assign n2583 = ~pi0221 & ~n2582;
  assign n2584 = ~n2457 & ~n2583;
  assign n2585 = ~pi0215 & ~n2584;
  assign n2586 = ~n2438 & n2572;
  assign n2587 = ~n2585 & n2586;
  assign n2588 = pi0055 & ~n2573;
  assign n2589 = ~n2587 & n2588;
  assign n2590 = pi0299 & n2460;
  assign n2591 = ~pi0224 & pi0833;
  assign n2592 = pi0222 & ~n2591;
  assign n2593 = ~pi0223 & ~n2592;
  assign n2594 = n2437 & ~n2593;
  assign n2595 = pi0224 & ~n2439;
  assign n2596 = ~pi0222 & ~n2595;
  assign n2597 = ~pi0332 & ~pi0929;
  assign n2598 = n2591 & n2597;
  assign n2599 = ~n2596 & ~n2598;
  assign n2600 = ~pi0223 & ~n2599;
  assign n2601 = ~n2594 & ~n2600;
  assign n2602 = ~pi0299 & ~n2601;
  assign n2603 = ~pi0222 & ~pi0224;
  assign n2604 = ~pi0223 & n2603;
  assign n2605 = ~n2444 & n2604;
  assign n2606 = n2602 & ~n2605;
  assign n2607 = ~n2590 & ~n2606;
  assign n2608 = ~pi0038 & ~pi0100;
  assign n2609 = ~pi0039 & ~pi0087;
  assign n2610 = n2608 & n2609;
  assign n2611 = n2569 & n2610;
  assign n2612 = n2607 & ~n2611;
  assign n2613 = ~n2525 & n2604;
  assign n2614 = ~n2601 & ~n2613;
  assign n2615 = ~pi0299 & ~n2614;
  assign n2616 = n2460 & ~n2528;
  assign n2617 = pi0299 & ~n2616;
  assign n2618 = ~n2615 & ~n2617;
  assign n2619 = ~pi0039 & ~n2618;
  assign n2620 = ~pi0038 & n2568;
  assign n2621 = n2569 & n2620;
  assign n2622 = n2619 & n2621;
  assign n2623 = ~n2612 & ~n2622;
  assign n2624 = pi0054 & n2623;
  assign n2625 = ~pi0039 & n2608;
  assign n2626 = ~n2607 & ~n2625;
  assign n2627 = pi0299 & ~n2560;
  assign n2628 = ~n2615 & ~n2627;
  assign n2629 = n2625 & n2628;
  assign n2630 = ~n2626 & ~n2629;
  assign n2631 = n2533 & ~n2630;
  assign n2632 = ~n2533 & ~n2607;
  assign n2633 = pi0092 & ~n2632;
  assign n2634 = ~n2631 & n2633;
  assign n2635 = pi0087 & ~n2630;
  assign n2636 = ~n2530 & ~n2607;
  assign n2637 = pi0095 & pi0234;
  assign n2638 = ~pi0152 & ~pi0161;
  assign n2639 = ~pi0166 & n2638;
  assign n2640 = ~pi0146 & ~n2639;
  assign n2641 = ~pi0210 & ~n2640;
  assign n2642 = ~pi0137 & ~n2637;
  assign n2643 = ~n2641 & n2642;
  assign n2644 = ~n2523 & ~n2643;
  assign n2645 = ~pi0332 & ~n2644;
  assign n2646 = pi0105 & ~n2645;
  assign n2647 = n2574 & ~n2646;
  assign n2648 = n2547 & n2640;
  assign n2649 = ~pi0137 & pi0210;
  assign n2650 = ~pi0252 & ~n2649;
  assign n2651 = ~n2640 & n2650;
  assign n2652 = n2549 & n2651;
  assign n2653 = n2446 & ~n2648;
  assign n2654 = ~n2652 & n2653;
  assign n2655 = pi0252 & ~n2640;
  assign n2656 = ~n2641 & ~n2655;
  assign n2657 = n2551 & n2656;
  assign n2658 = ~n2654 & ~n2657;
  assign n2659 = ~pi0228 & ~n2658;
  assign n2660 = ~pi0216 & ~n2659;
  assign n2661 = ~n2647 & n2660;
  assign n2662 = ~n2440 & ~n2661;
  assign n2663 = ~pi0221 & ~n2662;
  assign n2664 = ~n2457 & ~n2663;
  assign n2665 = ~pi0215 & ~n2664;
  assign n2666 = ~n2438 & ~n2665;
  assign n2667 = pi0299 & ~n2666;
  assign n2668 = ~pi0144 & ~pi0174;
  assign n2669 = ~pi0189 & n2668;
  assign n2670 = ~pi0223 & ~n2669;
  assign n2671 = pi0142 & ~pi0198;
  assign n2672 = ~pi0137 & ~n2671;
  assign n2673 = ~n2523 & ~n2672;
  assign n2674 = n2444 & ~n2673;
  assign n2675 = n2670 & ~n2674;
  assign n2676 = ~pi0234 & ~pi0332;
  assign n2677 = ~pi0137 & pi0198;
  assign n2678 = n2521 & ~n2677;
  assign n2679 = n2676 & ~n2678;
  assign n2680 = ~pi0223 & n2669;
  assign n2681 = pi0234 & ~pi0332;
  assign n2682 = ~pi0095 & n2677;
  assign n2683 = ~n2513 & ~n2682;
  assign n2684 = n2681 & ~n2683;
  assign n2685 = ~n2679 & n2680;
  assign n2686 = ~n2684 & n2685;
  assign n2687 = ~n2675 & ~n2686;
  assign n2688 = n2603 & ~n2687;
  assign n2689 = ~n2601 & ~n2688;
  assign n2690 = ~pi0299 & ~n2689;
  assign n2691 = n2530 & ~n2690;
  assign n2692 = ~n2667 & n2691;
  assign n2693 = pi0100 & ~n2636;
  assign n2694 = ~n2692 & n2693;
  assign n2695 = pi0039 & n2607;
  assign n2696 = pi0038 & ~n2695;
  assign n2697 = ~n2619 & n2696;
  assign n2698 = pi0039 & ~n2628;
  assign n2699 = n2491 & n2499;
  assign n2700 = ~pi0058 & ~pi0091;
  assign n2701 = ~pi0047 & n2700;
  assign n2702 = n2493 & n2701;
  assign n2703 = n2699 & n2702;
  assign n2704 = ~pi0090 & ~pi0093;
  assign n2705 = ~pi0070 & ~pi0096;
  assign n2706 = ~pi0035 & ~pi0051;
  assign n2707 = n2705 & n2706;
  assign n2708 = n2704 & n2707;
  assign n2709 = n2703 & n2708;
  assign n2710 = n2517 & n2709;
  assign n2711 = pi0225 & n2710;
  assign n2712 = pi0032 & ~n2711;
  assign n2713 = ~pi0095 & ~n2712;
  assign n2714 = ~pi0046 & n2493;
  assign n2715 = n2492 & n2496;
  assign n2716 = n2714 & n2715;
  assign n2717 = ~pi0058 & n2716;
  assign n2718 = pi0060 & n2491;
  assign n2719 = ~pi0053 & ~n2718;
  assign n2720 = ~pi0086 & ~pi0094;
  assign n2721 = ~pi0060 & n2491;
  assign n2722 = pi0053 & ~n2721;
  assign n2723 = n2720 & ~n2722;
  assign n2724 = ~n2719 & n2723;
  assign n2725 = n2704 & n2717;
  assign n2726 = n2724 & n2725;
  assign n2727 = ~pi0035 & ~n2726;
  assign n2728 = ~pi0093 & n2503;
  assign n2729 = pi0035 & ~n2728;
  assign n2730 = pi0035 & n2728;
  assign n2731 = ~pi0225 & n2730;
  assign n2732 = ~pi0070 & ~n2731;
  assign n2733 = ~pi0051 & n2732;
  assign n2734 = ~n2729 & n2733;
  assign n2735 = ~n2727 & n2734;
  assign n2736 = ~pi0040 & n2506;
  assign n2737 = n2735 & n2736;
  assign n2738 = ~pi0032 & ~n2737;
  assign n2739 = n2713 & ~n2738;
  assign n2740 = ~pi0137 & ~n2739;
  assign n2741 = pi0095 & ~n2511;
  assign n2742 = ~n2442 & ~n2741;
  assign n2743 = pi0040 & n2509;
  assign n2744 = ~pi0032 & ~n2743;
  assign n2745 = pi0072 & ~n2709;
  assign n2746 = ~pi0040 & ~n2745;
  assign n2747 = pi0051 & ~n2515;
  assign n2748 = ~pi0096 & ~n2747;
  assign n2749 = ~pi0051 & pi0070;
  assign n2750 = n2748 & ~n2749;
  assign n2751 = ~n2729 & ~n2731;
  assign n2752 = pi0093 & n2503;
  assign n2753 = ~pi0035 & ~n2752;
  assign n2754 = ~pi0047 & n2500;
  assign n2755 = n2491 & n2754;
  assign n2756 = pi0091 & n2755;
  assign n2757 = n2461 & ~n2756;
  assign n2758 = ~pi0109 & n2699;
  assign n2759 = pi0110 & ~n2758;
  assign n2760 = pi0047 & n2491;
  assign n2761 = n2500 & n2760;
  assign n2762 = pi0047 & ~n2761;
  assign n2763 = ~pi0091 & ~n2762;
  assign n2764 = ~n2759 & n2763;
  assign n2765 = ~pi0047 & ~pi0110;
  assign n2766 = pi0109 & ~n2699;
  assign n2767 = ~pi0102 & n2490;
  assign n2768 = n2462 & n2767;
  assign n2769 = ~pi0050 & n2494;
  assign n2770 = ~pi0077 & n2769;
  assign n2771 = n2720 & n2770;
  assign n2772 = n2768 & n2771;
  assign n2773 = ~pi0097 & n2772;
  assign n2774 = pi0108 & ~n2773;
  assign n2775 = ~pi0046 & ~n2774;
  assign n2776 = pi0097 & ~n2772;
  assign n2777 = n2463 & n2767;
  assign n2778 = n2769 & n2777;
  assign n2779 = ~pi0086 & pi0094;
  assign n2780 = n2778 & n2779;
  assign n2781 = ~pi0097 & ~n2780;
  assign n2782 = pi0086 & ~n2778;
  assign n2783 = ~pi0094 & ~n2782;
  assign n2784 = pi0077 & n2768;
  assign n2785 = ~pi0050 & ~n2784;
  assign n2786 = pi0081 & ~n2489;
  assign n2787 = pi0102 & ~n2490;
  assign n2788 = ~n2786 & ~n2787;
  assign n2789 = pi0064 & ~n2488;
  assign n2790 = pi0071 & ~n2485;
  assign n2791 = ~pi0065 & ~n2790;
  assign n2792 = ~pi0067 & n2483;
  assign n2793 = pi0069 & ~n2792;
  assign n2794 = pi0083 & ~n2484;
  assign n2795 = ~pi0103 & ~n2794;
  assign n2796 = ~n2793 & n2795;
  assign n2797 = ~pi0069 & ~pi0083;
  assign n2798 = pi0067 & ~n2483;
  assign n2799 = n2469 & n2477;
  assign n2800 = ~pi0084 & n2799;
  assign n2801 = ~pi0068 & n2800;
  assign n2802 = n2479 & n2801;
  assign n2803 = pi0036 & ~n2802;
  assign n2804 = ~pi0036 & ~pi0067;
  assign n2805 = ~pi0068 & ~pi0111;
  assign n2806 = pi0082 & n2805;
  assign n2807 = n2800 & n2806;
  assign n2808 = pi0111 & ~n2801;
  assign n2809 = ~pi0082 & ~n2808;
  assign n2810 = pi0068 & ~n2800;
  assign n2811 = pi0084 & ~n2799;
  assign n2812 = pi0104 & ~n2475;
  assign n2813 = pi0085 & pi0106;
  assign n2814 = n2470 & ~n2813;
  assign n2815 = pi0061 & pi0076;
  assign n2816 = n2471 & ~n2815;
  assign n2817 = ~n2814 & ~n2816;
  assign n2818 = ~pi0048 & ~n2817;
  assign n2819 = ~n2472 & ~n2818;
  assign n2820 = pi0089 & ~n2473;
  assign n2821 = ~pi0049 & ~n2820;
  assign n2822 = ~n2819 & n2821;
  assign n2823 = ~n2474 & ~n2822;
  assign n2824 = ~pi0045 & ~n2812;
  assign n2825 = ~n2823 & n2824;
  assign n2826 = ~n2476 & ~n2825;
  assign n2827 = ~n2477 & ~n2826;
  assign n2828 = n2469 & ~n2827;
  assign n2829 = pi0066 & pi0073;
  assign n2830 = ~n2469 & ~n2477;
  assign n2831 = ~n2829 & ~n2830;
  assign n2832 = ~n2828 & n2831;
  assign n2833 = ~pi0084 & ~n2832;
  assign n2834 = ~n2811 & ~n2833;
  assign n2835 = n2805 & ~n2834;
  assign n2836 = n2809 & ~n2810;
  assign n2837 = ~n2835 & n2836;
  assign n2838 = n2804 & ~n2807;
  assign n2839 = ~n2837 & n2838;
  assign n2840 = ~n2798 & ~n2803;
  assign n2841 = ~n2839 & n2840;
  assign n2842 = n2797 & ~n2841;
  assign n2843 = n2796 & ~n2842;
  assign n2844 = pi0103 & n2797;
  assign n2845 = n2792 & n2844;
  assign n2846 = ~pi0071 & ~n2845;
  assign n2847 = ~n2843 & n2846;
  assign n2848 = n2791 & ~n2847;
  assign n2849 = ~pi0107 & ~n2848;
  assign n2850 = pi0065 & ~pi0071;
  assign n2851 = n2485 & n2850;
  assign n2852 = n2849 & ~n2851;
  assign n2853 = pi0107 & ~n2486;
  assign n2854 = ~pi0063 & ~n2853;
  assign n2855 = ~n2852 & n2854;
  assign n2856 = ~pi0064 & ~n2855;
  assign n2857 = ~n2789 & ~n2856;
  assign n2858 = ~pi0081 & ~pi0102;
  assign n2859 = ~n2857 & n2858;
  assign n2860 = ~n2849 & n2854;
  assign n2861 = pi0063 & ~pi0107;
  assign n2862 = n2486 & n2861;
  assign n2863 = ~pi0064 & ~n2862;
  assign n2864 = ~n2860 & n2863;
  assign n2865 = ~n2789 & ~n2864;
  assign n2866 = n2859 & ~n2865;
  assign n2867 = n2788 & ~n2866;
  assign n2868 = n2462 & ~n2867;
  assign n2869 = pi0098 & ~n2767;
  assign n2870 = ~pi0098 & n2767;
  assign n2871 = pi0088 & ~n2870;
  assign n2872 = ~pi0077 & ~n2869;
  assign n2873 = ~n2871 & n2872;
  assign n2874 = ~n2868 & n2873;
  assign n2875 = n2785 & ~n2874;
  assign n2876 = pi0050 & ~n2777;
  assign n2877 = ~pi0060 & ~n2876;
  assign n2878 = ~n2875 & n2877;
  assign n2879 = n2719 & ~n2878;
  assign n2880 = ~n2722 & ~n2879;
  assign n2881 = ~pi0086 & ~n2880;
  assign n2882 = n2783 & ~n2881;
  assign n2883 = n2781 & ~n2882;
  assign n2884 = ~n2776 & ~n2883;
  assign n2885 = ~pi0108 & ~n2884;
  assign n2886 = n2775 & ~n2885;
  assign n2887 = pi0046 & n2496;
  assign n2888 = n2772 & n2887;
  assign n2889 = ~pi0109 & ~n2888;
  assign n2890 = ~n2886 & n2889;
  assign n2891 = ~n2766 & ~n2890;
  assign n2892 = n2765 & ~n2891;
  assign n2893 = n2764 & ~n2892;
  assign n2894 = n2757 & ~n2893;
  assign n2895 = pi0058 & ~n2502;
  assign n2896 = pi0090 & ~n2703;
  assign n2897 = ~pi0093 & ~n2896;
  assign n2898 = ~n2895 & n2897;
  assign n2899 = ~n2894 & n2898;
  assign n2900 = n2753 & ~n2899;
  assign n2901 = n2751 & ~n2900;
  assign n2902 = ~pi0051 & ~n2901;
  assign n2903 = n2750 & ~n2902;
  assign n2904 = ~pi0072 & ~n2903;
  assign n2905 = n2746 & ~n2904;
  assign n2906 = n2744 & ~n2905;
  assign n2907 = ~n2712 & ~n2906;
  assign n2908 = ~pi0095 & ~n2907;
  assign n2909 = n2742 & ~n2908;
  assign n2910 = pi0137 & ~n2909;
  assign n2911 = ~n2740 & ~n2910;
  assign n2912 = pi0210 & ~n2911;
  assign n2913 = ~pi0051 & ~pi0072;
  assign n2914 = pi0841 & n2503;
  assign n2915 = ~pi0093 & n2914;
  assign n2916 = n2913 & n2915;
  assign n2917 = ~pi0035 & ~pi0040;
  assign n2918 = pi0225 & n2917;
  assign n2919 = n2705 & n2918;
  assign n2920 = n2916 & n2919;
  assign n2921 = pi0032 & ~n2920;
  assign n2922 = ~pi0095 & ~n2921;
  assign n2923 = ~pi0833 & pi0957;
  assign n2924 = pi1091 & ~n2923;
  assign n2925 = pi0829 & pi0950;
  assign n2926 = pi1092 & pi1093;
  assign n2927 = n2925 & n2926;
  assign n2928 = n2924 & n2927;
  assign n2929 = ~n2727 & ~n2928;
  assign n2930 = pi1091 & pi1093;
  assign n2931 = ~n2923 & n2930;
  assign n2932 = pi0950 & pi1092;
  assign n2933 = pi0829 & n2932;
  assign n2934 = ~pi0046 & ~pi0109;
  assign n2935 = n2492 & n2934;
  assign n2936 = ~pi0108 & ~n2776;
  assign n2937 = ~pi0110 & n2936;
  assign n2938 = ~pi0093 & n2461;
  assign n2939 = ~pi0097 & ~n2724;
  assign n2940 = n2935 & n2938;
  assign n2941 = n2937 & n2940;
  assign n2942 = ~n2939 & n2941;
  assign n2943 = ~pi0035 & ~n2942;
  assign n2944 = n2931 & n2933;
  assign n2945 = ~n2943 & n2944;
  assign n2946 = ~n2929 & ~n2945;
  assign n2947 = n2734 & n2736;
  assign n2948 = ~n2946 & n2947;
  assign n2949 = ~pi0032 & ~n2948;
  assign n2950 = n2922 & ~n2949;
  assign n2951 = ~pi0137 & ~n2950;
  assign n2952 = ~n2906 & ~n2921;
  assign n2953 = ~pi0095 & ~n2952;
  assign n2954 = n2742 & ~n2953;
  assign n2955 = pi0137 & ~n2954;
  assign n2956 = ~n2951 & ~n2955;
  assign n2957 = ~pi0210 & ~n2956;
  assign n2958 = ~n2912 & ~n2957;
  assign n2959 = ~pi0234 & n2958;
  assign n2960 = ~pi0096 & ~n2735;
  assign n2961 = ~pi0035 & ~pi0070;
  assign n2962 = ~pi0051 & n2961;
  assign n2963 = ~pi0091 & n2938;
  assign n2964 = n2962 & n2963;
  assign n2965 = n2755 & n2964;
  assign n2966 = pi0096 & ~n2965;
  assign n2967 = n2517 & ~n2966;
  assign n2968 = ~n2960 & n2967;
  assign n2969 = ~pi0032 & ~n2968;
  assign n2970 = n2713 & ~n2969;
  assign n2971 = ~n2442 & ~n2970;
  assign n2972 = ~pi0137 & n2971;
  assign n2973 = pi0096 & n2965;
  assign n2974 = ~pi0040 & n2913;
  assign n2975 = n2505 & n2974;
  assign n2976 = n2973 & n2975;
  assign n2977 = n2906 & ~n2976;
  assign n2978 = ~n2712 & ~n2977;
  assign n2979 = ~pi0095 & ~n2978;
  assign n2980 = pi0479 & n2741;
  assign n2981 = ~n2979 & ~n2980;
  assign n2982 = pi0137 & ~n2981;
  assign n2983 = ~n2972 & ~n2982;
  assign n2984 = pi0210 & ~n2983;
  assign n2985 = ~n2921 & ~n2977;
  assign n2986 = ~pi0095 & ~n2985;
  assign n2987 = ~n2980 & ~n2986;
  assign n2988 = pi0137 & ~n2987;
  assign n2989 = pi0095 & pi0479;
  assign n2990 = ~n2921 & ~n2969;
  assign n2991 = ~pi0095 & ~n2990;
  assign n2992 = ~n2989 & ~n2991;
  assign n2993 = ~pi0137 & ~n2992;
  assign n2994 = ~n2988 & ~n2993;
  assign n2995 = ~n2924 & n2994;
  assign n2996 = n2734 & ~n2943;
  assign n2997 = ~pi0096 & ~n2996;
  assign n2998 = n2967 & ~n2997;
  assign n2999 = ~pi0032 & ~n2998;
  assign n3000 = ~n2921 & ~n2999;
  assign n3001 = ~pi0095 & ~n3000;
  assign n3002 = n2927 & ~n2989;
  assign n3003 = ~n3001 & n3002;
  assign n3004 = ~n2927 & n2992;
  assign n3005 = ~pi0137 & ~n3003;
  assign n3006 = ~n3004 & n3005;
  assign n3007 = n2924 & ~n3006;
  assign n3008 = ~n2988 & n3007;
  assign n3009 = ~n2995 & ~n3008;
  assign n3010 = ~pi0210 & n3009;
  assign n3011 = ~n2984 & ~n3010;
  assign n3012 = pi0234 & n3011;
  assign n3013 = ~pi0332 & ~n2959;
  assign n3014 = ~n3012 & n3013;
  assign n3015 = n2639 & ~n3014;
  assign n3016 = pi0146 & n3011;
  assign n3017 = ~pi0210 & ~n2994;
  assign n3018 = ~pi0146 & ~n2984;
  assign n3019 = ~n3017 & n3018;
  assign n3020 = n2681 & ~n3019;
  assign n3021 = ~n3016 & n3020;
  assign n3022 = pi0146 & n2958;
  assign n3023 = ~n2738 & n2922;
  assign n3024 = ~pi0137 & ~n3023;
  assign n3025 = ~n2955 & ~n3024;
  assign n3026 = ~pi0210 & ~n3025;
  assign n3027 = ~pi0146 & ~n2912;
  assign n3028 = ~n3026 & n3027;
  assign n3029 = n2676 & ~n3022;
  assign n3030 = ~n3028 & n3029;
  assign n3031 = ~n2639 & ~n3030;
  assign n3032 = ~n3021 & n3031;
  assign n3033 = ~n3015 & ~n3032;
  assign n3034 = pi0105 & ~n3033;
  assign n3035 = ~n2543 & ~n3034;
  assign n3036 = pi0228 & ~n3035;
  assign n3037 = ~pi0109 & ~n2886;
  assign n3038 = ~n2766 & ~n3037;
  assign n3039 = n2765 & ~n3038;
  assign n3040 = n2764 & ~n3039;
  assign n3041 = n2757 & ~n3040;
  assign n3042 = n2898 & ~n3041;
  assign n3043 = n2753 & ~n3042;
  assign n3044 = n2751 & ~n3043;
  assign n3045 = ~pi0051 & ~n3044;
  assign n3046 = n2750 & ~n3045;
  assign n3047 = ~pi0072 & ~n3046;
  assign n3048 = n2746 & ~n3047;
  assign n3049 = n2744 & ~n3048;
  assign n3050 = ~n2921 & ~n3049;
  assign n3051 = ~pi0095 & ~n3050;
  assign n3052 = n2742 & ~n3051;
  assign n3053 = pi0137 & ~n3052;
  assign n3054 = n2640 & n3024;
  assign n3055 = ~n2640 & n2951;
  assign n3056 = ~pi0210 & ~pi0234;
  assign n3057 = ~n3054 & n3056;
  assign n3058 = ~n3055 & n3057;
  assign n3059 = ~n3053 & n3058;
  assign n3060 = ~n2712 & ~n3049;
  assign n3061 = ~pi0095 & ~n3060;
  assign n3062 = n2742 & ~n3061;
  assign n3063 = pi0137 & ~n3062;
  assign n3064 = pi0210 & ~n2740;
  assign n3065 = ~n3063 & n3064;
  assign n3066 = ~n2976 & n3049;
  assign n3067 = ~n2921 & ~n3066;
  assign n3068 = ~pi0095 & ~n3067;
  assign n3069 = ~n2741 & ~n3068;
  assign n3070 = pi0137 & ~n3069;
  assign n3071 = ~n2640 & n2924;
  assign n3072 = ~n3004 & n3071;
  assign n3073 = ~n2741 & n2992;
  assign n3074 = ~n3072 & n3073;
  assign n3075 = ~n2741 & n3071;
  assign n3076 = n3003 & n3075;
  assign n3077 = ~pi0137 & ~n3076;
  assign n3078 = ~n3074 & n3077;
  assign n3079 = ~n3070 & ~n3078;
  assign n3080 = ~pi0210 & ~n3079;
  assign n3081 = pi0234 & ~n3080;
  assign n3082 = ~n3059 & ~n3065;
  assign n3083 = ~n3081 & n3082;
  assign n3084 = ~pi0137 & ~n2741;
  assign n3085 = ~n2971 & n3084;
  assign n3086 = ~n2712 & ~n3066;
  assign n3087 = ~pi0095 & ~n3086;
  assign n3088 = pi0137 & ~n2741;
  assign n3089 = ~n3087 & n3088;
  assign n3090 = pi0210 & pi0234;
  assign n3091 = ~n3085 & n3090;
  assign n3092 = ~n3089 & n3091;
  assign n3093 = ~n3083 & ~n3092;
  assign n3094 = n2446 & ~n3093;
  assign n3095 = pi0225 & pi0841;
  assign n3096 = n2710 & ~n3095;
  assign n3097 = pi0032 & ~n3096;
  assign n3098 = ~pi0095 & ~n3097;
  assign n3099 = pi0070 & ~n2505;
  assign n3100 = n2516 & ~n3099;
  assign n3101 = n2517 & n3100;
  assign n3102 = ~n2732 & n3101;
  assign n3103 = ~pi0032 & ~n3102;
  assign n3104 = n3098 & ~n3103;
  assign n3105 = pi0137 & ~n3104;
  assign n3106 = pi0093 & ~n2503;
  assign n3107 = ~pi0035 & ~n3106;
  assign n3108 = ~n2895 & ~n2896;
  assign n3109 = ~pi0053 & n2878;
  assign n3110 = ~pi0086 & ~n3109;
  assign n3111 = n2783 & ~n3110;
  assign n3112 = n2781 & ~n3111;
  assign n3113 = ~n2776 & ~n3112;
  assign n3114 = ~pi0108 & ~n3113;
  assign n3115 = n2775 & ~n3114;
  assign n3116 = ~pi0109 & ~n3115;
  assign n3117 = ~n2766 & ~n3116;
  assign n3118 = n2765 & ~n3117;
  assign n3119 = n2764 & ~n3118;
  assign n3120 = n2757 & ~n3119;
  assign n3121 = n3108 & ~n3120;
  assign n3122 = ~pi0093 & ~n3121;
  assign n3123 = n3107 & ~n3122;
  assign n3124 = n2733 & ~n3123;
  assign n3125 = n2748 & ~n3099;
  assign n3126 = ~n3124 & n3125;
  assign n3127 = ~pi0072 & ~n3126;
  assign n3128 = n2746 & ~n3127;
  assign n3129 = n2744 & ~n3128;
  assign n3130 = ~n2928 & n3129;
  assign n3131 = n2744 & n2928;
  assign n3132 = ~pi0097 & ~n3112;
  assign n3133 = ~pi0108 & ~n3132;
  assign n3134 = n2775 & ~n3133;
  assign n3135 = ~pi0109 & ~n3134;
  assign n3136 = ~n2766 & ~n3135;
  assign n3137 = n2765 & ~n3136;
  assign n3138 = n2764 & ~n3137;
  assign n3139 = n2757 & ~n3138;
  assign n3140 = n3108 & ~n3139;
  assign n3141 = ~pi0093 & ~n3140;
  assign n3142 = n3107 & ~n3141;
  assign n3143 = n2733 & ~n3142;
  assign n3144 = n3125 & ~n3143;
  assign n3145 = ~pi0072 & ~n3144;
  assign n3146 = n2746 & ~n3145;
  assign n3147 = n3131 & ~n3146;
  assign n3148 = ~n3097 & ~n3147;
  assign n3149 = ~n3130 & n3148;
  assign n3150 = ~pi0095 & ~n3149;
  assign n3151 = n2742 & ~n3150;
  assign n3152 = ~pi0137 & ~n3151;
  assign n3153 = ~n3105 & ~n3152;
  assign n3154 = ~pi0210 & ~n3153;
  assign n3155 = ~pi0225 & n2710;
  assign n3156 = pi0032 & ~n3155;
  assign n3157 = ~pi0095 & ~n3156;
  assign n3158 = pi0137 & n3157;
  assign n3159 = ~n3103 & n3158;
  assign n3160 = ~n3129 & ~n3156;
  assign n3161 = ~pi0095 & ~n3160;
  assign n3162 = ~pi0137 & n2742;
  assign n3163 = ~n3161 & n3162;
  assign n3164 = pi0210 & ~n3159;
  assign n3165 = ~n3163 & n3164;
  assign n3166 = n2681 & ~n3165;
  assign n3167 = ~n3154 & n3166;
  assign n3168 = ~pi0072 & ~n2973;
  assign n3169 = ~n3126 & n3168;
  assign n3170 = n2746 & ~n3169;
  assign n3171 = n2744 & ~n3170;
  assign n3172 = ~n2928 & n3171;
  assign n3173 = ~n3144 & n3168;
  assign n3174 = n2746 & ~n3173;
  assign n3175 = n3131 & ~n3174;
  assign n3176 = ~n3097 & ~n3175;
  assign n3177 = ~n3172 & n3176;
  assign n3178 = ~pi0095 & ~n3177;
  assign n3179 = ~n2741 & ~n3178;
  assign n3180 = ~pi0137 & ~n3179;
  assign n3181 = n2442 & n2511;
  assign n3182 = ~pi0072 & n2510;
  assign n3183 = n2973 & n3182;
  assign n3184 = n3103 & ~n3183;
  assign n3185 = n3098 & ~n3184;
  assign n3186 = pi0137 & ~n3181;
  assign n3187 = ~n3185 & n3186;
  assign n3188 = ~n3180 & ~n3187;
  assign n3189 = ~pi0210 & ~n3188;
  assign n3190 = ~n3156 & ~n3171;
  assign n3191 = ~pi0095 & ~n3190;
  assign n3192 = n3084 & ~n3191;
  assign n3193 = n3157 & ~n3184;
  assign n3194 = ~n3181 & ~n3193;
  assign n3195 = pi0137 & ~n3194;
  assign n3196 = pi0210 & ~n3195;
  assign n3197 = ~n3192 & n3196;
  assign n3198 = n2676 & ~n3197;
  assign n3199 = ~n3189 & n3198;
  assign n3200 = n2639 & ~n3167;
  assign n3201 = ~n3199 & n3200;
  assign n3202 = pi0146 & n3189;
  assign n3203 = ~pi0146 & ~pi0210;
  assign n3204 = ~n3097 & ~n3171;
  assign n3205 = ~pi0095 & ~n3204;
  assign n3206 = ~n2741 & ~n3205;
  assign n3207 = ~pi0137 & ~n3206;
  assign n3208 = ~n3187 & ~n3207;
  assign n3209 = n3203 & ~n3208;
  assign n3210 = n3198 & ~n3209;
  assign n3211 = ~n3202 & n3210;
  assign n3212 = ~n3097 & ~n3129;
  assign n3213 = ~pi0095 & ~n3212;
  assign n3214 = n2742 & ~n3213;
  assign n3215 = ~pi0137 & ~n3214;
  assign n3216 = ~n3105 & ~n3215;
  assign n3217 = n3203 & ~n3216;
  assign n3218 = pi0146 & n3154;
  assign n3219 = n3166 & ~n3217;
  assign n3220 = ~n3218 & n3219;
  assign n3221 = ~n2639 & ~n3211;
  assign n3222 = ~n3220 & n3221;
  assign n3223 = ~pi0153 & ~n3201;
  assign n3224 = ~n3222 & n3223;
  assign n3225 = ~pi0228 & ~n3094;
  assign n3226 = ~n3224 & n3225;
  assign n3227 = ~n3036 & ~n3226;
  assign n3228 = ~pi0216 & ~n3227;
  assign n3229 = ~n2440 & ~n3228;
  assign n3230 = ~pi0221 & ~n3229;
  assign n3231 = ~n2457 & ~n3230;
  assign n3232 = ~pi0215 & ~n3231;
  assign n3233 = pi0299 & ~n2438;
  assign n3234 = ~n3232 & n3233;
  assign n3235 = pi0198 & ~n2983;
  assign n3236 = ~pi0198 & n3009;
  assign n3237 = ~n3235 & ~n3236;
  assign n3238 = pi0142 & n3237;
  assign n3239 = ~pi0198 & ~n2994;
  assign n3240 = ~pi0142 & ~n3235;
  assign n3241 = ~n3239 & n3240;
  assign n3242 = n2681 & ~n3241;
  assign n3243 = ~n3238 & n3242;
  assign n3244 = pi0198 & ~n2911;
  assign n3245 = ~pi0198 & ~n2956;
  assign n3246 = ~n3244 & ~n3245;
  assign n3247 = pi0142 & n3246;
  assign n3248 = ~pi0198 & ~n3025;
  assign n3249 = ~pi0142 & ~n3244;
  assign n3250 = ~n3248 & n3249;
  assign n3251 = n2676 & ~n3247;
  assign n3252 = ~n3250 & n3251;
  assign n3253 = n2670 & ~n3252;
  assign n3254 = ~n3243 & n3253;
  assign n3255 = ~pi0234 & n3246;
  assign n3256 = pi0234 & n3237;
  assign n3257 = ~pi0332 & ~n3255;
  assign n3258 = ~n3256 & n3257;
  assign n3259 = n2680 & ~n3258;
  assign n3260 = ~n3254 & ~n3259;
  assign n3261 = n2603 & ~n3260;
  assign n3262 = n2602 & ~n3261;
  assign n3263 = ~pi0039 & ~n3262;
  assign n3264 = ~n3234 & n3263;
  assign n3265 = ~pi0038 & ~n2698;
  assign n3266 = ~n3264 & n3265;
  assign n3267 = ~pi0100 & ~n2697;
  assign n3268 = ~n3266 & n3267;
  assign n3269 = ~pi0087 & ~n2694;
  assign n3270 = ~n3268 & n3269;
  assign n3271 = ~pi0075 & ~n2635;
  assign n3272 = ~n3270 & n3271;
  assign n3273 = ~n2607 & ~n2610;
  assign n3274 = n2448 & ~n2647;
  assign n3275 = ~n2440 & ~n3274;
  assign n3276 = ~pi0221 & ~n3275;
  assign n3277 = ~n2457 & ~n3276;
  assign n3278 = ~pi0215 & ~n3277;
  assign n3279 = ~n2438 & ~n3278;
  assign n3280 = pi0299 & ~n3279;
  assign n3281 = n2610 & ~n2690;
  assign n3282 = ~n3280 & n3281;
  assign n3283 = pi0075 & ~n3273;
  assign n3284 = ~n3282 & n3283;
  assign n3285 = ~n3272 & ~n3284;
  assign n3286 = ~pi0092 & ~n3285;
  assign n3287 = ~pi0054 & ~n2634;
  assign n3288 = ~n3286 & n3287;
  assign n3289 = ~pi0074 & ~n2624;
  assign n3290 = ~n3288 & n3289;
  assign n3291 = pi0054 & ~n2607;
  assign n3292 = ~pi0054 & n2623;
  assign n3293 = pi0074 & ~n3291;
  assign n3294 = ~n3292 & n3293;
  assign n3295 = ~n3290 & ~n3294;
  assign n3296 = ~pi0055 & ~n3295;
  assign n3297 = ~pi0056 & ~n2589;
  assign n3298 = ~n3296 & n3297;
  assign n3299 = ~pi0062 & ~n2567;
  assign n3300 = ~n3298 & n3299;
  assign n3301 = ~pi0059 & ~n2566;
  assign n3302 = ~n3300 & n3301;
  assign n3303 = ~pi0057 & ~n2541;
  assign n3304 = ~n3302 & n3303;
  assign n3305 = ~pi0059 & n2539;
  assign n3306 = n2460 & ~n3305;
  assign n3307 = pi0057 & ~n3306;
  assign po0153 = n3304 | n3307;
  assign n3309 = pi0215 & pi1146;
  assign n3310 = pi0216 & ~pi0221;
  assign n3311 = pi0276 & n3310;
  assign n3312 = ~pi1146 & ~n2452;
  assign n3313 = ~pi0939 & n2452;
  assign n3314 = pi0221 & ~n3312;
  assign n3315 = ~n3313 & n3314;
  assign n3316 = ~n3311 & ~n3315;
  assign n3317 = ~pi0215 & ~n3316;
  assign n3318 = ~n3309 & ~n3317;
  assign n3319 = pi0154 & ~n3318;
  assign n3320 = ~pi0216 & ~n2441;
  assign n3321 = ~n3311 & ~n3320;
  assign n3322 = ~pi0221 & ~n3321;
  assign n3323 = ~n3315 & ~n3322;
  assign n3324 = ~pi0215 & ~n3323;
  assign n3325 = ~n3309 & ~n3324;
  assign n3326 = ~pi0154 & ~n3325;
  assign n3327 = ~n3319 & ~n3326;
  assign n3328 = ~pi0057 & ~pi0059;
  assign n3329 = n3327 & ~n3328;
  assign n3330 = ~pi0056 & n2536;
  assign n3331 = n2531 & n3330;
  assign n3332 = ~n3327 & ~n3331;
  assign n3333 = ~pi0055 & n2572;
  assign n3334 = ~n3309 & ~n3315;
  assign n3335 = ~pi0228 & n2521;
  assign n3336 = ~pi0216 & n3335;
  assign n3337 = n3334 & n3336;
  assign n3338 = ~n3319 & n3337;
  assign n3339 = ~n3327 & n3333;
  assign n3340 = ~n3338 & n3339;
  assign n3341 = ~n3332 & ~n3340;
  assign n3342 = pi0062 & ~n3341;
  assign n3343 = ~n2537 & ~n3327;
  assign n3344 = pi0056 & ~n3343;
  assign n3345 = ~n3340 & n3344;
  assign n3346 = n2572 & n3338;
  assign n3347 = pi0055 & ~n3327;
  assign n3348 = ~n3346 & n3347;
  assign n3349 = pi0299 & ~n3327;
  assign n3350 = pi0223 & ~pi1146;
  assign n3351 = ~pi0222 & pi0224;
  assign n3352 = pi0276 & n3351;
  assign n3353 = ~pi1146 & ~n2591;
  assign n3354 = ~pi0939 & n2591;
  assign n3355 = pi0222 & ~n3353;
  assign n3356 = ~n3354 & n3355;
  assign n3357 = ~pi0223 & ~n3352;
  assign n3358 = ~n3356 & n3357;
  assign n3359 = ~pi0299 & ~n3350;
  assign n3360 = ~n3358 & n3359;
  assign n3361 = ~n3349 & ~n3360;
  assign n3362 = ~n2532 & n3361;
  assign n3363 = pi0299 & ~n3318;
  assign n3364 = ~n3360 & ~n3363;
  assign n3365 = pi0154 & ~n3364;
  assign n3366 = pi0299 & ~n3325;
  assign n3367 = ~n3337 & n3366;
  assign n3368 = ~n3360 & ~n3367;
  assign n3369 = ~pi0154 & ~n3368;
  assign n3370 = n2625 & ~n3365;
  assign n3371 = ~n3369 & n3370;
  assign n3372 = n2533 & n3371;
  assign n3373 = n2531 & n2533;
  assign n3374 = n3361 & ~n3373;
  assign n3375 = pi0092 & ~n3374;
  assign n3376 = ~n3372 & n3375;
  assign n3377 = pi0075 & n3361;
  assign n3378 = ~n2625 & n3361;
  assign n3379 = ~n3371 & ~n3378;
  assign n3380 = pi0087 & ~n3379;
  assign n3381 = ~pi0038 & ~pi0216;
  assign n3382 = ~pi0228 & n3381;
  assign n3383 = ~pi0154 & pi0299;
  assign n3384 = ~pi0146 & ~n2521;
  assign n3385 = ~pi0252 & n2521;
  assign n3386 = pi0146 & ~n3385;
  assign n3387 = ~n3384 & ~n3386;
  assign n3388 = pi0152 & ~n3387;
  assign n3389 = ~pi0161 & ~pi0166;
  assign n3390 = n3385 & n3389;
  assign n3391 = n3387 & ~n3389;
  assign n3392 = ~pi0152 & ~n3390;
  assign n3393 = ~n3391 & n3392;
  assign n3394 = ~n3388 & ~n3393;
  assign n3395 = ~pi0039 & n3383;
  assign n3396 = n3382 & n3395;
  assign n3397 = n3334 & n3396;
  assign n3398 = n3394 & n3397;
  assign n3399 = pi0100 & ~n3361;
  assign n3400 = ~n3398 & n3399;
  assign n3401 = pi0038 & n3361;
  assign n3402 = pi0039 & ~n2521;
  assign n3403 = ~pi0070 & n3043;
  assign n3404 = ~n2729 & ~n3099;
  assign n3405 = ~n3403 & n3404;
  assign n3406 = ~pi0051 & ~n3405;
  assign n3407 = n2748 & ~n3406;
  assign n3408 = n3168 & ~n3407;
  assign n3409 = ~n2745 & ~n3408;
  assign n3410 = n2510 & ~n3409;
  assign n3411 = pi0040 & ~n2509;
  assign n3412 = pi0032 & ~n2710;
  assign n3413 = ~n3411 & ~n3412;
  assign n3414 = ~n3410 & n3413;
  assign n3415 = ~pi0095 & ~n3414;
  assign n3416 = ~n2741 & ~n3415;
  assign n3417 = ~pi0039 & ~n3416;
  assign n3418 = ~n3402 & ~n3417;
  assign n3419 = ~pi0216 & ~pi0228;
  assign n3420 = n3334 & n3419;
  assign n3421 = n3418 & n3420;
  assign n3422 = n3366 & ~n3421;
  assign n3423 = ~n3360 & ~n3422;
  assign n3424 = ~pi0154 & ~n3423;
  assign n3425 = ~pi0038 & ~n3365;
  assign n3426 = ~n3424 & n3425;
  assign n3427 = ~pi0100 & ~n3401;
  assign n3428 = ~n3426 & n3427;
  assign n3429 = ~pi0087 & ~n3400;
  assign n3430 = ~n3428 & n3429;
  assign n3431 = ~n3380 & ~n3430;
  assign n3432 = ~pi0075 & ~n3431;
  assign n3433 = ~pi0092 & ~n3377;
  assign n3434 = ~n3432 & n3433;
  assign n3435 = n2532 & ~n3376;
  assign n3436 = ~n3434 & n3435;
  assign n3437 = ~pi0055 & ~n3362;
  assign n3438 = ~n3436 & n3437;
  assign n3439 = ~pi0056 & ~n3348;
  assign n3440 = ~n3438 & n3439;
  assign n3441 = ~pi0062 & ~n3345;
  assign n3442 = ~n3440 & n3441;
  assign n3443 = n3328 & ~n3342;
  assign n3444 = ~n3442 & n3443;
  assign n3445 = ~pi0239 & ~n3329;
  assign n3446 = ~n3444 & n3445;
  assign n3447 = n2441 & n2442;
  assign n3448 = ~pi0216 & ~pi0221;
  assign n3449 = ~pi0215 & n3448;
  assign n3450 = n3447 & n3449;
  assign n3451 = n3318 & ~n3450;
  assign n3452 = ~pi0215 & ~n3451;
  assign n3453 = pi0154 & ~n3451;
  assign n3454 = ~n3326 & ~n3452;
  assign n3455 = ~n3453 & n3454;
  assign n3456 = ~n3328 & n3455;
  assign n3457 = ~n3331 & ~n3455;
  assign n3458 = n3337 & ~n3453;
  assign n3459 = ~n3455 & ~n3458;
  assign n3460 = n3333 & n3459;
  assign n3461 = ~pi0056 & n3460;
  assign n3462 = ~n3457 & ~n3461;
  assign n3463 = pi0062 & ~n3462;
  assign n3464 = ~n2537 & ~n3455;
  assign n3465 = pi0056 & ~n3464;
  assign n3466 = ~n3460 & n3465;
  assign n3467 = n2572 & n3458;
  assign n3468 = pi0055 & ~n3455;
  assign n3469 = ~n3467 & n3468;
  assign n3470 = ~pi0223 & ~pi0299;
  assign n3471 = n2603 & n3470;
  assign n3472 = n2442 & n3471;
  assign n3473 = pi0299 & ~n3455;
  assign n3474 = ~n3360 & ~n3472;
  assign n3475 = ~n3473 & n3474;
  assign n3476 = ~n2532 & n3475;
  assign n3477 = pi0299 & ~n3459;
  assign n3478 = n3373 & n3477;
  assign n3479 = pi0092 & ~n3475;
  assign n3480 = ~n3478 & n3479;
  assign n3481 = pi0075 & n3475;
  assign n3482 = n2625 & n3477;
  assign n3483 = pi0087 & ~n3475;
  assign n3484 = ~n3482 & n3483;
  assign n3485 = ~n3475 & ~n3477;
  assign n3486 = pi0039 & ~n3485;
  assign n3487 = n2519 & n2973;
  assign n3488 = ~n2442 & ~n3487;
  assign n3489 = ~pi0224 & n3488;
  assign n3490 = pi0224 & ~pi0276;
  assign n3491 = ~pi0222 & ~n3490;
  assign n3492 = ~n3489 & n3491;
  assign n3493 = ~pi0223 & ~n3356;
  assign n3494 = ~n3492 & n3493;
  assign n3495 = ~n3350 & ~n3494;
  assign n3496 = ~pi0299 & ~n3495;
  assign n3497 = pi0105 & ~n3488;
  assign n3498 = pi0228 & ~n3497;
  assign n3499 = ~n2741 & ~n3488;
  assign n3500 = ~pi0228 & ~n3499;
  assign n3501 = ~n3498 & ~n3500;
  assign n3502 = pi0154 & ~n3501;
  assign n3503 = ~pi0072 & ~n3407;
  assign n3504 = ~n2745 & ~n3503;
  assign n3505 = n2510 & ~n3504;
  assign n3506 = n3413 & ~n3505;
  assign n3507 = ~pi0095 & ~n3506;
  assign n3508 = n2742 & ~n3507;
  assign n3509 = ~pi0228 & n3508;
  assign n3510 = n2441 & n3488;
  assign n3511 = ~n3509 & ~n3510;
  assign n3512 = ~pi0154 & ~n3511;
  assign n3513 = n3449 & ~n3502;
  assign n3514 = ~n3512 & n3513;
  assign n3515 = pi0299 & n3318;
  assign n3516 = ~n3514 & n3515;
  assign n3517 = ~n3496 & ~n3516;
  assign n3518 = ~pi0039 & ~n3517;
  assign n3519 = n2608 & ~n3486;
  assign n3520 = ~n3518 & n3519;
  assign n3521 = pi0100 & n3398;
  assign n3522 = ~n2608 & ~n3475;
  assign n3523 = ~n3521 & n3522;
  assign n3524 = ~n3520 & ~n3523;
  assign n3525 = ~pi0087 & ~n3524;
  assign n3526 = ~pi0075 & ~n3484;
  assign n3527 = ~n3525 & n3526;
  assign n3528 = ~pi0092 & ~n3481;
  assign n3529 = ~n3527 & n3528;
  assign n3530 = n2532 & ~n3480;
  assign n3531 = ~n3529 & n3530;
  assign n3532 = ~pi0055 & ~n3476;
  assign n3533 = ~n3531 & n3532;
  assign n3534 = ~pi0056 & ~n3469;
  assign n3535 = ~n3533 & n3534;
  assign n3536 = ~pi0062 & ~n3466;
  assign n3537 = ~n3535 & n3536;
  assign n3538 = n3328 & ~n3463;
  assign n3539 = ~n3537 & n3538;
  assign n3540 = pi0239 & ~n3456;
  assign n3541 = ~n3539 & n3540;
  assign po0154 = n3446 | n3541;
  assign n3543 = pi0215 & pi1145;
  assign n3544 = pi0216 & pi0274;
  assign n3545 = ~pi0221 & ~n3544;
  assign n3546 = ~pi0151 & ~n2441;
  assign n3547 = ~pi0216 & ~n3546;
  assign n3548 = n3545 & ~n3547;
  assign n3549 = ~pi1145 & ~n2452;
  assign n3550 = ~pi0927 & n2452;
  assign n3551 = pi0221 & ~n3549;
  assign n3552 = ~n3550 & n3551;
  assign n3553 = ~n3548 & ~n3552;
  assign n3554 = ~pi0215 & ~n3553;
  assign n3555 = ~n3543 & ~n3554;
  assign n3556 = n2526 & n3447;
  assign n3557 = ~n3544 & n3556;
  assign n3558 = n3555 & ~n3557;
  assign n3559 = ~n3331 & n3558;
  assign n3560 = ~n3447 & ~n3546;
  assign n3561 = ~pi0151 & n3335;
  assign n3562 = ~n3560 & ~n3561;
  assign n3563 = ~pi0216 & ~n3562;
  assign n3564 = n3545 & ~n3563;
  assign n3565 = ~n3552 & ~n3564;
  assign n3566 = ~pi0215 & ~n3565;
  assign n3567 = ~n3543 & ~n3566;
  assign n3568 = n3331 & n3567;
  assign n3569 = pi0062 & ~n3559;
  assign n3570 = ~n3568 & n3569;
  assign n3571 = ~n2537 & ~n3558;
  assign n3572 = n2537 & ~n3567;
  assign n3573 = pi0056 & ~n3571;
  assign n3574 = ~n3572 & n3573;
  assign n3575 = ~n2572 & n3558;
  assign n3576 = n2572 & n3567;
  assign n3577 = pi0055 & ~n3575;
  assign n3578 = ~n3576 & n3577;
  assign n3579 = pi0223 & pi1145;
  assign n3580 = ~pi1145 & ~n2591;
  assign n3581 = ~pi0927 & n2591;
  assign n3582 = pi0222 & ~n3580;
  assign n3583 = ~n3581 & n3582;
  assign n3584 = pi0224 & pi0274;
  assign n3585 = n3351 & ~n3584;
  assign n3586 = ~n3583 & ~n3585;
  assign n3587 = ~pi0223 & ~n3586;
  assign n3588 = ~n3579 & ~n3587;
  assign n3589 = ~pi0299 & ~n3588;
  assign n3590 = ~n3472 & ~n3589;
  assign n3591 = pi0299 & ~n3558;
  assign n3592 = n3590 & ~n3591;
  assign n3593 = ~n2532 & n3592;
  assign n3594 = ~n2625 & n3592;
  assign n3595 = pi0299 & ~n3567;
  assign n3596 = n3590 & ~n3595;
  assign n3597 = n2625 & n3596;
  assign n3598 = ~n3594 & ~n3597;
  assign n3599 = n2533 & ~n3598;
  assign n3600 = ~n2533 & n3592;
  assign n3601 = pi0092 & ~n3600;
  assign n3602 = ~n3599 & n3601;
  assign n3603 = pi0075 & n3592;
  assign n3604 = pi0087 & n3598;
  assign n3605 = pi0038 & n3592;
  assign n3606 = pi0039 & ~n3596;
  assign n3607 = ~pi0222 & ~n3584;
  assign n3608 = ~n3489 & n3607;
  assign n3609 = ~n3583 & ~n3608;
  assign n3610 = ~pi0223 & ~n3609;
  assign n3611 = ~pi0299 & ~n3579;
  assign n3612 = ~n3610 & n3611;
  assign n3613 = ~pi0151 & n3511;
  assign n3614 = pi0151 & n3501;
  assign n3615 = ~pi0216 & ~n3614;
  assign n3616 = ~n3613 & n3615;
  assign n3617 = n3545 & ~n3616;
  assign n3618 = ~n3552 & ~n3617;
  assign n3619 = ~pi0215 & ~n3618;
  assign n3620 = pi0299 & ~n3543;
  assign n3621 = ~n3619 & n3620;
  assign n3622 = ~pi0039 & ~n3612;
  assign n3623 = ~n3621 & n3622;
  assign n3624 = ~pi0038 & ~n3606;
  assign n3625 = ~n3623 & n3624;
  assign n3626 = ~pi0100 & ~n3605;
  assign n3627 = ~n3625 & n3626;
  assign n3628 = ~n2530 & n3592;
  assign n3629 = ~pi0228 & n3394;
  assign n3630 = n2441 & ~n2442;
  assign n3631 = ~n3629 & ~n3630;
  assign n3632 = ~pi0151 & n3631;
  assign n3633 = n3563 & ~n3632;
  assign n3634 = n3545 & ~n3633;
  assign n3635 = ~n3552 & ~n3634;
  assign n3636 = ~pi0215 & ~n3635;
  assign n3637 = ~n3543 & ~n3636;
  assign n3638 = pi0299 & ~n3637;
  assign n3639 = n2530 & n3590;
  assign n3640 = ~n3638 & n3639;
  assign n3641 = pi0100 & ~n3628;
  assign n3642 = ~n3640 & n3641;
  assign n3643 = ~n3627 & ~n3642;
  assign n3644 = ~pi0087 & ~n3643;
  assign n3645 = ~pi0075 & ~n3604;
  assign n3646 = ~n3644 & n3645;
  assign n3647 = ~pi0092 & ~n3603;
  assign n3648 = ~n3646 & n3647;
  assign n3649 = n2532 & ~n3602;
  assign n3650 = ~n3648 & n3649;
  assign n3651 = ~pi0055 & ~n3593;
  assign n3652 = ~n3650 & n3651;
  assign n3653 = ~pi0056 & ~n3578;
  assign n3654 = ~n3652 & n3653;
  assign n3655 = ~pi0062 & ~n3574;
  assign n3656 = ~n3654 & n3655;
  assign n3657 = pi0235 & n3328;
  assign n3658 = ~n3570 & n3657;
  assign n3659 = ~n3656 & n3658;
  assign n3660 = ~n3543 & ~n3552;
  assign n3661 = n3336 & n3660;
  assign n3662 = n2537 & n3661;
  assign n3663 = ~pi0056 & n3662;
  assign n3664 = pi0062 & ~n3555;
  assign n3665 = ~n3663 & n3664;
  assign n3666 = ~n3555 & ~n3662;
  assign n3667 = pi0056 & ~n3666;
  assign n3668 = n2572 & n3661;
  assign n3669 = pi0055 & ~n3555;
  assign n3670 = ~n3668 & n3669;
  assign n3671 = pi0299 & ~n3555;
  assign n3672 = ~n3589 & ~n3671;
  assign n3673 = ~n2532 & n3672;
  assign n3674 = ~n3661 & n3671;
  assign n3675 = n2531 & ~n3589;
  assign n3676 = ~n3674 & n3675;
  assign n3677 = n2533 & n3676;
  assign n3678 = ~n3373 & n3672;
  assign n3679 = pi0092 & ~n3678;
  assign n3680 = ~n3677 & n3679;
  assign n3681 = pi0075 & n3672;
  assign n3682 = ~n2625 & n3672;
  assign n3683 = ~n3676 & ~n3682;
  assign n3684 = pi0087 & ~n3683;
  assign n3685 = ~pi0100 & n3418;
  assign n3686 = ~pi0039 & pi0100;
  assign n3687 = n3394 & n3686;
  assign n3688 = ~n3685 & ~n3687;
  assign n3689 = n3382 & n3660;
  assign n3690 = ~n3688 & n3689;
  assign n3691 = n3671 & ~n3690;
  assign n3692 = ~pi0087 & ~n3589;
  assign n3693 = ~n3691 & n3692;
  assign n3694 = ~n3684 & ~n3693;
  assign n3695 = ~pi0075 & ~n3694;
  assign n3696 = ~pi0092 & ~n3681;
  assign n3697 = ~n3695 & n3696;
  assign n3698 = n2532 & ~n3680;
  assign n3699 = ~n3697 & n3698;
  assign n3700 = ~pi0055 & ~n3673;
  assign n3701 = ~n3699 & n3700;
  assign n3702 = ~pi0056 & ~n3670;
  assign n3703 = ~n3701 & n3702;
  assign n3704 = ~pi0062 & ~n3667;
  assign n3705 = ~n3703 & n3704;
  assign n3706 = ~pi0235 & n3328;
  assign n3707 = ~n3665 & n3706;
  assign n3708 = ~n3705 & n3707;
  assign n3709 = pi0235 & n3557;
  assign n3710 = ~n3328 & ~n3709;
  assign n3711 = n3555 & n3710;
  assign n3712 = ~n3708 & ~n3711;
  assign po0155 = ~n3659 & n3712;
  assign n3714 = pi0215 & pi1143;
  assign n3715 = pi0216 & pi0264;
  assign n3716 = ~pi0221 & ~n3715;
  assign n3717 = ~pi0105 & pi0146;
  assign n3718 = pi0284 & ~n2442;
  assign n3719 = pi0105 & ~n3718;
  assign n3720 = pi0228 & ~n3717;
  assign n3721 = ~n3719 & n3720;
  assign n3722 = ~n3447 & ~n3721;
  assign n3723 = ~pi0146 & ~pi0228;
  assign n3724 = n3722 & ~n3723;
  assign n3725 = ~pi0216 & ~n3724;
  assign n3726 = n3716 & ~n3725;
  assign n3727 = ~pi1143 & ~n2452;
  assign n3728 = ~pi0944 & n2452;
  assign n3729 = pi0221 & ~n3727;
  assign n3730 = ~n3728 & n3729;
  assign n3731 = ~n3726 & ~n3730;
  assign n3732 = ~pi0215 & ~n3731;
  assign n3733 = ~n3714 & ~n3732;
  assign n3734 = ~n3331 & n3733;
  assign n3735 = pi0284 & n2521;
  assign n3736 = ~n3384 & ~n3735;
  assign n3737 = ~pi0228 & ~n3736;
  assign n3738 = n3722 & ~n3737;
  assign n3739 = ~pi0216 & ~n3738;
  assign n3740 = n3716 & ~n3739;
  assign n3741 = ~n3730 & ~n3740;
  assign n3742 = ~pi0215 & ~n3741;
  assign n3743 = ~n3714 & ~n3742;
  assign n3744 = n3331 & n3743;
  assign n3745 = pi0062 & ~n3734;
  assign n3746 = ~n3744 & n3745;
  assign n3747 = ~n2537 & ~n3733;
  assign n3748 = n2537 & ~n3743;
  assign n3749 = pi0056 & ~n3747;
  assign n3750 = ~n3748 & n3749;
  assign n3751 = ~n2572 & n3733;
  assign n3752 = n2572 & n3743;
  assign n3753 = pi0055 & ~n3751;
  assign n3754 = ~n3752 & n3753;
  assign n3755 = n2442 & n2604;
  assign n3756 = pi0223 & pi1143;
  assign n3757 = pi0224 & pi0264;
  assign n3758 = ~pi0222 & ~n3757;
  assign n3759 = ~pi0224 & n3718;
  assign n3760 = n3758 & ~n3759;
  assign n3761 = ~pi1143 & ~n2591;
  assign n3762 = ~pi0944 & n2591;
  assign n3763 = pi0222 & ~n3761;
  assign n3764 = ~n3762 & n3763;
  assign n3765 = ~n3760 & ~n3764;
  assign n3766 = ~pi0223 & ~n3765;
  assign n3767 = ~n3756 & ~n3766;
  assign n3768 = ~pi0299 & ~n3767;
  assign n3769 = ~n3755 & n3768;
  assign n3770 = pi0299 & ~n3733;
  assign n3771 = ~n3769 & ~n3770;
  assign n3772 = ~n2532 & n3771;
  assign n3773 = ~n2625 & n3771;
  assign n3774 = pi0299 & ~n3743;
  assign n3775 = ~n3769 & ~n3774;
  assign n3776 = n2625 & n3775;
  assign n3777 = ~n3773 & ~n3776;
  assign n3778 = n2533 & ~n3777;
  assign n3779 = ~n2533 & n3771;
  assign n3780 = pi0092 & ~n3779;
  assign n3781 = ~n3778 & n3780;
  assign n3782 = pi0075 & n3771;
  assign n3783 = pi0087 & n3777;
  assign n3784 = pi0038 & n3771;
  assign n3785 = pi0039 & ~n3775;
  assign n3786 = ~pi0299 & ~n3756;
  assign n3787 = ~pi0284 & n3488;
  assign n3788 = ~pi0224 & ~n3787;
  assign n3789 = n3758 & ~n3788;
  assign n3790 = ~n3764 & ~n3789;
  assign n3791 = n3786 & n3790;
  assign n3792 = pi0299 & ~n3714;
  assign n3793 = n2441 & ~n3488;
  assign n3794 = ~pi0146 & ~n3508;
  assign n3795 = pi0146 & n3499;
  assign n3796 = ~pi0284 & ~n3795;
  assign n3797 = pi0146 & pi0284;
  assign n3798 = ~n3416 & n3797;
  assign n3799 = ~n3796 & ~n3798;
  assign n3800 = ~n3794 & ~n3799;
  assign n3801 = ~pi0228 & ~n3800;
  assign n3802 = ~n3721 & ~n3793;
  assign n3803 = ~n3801 & n3802;
  assign n3804 = ~pi0216 & ~n3803;
  assign n3805 = n3716 & ~n3804;
  assign n3806 = ~n3730 & ~n3805;
  assign n3807 = ~pi0215 & ~n3806;
  assign n3808 = n3792 & ~n3807;
  assign n3809 = ~n3488 & n3758;
  assign n3810 = n3790 & ~n3809;
  assign n3811 = ~pi0223 & ~n3810;
  assign n3812 = n3786 & ~n3811;
  assign n3813 = ~pi0039 & ~n3812;
  assign n3814 = ~n3791 & n3813;
  assign n3815 = ~n3808 & n3814;
  assign n3816 = ~pi0038 & ~n3785;
  assign n3817 = ~n3815 & n3816;
  assign n3818 = ~pi0100 & ~n3784;
  assign n3819 = ~n3817 & n3818;
  assign n3820 = ~n2530 & n3771;
  assign n3821 = pi0252 & n2639;
  assign n3822 = ~pi0284 & ~n3821;
  assign n3823 = n2521 & n3822;
  assign n3824 = ~pi0228 & ~n3823;
  assign n3825 = ~n3386 & n3824;
  assign n3826 = n3722 & ~n3825;
  assign n3827 = ~pi0216 & ~n3826;
  assign n3828 = n3716 & ~n3827;
  assign n3829 = ~n3730 & ~n3828;
  assign n3830 = ~pi0215 & ~n3829;
  assign n3831 = ~n3714 & ~n3830;
  assign n3832 = pi0299 & ~n3831;
  assign n3833 = n2530 & ~n3769;
  assign n3834 = ~n3832 & n3833;
  assign n3835 = pi0100 & ~n3820;
  assign n3836 = ~n3834 & n3835;
  assign n3837 = ~n3819 & ~n3836;
  assign n3838 = ~pi0087 & ~n3837;
  assign n3839 = ~pi0075 & ~n3783;
  assign n3840 = ~n3838 & n3839;
  assign n3841 = ~pi0092 & ~n3782;
  assign n3842 = ~n3840 & n3841;
  assign n3843 = n2532 & ~n3781;
  assign n3844 = ~n3842 & n3843;
  assign n3845 = ~pi0055 & ~n3772;
  assign n3846 = ~n3844 & n3845;
  assign n3847 = ~pi0056 & ~n3754;
  assign n3848 = ~n3846 & n3847;
  assign n3849 = ~pi0062 & ~n3750;
  assign n3850 = ~n3848 & n3849;
  assign n3851 = ~pi0238 & n3328;
  assign n3852 = ~n3746 & n3851;
  assign n3853 = ~n3850 & n3852;
  assign n3854 = ~n3721 & ~n3737;
  assign n3855 = ~pi0216 & ~n3854;
  assign n3856 = n3716 & ~n3855;
  assign n3857 = ~n3730 & ~n3856;
  assign n3858 = ~pi0215 & ~n3857;
  assign n3859 = ~n3714 & ~n3858;
  assign n3860 = n3331 & n3859;
  assign n3861 = n3556 & ~n3715;
  assign n3862 = n3733 & ~n3861;
  assign n3863 = ~n3331 & n3862;
  assign n3864 = pi0062 & ~n3863;
  assign n3865 = ~n3860 & n3864;
  assign n3866 = ~n2537 & ~n3862;
  assign n3867 = n2537 & ~n3859;
  assign n3868 = pi0056 & ~n3866;
  assign n3869 = ~n3867 & n3868;
  assign n3870 = n2572 & n3859;
  assign n3871 = ~n2572 & n3862;
  assign n3872 = pi0055 & ~n3871;
  assign n3873 = ~n3870 & n3872;
  assign n3874 = pi0299 & ~n3862;
  assign n3875 = ~n3768 & ~n3874;
  assign n3876 = ~n2532 & n3875;
  assign n3877 = ~n2625 & n3875;
  assign n3878 = pi0299 & ~n3859;
  assign n3879 = ~n3768 & ~n3878;
  assign n3880 = n2625 & n3879;
  assign n3881 = ~n3877 & ~n3880;
  assign n3882 = n2533 & ~n3881;
  assign n3883 = ~n2533 & n3875;
  assign n3884 = pi0092 & ~n3883;
  assign n3885 = ~n3882 & n3884;
  assign n3886 = pi0075 & n3875;
  assign n3887 = pi0087 & n3881;
  assign n3888 = pi0038 & n3875;
  assign n3889 = pi0039 & ~n3879;
  assign n3890 = ~n3497 & n3721;
  assign n3891 = ~pi0146 & n3499;
  assign n3892 = pi0146 & ~n3508;
  assign n3893 = pi0284 & ~n3891;
  assign n3894 = ~n3892 & n3893;
  assign n3895 = ~pi0146 & ~pi0284;
  assign n3896 = ~n3416 & n3895;
  assign n3897 = ~n3894 & ~n3896;
  assign n3898 = ~pi0228 & ~n3897;
  assign n3899 = ~n3890 & ~n3898;
  assign n3900 = ~pi0216 & ~n3899;
  assign n3901 = n3716 & ~n3900;
  assign n3902 = ~n3730 & ~n3901;
  assign n3903 = ~pi0215 & ~n3902;
  assign n3904 = n3792 & ~n3903;
  assign n3905 = n3813 & ~n3904;
  assign n3906 = ~pi0038 & ~n3889;
  assign n3907 = ~n3905 & n3906;
  assign n3908 = ~pi0100 & ~n3888;
  assign n3909 = ~n3907 & n3908;
  assign n3910 = ~n2530 & n3875;
  assign n3911 = ~n3721 & ~n3825;
  assign n3912 = ~pi0216 & ~n3911;
  assign n3913 = n3716 & ~n3912;
  assign n3914 = ~n3730 & ~n3913;
  assign n3915 = ~pi0215 & ~n3914;
  assign n3916 = ~n3714 & ~n3915;
  assign n3917 = pi0299 & ~n3916;
  assign n3918 = n2530 & ~n3768;
  assign n3919 = ~n3917 & n3918;
  assign n3920 = pi0100 & ~n3910;
  assign n3921 = ~n3919 & n3920;
  assign n3922 = ~n3909 & ~n3921;
  assign n3923 = ~pi0087 & ~n3922;
  assign n3924 = ~pi0075 & ~n3887;
  assign n3925 = ~n3923 & n3924;
  assign n3926 = ~pi0092 & ~n3886;
  assign n3927 = ~n3925 & n3926;
  assign n3928 = n2532 & ~n3885;
  assign n3929 = ~n3927 & n3928;
  assign n3930 = ~pi0055 & ~n3876;
  assign n3931 = ~n3929 & n3930;
  assign n3932 = ~pi0056 & ~n3873;
  assign n3933 = ~n3931 & n3932;
  assign n3934 = ~pi0062 & ~n3869;
  assign n3935 = ~n3933 & n3934;
  assign n3936 = pi0238 & n3328;
  assign n3937 = ~n3865 & n3936;
  assign n3938 = ~n3935 & n3937;
  assign n3939 = pi0238 & n3861;
  assign n3940 = ~n3328 & ~n3939;
  assign n3941 = n3733 & n3940;
  assign n3942 = ~n3853 & ~n3941;
  assign po0156 = ~n3938 & n3942;
  assign n3944 = pi0215 & pi1142;
  assign n3945 = pi0216 & pi0277;
  assign n3946 = ~pi0221 & ~n3945;
  assign n3947 = pi0172 & ~pi0228;
  assign n3948 = ~pi0105 & pi0172;
  assign n3949 = pi0262 & ~n2442;
  assign n3950 = pi0105 & n3949;
  assign n3951 = ~n3948 & ~n3950;
  assign n3952 = pi0228 & ~n3951;
  assign n3953 = ~n3947 & ~n3952;
  assign n3954 = ~pi0216 & ~n3953;
  assign n3955 = n3946 & ~n3954;
  assign n3956 = ~pi1142 & ~n2452;
  assign n3957 = ~pi0932 & n2452;
  assign n3958 = pi0221 & ~n3956;
  assign n3959 = ~n3957 & n3958;
  assign n3960 = ~n3955 & ~n3959;
  assign n3961 = ~pi0215 & ~n3960;
  assign n3962 = ~n3944 & ~n3961;
  assign n3963 = ~n3450 & ~n3962;
  assign n3964 = ~n3328 & ~n3963;
  assign n3965 = ~n3331 & ~n3963;
  assign n3966 = ~pi0262 & n2521;
  assign n3967 = ~n3335 & ~n3947;
  assign n3968 = ~n3966 & ~n3967;
  assign n3969 = ~n3447 & ~n3952;
  assign n3970 = ~n3968 & n3969;
  assign n3971 = ~pi0216 & ~n3970;
  assign n3972 = n3946 & ~n3971;
  assign n3973 = ~n3959 & ~n3972;
  assign n3974 = ~pi0215 & ~n3973;
  assign n3975 = ~n3944 & ~n3974;
  assign n3976 = n3331 & n3975;
  assign n3977 = pi0062 & ~n3965;
  assign n3978 = ~n3976 & n3977;
  assign n3979 = n2537 & ~n3975;
  assign n3980 = ~n2537 & n3963;
  assign n3981 = pi0056 & ~n3980;
  assign n3982 = ~n3979 & n3981;
  assign n3983 = ~n2572 & ~n3963;
  assign n3984 = n2572 & n3975;
  assign n3985 = pi0055 & ~n3983;
  assign n3986 = ~n3984 & n3985;
  assign n3987 = pi0223 & pi1142;
  assign n3988 = pi0224 & pi0277;
  assign n3989 = ~pi0222 & ~n3988;
  assign n3990 = ~pi0224 & n3949;
  assign n3991 = n3989 & ~n3990;
  assign n3992 = ~pi1142 & ~n2591;
  assign n3993 = ~pi0932 & n2591;
  assign n3994 = pi0222 & ~n3992;
  assign n3995 = ~n3993 & n3994;
  assign n3996 = ~n3991 & ~n3995;
  assign n3997 = ~pi0223 & ~n3996;
  assign n3998 = ~n3987 & ~n3997;
  assign n3999 = ~pi0299 & ~n3998;
  assign n4000 = ~n3755 & n3999;
  assign n4001 = pi0299 & n3963;
  assign n4002 = ~n4000 & ~n4001;
  assign n4003 = ~n2532 & n4002;
  assign n4004 = ~n2625 & n4002;
  assign n4005 = pi0299 & ~n3975;
  assign n4006 = ~n4000 & ~n4005;
  assign n4007 = n2625 & n4006;
  assign n4008 = ~n4004 & ~n4007;
  assign n4009 = n2533 & ~n4008;
  assign n4010 = ~n2533 & n4002;
  assign n4011 = pi0092 & ~n4010;
  assign n4012 = ~n4009 & n4011;
  assign n4013 = pi0075 & n4002;
  assign n4014 = pi0087 & n4008;
  assign n4015 = pi0038 & n4002;
  assign n4016 = pi0039 & ~n4006;
  assign n4017 = ~pi0299 & ~n3987;
  assign n4018 = ~pi0262 & n3488;
  assign n4019 = ~pi0224 & ~n4018;
  assign n4020 = n3989 & ~n4019;
  assign n4021 = ~n3995 & ~n4020;
  assign n4022 = n4017 & n4021;
  assign n4023 = pi0299 & ~n3944;
  assign n4024 = pi0262 & n3416;
  assign n4025 = ~pi0262 & n3499;
  assign n4026 = ~pi0172 & ~n4025;
  assign n4027 = pi0172 & ~pi0262;
  assign n4028 = n3508 & n4027;
  assign n4029 = ~n4026 & ~n4028;
  assign n4030 = ~pi0228 & ~n4024;
  assign n4031 = ~n4029 & n4030;
  assign n4032 = ~n3487 & n3950;
  assign n4033 = pi0228 & ~n3948;
  assign n4034 = ~n4032 & n4033;
  assign n4035 = ~n3497 & n4034;
  assign n4036 = ~pi0216 & ~n4035;
  assign n4037 = ~n4031 & n4036;
  assign n4038 = n3946 & ~n4037;
  assign n4039 = ~n3959 & ~n4038;
  assign n4040 = ~pi0215 & ~n4039;
  assign n4041 = n4023 & ~n4040;
  assign n4042 = ~n3488 & n3989;
  assign n4043 = n4021 & ~n4042;
  assign n4044 = ~pi0223 & ~n4043;
  assign n4045 = n4017 & ~n4044;
  assign n4046 = ~pi0039 & ~n4045;
  assign n4047 = ~n4022 & n4046;
  assign n4048 = ~n4041 & n4047;
  assign n4049 = ~pi0038 & ~n4016;
  assign n4050 = ~n4048 & n4049;
  assign n4051 = ~pi0100 & ~n4015;
  assign n4052 = ~n4050 & n4051;
  assign n4053 = ~n2530 & n4002;
  assign n4054 = ~pi0262 & n3394;
  assign n4055 = ~n3629 & ~n3947;
  assign n4056 = ~n4054 & ~n4055;
  assign n4057 = n3969 & ~n4056;
  assign n4058 = ~pi0216 & ~n4057;
  assign n4059 = n3946 & ~n4058;
  assign n4060 = ~n3959 & ~n4059;
  assign n4061 = ~pi0215 & ~n4060;
  assign n4062 = ~n3944 & ~n4061;
  assign n4063 = pi0299 & ~n4062;
  assign n4064 = n2530 & ~n4000;
  assign n4065 = ~n4063 & n4064;
  assign n4066 = pi0100 & ~n4053;
  assign n4067 = ~n4065 & n4066;
  assign n4068 = ~n4052 & ~n4067;
  assign n4069 = ~pi0087 & ~n4068;
  assign n4070 = ~pi0075 & ~n4014;
  assign n4071 = ~n4069 & n4070;
  assign n4072 = ~pi0092 & ~n4013;
  assign n4073 = ~n4071 & n4072;
  assign n4074 = n2532 & ~n4012;
  assign n4075 = ~n4073 & n4074;
  assign n4076 = ~pi0055 & ~n4003;
  assign n4077 = ~n4075 & n4076;
  assign n4078 = ~pi0056 & ~n3986;
  assign n4079 = ~n4077 & n4078;
  assign n4080 = ~pi0062 & ~n3982;
  assign n4081 = ~n4079 & n4080;
  assign n4082 = n3328 & ~n3978;
  assign n4083 = ~n4081 & n4082;
  assign n4084 = ~pi0249 & ~n3964;
  assign n4085 = ~n4083 & n4084;
  assign n4086 = ~n3328 & n3962;
  assign n4087 = ~n3331 & n3962;
  assign n4088 = ~n3952 & ~n3968;
  assign n4089 = ~pi0216 & ~n4088;
  assign n4090 = n3946 & ~n4089;
  assign n4091 = ~n3959 & ~n4090;
  assign n4092 = ~pi0215 & ~n4091;
  assign n4093 = ~n3944 & ~n4092;
  assign n4094 = n3331 & n4093;
  assign n4095 = pi0062 & ~n4087;
  assign n4096 = ~n4094 & n4095;
  assign n4097 = ~n2537 & ~n3962;
  assign n4098 = n2537 & ~n4093;
  assign n4099 = pi0056 & ~n4097;
  assign n4100 = ~n4098 & n4099;
  assign n4101 = ~n2572 & n3962;
  assign n4102 = n2572 & n4093;
  assign n4103 = pi0055 & ~n4101;
  assign n4104 = ~n4102 & n4103;
  assign n4105 = pi0299 & ~n3962;
  assign n4106 = ~n3999 & ~n4105;
  assign n4107 = ~n2532 & n4106;
  assign n4108 = ~n2625 & n4106;
  assign n4109 = pi0299 & ~n4093;
  assign n4110 = ~n3999 & ~n4109;
  assign n4111 = n2625 & n4110;
  assign n4112 = ~n4108 & ~n4111;
  assign n4113 = n2533 & ~n4112;
  assign n4114 = ~n2533 & n4106;
  assign n4115 = pi0092 & ~n4114;
  assign n4116 = ~n4113 & n4115;
  assign n4117 = pi0075 & n4106;
  assign n4118 = pi0087 & n4112;
  assign n4119 = pi0038 & n4106;
  assign n4120 = pi0039 & ~n4110;
  assign n4121 = pi0262 & n3508;
  assign n4122 = ~pi0172 & ~n4121;
  assign n4123 = pi0262 & ~n3499;
  assign n4124 = ~pi0262 & ~n3416;
  assign n4125 = pi0172 & ~n4123;
  assign n4126 = ~n4124 & n4125;
  assign n4127 = ~n4122 & ~n4126;
  assign n4128 = ~pi0228 & ~n4127;
  assign n4129 = ~pi0216 & ~n4034;
  assign n4130 = ~n4128 & n4129;
  assign n4131 = n3946 & ~n4130;
  assign n4132 = ~n3959 & ~n4131;
  assign n4133 = ~pi0215 & ~n4132;
  assign n4134 = n4023 & ~n4133;
  assign n4135 = n4046 & ~n4134;
  assign n4136 = ~pi0038 & ~n4120;
  assign n4137 = ~n4135 & n4136;
  assign n4138 = ~pi0100 & ~n4119;
  assign n4139 = ~n4137 & n4138;
  assign n4140 = ~n2530 & n4106;
  assign n4141 = ~n3952 & ~n4056;
  assign n4142 = ~pi0216 & ~n4141;
  assign n4143 = n3946 & ~n4142;
  assign n4144 = ~n3959 & ~n4143;
  assign n4145 = ~pi0215 & ~n4144;
  assign n4146 = ~n3944 & ~n4145;
  assign n4147 = pi0299 & ~n4146;
  assign n4148 = n2530 & ~n3999;
  assign n4149 = ~n4147 & n4148;
  assign n4150 = pi0100 & ~n4140;
  assign n4151 = ~n4149 & n4150;
  assign n4152 = ~n4139 & ~n4151;
  assign n4153 = ~pi0087 & ~n4152;
  assign n4154 = ~pi0075 & ~n4118;
  assign n4155 = ~n4153 & n4154;
  assign n4156 = ~pi0092 & ~n4117;
  assign n4157 = ~n4155 & n4156;
  assign n4158 = n2532 & ~n4116;
  assign n4159 = ~n4157 & n4158;
  assign n4160 = ~pi0055 & ~n4107;
  assign n4161 = ~n4159 & n4160;
  assign n4162 = ~pi0056 & ~n4104;
  assign n4163 = ~n4161 & n4162;
  assign n4164 = ~pi0062 & ~n4100;
  assign n4165 = ~n4163 & n4164;
  assign n4166 = n3328 & ~n4096;
  assign n4167 = ~n4165 & n4166;
  assign n4168 = pi0249 & ~n4086;
  assign n4169 = ~n4167 & n4168;
  assign po0157 = n4085 | n4169;
  assign n4171 = pi0215 & pi1141;
  assign n4172 = pi0216 & pi0270;
  assign n4173 = ~pi0221 & ~n4172;
  assign n4174 = ~pi0105 & pi0171;
  assign n4175 = pi0861 & ~n2442;
  assign n4176 = pi0105 & ~n4175;
  assign n4177 = pi0228 & ~n4174;
  assign n4178 = ~n4176 & n4177;
  assign n4179 = ~pi0216 & ~n4178;
  assign n4180 = ~pi0171 & ~pi0228;
  assign n4181 = n4179 & ~n4180;
  assign n4182 = n4173 & ~n4181;
  assign n4183 = ~pi1141 & ~n2452;
  assign n4184 = ~pi0935 & n2452;
  assign n4185 = pi0221 & ~n4183;
  assign n4186 = ~n4184 & n4185;
  assign n4187 = ~n4182 & ~n4186;
  assign n4188 = ~pi0215 & ~n4187;
  assign n4189 = ~n4171 & ~n4188;
  assign n4190 = ~n3331 & n4189;
  assign n4191 = ~pi0861 & n2521;
  assign n4192 = pi0171 & ~n2521;
  assign n4193 = ~pi0228 & ~n4191;
  assign n4194 = ~n4192 & n4193;
  assign n4195 = n4179 & ~n4194;
  assign n4196 = n4173 & ~n4195;
  assign n4197 = ~n4186 & ~n4196;
  assign n4198 = ~pi0215 & ~n4197;
  assign n4199 = ~n4171 & ~n4198;
  assign n4200 = n3331 & n4199;
  assign n4201 = pi0062 & ~n4190;
  assign n4202 = ~n4200 & n4201;
  assign n4203 = ~n2537 & ~n4189;
  assign n4204 = n2537 & ~n4199;
  assign n4205 = pi0056 & ~n4203;
  assign n4206 = ~n4204 & n4205;
  assign n4207 = ~n2572 & n4189;
  assign n4208 = n2572 & n4199;
  assign n4209 = pi0055 & ~n4207;
  assign n4210 = ~n4208 & n4209;
  assign n4211 = pi0223 & pi1141;
  assign n4212 = pi0224 & pi0270;
  assign n4213 = ~pi0222 & ~n4212;
  assign n4214 = ~pi0224 & ~n4175;
  assign n4215 = n4213 & ~n4214;
  assign n4216 = ~pi1141 & ~n2591;
  assign n4217 = ~pi0935 & n2591;
  assign n4218 = pi0222 & ~n4216;
  assign n4219 = ~n4217 & n4218;
  assign n4220 = ~n4215 & ~n4219;
  assign n4221 = ~pi0223 & ~n4220;
  assign n4222 = ~n4211 & ~n4221;
  assign n4223 = ~pi0299 & ~n4222;
  assign n4224 = pi0299 & ~n4189;
  assign n4225 = ~n4223 & ~n4224;
  assign n4226 = ~n2532 & n4225;
  assign n4227 = ~n2625 & n4225;
  assign n4228 = pi0299 & ~n4199;
  assign n4229 = ~n4223 & ~n4228;
  assign n4230 = n2625 & n4229;
  assign n4231 = ~n4227 & ~n4230;
  assign n4232 = n2533 & ~n4231;
  assign n4233 = ~n2533 & n4225;
  assign n4234 = pi0092 & ~n4233;
  assign n4235 = ~n4232 & n4234;
  assign n4236 = pi0075 & n4225;
  assign n4237 = pi0087 & n4231;
  assign n4238 = pi0038 & n4225;
  assign n4239 = pi0039 & ~n4229;
  assign n4240 = ~pi0299 & ~n4211;
  assign n4241 = pi0861 & n3488;
  assign n4242 = ~pi0224 & ~n4241;
  assign n4243 = n4213 & ~n4242;
  assign n4244 = ~n4219 & ~n4243;
  assign n4245 = n4240 & n4244;
  assign n4246 = pi0299 & ~n4171;
  assign n4247 = pi0861 & n3499;
  assign n4248 = ~pi0171 & ~n4247;
  assign n4249 = pi0171 & n3508;
  assign n4250 = ~n4248 & ~n4249;
  assign n4251 = pi0861 & ~n4250;
  assign n4252 = ~n3416 & n4248;
  assign n4253 = ~n4251 & ~n4252;
  assign n4254 = ~pi0228 & ~n4253;
  assign n4255 = ~n3497 & n4178;
  assign n4256 = ~pi0216 & ~n4255;
  assign n4257 = ~n4254 & n4256;
  assign n4258 = n4173 & ~n4257;
  assign n4259 = ~n4186 & ~n4258;
  assign n4260 = ~pi0215 & ~n4259;
  assign n4261 = n4246 & ~n4260;
  assign n4262 = ~n3488 & n4213;
  assign n4263 = n4244 & ~n4262;
  assign n4264 = ~pi0223 & ~n4263;
  assign n4265 = n4240 & ~n4264;
  assign n4266 = ~pi0039 & ~n4265;
  assign n4267 = ~n4245 & n4266;
  assign n4268 = ~n4261 & n4267;
  assign n4269 = ~pi0038 & ~n4239;
  assign n4270 = ~n4268 & n4269;
  assign n4271 = ~pi0100 & ~n4238;
  assign n4272 = ~n4270 & n4271;
  assign n4273 = ~n2530 & n4225;
  assign n4274 = ~pi0861 & n3394;
  assign n4275 = pi0171 & ~n3394;
  assign n4276 = ~pi0228 & ~n4274;
  assign n4277 = ~n4275 & n4276;
  assign n4278 = n4179 & ~n4277;
  assign n4279 = n4173 & ~n4278;
  assign n4280 = ~n4186 & ~n4279;
  assign n4281 = ~pi0215 & ~n4280;
  assign n4282 = ~n4171 & ~n4281;
  assign n4283 = pi0299 & ~n4282;
  assign n4284 = n2530 & ~n4223;
  assign n4285 = ~n4283 & n4284;
  assign n4286 = pi0100 & ~n4273;
  assign n4287 = ~n4285 & n4286;
  assign n4288 = ~n4272 & ~n4287;
  assign n4289 = ~pi0087 & ~n4288;
  assign n4290 = ~pi0075 & ~n4237;
  assign n4291 = ~n4289 & n4290;
  assign n4292 = ~pi0092 & ~n4236;
  assign n4293 = ~n4291 & n4292;
  assign n4294 = n2532 & ~n4235;
  assign n4295 = ~n4293 & n4294;
  assign n4296 = ~pi0055 & ~n4226;
  assign n4297 = ~n4295 & n4296;
  assign n4298 = ~pi0056 & ~n4210;
  assign n4299 = ~n4297 & n4298;
  assign n4300 = ~pi0062 & ~n4206;
  assign n4301 = ~n4299 & n4300;
  assign n4302 = ~pi0241 & n3328;
  assign n4303 = ~n4202 & n4302;
  assign n4304 = ~n4301 & n4303;
  assign n4305 = ~n3447 & n4179;
  assign n4306 = ~n4194 & n4305;
  assign n4307 = n4173 & ~n4306;
  assign n4308 = ~n4186 & ~n4307;
  assign n4309 = ~pi0215 & ~n4308;
  assign n4310 = ~n4171 & ~n4309;
  assign n4311 = n3331 & n4310;
  assign n4312 = n3556 & ~n4172;
  assign n4313 = n4189 & ~n4312;
  assign n4314 = ~n3331 & n4313;
  assign n4315 = pi0062 & ~n4314;
  assign n4316 = ~n4311 & n4315;
  assign n4317 = ~n2537 & ~n4313;
  assign n4318 = n2537 & ~n4310;
  assign n4319 = pi0056 & ~n4317;
  assign n4320 = ~n4318 & n4319;
  assign n4321 = n2572 & n4310;
  assign n4322 = ~n2572 & n4313;
  assign n4323 = pi0055 & ~n4322;
  assign n4324 = ~n4321 & n4323;
  assign n4325 = ~n3472 & ~n4223;
  assign n4326 = pi0299 & ~n4313;
  assign n4327 = n4325 & ~n4326;
  assign n4328 = ~n2532 & n4327;
  assign n4329 = ~n2625 & n4327;
  assign n4330 = pi0299 & ~n4310;
  assign n4331 = n4325 & ~n4330;
  assign n4332 = n2625 & n4331;
  assign n4333 = ~n4329 & ~n4332;
  assign n4334 = n2533 & ~n4333;
  assign n4335 = ~n2533 & n4327;
  assign n4336 = pi0092 & ~n4335;
  assign n4337 = ~n4334 & n4336;
  assign n4338 = pi0075 & n4327;
  assign n4339 = pi0087 & n4333;
  assign n4340 = pi0038 & n4327;
  assign n4341 = pi0039 & ~n4331;
  assign n4342 = ~pi0861 & n3508;
  assign n4343 = ~pi0171 & ~n4342;
  assign n4344 = ~pi0861 & ~n3499;
  assign n4345 = pi0861 & ~n3416;
  assign n4346 = pi0171 & ~n4344;
  assign n4347 = ~n4345 & n4346;
  assign n4348 = ~n4343 & ~n4347;
  assign n4349 = ~pi0228 & ~n4348;
  assign n4350 = ~n3793 & n4179;
  assign n4351 = ~n4349 & n4350;
  assign n4352 = n4173 & ~n4351;
  assign n4353 = ~n4186 & ~n4352;
  assign n4354 = ~pi0215 & ~n4353;
  assign n4355 = n4246 & ~n4354;
  assign n4356 = n4266 & ~n4355;
  assign n4357 = ~pi0038 & ~n4341;
  assign n4358 = ~n4356 & n4357;
  assign n4359 = ~pi0100 & ~n4340;
  assign n4360 = ~n4358 & n4359;
  assign n4361 = ~n2530 & n4327;
  assign n4362 = ~n4277 & n4305;
  assign n4363 = n4173 & ~n4362;
  assign n4364 = ~n4186 & ~n4363;
  assign n4365 = ~pi0215 & ~n4364;
  assign n4366 = ~n4171 & ~n4365;
  assign n4367 = pi0299 & ~n4366;
  assign n4368 = n2530 & n4325;
  assign n4369 = ~n4367 & n4368;
  assign n4370 = pi0100 & ~n4361;
  assign n4371 = ~n4369 & n4370;
  assign n4372 = ~n4360 & ~n4371;
  assign n4373 = ~pi0087 & ~n4372;
  assign n4374 = ~pi0075 & ~n4339;
  assign n4375 = ~n4373 & n4374;
  assign n4376 = ~pi0092 & ~n4338;
  assign n4377 = ~n4375 & n4376;
  assign n4378 = n2532 & ~n4337;
  assign n4379 = ~n4377 & n4378;
  assign n4380 = ~pi0055 & ~n4328;
  assign n4381 = ~n4379 & n4380;
  assign n4382 = ~pi0056 & ~n4324;
  assign n4383 = ~n4381 & n4382;
  assign n4384 = ~pi0062 & ~n4320;
  assign n4385 = ~n4383 & n4384;
  assign n4386 = pi0241 & n3328;
  assign n4387 = ~n4316 & n4386;
  assign n4388 = ~n4385 & n4387;
  assign n4389 = pi0241 & n4312;
  assign n4390 = ~n3328 & ~n4389;
  assign n4391 = n4189 & n4390;
  assign n4392 = ~n4388 & ~n4391;
  assign po0158 = ~n4304 & n4392;
  assign n4394 = pi0215 & pi1140;
  assign n4395 = pi0216 & pi0282;
  assign n4396 = ~pi0221 & ~n4395;
  assign n4397 = ~pi0105 & pi0170;
  assign n4398 = pi0869 & ~n2442;
  assign n4399 = pi0105 & ~n4398;
  assign n4400 = pi0228 & ~n4397;
  assign n4401 = ~n4399 & n4400;
  assign n4402 = ~pi0216 & ~n4401;
  assign n4403 = ~pi0170 & ~pi0228;
  assign n4404 = n4402 & ~n4403;
  assign n4405 = n4396 & ~n4404;
  assign n4406 = ~pi1140 & ~n2452;
  assign n4407 = ~pi0921 & n2452;
  assign n4408 = pi0221 & ~n4406;
  assign n4409 = ~n4407 & n4408;
  assign n4410 = ~n4405 & ~n4409;
  assign n4411 = ~pi0215 & ~n4410;
  assign n4412 = ~n4394 & ~n4411;
  assign n4413 = ~n3331 & n4412;
  assign n4414 = ~pi0869 & n2521;
  assign n4415 = pi0170 & ~n2521;
  assign n4416 = ~pi0228 & ~n4414;
  assign n4417 = ~n4415 & n4416;
  assign n4418 = n4402 & ~n4417;
  assign n4419 = n4396 & ~n4418;
  assign n4420 = ~n4409 & ~n4419;
  assign n4421 = ~pi0215 & ~n4420;
  assign n4422 = ~n4394 & ~n4421;
  assign n4423 = n3331 & n4422;
  assign n4424 = pi0062 & ~n4413;
  assign n4425 = ~n4423 & n4424;
  assign n4426 = ~n2537 & ~n4412;
  assign n4427 = n2537 & ~n4422;
  assign n4428 = pi0056 & ~n4426;
  assign n4429 = ~n4427 & n4428;
  assign n4430 = ~n2572 & n4412;
  assign n4431 = n2572 & n4422;
  assign n4432 = pi0055 & ~n4430;
  assign n4433 = ~n4431 & n4432;
  assign n4434 = pi0223 & pi1140;
  assign n4435 = pi0224 & pi0282;
  assign n4436 = ~pi0222 & ~n4435;
  assign n4437 = ~pi0224 & ~n4398;
  assign n4438 = n4436 & ~n4437;
  assign n4439 = ~pi1140 & ~n2591;
  assign n4440 = ~pi0921 & n2591;
  assign n4441 = pi0222 & ~n4439;
  assign n4442 = ~n4440 & n4441;
  assign n4443 = ~n4438 & ~n4442;
  assign n4444 = ~pi0223 & ~n4443;
  assign n4445 = ~n4434 & ~n4444;
  assign n4446 = ~pi0299 & ~n4445;
  assign n4447 = pi0299 & ~n4412;
  assign n4448 = ~n4446 & ~n4447;
  assign n4449 = ~n2532 & n4448;
  assign n4450 = ~n2625 & n4448;
  assign n4451 = pi0299 & ~n4422;
  assign n4452 = ~n4446 & ~n4451;
  assign n4453 = n2625 & n4452;
  assign n4454 = ~n4450 & ~n4453;
  assign n4455 = n2533 & ~n4454;
  assign n4456 = ~n2533 & n4448;
  assign n4457 = pi0092 & ~n4456;
  assign n4458 = ~n4455 & n4457;
  assign n4459 = pi0075 & n4448;
  assign n4460 = pi0087 & n4454;
  assign n4461 = pi0038 & n4448;
  assign n4462 = pi0039 & ~n4452;
  assign n4463 = ~pi0299 & ~n4434;
  assign n4464 = pi0869 & n3488;
  assign n4465 = ~pi0224 & ~n4464;
  assign n4466 = n4436 & ~n4465;
  assign n4467 = ~n4442 & ~n4466;
  assign n4468 = n4463 & n4467;
  assign n4469 = pi0299 & ~n4394;
  assign n4470 = pi0869 & n3499;
  assign n4471 = ~pi0170 & ~n4470;
  assign n4472 = pi0170 & n3508;
  assign n4473 = ~n4471 & ~n4472;
  assign n4474 = pi0869 & ~n4473;
  assign n4475 = ~n3416 & n4471;
  assign n4476 = ~n4474 & ~n4475;
  assign n4477 = ~pi0228 & ~n4476;
  assign n4478 = ~n3497 & n4401;
  assign n4479 = ~pi0216 & ~n4478;
  assign n4480 = ~n4477 & n4479;
  assign n4481 = n4396 & ~n4480;
  assign n4482 = ~n4409 & ~n4481;
  assign n4483 = ~pi0215 & ~n4482;
  assign n4484 = n4469 & ~n4483;
  assign n4485 = ~n3488 & n4436;
  assign n4486 = n4467 & ~n4485;
  assign n4487 = ~pi0223 & ~n4486;
  assign n4488 = n4463 & ~n4487;
  assign n4489 = ~pi0039 & ~n4488;
  assign n4490 = ~n4468 & n4489;
  assign n4491 = ~n4484 & n4490;
  assign n4492 = ~pi0038 & ~n4462;
  assign n4493 = ~n4491 & n4492;
  assign n4494 = ~pi0100 & ~n4461;
  assign n4495 = ~n4493 & n4494;
  assign n4496 = ~n2530 & n4448;
  assign n4497 = ~pi0869 & n3394;
  assign n4498 = pi0170 & ~n3394;
  assign n4499 = ~pi0228 & ~n4497;
  assign n4500 = ~n4498 & n4499;
  assign n4501 = n4402 & ~n4500;
  assign n4502 = n4396 & ~n4501;
  assign n4503 = ~n4409 & ~n4502;
  assign n4504 = ~pi0215 & ~n4503;
  assign n4505 = ~n4394 & ~n4504;
  assign n4506 = pi0299 & ~n4505;
  assign n4507 = n2530 & ~n4446;
  assign n4508 = ~n4506 & n4507;
  assign n4509 = pi0100 & ~n4496;
  assign n4510 = ~n4508 & n4509;
  assign n4511 = ~n4495 & ~n4510;
  assign n4512 = ~pi0087 & ~n4511;
  assign n4513 = ~pi0075 & ~n4460;
  assign n4514 = ~n4512 & n4513;
  assign n4515 = ~pi0092 & ~n4459;
  assign n4516 = ~n4514 & n4515;
  assign n4517 = n2532 & ~n4458;
  assign n4518 = ~n4516 & n4517;
  assign n4519 = ~pi0055 & ~n4449;
  assign n4520 = ~n4518 & n4519;
  assign n4521 = ~pi0056 & ~n4433;
  assign n4522 = ~n4520 & n4521;
  assign n4523 = ~pi0062 & ~n4429;
  assign n4524 = ~n4522 & n4523;
  assign n4525 = ~pi0248 & n3328;
  assign n4526 = ~n4425 & n4525;
  assign n4527 = ~n4524 & n4526;
  assign n4528 = ~n3447 & n4402;
  assign n4529 = ~n4417 & n4528;
  assign n4530 = n4396 & ~n4529;
  assign n4531 = ~n4409 & ~n4530;
  assign n4532 = ~pi0215 & ~n4531;
  assign n4533 = ~n4394 & ~n4532;
  assign n4534 = n3331 & n4533;
  assign n4535 = n3556 & ~n4395;
  assign n4536 = n4412 & ~n4535;
  assign n4537 = ~n3331 & n4536;
  assign n4538 = pi0062 & ~n4537;
  assign n4539 = ~n4534 & n4538;
  assign n4540 = ~n2537 & ~n4536;
  assign n4541 = n2537 & ~n4533;
  assign n4542 = pi0056 & ~n4540;
  assign n4543 = ~n4541 & n4542;
  assign n4544 = n2572 & n4533;
  assign n4545 = ~n2572 & n4536;
  assign n4546 = pi0055 & ~n4545;
  assign n4547 = ~n4544 & n4546;
  assign n4548 = ~n3472 & ~n4446;
  assign n4549 = pi0299 & ~n4536;
  assign n4550 = n4548 & ~n4549;
  assign n4551 = ~n2532 & n4550;
  assign n4552 = ~n2625 & n4550;
  assign n4553 = pi0299 & ~n4533;
  assign n4554 = n4548 & ~n4553;
  assign n4555 = n2625 & n4554;
  assign n4556 = ~n4552 & ~n4555;
  assign n4557 = n2533 & ~n4556;
  assign n4558 = ~n2533 & n4550;
  assign n4559 = pi0092 & ~n4558;
  assign n4560 = ~n4557 & n4559;
  assign n4561 = pi0075 & n4550;
  assign n4562 = pi0087 & n4556;
  assign n4563 = pi0038 & n4550;
  assign n4564 = pi0039 & ~n4554;
  assign n4565 = ~pi0869 & n3508;
  assign n4566 = ~pi0170 & ~n4565;
  assign n4567 = ~pi0869 & ~n3499;
  assign n4568 = pi0869 & ~n3416;
  assign n4569 = pi0170 & ~n4567;
  assign n4570 = ~n4568 & n4569;
  assign n4571 = ~n4566 & ~n4570;
  assign n4572 = ~pi0228 & ~n4571;
  assign n4573 = ~n3793 & n4402;
  assign n4574 = ~n4572 & n4573;
  assign n4575 = n4396 & ~n4574;
  assign n4576 = ~n4409 & ~n4575;
  assign n4577 = ~pi0215 & ~n4576;
  assign n4578 = n4469 & ~n4577;
  assign n4579 = n4489 & ~n4578;
  assign n4580 = ~pi0038 & ~n4564;
  assign n4581 = ~n4579 & n4580;
  assign n4582 = ~pi0100 & ~n4563;
  assign n4583 = ~n4581 & n4582;
  assign n4584 = ~n2530 & n4550;
  assign n4585 = ~n4500 & n4528;
  assign n4586 = n4396 & ~n4585;
  assign n4587 = ~n4409 & ~n4586;
  assign n4588 = ~pi0215 & ~n4587;
  assign n4589 = ~n4394 & ~n4588;
  assign n4590 = pi0299 & ~n4589;
  assign n4591 = n2530 & n4548;
  assign n4592 = ~n4590 & n4591;
  assign n4593 = pi0100 & ~n4584;
  assign n4594 = ~n4592 & n4593;
  assign n4595 = ~n4583 & ~n4594;
  assign n4596 = ~pi0087 & ~n4595;
  assign n4597 = ~pi0075 & ~n4562;
  assign n4598 = ~n4596 & n4597;
  assign n4599 = ~pi0092 & ~n4561;
  assign n4600 = ~n4598 & n4599;
  assign n4601 = n2532 & ~n4560;
  assign n4602 = ~n4600 & n4601;
  assign n4603 = ~pi0055 & ~n4551;
  assign n4604 = ~n4602 & n4603;
  assign n4605 = ~pi0056 & ~n4547;
  assign n4606 = ~n4604 & n4605;
  assign n4607 = ~pi0062 & ~n4543;
  assign n4608 = ~n4606 & n4607;
  assign n4609 = pi0248 & n3328;
  assign n4610 = ~n4539 & n4609;
  assign n4611 = ~n4608 & n4610;
  assign n4612 = pi0248 & n4535;
  assign n4613 = ~n3328 & ~n4612;
  assign n4614 = n4412 & n4613;
  assign n4615 = ~n4611 & ~n4614;
  assign po0159 = ~n4527 & n4615;
  assign n4617 = pi0215 & pi1139;
  assign n4618 = pi0216 & ~pi1139;
  assign n4619 = pi0833 & pi0920;
  assign n4620 = ~pi0833 & pi1139;
  assign n4621 = ~pi0216 & ~n4619;
  assign n4622 = ~n4620 & n4621;
  assign n4623 = pi0221 & ~n4622;
  assign n4624 = ~n4618 & n4623;
  assign n4625 = pi0216 & pi0281;
  assign n4626 = ~pi0221 & ~n4625;
  assign n4627 = ~pi0216 & ~pi0862;
  assign n4628 = n3630 & n4627;
  assign n4629 = n4626 & ~n4628;
  assign n4630 = ~n4624 & ~n4629;
  assign n4631 = ~pi0216 & ~n4623;
  assign n4632 = pi0148 & ~n2441;
  assign n4633 = n4631 & n4632;
  assign n4634 = ~pi0215 & ~n4633;
  assign n4635 = ~n4630 & n4634;
  assign n4636 = ~n4617 & ~n4635;
  assign n4637 = ~n3450 & ~n4636;
  assign n4638 = ~n3328 & ~n4637;
  assign n4639 = ~n3331 & ~n4637;
  assign n4640 = ~pi0148 & ~pi0215;
  assign n4641 = pi0862 & ~n3447;
  assign n4642 = ~n2441 & ~n3335;
  assign n4643 = ~pi0216 & ~n4641;
  assign n4644 = ~n4642 & n4643;
  assign n4645 = n4626 & ~n4644;
  assign n4646 = ~n4624 & ~n4645;
  assign n4647 = n4640 & ~n4646;
  assign n4648 = pi0148 & ~pi0215;
  assign n4649 = ~n3335 & ~n3630;
  assign n4650 = n4627 & ~n4649;
  assign n4651 = n4626 & ~n4650;
  assign n4652 = ~n4624 & ~n4651;
  assign n4653 = n4631 & n4649;
  assign n4654 = n4648 & ~n4653;
  assign n4655 = ~n4652 & n4654;
  assign n4656 = ~n4617 & ~n4655;
  assign n4657 = ~n4647 & n4656;
  assign n4658 = n3331 & n4657;
  assign n4659 = pi0062 & ~n4639;
  assign n4660 = ~n4658 & n4659;
  assign n4661 = n2537 & ~n4657;
  assign n4662 = ~n2537 & n4637;
  assign n4663 = pi0056 & ~n4662;
  assign n4664 = ~n4661 & n4663;
  assign n4665 = ~n2572 & ~n4637;
  assign n4666 = n2572 & n4657;
  assign n4667 = pi0055 & ~n4665;
  assign n4668 = ~n4666 & n4667;
  assign n4669 = pi0223 & pi1139;
  assign n4670 = ~pi1139 & ~n2591;
  assign n4671 = ~pi0920 & n2591;
  assign n4672 = pi0222 & ~n4670;
  assign n4673 = ~n4671 & n4672;
  assign n4674 = ~pi0224 & ~n4669;
  assign n4675 = ~n4673 & n4674;
  assign n4676 = n2442 & n4675;
  assign n4677 = ~pi0862 & n4675;
  assign n4678 = pi0224 & pi0281;
  assign n4679 = ~pi0222 & ~n4678;
  assign n4680 = ~n4673 & ~n4679;
  assign n4681 = ~pi0223 & ~n4680;
  assign n4682 = ~n4669 & ~n4681;
  assign n4683 = ~pi0299 & ~n4682;
  assign n4684 = ~n4677 & n4683;
  assign n4685 = ~n4676 & n4684;
  assign n4686 = pi0299 & n4637;
  assign n4687 = ~n4685 & ~n4686;
  assign n4688 = ~n2532 & n4687;
  assign n4689 = ~n2625 & n4687;
  assign n4690 = pi0299 & ~n4657;
  assign n4691 = ~n4685 & ~n4690;
  assign n4692 = n2625 & n4691;
  assign n4693 = ~n4689 & ~n4692;
  assign n4694 = n2533 & ~n4693;
  assign n4695 = ~n2533 & n4687;
  assign n4696 = pi0092 & ~n4695;
  assign n4697 = ~n4694 & n4696;
  assign n4698 = pi0075 & n4687;
  assign n4699 = pi0087 & n4693;
  assign n4700 = ~n2530 & n4687;
  assign n4701 = ~n2441 & ~n3629;
  assign n4702 = n4626 & n4701;
  assign n4703 = n4646 & ~n4702;
  assign n4704 = n4640 & ~n4703;
  assign n4705 = n3631 & n4626;
  assign n4706 = n4652 & ~n4705;
  assign n4707 = n3631 & n4631;
  assign n4708 = n4648 & ~n4707;
  assign n4709 = ~n4706 & n4708;
  assign n4710 = ~n4617 & ~n4704;
  assign n4711 = ~n4709 & n4710;
  assign n4712 = pi0299 & ~n4711;
  assign n4713 = n2530 & ~n4685;
  assign n4714 = ~n4712 & n4713;
  assign n4715 = pi0100 & ~n4700;
  assign n4716 = ~n4714 & n4715;
  assign n4717 = pi0038 & n4687;
  assign n4718 = pi0039 & ~n4691;
  assign n4719 = ~n3488 & n4675;
  assign n4720 = ~n4677 & ~n4682;
  assign n4721 = ~n4719 & n4720;
  assign n4722 = ~pi0299 & ~n4721;
  assign n4723 = ~n3511 & n4627;
  assign n4724 = n4626 & ~n4723;
  assign n4725 = ~n4624 & ~n4724;
  assign n4726 = n3511 & n4631;
  assign n4727 = n4648 & ~n4726;
  assign n4728 = ~n4725 & n4727;
  assign n4729 = pi0862 & ~n3501;
  assign n4730 = ~pi0228 & n3416;
  assign n4731 = ~n2441 & ~n4730;
  assign n4732 = ~pi0862 & n4731;
  assign n4733 = ~pi0216 & ~n4729;
  assign n4734 = ~n4732 & n4733;
  assign n4735 = n4626 & ~n4734;
  assign n4736 = ~n4624 & ~n4735;
  assign n4737 = n4640 & ~n4736;
  assign n4738 = pi0299 & ~n4617;
  assign n4739 = ~n4728 & n4738;
  assign n4740 = ~n4737 & n4739;
  assign n4741 = ~pi0039 & ~n4722;
  assign n4742 = ~n4740 & n4741;
  assign n4743 = ~pi0038 & ~n4718;
  assign n4744 = ~n4742 & n4743;
  assign n4745 = ~pi0100 & ~n4717;
  assign n4746 = ~n4744 & n4745;
  assign n4747 = ~n4716 & ~n4746;
  assign n4748 = ~pi0087 & ~n4747;
  assign n4749 = ~pi0075 & ~n4699;
  assign n4750 = ~n4748 & n4749;
  assign n4751 = ~pi0092 & ~n4698;
  assign n4752 = ~n4750 & n4751;
  assign n4753 = n2532 & ~n4697;
  assign n4754 = ~n4752 & n4753;
  assign n4755 = ~pi0055 & ~n4688;
  assign n4756 = ~n4754 & n4755;
  assign n4757 = ~pi0056 & ~n4668;
  assign n4758 = ~n4756 & n4757;
  assign n4759 = ~pi0062 & ~n4664;
  assign n4760 = ~n4758 & n4759;
  assign n4761 = n3328 & ~n4660;
  assign n4762 = ~n4760 & n4761;
  assign n4763 = ~pi0247 & ~n4638;
  assign n4764 = ~n4762 & n4763;
  assign n4765 = ~n3328 & n4636;
  assign n4766 = ~n3331 & n4636;
  assign n4767 = n4634 & ~n4652;
  assign n4768 = n4656 & ~n4767;
  assign n4769 = n3331 & n4768;
  assign n4770 = pi0062 & ~n4766;
  assign n4771 = ~n4769 & n4770;
  assign n4772 = ~n2537 & ~n4636;
  assign n4773 = n2537 & ~n4768;
  assign n4774 = pi0056 & ~n4772;
  assign n4775 = ~n4773 & n4774;
  assign n4776 = ~n2572 & n4636;
  assign n4777 = n2572 & n4768;
  assign n4778 = pi0055 & ~n4776;
  assign n4779 = ~n4777 & n4778;
  assign n4780 = ~n3472 & ~n4684;
  assign n4781 = pi0299 & ~n4636;
  assign n4782 = n4780 & ~n4781;
  assign n4783 = ~n2532 & n4782;
  assign n4784 = ~n2625 & n4782;
  assign n4785 = pi0299 & ~n4768;
  assign n4786 = n4780 & ~n4785;
  assign n4787 = n2625 & n4786;
  assign n4788 = ~n4784 & ~n4787;
  assign n4789 = n2533 & ~n4788;
  assign n4790 = ~n2533 & n4782;
  assign n4791 = pi0092 & ~n4790;
  assign n4792 = ~n4789 & n4791;
  assign n4793 = pi0075 & n4782;
  assign n4794 = pi0087 & n4788;
  assign n4795 = ~n2530 & n4782;
  assign n4796 = n4640 & ~n4706;
  assign n4797 = ~pi0216 & ~n4624;
  assign n4798 = n4701 & n4797;
  assign n4799 = n4648 & ~n4652;
  assign n4800 = ~n4798 & n4799;
  assign n4801 = ~n4617 & ~n4800;
  assign n4802 = ~n4796 & n4801;
  assign n4803 = pi0299 & ~n4802;
  assign n4804 = n2530 & n4780;
  assign n4805 = ~n4803 & n4804;
  assign n4806 = pi0100 & ~n4795;
  assign n4807 = ~n4805 & n4806;
  assign n4808 = pi0038 & n4782;
  assign n4809 = pi0039 & ~n4786;
  assign n4810 = n3488 & n4677;
  assign n4811 = n4683 & ~n4810;
  assign n4812 = pi0862 & ~n4731;
  assign n4813 = ~pi0862 & n3501;
  assign n4814 = ~pi0216 & ~n4813;
  assign n4815 = ~n4812 & n4814;
  assign n4816 = n4626 & ~n4815;
  assign n4817 = ~n4624 & ~n4816;
  assign n4818 = n4648 & ~n4817;
  assign n4819 = n4640 & ~n4725;
  assign n4820 = ~n4617 & ~n4819;
  assign n4821 = ~n4818 & n4820;
  assign n4822 = pi0299 & ~n4821;
  assign n4823 = ~n4811 & ~n4822;
  assign n4824 = ~pi0039 & ~n4823;
  assign n4825 = ~pi0038 & ~n4809;
  assign n4826 = ~n4824 & n4825;
  assign n4827 = ~pi0100 & ~n4808;
  assign n4828 = ~n4826 & n4827;
  assign n4829 = ~n4807 & ~n4828;
  assign n4830 = ~pi0087 & ~n4829;
  assign n4831 = ~pi0075 & ~n4794;
  assign n4832 = ~n4830 & n4831;
  assign n4833 = ~pi0092 & ~n4793;
  assign n4834 = ~n4832 & n4833;
  assign n4835 = n2532 & ~n4792;
  assign n4836 = ~n4834 & n4835;
  assign n4837 = ~pi0055 & ~n4783;
  assign n4838 = ~n4836 & n4837;
  assign n4839 = ~pi0056 & ~n4779;
  assign n4840 = ~n4838 & n4839;
  assign n4841 = ~pi0062 & ~n4775;
  assign n4842 = ~n4840 & n4841;
  assign n4843 = n3328 & ~n4771;
  assign n4844 = ~n4842 & n4843;
  assign n4845 = pi0247 & ~n4765;
  assign n4846 = ~n4844 & n4845;
  assign po0160 = n4764 | n4846;
  assign n4848 = pi0215 & pi1138;
  assign n4849 = pi0216 & pi0269;
  assign n4850 = ~pi0221 & ~n4849;
  assign n4851 = ~pi0105 & pi0169;
  assign n4852 = pi0877 & ~n2442;
  assign n4853 = pi0105 & ~n4852;
  assign n4854 = pi0228 & ~n4851;
  assign n4855 = ~n4853 & n4854;
  assign n4856 = ~pi0216 & ~n4855;
  assign n4857 = ~pi0169 & ~pi0228;
  assign n4858 = n4856 & ~n4857;
  assign n4859 = n4850 & ~n4858;
  assign n4860 = ~pi1138 & ~n2452;
  assign n4861 = ~pi0940 & n2452;
  assign n4862 = pi0221 & ~n4860;
  assign n4863 = ~n4861 & n4862;
  assign n4864 = ~n4859 & ~n4863;
  assign n4865 = ~pi0215 & ~n4864;
  assign n4866 = ~n4848 & ~n4865;
  assign n4867 = ~n3331 & n4866;
  assign n4868 = ~pi0877 & n2521;
  assign n4869 = pi0169 & ~n2521;
  assign n4870 = ~pi0228 & ~n4868;
  assign n4871 = ~n4869 & n4870;
  assign n4872 = n4856 & ~n4871;
  assign n4873 = n4850 & ~n4872;
  assign n4874 = ~n4863 & ~n4873;
  assign n4875 = ~pi0215 & ~n4874;
  assign n4876 = ~n4848 & ~n4875;
  assign n4877 = n3331 & n4876;
  assign n4878 = pi0062 & ~n4867;
  assign n4879 = ~n4877 & n4878;
  assign n4880 = ~n2537 & ~n4866;
  assign n4881 = n2537 & ~n4876;
  assign n4882 = pi0056 & ~n4880;
  assign n4883 = ~n4881 & n4882;
  assign n4884 = ~n2572 & n4866;
  assign n4885 = n2572 & n4876;
  assign n4886 = pi0055 & ~n4884;
  assign n4887 = ~n4885 & n4886;
  assign n4888 = pi0223 & pi1138;
  assign n4889 = pi0224 & pi0269;
  assign n4890 = ~pi0222 & ~n4889;
  assign n4891 = ~pi0224 & ~n4852;
  assign n4892 = n4890 & ~n4891;
  assign n4893 = ~pi1138 & ~n2591;
  assign n4894 = ~pi0940 & n2591;
  assign n4895 = pi0222 & ~n4893;
  assign n4896 = ~n4894 & n4895;
  assign n4897 = ~n4892 & ~n4896;
  assign n4898 = ~pi0223 & ~n4897;
  assign n4899 = ~n4888 & ~n4898;
  assign n4900 = ~pi0299 & ~n4899;
  assign n4901 = pi0299 & ~n4866;
  assign n4902 = ~n4900 & ~n4901;
  assign n4903 = ~n2532 & n4902;
  assign n4904 = ~n2625 & n4902;
  assign n4905 = pi0299 & ~n4876;
  assign n4906 = ~n4900 & ~n4905;
  assign n4907 = n2625 & n4906;
  assign n4908 = ~n4904 & ~n4907;
  assign n4909 = n2533 & ~n4908;
  assign n4910 = ~n2533 & n4902;
  assign n4911 = pi0092 & ~n4910;
  assign n4912 = ~n4909 & n4911;
  assign n4913 = pi0075 & n4902;
  assign n4914 = pi0087 & n4908;
  assign n4915 = pi0038 & n4902;
  assign n4916 = pi0039 & ~n4906;
  assign n4917 = ~pi0299 & ~n4888;
  assign n4918 = pi0877 & n3488;
  assign n4919 = ~pi0224 & ~n4918;
  assign n4920 = n4890 & ~n4919;
  assign n4921 = ~n4896 & ~n4920;
  assign n4922 = n4917 & n4921;
  assign n4923 = pi0299 & ~n4848;
  assign n4924 = pi0877 & n3499;
  assign n4925 = ~pi0169 & ~n4924;
  assign n4926 = pi0169 & n3508;
  assign n4927 = ~n4925 & ~n4926;
  assign n4928 = pi0877 & ~n4927;
  assign n4929 = ~n3416 & n4925;
  assign n4930 = ~n4928 & ~n4929;
  assign n4931 = ~pi0228 & ~n4930;
  assign n4932 = ~n3497 & n4855;
  assign n4933 = ~pi0216 & ~n4932;
  assign n4934 = ~n4931 & n4933;
  assign n4935 = n4850 & ~n4934;
  assign n4936 = ~n4863 & ~n4935;
  assign n4937 = ~pi0215 & ~n4936;
  assign n4938 = n4923 & ~n4937;
  assign n4939 = ~n3488 & n4890;
  assign n4940 = n4921 & ~n4939;
  assign n4941 = ~pi0223 & ~n4940;
  assign n4942 = n4917 & ~n4941;
  assign n4943 = ~pi0039 & ~n4942;
  assign n4944 = ~n4922 & n4943;
  assign n4945 = ~n4938 & n4944;
  assign n4946 = ~pi0038 & ~n4916;
  assign n4947 = ~n4945 & n4946;
  assign n4948 = ~pi0100 & ~n4915;
  assign n4949 = ~n4947 & n4948;
  assign n4950 = ~n2530 & n4902;
  assign n4951 = ~pi0877 & n3394;
  assign n4952 = pi0169 & ~n3394;
  assign n4953 = ~pi0228 & ~n4951;
  assign n4954 = ~n4952 & n4953;
  assign n4955 = n4856 & ~n4954;
  assign n4956 = n4850 & ~n4955;
  assign n4957 = ~n4863 & ~n4956;
  assign n4958 = ~pi0215 & ~n4957;
  assign n4959 = ~n4848 & ~n4958;
  assign n4960 = pi0299 & ~n4959;
  assign n4961 = n2530 & ~n4900;
  assign n4962 = ~n4960 & n4961;
  assign n4963 = pi0100 & ~n4950;
  assign n4964 = ~n4962 & n4963;
  assign n4965 = ~n4949 & ~n4964;
  assign n4966 = ~pi0087 & ~n4965;
  assign n4967 = ~pi0075 & ~n4914;
  assign n4968 = ~n4966 & n4967;
  assign n4969 = ~pi0092 & ~n4913;
  assign n4970 = ~n4968 & n4969;
  assign n4971 = n2532 & ~n4912;
  assign n4972 = ~n4970 & n4971;
  assign n4973 = ~pi0055 & ~n4903;
  assign n4974 = ~n4972 & n4973;
  assign n4975 = ~pi0056 & ~n4887;
  assign n4976 = ~n4974 & n4975;
  assign n4977 = ~pi0062 & ~n4883;
  assign n4978 = ~n4976 & n4977;
  assign n4979 = ~pi0246 & n3328;
  assign n4980 = ~n4879 & n4979;
  assign n4981 = ~n4978 & n4980;
  assign n4982 = ~n3447 & n4856;
  assign n4983 = ~n4871 & n4982;
  assign n4984 = n4850 & ~n4983;
  assign n4985 = ~n4863 & ~n4984;
  assign n4986 = ~pi0215 & ~n4985;
  assign n4987 = ~n4848 & ~n4986;
  assign n4988 = n3331 & n4987;
  assign n4989 = n3556 & ~n4849;
  assign n4990 = n4866 & ~n4989;
  assign n4991 = ~n3331 & n4990;
  assign n4992 = pi0062 & ~n4991;
  assign n4993 = ~n4988 & n4992;
  assign n4994 = ~n2537 & ~n4990;
  assign n4995 = n2537 & ~n4987;
  assign n4996 = pi0056 & ~n4994;
  assign n4997 = ~n4995 & n4996;
  assign n4998 = n2572 & n4987;
  assign n4999 = ~n2572 & n4990;
  assign n5000 = pi0055 & ~n4999;
  assign n5001 = ~n4998 & n5000;
  assign n5002 = ~n3472 & ~n4900;
  assign n5003 = pi0299 & ~n4990;
  assign n5004 = n5002 & ~n5003;
  assign n5005 = ~n2532 & n5004;
  assign n5006 = ~n2625 & n5004;
  assign n5007 = pi0299 & ~n4987;
  assign n5008 = n5002 & ~n5007;
  assign n5009 = n2625 & n5008;
  assign n5010 = ~n5006 & ~n5009;
  assign n5011 = n2533 & ~n5010;
  assign n5012 = ~n2533 & n5004;
  assign n5013 = pi0092 & ~n5012;
  assign n5014 = ~n5011 & n5013;
  assign n5015 = pi0075 & n5004;
  assign n5016 = pi0087 & n5010;
  assign n5017 = pi0038 & n5004;
  assign n5018 = pi0039 & ~n5008;
  assign n5019 = ~pi0877 & n3508;
  assign n5020 = ~pi0169 & ~n5019;
  assign n5021 = ~pi0877 & ~n3499;
  assign n5022 = pi0877 & ~n3416;
  assign n5023 = pi0169 & ~n5021;
  assign n5024 = ~n5022 & n5023;
  assign n5025 = ~n5020 & ~n5024;
  assign n5026 = ~pi0228 & ~n5025;
  assign n5027 = ~n3793 & n4856;
  assign n5028 = ~n5026 & n5027;
  assign n5029 = n4850 & ~n5028;
  assign n5030 = ~n4863 & ~n5029;
  assign n5031 = ~pi0215 & ~n5030;
  assign n5032 = n4923 & ~n5031;
  assign n5033 = n4943 & ~n5032;
  assign n5034 = ~pi0038 & ~n5018;
  assign n5035 = ~n5033 & n5034;
  assign n5036 = ~pi0100 & ~n5017;
  assign n5037 = ~n5035 & n5036;
  assign n5038 = ~n2530 & n5004;
  assign n5039 = ~n4954 & n4982;
  assign n5040 = n4850 & ~n5039;
  assign n5041 = ~n4863 & ~n5040;
  assign n5042 = ~pi0215 & ~n5041;
  assign n5043 = ~n4848 & ~n5042;
  assign n5044 = pi0299 & ~n5043;
  assign n5045 = n2530 & n5002;
  assign n5046 = ~n5044 & n5045;
  assign n5047 = pi0100 & ~n5038;
  assign n5048 = ~n5046 & n5047;
  assign n5049 = ~n5037 & ~n5048;
  assign n5050 = ~pi0087 & ~n5049;
  assign n5051 = ~pi0075 & ~n5016;
  assign n5052 = ~n5050 & n5051;
  assign n5053 = ~pi0092 & ~n5015;
  assign n5054 = ~n5052 & n5053;
  assign n5055 = n2532 & ~n5014;
  assign n5056 = ~n5054 & n5055;
  assign n5057 = ~pi0055 & ~n5005;
  assign n5058 = ~n5056 & n5057;
  assign n5059 = ~pi0056 & ~n5001;
  assign n5060 = ~n5058 & n5059;
  assign n5061 = ~pi0062 & ~n4997;
  assign n5062 = ~n5060 & n5061;
  assign n5063 = pi0246 & n3328;
  assign n5064 = ~n4993 & n5063;
  assign n5065 = ~n5062 & n5064;
  assign n5066 = pi0246 & n4989;
  assign n5067 = ~n3328 & ~n5066;
  assign n5068 = n4866 & n5067;
  assign n5069 = ~n5065 & ~n5068;
  assign po0161 = ~n4981 & n5069;
  assign n5071 = pi0215 & pi1137;
  assign n5072 = pi0216 & pi0280;
  assign n5073 = ~pi0221 & ~n5072;
  assign n5074 = ~pi0105 & pi0168;
  assign n5075 = pi0878 & ~n2442;
  assign n5076 = pi0105 & ~n5075;
  assign n5077 = pi0228 & ~n5074;
  assign n5078 = ~n5076 & n5077;
  assign n5079 = ~pi0216 & ~n5078;
  assign n5080 = ~pi0168 & ~pi0228;
  assign n5081 = n5079 & ~n5080;
  assign n5082 = n5073 & ~n5081;
  assign n5083 = ~pi1137 & ~n2452;
  assign n5084 = ~pi0933 & n2452;
  assign n5085 = pi0221 & ~n5083;
  assign n5086 = ~n5084 & n5085;
  assign n5087 = ~n5082 & ~n5086;
  assign n5088 = ~pi0215 & ~n5087;
  assign n5089 = ~n5071 & ~n5088;
  assign n5090 = ~n3331 & n5089;
  assign n5091 = ~pi0878 & n2521;
  assign n5092 = pi0168 & ~n2521;
  assign n5093 = ~pi0228 & ~n5091;
  assign n5094 = ~n5092 & n5093;
  assign n5095 = n5079 & ~n5094;
  assign n5096 = n5073 & ~n5095;
  assign n5097 = ~n5086 & ~n5096;
  assign n5098 = ~pi0215 & ~n5097;
  assign n5099 = ~n5071 & ~n5098;
  assign n5100 = n3331 & n5099;
  assign n5101 = pi0062 & ~n5090;
  assign n5102 = ~n5100 & n5101;
  assign n5103 = ~n2537 & ~n5089;
  assign n5104 = n2537 & ~n5099;
  assign n5105 = pi0056 & ~n5103;
  assign n5106 = ~n5104 & n5105;
  assign n5107 = ~n2572 & n5089;
  assign n5108 = n2572 & n5099;
  assign n5109 = pi0055 & ~n5107;
  assign n5110 = ~n5108 & n5109;
  assign n5111 = pi0223 & pi1137;
  assign n5112 = pi0224 & pi0280;
  assign n5113 = ~pi0222 & ~n5112;
  assign n5114 = ~pi0224 & ~n5075;
  assign n5115 = n5113 & ~n5114;
  assign n5116 = ~pi1137 & ~n2591;
  assign n5117 = ~pi0933 & n2591;
  assign n5118 = pi0222 & ~n5116;
  assign n5119 = ~n5117 & n5118;
  assign n5120 = ~n5115 & ~n5119;
  assign n5121 = ~pi0223 & ~n5120;
  assign n5122 = ~n5111 & ~n5121;
  assign n5123 = ~pi0299 & ~n5122;
  assign n5124 = pi0299 & ~n5089;
  assign n5125 = ~n5123 & ~n5124;
  assign n5126 = ~n2532 & n5125;
  assign n5127 = ~n2625 & n5125;
  assign n5128 = pi0299 & ~n5099;
  assign n5129 = ~n5123 & ~n5128;
  assign n5130 = n2625 & n5129;
  assign n5131 = ~n5127 & ~n5130;
  assign n5132 = n2533 & ~n5131;
  assign n5133 = ~n2533 & n5125;
  assign n5134 = pi0092 & ~n5133;
  assign n5135 = ~n5132 & n5134;
  assign n5136 = pi0075 & n5125;
  assign n5137 = pi0087 & n5131;
  assign n5138 = pi0038 & n5125;
  assign n5139 = pi0039 & ~n5129;
  assign n5140 = ~pi0299 & ~n5111;
  assign n5141 = pi0878 & n3488;
  assign n5142 = ~pi0224 & ~n5141;
  assign n5143 = n5113 & ~n5142;
  assign n5144 = ~n5119 & ~n5143;
  assign n5145 = n5140 & n5144;
  assign n5146 = pi0299 & ~n5071;
  assign n5147 = pi0878 & n3499;
  assign n5148 = ~pi0168 & ~n5147;
  assign n5149 = pi0168 & n3508;
  assign n5150 = ~n5148 & ~n5149;
  assign n5151 = pi0878 & ~n5150;
  assign n5152 = ~n3416 & n5148;
  assign n5153 = ~n5151 & ~n5152;
  assign n5154 = ~pi0228 & ~n5153;
  assign n5155 = ~n3497 & n5078;
  assign n5156 = ~pi0216 & ~n5155;
  assign n5157 = ~n5154 & n5156;
  assign n5158 = n5073 & ~n5157;
  assign n5159 = ~n5086 & ~n5158;
  assign n5160 = ~pi0215 & ~n5159;
  assign n5161 = n5146 & ~n5160;
  assign n5162 = ~n3488 & n5113;
  assign n5163 = n5144 & ~n5162;
  assign n5164 = ~pi0223 & ~n5163;
  assign n5165 = n5140 & ~n5164;
  assign n5166 = ~pi0039 & ~n5165;
  assign n5167 = ~n5145 & n5166;
  assign n5168 = ~n5161 & n5167;
  assign n5169 = ~pi0038 & ~n5139;
  assign n5170 = ~n5168 & n5169;
  assign n5171 = ~pi0100 & ~n5138;
  assign n5172 = ~n5170 & n5171;
  assign n5173 = ~n2530 & n5125;
  assign n5174 = ~pi0878 & n3394;
  assign n5175 = pi0168 & ~n3394;
  assign n5176 = ~pi0228 & ~n5174;
  assign n5177 = ~n5175 & n5176;
  assign n5178 = n5079 & ~n5177;
  assign n5179 = n5073 & ~n5178;
  assign n5180 = ~n5086 & ~n5179;
  assign n5181 = ~pi0215 & ~n5180;
  assign n5182 = ~n5071 & ~n5181;
  assign n5183 = pi0299 & ~n5182;
  assign n5184 = n2530 & ~n5123;
  assign n5185 = ~n5183 & n5184;
  assign n5186 = pi0100 & ~n5173;
  assign n5187 = ~n5185 & n5186;
  assign n5188 = ~n5172 & ~n5187;
  assign n5189 = ~pi0087 & ~n5188;
  assign n5190 = ~pi0075 & ~n5137;
  assign n5191 = ~n5189 & n5190;
  assign n5192 = ~pi0092 & ~n5136;
  assign n5193 = ~n5191 & n5192;
  assign n5194 = n2532 & ~n5135;
  assign n5195 = ~n5193 & n5194;
  assign n5196 = ~pi0055 & ~n5126;
  assign n5197 = ~n5195 & n5196;
  assign n5198 = ~pi0056 & ~n5110;
  assign n5199 = ~n5197 & n5198;
  assign n5200 = ~pi0062 & ~n5106;
  assign n5201 = ~n5199 & n5200;
  assign n5202 = ~pi0240 & n3328;
  assign n5203 = ~n5102 & n5202;
  assign n5204 = ~n5201 & n5203;
  assign n5205 = ~n3447 & n5079;
  assign n5206 = ~n5094 & n5205;
  assign n5207 = n5073 & ~n5206;
  assign n5208 = ~n5086 & ~n5207;
  assign n5209 = ~pi0215 & ~n5208;
  assign n5210 = ~n5071 & ~n5209;
  assign n5211 = n3331 & n5210;
  assign n5212 = n3556 & ~n5072;
  assign n5213 = n5089 & ~n5212;
  assign n5214 = ~n3331 & n5213;
  assign n5215 = pi0062 & ~n5214;
  assign n5216 = ~n5211 & n5215;
  assign n5217 = ~n2537 & ~n5213;
  assign n5218 = n2537 & ~n5210;
  assign n5219 = pi0056 & ~n5217;
  assign n5220 = ~n5218 & n5219;
  assign n5221 = n2572 & n5210;
  assign n5222 = ~n2572 & n5213;
  assign n5223 = pi0055 & ~n5222;
  assign n5224 = ~n5221 & n5223;
  assign n5225 = ~n3472 & ~n5123;
  assign n5226 = pi0299 & ~n5213;
  assign n5227 = n5225 & ~n5226;
  assign n5228 = ~n2532 & n5227;
  assign n5229 = ~n2625 & n5227;
  assign n5230 = pi0299 & ~n5210;
  assign n5231 = n5225 & ~n5230;
  assign n5232 = n2625 & n5231;
  assign n5233 = ~n5229 & ~n5232;
  assign n5234 = n2533 & ~n5233;
  assign n5235 = ~n2533 & n5227;
  assign n5236 = pi0092 & ~n5235;
  assign n5237 = ~n5234 & n5236;
  assign n5238 = pi0075 & n5227;
  assign n5239 = pi0087 & n5233;
  assign n5240 = pi0038 & n5227;
  assign n5241 = pi0039 & ~n5231;
  assign n5242 = ~pi0878 & n3508;
  assign n5243 = ~pi0168 & ~n5242;
  assign n5244 = ~pi0878 & ~n3499;
  assign n5245 = pi0878 & ~n3416;
  assign n5246 = pi0168 & ~n5244;
  assign n5247 = ~n5245 & n5246;
  assign n5248 = ~n5243 & ~n5247;
  assign n5249 = ~pi0228 & ~n5248;
  assign n5250 = ~n3793 & n5079;
  assign n5251 = ~n5249 & n5250;
  assign n5252 = n5073 & ~n5251;
  assign n5253 = ~n5086 & ~n5252;
  assign n5254 = ~pi0215 & ~n5253;
  assign n5255 = n5146 & ~n5254;
  assign n5256 = n5166 & ~n5255;
  assign n5257 = ~pi0038 & ~n5241;
  assign n5258 = ~n5256 & n5257;
  assign n5259 = ~pi0100 & ~n5240;
  assign n5260 = ~n5258 & n5259;
  assign n5261 = ~n2530 & n5227;
  assign n5262 = ~n5177 & n5205;
  assign n5263 = n5073 & ~n5262;
  assign n5264 = ~n5086 & ~n5263;
  assign n5265 = ~pi0215 & ~n5264;
  assign n5266 = ~n5071 & ~n5265;
  assign n5267 = pi0299 & ~n5266;
  assign n5268 = n2530 & n5225;
  assign n5269 = ~n5267 & n5268;
  assign n5270 = pi0100 & ~n5261;
  assign n5271 = ~n5269 & n5270;
  assign n5272 = ~n5260 & ~n5271;
  assign n5273 = ~pi0087 & ~n5272;
  assign n5274 = ~pi0075 & ~n5239;
  assign n5275 = ~n5273 & n5274;
  assign n5276 = ~pi0092 & ~n5238;
  assign n5277 = ~n5275 & n5276;
  assign n5278 = n2532 & ~n5237;
  assign n5279 = ~n5277 & n5278;
  assign n5280 = ~pi0055 & ~n5228;
  assign n5281 = ~n5279 & n5280;
  assign n5282 = ~pi0056 & ~n5224;
  assign n5283 = ~n5281 & n5282;
  assign n5284 = ~pi0062 & ~n5220;
  assign n5285 = ~n5283 & n5284;
  assign n5286 = pi0240 & n3328;
  assign n5287 = ~n5216 & n5286;
  assign n5288 = ~n5285 & n5287;
  assign n5289 = pi0240 & n5212;
  assign n5290 = ~n3328 & ~n5289;
  assign n5291 = n5089 & n5290;
  assign n5292 = ~n5288 & ~n5291;
  assign po0162 = ~n5204 & n5292;
  assign n5294 = pi0215 & pi1136;
  assign n5295 = pi0216 & pi0266;
  assign n5296 = pi0875 & ~n2442;
  assign n5297 = pi0105 & ~n5296;
  assign n5298 = ~pi0105 & ~pi0166;
  assign n5299 = ~n5297 & ~n5298;
  assign n5300 = pi0228 & n5299;
  assign n5301 = pi0166 & ~pi0228;
  assign n5302 = ~n5300 & ~n5301;
  assign n5303 = ~pi0216 & ~n5302;
  assign n5304 = ~n5295 & ~n5303;
  assign n5305 = ~pi0221 & ~n5304;
  assign n5306 = ~pi1136 & ~n2452;
  assign n5307 = ~pi0928 & n2452;
  assign n5308 = pi0221 & ~n5306;
  assign n5309 = ~n5307 & n5308;
  assign n5310 = ~n5305 & ~n5309;
  assign n5311 = ~pi0215 & ~n5310;
  assign n5312 = ~n5294 & ~n5311;
  assign n5313 = ~n3328 & n5312;
  assign n5314 = ~n3331 & n5312;
  assign n5315 = ~pi0166 & ~n2521;
  assign n5316 = ~pi0875 & n2521;
  assign n5317 = ~pi0228 & ~n5315;
  assign n5318 = ~n5316 & n5317;
  assign n5319 = ~n5300 & ~n5318;
  assign n5320 = ~pi0216 & ~n5319;
  assign n5321 = ~n5295 & ~n5320;
  assign n5322 = ~pi0221 & ~n5321;
  assign n5323 = ~n5309 & ~n5322;
  assign n5324 = ~pi0215 & ~n5323;
  assign n5325 = ~n5294 & ~n5324;
  assign n5326 = n3331 & n5325;
  assign n5327 = pi0062 & ~n5314;
  assign n5328 = ~n5326 & n5327;
  assign n5329 = ~n2537 & ~n5312;
  assign n5330 = n2537 & ~n5325;
  assign n5331 = pi0056 & ~n5329;
  assign n5332 = ~n5330 & n5331;
  assign n5333 = ~n2572 & n5312;
  assign n5334 = n2572 & n5325;
  assign n5335 = pi0055 & ~n5333;
  assign n5336 = ~n5334 & n5335;
  assign n5337 = pi0223 & pi1136;
  assign n5338 = pi0224 & ~pi0266;
  assign n5339 = ~pi0224 & ~pi0875;
  assign n5340 = ~n2442 & n5339;
  assign n5341 = ~pi0222 & ~n5338;
  assign n5342 = ~n5340 & n5341;
  assign n5343 = ~pi1136 & ~n2591;
  assign n5344 = ~pi0928 & n2591;
  assign n5345 = pi0222 & ~n5343;
  assign n5346 = ~n5344 & n5345;
  assign n5347 = ~n5342 & ~n5346;
  assign n5348 = ~pi0223 & ~n5347;
  assign n5349 = ~n5337 & ~n5348;
  assign n5350 = ~pi0299 & ~n5349;
  assign n5351 = n2604 & ~n5296;
  assign n5352 = n5350 & ~n5351;
  assign n5353 = pi0299 & ~n5312;
  assign n5354 = ~n5352 & ~n5353;
  assign n5355 = ~n2532 & n5354;
  assign n5356 = ~n2625 & n5354;
  assign n5357 = pi0299 & ~n5325;
  assign n5358 = ~n5352 & ~n5357;
  assign n5359 = n2625 & n5358;
  assign n5360 = ~n5356 & ~n5359;
  assign n5361 = n2533 & ~n5360;
  assign n5362 = ~n2533 & n5354;
  assign n5363 = pi0092 & ~n5362;
  assign n5364 = ~n5361 & n5363;
  assign n5365 = pi0075 & n5354;
  assign n5366 = pi0087 & n5360;
  assign n5367 = pi0038 & n5354;
  assign n5368 = pi0039 & ~n5358;
  assign n5369 = n2603 & ~n3488;
  assign n5370 = n5342 & ~n5369;
  assign n5371 = ~pi0299 & ~n5337;
  assign n5372 = ~n5346 & n5371;
  assign n5373 = ~n5370 & n5372;
  assign n5374 = n3498 & ~n5299;
  assign n5375 = ~pi0216 & ~n5374;
  assign n5376 = pi0166 & n3499;
  assign n5377 = ~pi0166 & ~n3508;
  assign n5378 = pi0875 & ~n5376;
  assign n5379 = ~n5377 & n5378;
  assign n5380 = pi0166 & ~pi0875;
  assign n5381 = ~n3416 & n5380;
  assign n5382 = ~n5379 & ~n5381;
  assign n5383 = ~pi0228 & ~n5382;
  assign n5384 = ~n3498 & ~n5383;
  assign n5385 = n5375 & ~n5384;
  assign n5386 = ~n5295 & ~n5385;
  assign n5387 = ~pi0221 & ~n5386;
  assign n5388 = ~n5309 & ~n5387;
  assign n5389 = ~pi0215 & ~n5388;
  assign n5390 = pi0299 & ~n5294;
  assign n5391 = ~n5389 & n5390;
  assign n5392 = n5347 & ~n5369;
  assign n5393 = ~pi0223 & ~n5392;
  assign n5394 = n5371 & ~n5393;
  assign n5395 = ~pi0039 & ~n5394;
  assign n5396 = ~n5373 & n5395;
  assign n5397 = ~n5391 & n5396;
  assign n5398 = ~pi0038 & ~n5368;
  assign n5399 = ~n5397 & n5398;
  assign n5400 = ~pi0100 & ~n5367;
  assign n5401 = ~n5399 & n5400;
  assign n5402 = ~n2530 & n5354;
  assign n5403 = ~pi0875 & n3387;
  assign n5404 = pi0166 & ~n5403;
  assign n5405 = ~n2638 & ~n3387;
  assign n5406 = n2638 & ~n3385;
  assign n5407 = pi0875 & ~n5406;
  assign n5408 = ~n5405 & n5407;
  assign n5409 = ~n5404 & ~n5408;
  assign n5410 = ~pi0228 & ~n5409;
  assign n5411 = ~n5300 & ~n5410;
  assign n5412 = ~pi0216 & ~n5411;
  assign n5413 = ~n5295 & ~n5412;
  assign n5414 = ~pi0221 & ~n5413;
  assign n5415 = ~n5309 & ~n5414;
  assign n5416 = ~pi0215 & ~n5415;
  assign n5417 = ~n5294 & ~n5416;
  assign n5418 = pi0299 & ~n5417;
  assign n5419 = n2530 & ~n5352;
  assign n5420 = ~n5418 & n5419;
  assign n5421 = pi0100 & ~n5402;
  assign n5422 = ~n5420 & n5421;
  assign n5423 = ~n5401 & ~n5422;
  assign n5424 = ~pi0087 & ~n5423;
  assign n5425 = ~pi0075 & ~n5366;
  assign n5426 = ~n5424 & n5425;
  assign n5427 = ~pi0092 & ~n5365;
  assign n5428 = ~n5426 & n5427;
  assign n5429 = n2532 & ~n5364;
  assign n5430 = ~n5428 & n5429;
  assign n5431 = ~pi0055 & ~n5355;
  assign n5432 = ~n5430 & n5431;
  assign n5433 = ~pi0056 & ~n5336;
  assign n5434 = ~n5432 & n5433;
  assign n5435 = ~pi0062 & ~n5332;
  assign n5436 = ~n5434 & n5435;
  assign n5437 = n3328 & ~n5328;
  assign n5438 = ~n5436 & n5437;
  assign n5439 = ~pi0245 & ~n5313;
  assign n5440 = ~n5438 & n5439;
  assign n5441 = ~n3450 & n5312;
  assign n5442 = ~n3328 & n5441;
  assign n5443 = ~n3447 & ~n5300;
  assign n5444 = ~n5318 & n5443;
  assign n5445 = ~pi0216 & ~n5444;
  assign n5446 = ~n5295 & ~n5445;
  assign n5447 = ~pi0221 & ~n5446;
  assign n5448 = ~n5309 & ~n5447;
  assign n5449 = ~pi0215 & ~n5448;
  assign n5450 = ~n5294 & ~n5449;
  assign n5451 = n3331 & n5450;
  assign n5452 = ~n3331 & n5441;
  assign n5453 = pi0062 & ~n5452;
  assign n5454 = ~n5451 & n5453;
  assign n5455 = ~n2537 & ~n5441;
  assign n5456 = n2537 & ~n5450;
  assign n5457 = pi0056 & ~n5455;
  assign n5458 = ~n5456 & n5457;
  assign n5459 = n2572 & n5450;
  assign n5460 = ~n2572 & n5441;
  assign n5461 = pi0055 & ~n5460;
  assign n5462 = ~n5459 & n5461;
  assign n5463 = pi0299 & ~n5441;
  assign n5464 = ~n5350 & ~n5463;
  assign n5465 = ~n2532 & n5464;
  assign n5466 = ~n2625 & n5464;
  assign n5467 = pi0299 & ~n5450;
  assign n5468 = ~n5350 & ~n5467;
  assign n5469 = n2625 & n5468;
  assign n5470 = ~n5466 & ~n5469;
  assign n5471 = n2533 & ~n5470;
  assign n5472 = ~n2533 & n5464;
  assign n5473 = pi0092 & ~n5472;
  assign n5474 = ~n5471 & n5473;
  assign n5475 = pi0075 & n5464;
  assign n5476 = pi0087 & n5470;
  assign n5477 = pi0038 & n5464;
  assign n5478 = pi0039 & ~n5468;
  assign n5479 = ~pi0166 & ~n3499;
  assign n5480 = pi0166 & n3508;
  assign n5481 = ~pi0875 & ~n5479;
  assign n5482 = ~n5480 & n5481;
  assign n5483 = ~pi0166 & ~n3416;
  assign n5484 = pi0875 & ~n5483;
  assign n5485 = ~pi0228 & ~n5482;
  assign n5486 = ~n5484 & n5485;
  assign n5487 = n5375 & ~n5486;
  assign n5488 = ~n5295 & ~n5487;
  assign n5489 = ~pi0221 & ~n5488;
  assign n5490 = ~n5309 & ~n5489;
  assign n5491 = ~pi0215 & ~n5490;
  assign n5492 = n5390 & ~n5491;
  assign n5493 = n5395 & ~n5492;
  assign n5494 = ~pi0038 & ~n5478;
  assign n5495 = ~n5493 & n5494;
  assign n5496 = ~pi0100 & ~n5477;
  assign n5497 = ~n5495 & n5496;
  assign n5498 = ~n2530 & n5464;
  assign n5499 = ~n5410 & n5443;
  assign n5500 = ~pi0216 & ~n5499;
  assign n5501 = ~n5295 & ~n5500;
  assign n5502 = ~pi0221 & ~n5501;
  assign n5503 = ~n5309 & ~n5502;
  assign n5504 = ~pi0215 & ~n5503;
  assign n5505 = ~n5294 & ~n5504;
  assign n5506 = pi0299 & ~n5505;
  assign n5507 = n2530 & ~n5350;
  assign n5508 = ~n5506 & n5507;
  assign n5509 = pi0100 & ~n5498;
  assign n5510 = ~n5508 & n5509;
  assign n5511 = ~n5497 & ~n5510;
  assign n5512 = ~pi0087 & ~n5511;
  assign n5513 = ~pi0075 & ~n5476;
  assign n5514 = ~n5512 & n5513;
  assign n5515 = ~pi0092 & ~n5475;
  assign n5516 = ~n5514 & n5515;
  assign n5517 = n2532 & ~n5474;
  assign n5518 = ~n5516 & n5517;
  assign n5519 = ~pi0055 & ~n5465;
  assign n5520 = ~n5518 & n5519;
  assign n5521 = ~pi0056 & ~n5462;
  assign n5522 = ~n5520 & n5521;
  assign n5523 = ~pi0062 & ~n5458;
  assign n5524 = ~n5522 & n5523;
  assign n5525 = n3328 & ~n5454;
  assign n5526 = ~n5524 & n5525;
  assign n5527 = pi0245 & ~n5442;
  assign n5528 = ~n5526 & n5527;
  assign po0163 = n5440 | n5528;
  assign n5530 = pi0215 & pi1135;
  assign n5531 = pi0216 & pi0279;
  assign n5532 = pi0879 & ~n2442;
  assign n5533 = pi0105 & ~n5532;
  assign n5534 = ~pi0105 & ~pi0161;
  assign n5535 = ~n5533 & ~n5534;
  assign n5536 = pi0228 & n5535;
  assign n5537 = pi0161 & ~pi0228;
  assign n5538 = ~n5536 & ~n5537;
  assign n5539 = ~pi0216 & ~n5538;
  assign n5540 = ~n5531 & ~n5539;
  assign n5541 = ~pi0221 & ~n5540;
  assign n5542 = ~pi1135 & ~n2452;
  assign n5543 = ~pi0938 & n2452;
  assign n5544 = pi0221 & ~n5542;
  assign n5545 = ~n5543 & n5544;
  assign n5546 = ~n5541 & ~n5545;
  assign n5547 = ~pi0215 & ~n5546;
  assign n5548 = ~n5530 & ~n5547;
  assign n5549 = ~n3328 & n5548;
  assign n5550 = ~n3331 & n5548;
  assign n5551 = ~pi0879 & n2521;
  assign n5552 = ~n3335 & ~n5537;
  assign n5553 = ~n5551 & ~n5552;
  assign n5554 = ~n5536 & ~n5553;
  assign n5555 = ~pi0216 & ~n5554;
  assign n5556 = ~n5531 & ~n5555;
  assign n5557 = ~pi0221 & ~n5556;
  assign n5558 = ~n5545 & ~n5557;
  assign n5559 = ~pi0215 & ~n5558;
  assign n5560 = ~n5530 & ~n5559;
  assign n5561 = n3331 & n5560;
  assign n5562 = pi0062 & ~n5550;
  assign n5563 = ~n5561 & n5562;
  assign n5564 = ~n2537 & ~n5548;
  assign n5565 = n2537 & ~n5560;
  assign n5566 = pi0056 & ~n5564;
  assign n5567 = ~n5565 & n5566;
  assign n5568 = ~n2572 & n5548;
  assign n5569 = n2572 & n5560;
  assign n5570 = pi0055 & ~n5568;
  assign n5571 = ~n5569 & n5570;
  assign n5572 = pi0223 & pi1135;
  assign n5573 = ~pi1135 & ~n2591;
  assign n5574 = ~pi0938 & n2591;
  assign n5575 = pi0222 & ~n5573;
  assign n5576 = ~n5574 & n5575;
  assign n5577 = pi0224 & ~pi0279;
  assign n5578 = ~pi0224 & ~pi0879;
  assign n5579 = ~n2442 & n5578;
  assign n5580 = ~pi0222 & ~n5577;
  assign n5581 = ~n5579 & n5580;
  assign n5582 = ~n5576 & ~n5581;
  assign n5583 = ~pi0223 & ~n5582;
  assign n5584 = ~n5572 & ~n5583;
  assign n5585 = ~pi0299 & ~n5584;
  assign n5586 = n2604 & ~n5532;
  assign n5587 = n5585 & ~n5586;
  assign n5588 = pi0299 & ~n5548;
  assign n5589 = ~n5587 & ~n5588;
  assign n5590 = ~n2532 & n5589;
  assign n5591 = ~n2625 & n5589;
  assign n5592 = pi0299 & ~n5560;
  assign n5593 = ~n5587 & ~n5592;
  assign n5594 = n2625 & n5593;
  assign n5595 = ~n5591 & ~n5594;
  assign n5596 = n2533 & ~n5595;
  assign n5597 = ~n2533 & n5589;
  assign n5598 = pi0092 & ~n5597;
  assign n5599 = ~n5596 & n5598;
  assign n5600 = pi0075 & n5589;
  assign n5601 = pi0087 & n5595;
  assign n5602 = pi0038 & n5589;
  assign n5603 = pi0039 & ~n5593;
  assign n5604 = ~pi0299 & ~n5572;
  assign n5605 = n5369 & ~n5576;
  assign n5606 = n5583 & ~n5605;
  assign n5607 = n5604 & ~n5606;
  assign n5608 = n3498 & ~n5535;
  assign n5609 = ~pi0216 & ~n5608;
  assign n5610 = pi0161 & n3499;
  assign n5611 = ~pi0161 & ~n3508;
  assign n5612 = pi0879 & ~n5610;
  assign n5613 = ~n5611 & n5612;
  assign n5614 = pi0161 & ~pi0879;
  assign n5615 = ~n3416 & n5614;
  assign n5616 = ~n5613 & ~n5615;
  assign n5617 = ~pi0228 & ~n5616;
  assign n5618 = ~n3498 & ~n5617;
  assign n5619 = n5609 & ~n5618;
  assign n5620 = ~n5531 & ~n5619;
  assign n5621 = ~pi0221 & ~n5620;
  assign n5622 = ~n5545 & ~n5621;
  assign n5623 = ~pi0215 & ~n5622;
  assign n5624 = pi0299 & ~n5530;
  assign n5625 = ~n5623 & n5624;
  assign n5626 = ~pi0039 & ~n5607;
  assign n5627 = ~n5625 & n5626;
  assign n5628 = ~pi0038 & ~n5603;
  assign n5629 = ~n5627 & n5628;
  assign n5630 = ~pi0100 & ~n5602;
  assign n5631 = ~n5629 & n5630;
  assign n5632 = ~n2530 & n5589;
  assign n5633 = ~pi0879 & n3387;
  assign n5634 = pi0161 & ~n5633;
  assign n5635 = ~pi0152 & ~pi0166;
  assign n5636 = ~n3385 & n5635;
  assign n5637 = ~n3387 & ~n5635;
  assign n5638 = pi0879 & ~n5636;
  assign n5639 = ~n5637 & n5638;
  assign n5640 = ~n5634 & ~n5639;
  assign n5641 = ~pi0228 & ~n5640;
  assign n5642 = ~n5536 & ~n5641;
  assign n5643 = ~pi0216 & ~n5642;
  assign n5644 = ~n5531 & ~n5643;
  assign n5645 = ~pi0221 & ~n5644;
  assign n5646 = ~n5545 & ~n5645;
  assign n5647 = ~pi0215 & ~n5646;
  assign n5648 = ~n5530 & ~n5647;
  assign n5649 = pi0299 & ~n5648;
  assign n5650 = n2530 & ~n5587;
  assign n5651 = ~n5649 & n5650;
  assign n5652 = pi0100 & ~n5632;
  assign n5653 = ~n5651 & n5652;
  assign n5654 = ~n5631 & ~n5653;
  assign n5655 = ~pi0087 & ~n5654;
  assign n5656 = ~pi0075 & ~n5601;
  assign n5657 = ~n5655 & n5656;
  assign n5658 = ~pi0092 & ~n5600;
  assign n5659 = ~n5657 & n5658;
  assign n5660 = n2532 & ~n5599;
  assign n5661 = ~n5659 & n5660;
  assign n5662 = ~pi0055 & ~n5590;
  assign n5663 = ~n5661 & n5662;
  assign n5664 = ~pi0056 & ~n5571;
  assign n5665 = ~n5663 & n5664;
  assign n5666 = ~pi0062 & ~n5567;
  assign n5667 = ~n5665 & n5666;
  assign n5668 = n3328 & ~n5563;
  assign n5669 = ~n5667 & n5668;
  assign n5670 = ~pi0244 & ~n5549;
  assign n5671 = ~n5669 & n5670;
  assign n5672 = ~n3450 & n5548;
  assign n5673 = ~n3328 & n5672;
  assign n5674 = ~n3447 & ~n5536;
  assign n5675 = ~n5553 & n5674;
  assign n5676 = ~pi0216 & ~n5675;
  assign n5677 = ~n5531 & ~n5676;
  assign n5678 = ~pi0221 & ~n5677;
  assign n5679 = ~n5545 & ~n5678;
  assign n5680 = ~pi0215 & ~n5679;
  assign n5681 = ~n5530 & ~n5680;
  assign n5682 = n3331 & n5681;
  assign n5683 = ~n3331 & n5672;
  assign n5684 = pi0062 & ~n5683;
  assign n5685 = ~n5682 & n5684;
  assign n5686 = ~n2537 & ~n5672;
  assign n5687 = n2537 & ~n5681;
  assign n5688 = pi0056 & ~n5686;
  assign n5689 = ~n5687 & n5688;
  assign n5690 = n2572 & n5681;
  assign n5691 = ~n2572 & n5672;
  assign n5692 = pi0055 & ~n5691;
  assign n5693 = ~n5690 & n5692;
  assign n5694 = pi0299 & ~n5672;
  assign n5695 = ~n5585 & ~n5694;
  assign n5696 = ~n2532 & n5695;
  assign n5697 = ~n2625 & n5695;
  assign n5698 = pi0299 & ~n5681;
  assign n5699 = ~n5585 & ~n5698;
  assign n5700 = n2625 & n5699;
  assign n5701 = ~n5697 & ~n5700;
  assign n5702 = n2533 & ~n5701;
  assign n5703 = ~n2533 & n5695;
  assign n5704 = pi0092 & ~n5703;
  assign n5705 = ~n5702 & n5704;
  assign n5706 = pi0075 & n5695;
  assign n5707 = pi0087 & n5701;
  assign n5708 = pi0038 & n5695;
  assign n5709 = pi0039 & ~n5699;
  assign n5710 = ~n5369 & n5582;
  assign n5711 = ~pi0223 & ~n5710;
  assign n5712 = n5604 & ~n5711;
  assign n5713 = ~pi0161 & ~n3499;
  assign n5714 = pi0161 & n3508;
  assign n5715 = ~pi0879 & ~n5713;
  assign n5716 = ~n5714 & n5715;
  assign n5717 = ~pi0161 & ~n3416;
  assign n5718 = pi0879 & ~n5717;
  assign n5719 = ~pi0228 & ~n5716;
  assign n5720 = ~n5718 & n5719;
  assign n5721 = n5609 & ~n5720;
  assign n5722 = ~n5531 & ~n5721;
  assign n5723 = ~pi0221 & ~n5722;
  assign n5724 = ~n5545 & ~n5723;
  assign n5725 = ~pi0215 & ~n5724;
  assign n5726 = n5624 & ~n5725;
  assign n5727 = ~pi0039 & ~n5712;
  assign n5728 = ~n5726 & n5727;
  assign n5729 = ~pi0038 & ~n5709;
  assign n5730 = ~n5728 & n5729;
  assign n5731 = ~pi0100 & ~n5708;
  assign n5732 = ~n5730 & n5731;
  assign n5733 = ~n2530 & n5695;
  assign n5734 = ~n5641 & n5674;
  assign n5735 = ~pi0216 & ~n5734;
  assign n5736 = ~n5531 & ~n5735;
  assign n5737 = ~pi0221 & ~n5736;
  assign n5738 = ~n5545 & ~n5737;
  assign n5739 = ~pi0215 & ~n5738;
  assign n5740 = ~n5530 & ~n5739;
  assign n5741 = pi0299 & ~n5740;
  assign n5742 = n2530 & ~n5585;
  assign n5743 = ~n5741 & n5742;
  assign n5744 = pi0100 & ~n5733;
  assign n5745 = ~n5743 & n5744;
  assign n5746 = ~n5732 & ~n5745;
  assign n5747 = ~pi0087 & ~n5746;
  assign n5748 = ~pi0075 & ~n5707;
  assign n5749 = ~n5747 & n5748;
  assign n5750 = ~pi0092 & ~n5706;
  assign n5751 = ~n5749 & n5750;
  assign n5752 = n2532 & ~n5705;
  assign n5753 = ~n5751 & n5752;
  assign n5754 = ~pi0055 & ~n5696;
  assign n5755 = ~n5753 & n5754;
  assign n5756 = ~pi0056 & ~n5693;
  assign n5757 = ~n5755 & n5756;
  assign n5758 = ~pi0062 & ~n5689;
  assign n5759 = ~n5757 & n5758;
  assign n5760 = n3328 & ~n5685;
  assign n5761 = ~n5759 & n5760;
  assign n5762 = pi0244 & ~n5673;
  assign n5763 = ~n5761 & n5762;
  assign po0164 = n5671 | n5763;
  assign n5765 = pi0216 & pi0278;
  assign n5766 = ~pi0221 & ~n5765;
  assign n5767 = ~pi0105 & pi0152;
  assign n5768 = pi0846 & ~n2442;
  assign n5769 = pi0105 & n5768;
  assign n5770 = ~n5767 & ~n5769;
  assign n5771 = pi0228 & ~n5770;
  assign n5772 = pi0152 & ~pi0228;
  assign n5773 = ~n5771 & ~n5772;
  assign n5774 = ~pi0216 & ~n5773;
  assign n5775 = n5766 & ~n5774;
  assign n5776 = pi0833 & ~pi0930;
  assign n5777 = ~pi0216 & pi0221;
  assign n5778 = n5776 & n5777;
  assign n5779 = pi0221 & ~n2452;
  assign n5780 = ~pi0215 & ~n5779;
  assign n5781 = ~n5778 & n5780;
  assign n5782 = ~n5775 & n5781;
  assign n5783 = ~n3450 & ~n5782;
  assign n5784 = ~n3328 & ~n5783;
  assign n5785 = ~n3331 & ~n5783;
  assign n5786 = ~n3447 & ~n5771;
  assign n5787 = ~pi0152 & ~n2521;
  assign n5788 = ~pi0846 & n2521;
  assign n5789 = ~pi0228 & ~n5787;
  assign n5790 = ~n5788 & n5789;
  assign n5791 = n5786 & ~n5790;
  assign n5792 = ~pi0216 & ~n5791;
  assign n5793 = n5766 & ~n5792;
  assign n5794 = n5781 & ~n5793;
  assign n5795 = n3331 & n5794;
  assign n5796 = pi0062 & ~n5785;
  assign n5797 = ~n5795 & n5796;
  assign n5798 = n2537 & ~n5794;
  assign n5799 = ~n2537 & n5783;
  assign n5800 = pi0056 & ~n5799;
  assign n5801 = ~n5798 & n5800;
  assign n5802 = ~n2572 & ~n5783;
  assign n5803 = n2572 & n5794;
  assign n5804 = pi0055 & ~n5802;
  assign n5805 = ~n5803 & n5804;
  assign n5806 = pi0224 & pi0278;
  assign n5807 = ~pi0222 & ~n5806;
  assign n5808 = ~pi0224 & n5768;
  assign n5809 = n5807 & ~n5808;
  assign n5810 = pi0222 & ~pi0224;
  assign n5811 = n5776 & n5810;
  assign n5812 = n2593 & ~n5811;
  assign n5813 = ~n5809 & n5812;
  assign n5814 = ~pi0299 & ~n5813;
  assign n5815 = ~n3755 & n5814;
  assign n5816 = pi0299 & n5783;
  assign n5817 = ~n5815 & ~n5816;
  assign n5818 = ~n2532 & n5817;
  assign n5819 = ~n2625 & n5817;
  assign n5820 = pi0299 & ~n5794;
  assign n5821 = ~n5815 & ~n5820;
  assign n5822 = n2625 & n5821;
  assign n5823 = ~n5819 & ~n5822;
  assign n5824 = n2533 & ~n5823;
  assign n5825 = ~n2533 & n5817;
  assign n5826 = pi0092 & ~n5825;
  assign n5827 = ~n5824 & n5826;
  assign n5828 = pi0075 & n5817;
  assign n5829 = pi0087 & n5823;
  assign n5830 = pi0038 & n5817;
  assign n5831 = pi0039 & ~n5821;
  assign n5832 = ~pi0846 & n3488;
  assign n5833 = ~pi0224 & ~n5832;
  assign n5834 = n5807 & ~n5833;
  assign n5835 = ~n5811 & ~n5834;
  assign n5836 = ~n2592 & n3470;
  assign n5837 = n5835 & n5836;
  assign n5838 = pi0228 & ~n5767;
  assign n5839 = pi0105 & ~n5832;
  assign n5840 = n5838 & ~n5839;
  assign n5841 = ~pi0216 & ~n5840;
  assign n5842 = ~pi0152 & n3499;
  assign n5843 = pi0152 & ~n3508;
  assign n5844 = ~pi0846 & ~n5842;
  assign n5845 = ~n5843 & n5844;
  assign n5846 = ~pi0152 & pi0846;
  assign n5847 = ~n3416 & n5846;
  assign n5848 = ~n5845 & ~n5847;
  assign n5849 = ~pi0228 & ~n5848;
  assign n5850 = n5841 & ~n5849;
  assign n5851 = n5766 & ~n5850;
  assign n5852 = ~n5778 & ~n5851;
  assign n5853 = ~pi0215 & pi0299;
  assign n5854 = ~n5779 & n5853;
  assign n5855 = n5852 & n5854;
  assign n5856 = ~pi0039 & ~n5837;
  assign n5857 = ~n5855 & n5856;
  assign n5858 = ~pi0038 & ~n5831;
  assign n5859 = ~n5857 & n5858;
  assign n5860 = ~pi0100 & ~n5830;
  assign n5861 = ~n5859 & n5860;
  assign n5862 = ~n2530 & n5817;
  assign n5863 = pi0846 & ~n3393;
  assign n5864 = ~n3388 & ~n5863;
  assign n5865 = ~pi0228 & ~n5864;
  assign n5866 = n5786 & ~n5865;
  assign n5867 = ~pi0216 & ~n5866;
  assign n5868 = n5766 & ~n5867;
  assign n5869 = n5781 & ~n5868;
  assign n5870 = pi0299 & ~n5869;
  assign n5871 = n2530 & ~n5815;
  assign n5872 = ~n5870 & n5871;
  assign n5873 = pi0100 & ~n5862;
  assign n5874 = ~n5872 & n5873;
  assign n5875 = ~n5861 & ~n5874;
  assign n5876 = ~pi0087 & ~n5875;
  assign n5877 = ~pi0075 & ~n5829;
  assign n5878 = ~n5876 & n5877;
  assign n5879 = ~pi0092 & ~n5828;
  assign n5880 = ~n5878 & n5879;
  assign n5881 = n2532 & ~n5827;
  assign n5882 = ~n5880 & n5881;
  assign n5883 = ~pi0055 & ~n5818;
  assign n5884 = ~n5882 & n5883;
  assign n5885 = ~pi0056 & ~n5805;
  assign n5886 = ~n5884 & n5885;
  assign n5887 = ~pi0062 & ~n5801;
  assign n5888 = ~n5886 & n5887;
  assign n5889 = n3328 & ~n5797;
  assign n5890 = ~n5888 & n5889;
  assign n5891 = pi0242 & ~n5784;
  assign n5892 = ~n5890 & n5891;
  assign n5893 = ~n3328 & n5782;
  assign n5894 = ~n3331 & n5782;
  assign n5895 = ~n5771 & ~n5790;
  assign n5896 = ~pi0216 & ~n5895;
  assign n5897 = n5766 & ~n5896;
  assign n5898 = n5781 & ~n5897;
  assign n5899 = n3331 & n5898;
  assign n5900 = pi0062 & ~n5894;
  assign n5901 = ~n5899 & n5900;
  assign n5902 = ~n2537 & ~n5782;
  assign n5903 = n2537 & ~n5898;
  assign n5904 = pi0056 & ~n5902;
  assign n5905 = ~n5903 & n5904;
  assign n5906 = ~n2572 & n5782;
  assign n5907 = n2572 & n5898;
  assign n5908 = pi0055 & ~n5906;
  assign n5909 = ~n5907 & n5908;
  assign n5910 = pi0299 & ~n5782;
  assign n5911 = ~n5814 & ~n5910;
  assign n5912 = ~n2532 & n5911;
  assign n5913 = ~n2625 & n5911;
  assign n5914 = pi0299 & ~n5898;
  assign n5915 = ~n5814 & ~n5914;
  assign n5916 = n2625 & n5915;
  assign n5917 = ~n5913 & ~n5916;
  assign n5918 = n2533 & ~n5917;
  assign n5919 = ~n2533 & n5911;
  assign n5920 = pi0092 & ~n5919;
  assign n5921 = ~n5918 & n5920;
  assign n5922 = pi0075 & n5911;
  assign n5923 = pi0087 & n5917;
  assign n5924 = pi0038 & n5911;
  assign n5925 = pi0039 & ~n5915;
  assign n5926 = ~n3487 & n5808;
  assign n5927 = n5807 & ~n5926;
  assign n5928 = ~n5811 & n5836;
  assign n5929 = ~n5927 & n5928;
  assign n5930 = ~n3488 & n5838;
  assign n5931 = pi0152 & ~pi0846;
  assign n5932 = ~n3416 & n5931;
  assign n5933 = pi0152 & n3499;
  assign n5934 = ~pi0152 & ~n3508;
  assign n5935 = pi0846 & ~n5933;
  assign n5936 = ~n5934 & n5935;
  assign n5937 = ~pi0228 & ~n5932;
  assign n5938 = ~n5936 & n5937;
  assign n5939 = n5841 & ~n5930;
  assign n5940 = ~n5938 & n5939;
  assign n5941 = n5766 & ~n5940;
  assign n5942 = ~n5778 & ~n5941;
  assign n5943 = n5854 & n5942;
  assign n5944 = ~pi0039 & ~n5929;
  assign n5945 = ~n5943 & n5944;
  assign n5946 = ~pi0038 & ~n5925;
  assign n5947 = ~n5945 & n5946;
  assign n5948 = ~pi0100 & ~n5924;
  assign n5949 = ~n5947 & n5948;
  assign n5950 = ~n2530 & n5911;
  assign n5951 = ~n5771 & ~n5865;
  assign n5952 = ~pi0216 & ~n5951;
  assign n5953 = n5766 & ~n5952;
  assign n5954 = n5781 & ~n5953;
  assign n5955 = pi0299 & ~n5954;
  assign n5956 = n2530 & ~n5814;
  assign n5957 = ~n5955 & n5956;
  assign n5958 = pi0100 & ~n5950;
  assign n5959 = ~n5957 & n5958;
  assign n5960 = ~n5949 & ~n5959;
  assign n5961 = ~pi0087 & ~n5960;
  assign n5962 = ~pi0075 & ~n5923;
  assign n5963 = ~n5961 & n5962;
  assign n5964 = ~pi0092 & ~n5922;
  assign n5965 = ~n5963 & n5964;
  assign n5966 = n2532 & ~n5921;
  assign n5967 = ~n5965 & n5966;
  assign n5968 = ~pi0055 & ~n5912;
  assign n5969 = ~n5967 & n5968;
  assign n5970 = ~pi0056 & ~n5909;
  assign n5971 = ~n5969 & n5970;
  assign n5972 = ~pi0062 & ~n5905;
  assign n5973 = ~n5971 & n5972;
  assign n5974 = n3328 & ~n5901;
  assign n5975 = ~n5973 & n5974;
  assign n5976 = ~pi0242 & ~n5893;
  assign n5977 = ~n5975 & n5976;
  assign n5978 = ~n5892 & ~n5977;
  assign n5979 = ~pi1134 & ~n5978;
  assign n5980 = ~n5775 & ~n5778;
  assign n5981 = ~pi0215 & ~n5980;
  assign n5982 = ~n3328 & n5981;
  assign n5983 = ~n3331 & n5981;
  assign n5984 = ~n5778 & ~n5897;
  assign n5985 = ~pi0215 & ~n5984;
  assign n5986 = n3331 & n5985;
  assign n5987 = pi0062 & ~n5983;
  assign n5988 = ~n5986 & n5987;
  assign n5989 = ~n2537 & ~n5981;
  assign n5990 = n2537 & ~n5985;
  assign n5991 = pi0056 & ~n5989;
  assign n5992 = ~n5990 & n5991;
  assign n5993 = ~n2572 & n5981;
  assign n5994 = n2572 & n5985;
  assign n5995 = pi0055 & ~n5993;
  assign n5996 = ~n5994 & n5995;
  assign n5997 = n2593 & n5815;
  assign n5998 = ~pi0299 & ~n5997;
  assign n5999 = ~pi0223 & n5809;
  assign n6000 = n5998 & ~n5999;
  assign n6001 = pi0299 & ~n5981;
  assign n6002 = ~n6000 & ~n6001;
  assign n6003 = ~n2532 & n6002;
  assign n6004 = ~n2625 & n6002;
  assign n6005 = pi0299 & ~n5985;
  assign n6006 = ~n6000 & ~n6005;
  assign n6007 = n2625 & n6006;
  assign n6008 = ~n6004 & ~n6007;
  assign n6009 = n2533 & ~n6008;
  assign n6010 = ~n2533 & n6002;
  assign n6011 = pi0092 & ~n6010;
  assign n6012 = ~n6009 & n6011;
  assign n6013 = pi0075 & n6002;
  assign n6014 = pi0087 & n6008;
  assign n6015 = pi0038 & n6002;
  assign n6016 = pi0039 & ~n6006;
  assign n6017 = n3470 & n5927;
  assign n6018 = n5853 & ~n5942;
  assign n6019 = n3470 & ~n5835;
  assign n6020 = ~pi0039 & ~n6019;
  assign n6021 = ~n6017 & n6020;
  assign n6022 = ~n6018 & n6021;
  assign n6023 = ~pi0038 & ~n6016;
  assign n6024 = ~n6022 & n6023;
  assign n6025 = ~pi0100 & ~n6015;
  assign n6026 = ~n6024 & n6025;
  assign n6027 = ~n2530 & n6002;
  assign n6028 = ~n5778 & ~n5953;
  assign n6029 = ~pi0215 & ~n6028;
  assign n6030 = pi0299 & ~n6029;
  assign n6031 = n2530 & ~n6000;
  assign n6032 = ~n6030 & n6031;
  assign n6033 = pi0100 & ~n6027;
  assign n6034 = ~n6032 & n6033;
  assign n6035 = ~n6026 & ~n6034;
  assign n6036 = ~pi0087 & ~n6035;
  assign n6037 = ~pi0075 & ~n6014;
  assign n6038 = ~n6036 & n6037;
  assign n6039 = ~pi0092 & ~n6013;
  assign n6040 = ~n6038 & n6039;
  assign n6041 = n2532 & ~n6012;
  assign n6042 = ~n6040 & n6041;
  assign n6043 = ~pi0055 & ~n6003;
  assign n6044 = ~n6042 & n6043;
  assign n6045 = ~pi0056 & ~n5996;
  assign n6046 = ~n6044 & n6045;
  assign n6047 = ~pi0062 & ~n5992;
  assign n6048 = ~n6046 & n6047;
  assign n6049 = n3328 & ~n5988;
  assign n6050 = ~n6048 & n6049;
  assign n6051 = ~pi0242 & ~n5982;
  assign n6052 = ~n6050 & n6051;
  assign n6053 = ~n3450 & n5981;
  assign n6054 = ~n3328 & n6053;
  assign n6055 = ~n5778 & ~n5793;
  assign n6056 = ~pi0215 & ~n6055;
  assign n6057 = n3331 & n6056;
  assign n6058 = ~n3331 & n6053;
  assign n6059 = pi0062 & ~n6058;
  assign n6060 = ~n6057 & n6059;
  assign n6061 = ~n2537 & ~n6053;
  assign n6062 = n2537 & ~n6056;
  assign n6063 = pi0056 & ~n6061;
  assign n6064 = ~n6062 & n6063;
  assign n6065 = n2572 & n6056;
  assign n6066 = ~n2572 & n6053;
  assign n6067 = pi0055 & ~n6066;
  assign n6068 = ~n6065 & n6067;
  assign n6069 = pi0299 & ~n6053;
  assign n6070 = ~n5998 & ~n6069;
  assign n6071 = ~n2532 & n6070;
  assign n6072 = ~n2625 & n6070;
  assign n6073 = pi0299 & ~n6056;
  assign n6074 = ~n5998 & ~n6073;
  assign n6075 = n2625 & n6074;
  assign n6076 = ~n6072 & ~n6075;
  assign n6077 = n2533 & ~n6076;
  assign n6078 = ~n2533 & n6070;
  assign n6079 = pi0092 & ~n6078;
  assign n6080 = ~n6077 & n6079;
  assign n6081 = pi0075 & n6070;
  assign n6082 = pi0087 & n6076;
  assign n6083 = pi0038 & n6070;
  assign n6084 = pi0039 & ~n6074;
  assign n6085 = ~n5852 & n5853;
  assign n6086 = n6020 & ~n6085;
  assign n6087 = ~pi0038 & ~n6084;
  assign n6088 = ~n6086 & n6087;
  assign n6089 = ~pi0100 & ~n6083;
  assign n6090 = ~n6088 & n6089;
  assign n6091 = ~n2530 & n6070;
  assign n6092 = ~n5778 & ~n5868;
  assign n6093 = ~pi0215 & ~n6092;
  assign n6094 = pi0299 & ~n6093;
  assign n6095 = n2530 & ~n5998;
  assign n6096 = ~n6094 & n6095;
  assign n6097 = pi0100 & ~n6091;
  assign n6098 = ~n6096 & n6097;
  assign n6099 = ~n6090 & ~n6098;
  assign n6100 = ~pi0087 & ~n6099;
  assign n6101 = ~pi0075 & ~n6082;
  assign n6102 = ~n6100 & n6101;
  assign n6103 = ~pi0092 & ~n6081;
  assign n6104 = ~n6102 & n6103;
  assign n6105 = n2532 & ~n6080;
  assign n6106 = ~n6104 & n6105;
  assign n6107 = ~pi0055 & ~n6071;
  assign n6108 = ~n6106 & n6107;
  assign n6109 = ~pi0056 & ~n6068;
  assign n6110 = ~n6108 & n6109;
  assign n6111 = ~pi0062 & ~n6064;
  assign n6112 = ~n6110 & n6111;
  assign n6113 = n3328 & ~n6060;
  assign n6114 = ~n6112 & n6113;
  assign n6115 = pi0242 & ~n6054;
  assign n6116 = ~n6114 & n6115;
  assign n6117 = pi1134 & ~n6052;
  assign n6118 = ~n6116 & n6117;
  assign po0165 = ~n5979 & ~n6118;
  assign n6120 = pi0057 & pi0059;
  assign n6121 = n2521 & n2538;
  assign n6122 = ~n3328 & ~n6121;
  assign n6123 = ~n6120 & ~n6122;
  assign n6124 = pi0057 & ~n6123;
  assign n6125 = n2512 & n2625;
  assign n6126 = n2536 & n6125;
  assign n6127 = pi0056 & ~n6126;
  assign n6128 = ~pi0054 & n2534;
  assign n6129 = n6125 & n6128;
  assign n6130 = pi0074 & ~n6129;
  assign n6131 = ~pi0055 & ~n6130;
  assign n6132 = pi0087 & ~n6125;
  assign n6133 = ~pi0075 & ~n6132;
  assign n6134 = ~pi0054 & ~pi0092;
  assign n6135 = ~pi0039 & n2512;
  assign n6136 = pi0038 & ~n6135;
  assign n6137 = ~pi0100 & ~n6136;
  assign n6138 = pi0058 & n2502;
  assign n6139 = ~pi0090 & ~n6138;
  assign n6140 = n2720 & n2769;
  assign n6141 = n2874 & n6140;
  assign n6142 = n2781 & ~n6141;
  assign n6143 = ~n2776 & ~n6142;
  assign n6144 = ~pi0108 & ~n6143;
  assign n6145 = n2775 & ~n6144;
  assign n6146 = ~pi0110 & n2889;
  assign n6147 = ~n6145 & n6146;
  assign n6148 = ~n2759 & ~n2766;
  assign n6149 = ~n6147 & n6148;
  assign n6150 = ~pi0047 & ~n6149;
  assign n6151 = n2700 & ~n2762;
  assign n6152 = ~n6150 & n6151;
  assign n6153 = n6139 & ~n6152;
  assign n6154 = ~n2896 & ~n6153;
  assign n6155 = ~pi0093 & ~n6154;
  assign n6156 = ~pi0841 & n2503;
  assign n6157 = pi0093 & ~n6156;
  assign n6158 = ~n6155 & ~n6157;
  assign n6159 = ~pi0035 & ~n6158;
  assign n6160 = ~pi0070 & ~n2729;
  assign n6161 = ~n6159 & n6160;
  assign n6162 = ~pi0051 & ~n6161;
  assign n6163 = n2748 & ~n6162;
  assign n6164 = n3168 & ~n6163;
  assign n6165 = n2746 & ~n6164;
  assign n6166 = n2744 & ~n6165;
  assign n6167 = ~pi0198 & ~pi0299;
  assign n6168 = ~pi0210 & pi0299;
  assign n6169 = ~n6167 & ~n6168;
  assign n6170 = ~pi0035 & n2508;
  assign n6171 = ~pi0040 & n6170;
  assign n6172 = n2915 & n6171;
  assign n6173 = pi0032 & ~n6172;
  assign n6174 = ~n6169 & ~n6173;
  assign n6175 = ~n3412 & n6169;
  assign n6176 = ~n6174 & ~n6175;
  assign n6177 = ~n6166 & ~n6176;
  assign n6178 = ~pi0095 & ~n6177;
  assign n6179 = ~n2741 & ~n6178;
  assign n6180 = ~pi0039 & ~n6179;
  assign n6181 = pi0835 & pi0984;
  assign n6182 = ~pi0252 & ~pi1001;
  assign n6183 = ~pi0979 & ~n6182;
  assign n6184 = ~n6181 & n6183;
  assign n6185 = ~pi0287 & n6184;
  assign n6186 = pi0835 & pi0950;
  assign n6187 = n6185 & n6186;
  assign n6188 = n2928 & n6187;
  assign n6189 = pi0222 & pi0224;
  assign n6190 = pi0603 & ~pi0642;
  assign n6191 = ~pi0614 & ~pi0616;
  assign n6192 = n6190 & n6191;
  assign n6193 = ~pi0662 & pi0680;
  assign n6194 = ~pi0661 & n6193;
  assign n6195 = ~pi0681 & n6194;
  assign po1101 = n6192 | n6195;
  assign n6197 = ~pi0332 & ~pi0468;
  assign n6198 = po1101 & ~n6197;
  assign n6199 = ~pi0587 & ~pi0602;
  assign n6200 = ~pi0961 & ~pi0967;
  assign n6201 = ~pi0969 & ~pi0971;
  assign n6202 = ~pi0974 & ~pi0977;
  assign n6203 = n6201 & n6202;
  assign n6204 = n6199 & n6200;
  assign n6205 = n6203 & n6204;
  assign n6206 = n6197 & ~n6205;
  assign n6207 = ~n6198 & ~n6206;
  assign n6208 = n6188 & n6189;
  assign n6209 = ~n6207 & n6208;
  assign n6210 = n2521 & ~n6209;
  assign n6211 = ~pi0223 & ~n6210;
  assign n6212 = pi1092 & n6187;
  assign n6213 = ~pi0824 & ~pi0829;
  assign n6214 = pi0824 & ~pi1091;
  assign n6215 = pi1093 & ~n2924;
  assign n6216 = ~n6214 & n6215;
  assign n6217 = ~n6213 & ~n6216;
  assign n6218 = n6212 & n6217;
  assign n6219 = ~n6197 & ~n6218;
  assign n6220 = po1101 & ~n6219;
  assign n6221 = n2521 & ~n6220;
  assign n6222 = n2512 & n6197;
  assign n6223 = po1101 & n6222;
  assign n6224 = ~n6221 & ~n6223;
  assign n6225 = n6205 & ~n6224;
  assign n6226 = ~n6192 & ~n6197;
  assign n6227 = ~n6195 & n6226;
  assign n6228 = n6218 & ~n6227;
  assign n6229 = n2521 & ~n6228;
  assign n6230 = ~n6205 & n6229;
  assign n6231 = pi0223 & ~n6230;
  assign n6232 = ~n6225 & n6231;
  assign n6233 = ~pi0299 & ~n6211;
  assign n6234 = ~n6232 & n6233;
  assign n6235 = pi0216 & pi0221;
  assign n6236 = ~pi0907 & ~pi0947;
  assign n6237 = ~pi0960 & ~pi0963;
  assign n6238 = ~pi0970 & ~pi0972;
  assign n6239 = ~pi0975 & ~pi0978;
  assign n6240 = n6238 & n6239;
  assign n6241 = n6237 & n6240;
  assign n6242 = n6236 & n6241;
  assign n6243 = n6197 & ~n6242;
  assign n6244 = ~n6198 & ~n6243;
  assign n6245 = n6188 & n6235;
  assign n6246 = ~n6244 & n6245;
  assign n6247 = n2521 & ~n6246;
  assign n6248 = ~pi0215 & ~n6247;
  assign n6249 = n6229 & ~n6242;
  assign n6250 = ~n6224 & n6242;
  assign n6251 = pi0215 & ~n6249;
  assign n6252 = ~n6250 & n6251;
  assign n6253 = pi0299 & ~n6248;
  assign n6254 = ~n6252 & n6253;
  assign n6255 = pi0039 & ~n6234;
  assign n6256 = ~n6254 & n6255;
  assign n6257 = ~n6180 & ~n6256;
  assign n6258 = ~pi0038 & ~n6257;
  assign n6259 = n6137 & ~n6258;
  assign n6260 = ~pi0142 & ~n2669;
  assign n6261 = ~pi0299 & n6260;
  assign n6262 = pi0299 & n2640;
  assign n6263 = ~n6261 & ~n6262;
  assign n6264 = ~n3385 & n6263;
  assign n6265 = ~pi0041 & ~pi0099;
  assign n6266 = ~pi0101 & n6265;
  assign n6267 = ~pi0042 & ~pi0043;
  assign n6268 = ~pi0052 & n6267;
  assign n6269 = ~pi0113 & ~pi0116;
  assign n6270 = ~pi0114 & ~pi0115;
  assign n6271 = n6269 & n6270;
  assign n6272 = n6268 & n6271;
  assign n6273 = n6266 & n6272;
  assign po1057 = pi0044 | ~n6273;
  assign n6275 = ~pi0683 & po1057;
  assign n6276 = pi0129 & pi0250;
  assign n6277 = n2932 & ~n6213;
  assign po0740 = ~pi1093 & n6277;
  assign n6279 = ~pi0250 & ~po0740;
  assign n6280 = ~n6276 & ~n6279;
  assign n6281 = ~n6275 & ~n6280;
  assign n6282 = ~n6263 & po1057;
  assign n6283 = n6281 & n6282;
  assign n6284 = ~pi0039 & n2521;
  assign n6285 = ~pi0038 & pi0100;
  assign n6286 = n6284 & n6285;
  assign n6287 = ~n6264 & ~n6283;
  assign n6288 = n6286 & n6287;
  assign n6289 = ~pi0087 & ~n6288;
  assign n6290 = ~n6259 & n6289;
  assign n6291 = n6133 & n6134;
  assign n6292 = ~n6290 & n6291;
  assign n6293 = ~pi0074 & ~n6292;
  assign n6294 = n6131 & ~n6293;
  assign n6295 = ~pi0056 & ~n6294;
  assign n6296 = ~n6127 & ~n6295;
  assign n6297 = ~pi0062 & ~n6296;
  assign n6298 = n3330 & n6125;
  assign n6299 = pi0062 & ~n6298;
  assign n6300 = ~pi0059 & ~n6299;
  assign n6301 = ~n6297 & n6300;
  assign n6302 = ~pi0057 & ~n6301;
  assign po0167 = ~n6124 & ~n6302;
  assign n6304 = ~pi0055 & n2529;
  assign n6305 = ~pi0059 & n6304;
  assign n6306 = ~pi0228 & ~n6305;
  assign n6307 = pi0057 & ~n6306;
  assign n6308 = ~n6195 & ~n6197;
  assign n6309 = ~pi0907 & n6197;
  assign n6310 = ~n6308 & ~n6309;
  assign n6311 = ~pi0228 & ~n2572;
  assign n6312 = pi0030 & pi0228;
  assign n6313 = ~n3335 & ~n6312;
  assign n6314 = ~n6311 & ~n6313;
  assign n6315 = n6310 & n6314;
  assign n6316 = n6307 & n6315;
  assign n6317 = ~pi0228 & ~n6304;
  assign n6318 = n6315 & ~n6317;
  assign n6319 = pi0059 & ~n6318;
  assign n6320 = n6310 & n6312;
  assign n6321 = ~n2529 & n6320;
  assign n6322 = pi0055 & ~n6315;
  assign n6323 = ~pi0054 & n2569;
  assign n6324 = pi0299 & n6310;
  assign n6325 = ~pi0602 & n6197;
  assign n6326 = ~n6308 & ~n6325;
  assign n6327 = ~pi0299 & n6326;
  assign n6328 = ~n6324 & ~n6327;
  assign n6329 = n6312 & ~n6328;
  assign n6330 = ~n6323 & ~n6329;
  assign n6331 = ~n2610 & n6329;
  assign n6332 = ~pi0039 & ~n6313;
  assign n6333 = ~n6328 & n6332;
  assign n6334 = n2620 & n6333;
  assign n6335 = ~n6331 & ~n6334;
  assign n6336 = n2569 & n6335;
  assign n6337 = ~pi0054 & n6336;
  assign n6338 = pi0074 & ~n6330;
  assign n6339 = ~n6337 & n6338;
  assign n6340 = ~n2569 & ~n6329;
  assign n6341 = ~n6336 & ~n6340;
  assign n6342 = pi0054 & ~n6341;
  assign n6343 = ~pi0075 & n6335;
  assign n6344 = pi0075 & ~n6329;
  assign n6345 = pi0092 & ~n6344;
  assign n6346 = ~n6343 & n6345;
  assign n6347 = pi0075 & n6335;
  assign n6348 = pi0087 & n6329;
  assign n6349 = ~n2530 & n6329;
  assign n6350 = n6312 & n6326;
  assign n6351 = n2521 & ~n6280;
  assign n6352 = pi0683 & po1057;
  assign n6353 = n6351 & n6352;
  assign n6354 = ~n6308 & n6353;
  assign n6355 = n6260 & n6354;
  assign n6356 = pi0252 & ~n6260;
  assign n6357 = pi0252 & n6222;
  assign n6358 = ~n6195 & n6357;
  assign n6359 = pi0252 & n2521;
  assign n6360 = n6195 & n6359;
  assign n6361 = ~n6358 & ~n6360;
  assign n6362 = n6356 & ~n6361;
  assign n6363 = ~n6355 & ~n6362;
  assign n6364 = ~pi0228 & ~n6325;
  assign n6365 = ~n6363 & n6364;
  assign n6366 = ~pi0299 & ~n6350;
  assign n6367 = ~n6365 & n6366;
  assign n6368 = pi0299 & ~n6320;
  assign n6369 = n2640 & ~n6354;
  assign n6370 = ~n2640 & n6361;
  assign n6371 = ~pi0228 & ~n6309;
  assign n6372 = ~n6369 & n6371;
  assign n6373 = ~n6370 & n6372;
  assign n6374 = n6368 & ~n6373;
  assign n6375 = n2530 & ~n6374;
  assign n6376 = ~n6367 & n6375;
  assign n6377 = pi0100 & ~n6349;
  assign n6378 = ~n6376 & n6377;
  assign n6379 = ~pi0215 & pi0221;
  assign n6380 = ~pi0287 & n2521;
  assign n6381 = pi0835 & n6184;
  assign n6382 = n6380 & n6381;
  assign n6383 = pi0824 & pi1093;
  assign n6384 = n2932 & n6383;
  assign n6385 = n6382 & n6384;
  assign n6386 = ~pi1091 & n6385;
  assign n6387 = pi1091 & n2923;
  assign n6388 = n6384 & ~n6387;
  assign n6389 = ~n2928 & ~n6388;
  assign n6390 = pi1091 & ~n6389;
  assign n6391 = n6382 & n6390;
  assign n6392 = ~n6386 & ~n6391;
  assign n6393 = pi0216 & ~n6392;
  assign n6394 = ~pi0829 & ~n2923;
  assign n6395 = pi1091 & ~n6394;
  assign n6396 = n6385 & ~n6395;
  assign n6397 = ~pi0216 & n6396;
  assign n6398 = ~n6393 & ~n6397;
  assign n6399 = ~pi0228 & ~n6398;
  assign n6400 = ~n6312 & ~n6399;
  assign n6401 = n6379 & ~n6400;
  assign n6402 = ~n6312 & ~n6401;
  assign n6403 = n6310 & ~n6402;
  assign n6404 = pi0299 & ~n6403;
  assign n6405 = pi0222 & ~pi0223;
  assign n6406 = ~pi0224 & ~n6396;
  assign n6407 = pi0224 & n6392;
  assign n6408 = n6405 & ~n6406;
  assign n6409 = ~n6407 & n6408;
  assign n6410 = ~pi0228 & n6409;
  assign n6411 = ~n6312 & ~n6410;
  assign n6412 = n6326 & ~n6411;
  assign n6413 = ~pi0299 & ~n6412;
  assign n6414 = pi0039 & ~n6413;
  assign n6415 = ~n6404 & n6414;
  assign n6416 = pi0158 & pi0159;
  assign n6417 = pi0160 & pi0197;
  assign n6418 = n6416 & n6417;
  assign n6419 = pi0091 & ~n2755;
  assign n6420 = ~pi0058 & ~n6419;
  assign n6421 = ~pi0091 & ~pi0314;
  assign n6422 = n2765 & ~n2766;
  assign n6423 = pi0067 & n2483;
  assign n6424 = pi0085 & n2827;
  assign n6425 = n2469 & ~n6424;
  assign n6426 = n2831 & ~n6425;
  assign n6427 = n2478 & ~n6426;
  assign n6428 = ~n2810 & ~n2811;
  assign n6429 = ~n6427 & n6428;
  assign n6430 = n2479 & n6429;
  assign n6431 = ~n2807 & ~n6430;
  assign n6432 = n2804 & ~n6431;
  assign n6433 = n2797 & ~n6423;
  assign n6434 = ~n6432 & n6433;
  assign n6435 = n2796 & ~n6434;
  assign n6436 = ~pi0071 & ~n6435;
  assign po1049 = pi0064 | ~n2487;
  assign n6438 = n2791 & ~po1049;
  assign n6439 = ~n6436 & n6438;
  assign n6440 = ~pi0081 & ~n6439;
  assign n6441 = n2845 & n6438;
  assign n6442 = n6440 & ~n6441;
  assign n6443 = ~pi0102 & ~n2786;
  assign n6444 = n2463 & n6443;
  assign n6445 = ~n6442 & n6444;
  assign n6446 = n2785 & ~n6445;
  assign n6447 = n2877 & ~n6446;
  assign n6448 = n2719 & ~n6447;
  assign n6449 = ~n2722 & ~n6448;
  assign n6450 = ~pi0086 & ~n6449;
  assign n6451 = ~pi0046 & n2496;
  assign n6452 = n2783 & n6451;
  assign n6453 = ~n6450 & n6452;
  assign n6454 = n2889 & ~n6453;
  assign n6455 = n6422 & ~n6454;
  assign n6456 = n6421 & ~n6455;
  assign n6457 = ~pi0091 & pi0314;
  assign n6458 = ~n6440 & n6444;
  assign n6459 = n2785 & ~n6458;
  assign n6460 = n2877 & ~n6459;
  assign n6461 = n2719 & ~n6460;
  assign n6462 = ~n2722 & ~n6461;
  assign n6463 = ~pi0086 & ~n6462;
  assign n6464 = n6452 & ~n6463;
  assign n6465 = n2889 & ~n6464;
  assign n6466 = n6422 & ~n6465;
  assign n6467 = n6457 & ~n6466;
  assign n6468 = n6420 & ~n6467;
  assign n6469 = ~n6456 & n6468;
  assign n6470 = ~pi0090 & ~n6469;
  assign n6471 = ~n2896 & ~n6470;
  assign n6472 = ~pi0093 & ~n6471;
  assign n6473 = pi0093 & ~n2914;
  assign n6474 = ~pi0035 & ~n6473;
  assign n6475 = ~n6472 & n6474;
  assign n6476 = ~pi0070 & ~n6475;
  assign n6477 = n3100 & ~n6476;
  assign n6478 = ~pi0072 & ~n6477;
  assign n6479 = ~pi0095 & n2510;
  assign n6480 = ~n2745 & n6479;
  assign n6481 = ~n6478 & n6480;
  assign n6482 = ~n3181 & ~n6481;
  assign n6483 = ~pi0841 & n2728;
  assign n6484 = n2962 & n6483;
  assign n6485 = n2736 & n6484;
  assign n6486 = pi0032 & n6485;
  assign n6487 = ~pi0095 & n6486;
  assign n6488 = ~pi0210 & n6487;
  assign n6489 = n6482 & ~n6488;
  assign n6490 = ~n6197 & ~n6489;
  assign n6491 = ~pi0047 & n2493;
  assign n6492 = ~n2888 & ~n6453;
  assign n6493 = n6491 & ~n6492;
  assign n6494 = n6421 & ~n6493;
  assign n6495 = ~n2888 & ~n6464;
  assign n6496 = n6491 & ~n6495;
  assign n6497 = n6457 & ~n6496;
  assign n6498 = n6420 & ~n6497;
  assign n6499 = ~n6494 & n6498;
  assign n6500 = ~pi0090 & ~n6499;
  assign n6501 = ~n2896 & ~n6500;
  assign n6502 = ~pi0093 & ~n6501;
  assign n6503 = n6474 & ~n6502;
  assign n6504 = ~pi0070 & ~n6503;
  assign n6505 = n3100 & ~n6504;
  assign n6506 = ~pi0072 & ~n6505;
  assign n6507 = n6480 & ~n6506;
  assign n6508 = ~n3181 & ~n6507;
  assign n6509 = ~n6488 & n6508;
  assign n6510 = n6197 & ~n6509;
  assign n6511 = ~n6490 & ~n6510;
  assign n6512 = n6310 & ~n6511;
  assign n6513 = n6418 & ~n6512;
  assign n6514 = n6310 & ~n6489;
  assign n6515 = ~n6418 & ~n6514;
  assign n6516 = ~pi0228 & ~n6515;
  assign n6517 = ~n6513 & n6516;
  assign n6518 = n6368 & ~n6517;
  assign n6519 = ~pi0198 & n6487;
  assign n6520 = n6482 & ~n6519;
  assign n6521 = ~pi0228 & ~n6520;
  assign n6522 = ~n6312 & ~n6521;
  assign n6523 = n6326 & ~n6522;
  assign n6524 = ~pi0299 & ~n6523;
  assign n6525 = pi0145 & pi0180;
  assign n6526 = pi0181 & pi0182;
  assign n6527 = n6525 & n6526;
  assign n6528 = ~pi0299 & n6527;
  assign n6529 = ~n6524 & ~n6528;
  assign n6530 = ~n6197 & ~n6520;
  assign n6531 = n6508 & ~n6519;
  assign n6532 = n6197 & ~n6531;
  assign n6533 = ~n6530 & ~n6532;
  assign n6534 = ~pi0228 & n6326;
  assign n6535 = ~n6533 & n6534;
  assign n6536 = ~n6350 & ~n6535;
  assign n6537 = n6527 & ~n6536;
  assign n6538 = ~n6529 & ~n6537;
  assign n6539 = pi0232 & ~n6518;
  assign n6540 = ~n6538 & n6539;
  assign n6541 = ~pi0228 & n6514;
  assign n6542 = n6368 & ~n6541;
  assign n6543 = ~pi0232 & ~n6542;
  assign n6544 = ~n6524 & n6543;
  assign n6545 = ~n6540 & ~n6544;
  assign n6546 = ~pi0039 & ~n6545;
  assign n6547 = ~pi0038 & ~n6415;
  assign n6548 = ~n6546 & n6547;
  assign n6549 = pi0038 & ~n6329;
  assign n6550 = ~n6333 & n6549;
  assign n6551 = ~n6548 & ~n6550;
  assign n6552 = ~pi0100 & ~n6551;
  assign n6553 = ~pi0087 & ~n6378;
  assign n6554 = ~n6552 & n6553;
  assign n6555 = ~pi0075 & ~n6348;
  assign n6556 = ~n6554 & n6555;
  assign n6557 = ~pi0092 & ~n6347;
  assign n6558 = ~n6556 & n6557;
  assign n6559 = ~pi0054 & ~n6346;
  assign n6560 = ~n6558 & n6559;
  assign n6561 = ~pi0074 & ~n6342;
  assign n6562 = ~n6560 & n6561;
  assign n6563 = ~pi0055 & ~n6339;
  assign n6564 = ~n6562 & n6563;
  assign n6565 = n2529 & ~n6322;
  assign n6566 = ~n6564 & n6565;
  assign n6567 = ~pi0059 & ~n6321;
  assign n6568 = ~n6566 & n6567;
  assign n6569 = ~pi0057 & ~n6319;
  assign n6570 = ~n6568 & n6569;
  assign po0171 = ~n6316 & ~n6570;
  assign n6572 = ~pi0947 & n6197;
  assign n6573 = ~n6226 & ~n6572;
  assign n6574 = n6314 & n6573;
  assign n6575 = n6307 & n6574;
  assign n6576 = ~n6317 & n6574;
  assign n6577 = pi0059 & ~n6576;
  assign n6578 = n6312 & n6573;
  assign n6579 = ~n2529 & n6578;
  assign n6580 = pi0055 & ~n6574;
  assign n6581 = pi0299 & ~n6573;
  assign n6582 = ~pi0587 & n6197;
  assign n6583 = ~n6226 & ~n6582;
  assign n6584 = ~pi0299 & ~n6583;
  assign n6585 = ~n6581 & ~n6584;
  assign n6586 = n6312 & n6585;
  assign n6587 = ~n6323 & ~n6586;
  assign n6588 = ~n2610 & n6586;
  assign n6589 = n6332 & n6585;
  assign n6590 = n2620 & n6589;
  assign n6591 = ~n6588 & ~n6590;
  assign n6592 = n2569 & n6591;
  assign n6593 = ~pi0054 & n6592;
  assign n6594 = pi0074 & ~n6587;
  assign n6595 = ~n6593 & n6594;
  assign n6596 = ~n2569 & ~n6586;
  assign n6597 = ~n6592 & ~n6596;
  assign n6598 = pi0054 & ~n6597;
  assign n6599 = ~pi0075 & n6591;
  assign n6600 = pi0075 & ~n6586;
  assign n6601 = pi0092 & ~n6600;
  assign n6602 = ~n6599 & n6601;
  assign n6603 = pi0075 & n6591;
  assign n6604 = pi0087 & n6586;
  assign n6605 = ~n2530 & n6586;
  assign n6606 = pi0299 & ~n6578;
  assign n6607 = ~n6226 & n6353;
  assign n6608 = n2640 & ~n6572;
  assign n6609 = n6607 & n6608;
  assign n6610 = ~n6192 & ~n6357;
  assign n6611 = n6192 & ~n6359;
  assign n6612 = ~n6610 & ~n6611;
  assign n6613 = n6192 & ~n6197;
  assign n6614 = ~pi0947 & ~n6613;
  assign n6615 = ~n2640 & ~n6614;
  assign n6616 = n6612 & n6615;
  assign n6617 = ~n6609 & ~n6616;
  assign n6618 = ~pi0228 & ~n6617;
  assign n6619 = n6606 & ~n6618;
  assign n6620 = ~pi0228 & n2669;
  assign n6621 = ~n6582 & n6612;
  assign n6622 = n6620 & ~n6621;
  assign n6623 = ~pi0587 & ~n6613;
  assign n6624 = pi0142 & ~n6612;
  assign n6625 = ~pi0142 & ~n6607;
  assign n6626 = ~pi0228 & ~n6623;
  assign n6627 = ~n6625 & n6626;
  assign n6628 = ~n6624 & n6627;
  assign n6629 = n6312 & n6583;
  assign n6630 = ~n6620 & ~n6629;
  assign n6631 = ~n6628 & n6630;
  assign n6632 = ~n6622 & ~n6631;
  assign n6633 = ~pi0299 & ~n6632;
  assign n6634 = n2530 & ~n6619;
  assign n6635 = ~n6633 & n6634;
  assign n6636 = pi0100 & ~n6605;
  assign n6637 = ~n6635 & n6636;
  assign n6638 = ~n6411 & n6583;
  assign n6639 = ~pi0299 & ~n6638;
  assign n6640 = pi0299 & n6379;
  assign n6641 = ~n6606 & ~n6640;
  assign n6642 = n6401 & n6573;
  assign n6643 = ~n6641 & ~n6642;
  assign n6644 = pi0039 & ~n6639;
  assign n6645 = ~n6643 & n6644;
  assign n6646 = ~n6511 & n6573;
  assign n6647 = n6418 & ~n6646;
  assign n6648 = ~n6489 & n6573;
  assign n6649 = ~n6418 & ~n6648;
  assign n6650 = ~pi0228 & ~n6649;
  assign n6651 = ~n6647 & n6650;
  assign n6652 = n6606 & ~n6651;
  assign n6653 = ~n6522 & n6583;
  assign n6654 = ~n6527 & n6653;
  assign n6655 = ~pi0228 & n6583;
  assign n6656 = ~n6533 & n6655;
  assign n6657 = ~n6629 & ~n6656;
  assign n6658 = n6527 & ~n6657;
  assign n6659 = ~pi0299 & ~n6654;
  assign n6660 = ~n6658 & n6659;
  assign n6661 = pi0232 & ~n6652;
  assign n6662 = ~n6660 & n6661;
  assign n6663 = ~pi0228 & n6648;
  assign n6664 = n6606 & ~n6663;
  assign n6665 = ~pi0299 & ~n6653;
  assign n6666 = ~pi0232 & ~n6664;
  assign n6667 = ~n6665 & n6666;
  assign n6668 = ~n6662 & ~n6667;
  assign n6669 = ~pi0039 & ~n6668;
  assign n6670 = ~pi0038 & ~n6645;
  assign n6671 = ~n6669 & n6670;
  assign n6672 = pi0038 & ~n6586;
  assign n6673 = ~n6589 & n6672;
  assign n6674 = ~n6671 & ~n6673;
  assign n6675 = ~pi0100 & ~n6674;
  assign n6676 = ~pi0087 & ~n6637;
  assign n6677 = ~n6675 & n6676;
  assign n6678 = ~pi0075 & ~n6604;
  assign n6679 = ~n6677 & n6678;
  assign n6680 = ~pi0092 & ~n6603;
  assign n6681 = ~n6679 & n6680;
  assign n6682 = ~pi0054 & ~n6602;
  assign n6683 = ~n6681 & n6682;
  assign n6684 = ~pi0074 & ~n6598;
  assign n6685 = ~n6683 & n6684;
  assign n6686 = ~pi0055 & ~n6595;
  assign n6687 = ~n6685 & n6686;
  assign n6688 = n2529 & ~n6580;
  assign n6689 = ~n6687 & n6688;
  assign n6690 = ~pi0059 & ~n6579;
  assign n6691 = ~n6689 & n6690;
  assign n6692 = ~pi0057 & ~n6577;
  assign n6693 = ~n6691 & n6692;
  assign po0172 = ~n6575 & ~n6693;
  assign n6695 = pi0030 & n6197;
  assign n6696 = pi0228 & n6695;
  assign n6697 = pi0970 & n6696;
  assign n6698 = ~pi0228 & pi0970;
  assign n6699 = n6222 & n6698;
  assign n6700 = n2572 & n6699;
  assign n6701 = n6305 & n6700;
  assign n6702 = ~n6697 & ~n6701;
  assign n6703 = pi0057 & ~n6702;
  assign n6704 = n6304 & n6700;
  assign n6705 = pi0059 & ~n6697;
  assign n6706 = ~n6704 & n6705;
  assign n6707 = ~n2529 & n6697;
  assign n6708 = pi0055 & ~n6697;
  assign n6709 = ~n6700 & n6708;
  assign n6710 = pi0299 & pi0970;
  assign n6711 = ~pi0299 & pi0967;
  assign n6712 = ~n6710 & ~n6711;
  assign n6713 = n6696 & ~n6712;
  assign n6714 = ~n6323 & ~n6713;
  assign n6715 = ~n2610 & n6713;
  assign n6716 = pi0299 & ~n6697;
  assign n6717 = ~n6699 & n6716;
  assign n6718 = pi0228 & ~n6695;
  assign n6719 = ~pi0228 & ~n6222;
  assign n6720 = ~n6718 & ~n6719;
  assign n6721 = pi0967 & n6720;
  assign n6722 = ~pi0299 & ~n6721;
  assign n6723 = ~pi0039 & ~n6717;
  assign n6724 = ~n6722 & n6723;
  assign n6725 = n2620 & n6724;
  assign n6726 = ~n6715 & ~n6725;
  assign n6727 = n2569 & n6726;
  assign n6728 = ~pi0054 & n6727;
  assign n6729 = pi0074 & ~n6714;
  assign n6730 = ~n6728 & n6729;
  assign n6731 = ~n2569 & ~n6713;
  assign n6732 = ~n6727 & ~n6731;
  assign n6733 = pi0054 & ~n6732;
  assign n6734 = ~pi0075 & n6726;
  assign n6735 = pi0075 & ~n6713;
  assign n6736 = pi0092 & ~n6735;
  assign n6737 = ~n6734 & n6736;
  assign n6738 = pi0075 & n6726;
  assign n6739 = pi0087 & n6713;
  assign n6740 = ~n2530 & n6713;
  assign n6741 = ~n2640 & ~n6357;
  assign n6742 = n6197 & n6353;
  assign n6743 = n2640 & ~n6742;
  assign n6744 = ~pi0228 & ~n6741;
  assign n6745 = ~n6743 & n6744;
  assign n6746 = pi0970 & n6745;
  assign n6747 = n6716 & ~n6746;
  assign n6748 = ~n6260 & n6357;
  assign n6749 = n6260 & n6742;
  assign n6750 = ~pi0228 & ~n6748;
  assign n6751 = ~n6749 & n6750;
  assign n6752 = ~n6718 & ~n6751;
  assign n6753 = pi0967 & n6752;
  assign n6754 = ~pi0299 & ~n6753;
  assign n6755 = n2530 & ~n6747;
  assign n6756 = ~n6754 & n6755;
  assign n6757 = pi0100 & ~n6740;
  assign n6758 = ~n6756 & n6757;
  assign n6759 = n6379 & ~n6398;
  assign n6760 = n6197 & n6759;
  assign n6761 = ~pi0228 & ~n6760;
  assign n6762 = n6710 & ~n6761;
  assign n6763 = n6197 & n6409;
  assign n6764 = ~pi0228 & ~n6763;
  assign n6765 = n6711 & ~n6764;
  assign n6766 = ~n6762 & ~n6765;
  assign n6767 = pi0039 & ~n6718;
  assign n6768 = ~n6766 & n6767;
  assign n6769 = n6197 & ~n6522;
  assign n6770 = ~n6527 & ~n6769;
  assign n6771 = ~n6520 & ~n6527;
  assign n6772 = ~pi0228 & n6532;
  assign n6773 = ~n6696 & ~n6771;
  assign n6774 = ~n6772 & n6773;
  assign n6775 = ~n6770 & ~n6774;
  assign n6776 = pi0967 & n6775;
  assign n6777 = ~pi0299 & ~n6776;
  assign n6778 = n6197 & ~n6489;
  assign n6779 = n6698 & n6778;
  assign n6780 = n6716 & ~n6779;
  assign n6781 = pi0299 & n6416;
  assign n6782 = ~n6780 & ~n6781;
  assign n6783 = n6417 & ~n6510;
  assign n6784 = ~n6417 & n6489;
  assign n6785 = ~n6783 & ~n6784;
  assign n6786 = n6197 & n6785;
  assign n6787 = n6698 & n6786;
  assign n6788 = ~n6697 & ~n6787;
  assign n6789 = n6416 & ~n6788;
  assign n6790 = ~n6782 & ~n6789;
  assign n6791 = pi0232 & ~n6777;
  assign n6792 = ~n6790 & n6791;
  assign n6793 = pi0967 & n6769;
  assign n6794 = ~pi0299 & ~n6793;
  assign n6795 = ~pi0232 & ~n6780;
  assign n6796 = ~n6794 & n6795;
  assign n6797 = ~n6792 & ~n6796;
  assign n6798 = ~pi0039 & ~n6797;
  assign n6799 = ~pi0038 & ~n6768;
  assign n6800 = ~n6798 & n6799;
  assign n6801 = pi0039 & n6713;
  assign n6802 = pi0038 & ~n6801;
  assign n6803 = ~n6724 & n6802;
  assign n6804 = ~n6800 & ~n6803;
  assign n6805 = ~pi0100 & ~n6804;
  assign n6806 = ~pi0087 & ~n6758;
  assign n6807 = ~n6805 & n6806;
  assign n6808 = ~pi0075 & ~n6739;
  assign n6809 = ~n6807 & n6808;
  assign n6810 = ~pi0092 & ~n6738;
  assign n6811 = ~n6809 & n6810;
  assign n6812 = ~pi0054 & ~n6737;
  assign n6813 = ~n6811 & n6812;
  assign n6814 = ~pi0074 & ~n6733;
  assign n6815 = ~n6813 & n6814;
  assign n6816 = ~pi0055 & ~n6730;
  assign n6817 = ~n6815 & n6816;
  assign n6818 = n2529 & ~n6709;
  assign n6819 = ~n6817 & n6818;
  assign n6820 = ~pi0059 & ~n6707;
  assign n6821 = ~n6819 & n6820;
  assign n6822 = ~pi0057 & ~n6706;
  assign n6823 = ~n6821 & n6822;
  assign po0173 = ~n6703 & ~n6823;
  assign n6825 = pi0972 & n6696;
  assign n6826 = ~pi0228 & pi0972;
  assign n6827 = n6222 & n6826;
  assign n6828 = n2572 & n6827;
  assign n6829 = n6305 & n6828;
  assign n6830 = ~n6825 & ~n6829;
  assign n6831 = pi0057 & ~n6830;
  assign n6832 = n6304 & n6828;
  assign n6833 = pi0059 & ~n6825;
  assign n6834 = ~n6832 & n6833;
  assign n6835 = ~n2529 & n6825;
  assign n6836 = pi0055 & ~n6825;
  assign n6837 = ~n6828 & n6836;
  assign n6838 = ~pi0299 & pi0961;
  assign n6839 = pi0299 & pi0972;
  assign n6840 = ~n6838 & ~n6839;
  assign n6841 = n6696 & ~n6840;
  assign n6842 = ~n6323 & ~n6841;
  assign n6843 = ~n2610 & n6841;
  assign n6844 = pi0299 & ~n6825;
  assign n6845 = ~n6827 & n6844;
  assign n6846 = pi0961 & n6720;
  assign n6847 = ~pi0299 & ~n6846;
  assign n6848 = ~pi0039 & ~n6845;
  assign n6849 = ~n6847 & n6848;
  assign n6850 = n2620 & n6849;
  assign n6851 = ~n6843 & ~n6850;
  assign n6852 = n2569 & n6851;
  assign n6853 = ~pi0054 & n6852;
  assign n6854 = pi0074 & ~n6842;
  assign n6855 = ~n6853 & n6854;
  assign n6856 = ~n2569 & ~n6841;
  assign n6857 = ~n6852 & ~n6856;
  assign n6858 = pi0054 & ~n6857;
  assign n6859 = ~pi0075 & n6851;
  assign n6860 = pi0075 & ~n6841;
  assign n6861 = pi0092 & ~n6860;
  assign n6862 = ~n6859 & n6861;
  assign n6863 = pi0075 & n6851;
  assign n6864 = pi0087 & n6841;
  assign n6865 = ~n2530 & n6841;
  assign n6866 = pi0972 & n6745;
  assign n6867 = n6844 & ~n6866;
  assign n6868 = pi0961 & n6752;
  assign n6869 = ~pi0299 & ~n6868;
  assign n6870 = n2530 & ~n6867;
  assign n6871 = ~n6869 & n6870;
  assign n6872 = pi0100 & ~n6865;
  assign n6873 = ~n6871 & n6872;
  assign n6874 = ~n6764 & n6838;
  assign n6875 = ~n6761 & n6839;
  assign n6876 = ~n6874 & ~n6875;
  assign n6877 = n6767 & ~n6876;
  assign n6878 = pi0961 & n6775;
  assign n6879 = ~pi0299 & ~n6878;
  assign n6880 = n6778 & n6826;
  assign n6881 = n6844 & ~n6880;
  assign n6882 = ~n6781 & ~n6881;
  assign n6883 = n6786 & n6826;
  assign n6884 = ~n6825 & ~n6883;
  assign n6885 = n6416 & ~n6884;
  assign n6886 = ~n6882 & ~n6885;
  assign n6887 = pi0232 & ~n6879;
  assign n6888 = ~n6886 & n6887;
  assign n6889 = pi0961 & n6769;
  assign n6890 = ~pi0299 & ~n6889;
  assign n6891 = ~pi0232 & ~n6881;
  assign n6892 = ~n6890 & n6891;
  assign n6893 = ~n6888 & ~n6892;
  assign n6894 = ~pi0039 & ~n6893;
  assign n6895 = ~pi0038 & ~n6877;
  assign n6896 = ~n6894 & n6895;
  assign n6897 = pi0039 & n6841;
  assign n6898 = pi0038 & ~n6897;
  assign n6899 = ~n6849 & n6898;
  assign n6900 = ~n6896 & ~n6899;
  assign n6901 = ~pi0100 & ~n6900;
  assign n6902 = ~pi0087 & ~n6873;
  assign n6903 = ~n6901 & n6902;
  assign n6904 = ~pi0075 & ~n6864;
  assign n6905 = ~n6903 & n6904;
  assign n6906 = ~pi0092 & ~n6863;
  assign n6907 = ~n6905 & n6906;
  assign n6908 = ~pi0054 & ~n6862;
  assign n6909 = ~n6907 & n6908;
  assign n6910 = ~pi0074 & ~n6858;
  assign n6911 = ~n6909 & n6910;
  assign n6912 = ~pi0055 & ~n6855;
  assign n6913 = ~n6911 & n6912;
  assign n6914 = n2529 & ~n6837;
  assign n6915 = ~n6913 & n6914;
  assign n6916 = ~pi0059 & ~n6835;
  assign n6917 = ~n6915 & n6916;
  assign n6918 = ~pi0057 & ~n6834;
  assign n6919 = ~n6917 & n6918;
  assign po0174 = ~n6831 & ~n6919;
  assign n6921 = pi0960 & n6696;
  assign n6922 = ~pi0228 & pi0960;
  assign n6923 = n6222 & n6922;
  assign n6924 = n2572 & n6923;
  assign n6925 = n6305 & n6924;
  assign n6926 = ~n6921 & ~n6925;
  assign n6927 = pi0057 & ~n6926;
  assign n6928 = n6304 & n6924;
  assign n6929 = pi0059 & ~n6921;
  assign n6930 = ~n6928 & n6929;
  assign n6931 = ~n2529 & n6921;
  assign n6932 = pi0055 & ~n6921;
  assign n6933 = ~n6924 & n6932;
  assign n6934 = ~pi0299 & pi0977;
  assign n6935 = pi0299 & pi0960;
  assign n6936 = ~n6934 & ~n6935;
  assign n6937 = n6696 & ~n6936;
  assign n6938 = ~n6323 & ~n6937;
  assign n6939 = ~n2610 & n6937;
  assign n6940 = pi0299 & ~n6921;
  assign n6941 = ~n6923 & n6940;
  assign n6942 = pi0977 & n6720;
  assign n6943 = ~pi0299 & ~n6942;
  assign n6944 = ~pi0039 & ~n6941;
  assign n6945 = ~n6943 & n6944;
  assign n6946 = n2620 & n6945;
  assign n6947 = ~n6939 & ~n6946;
  assign n6948 = n2569 & n6947;
  assign n6949 = ~pi0054 & n6948;
  assign n6950 = pi0074 & ~n6938;
  assign n6951 = ~n6949 & n6950;
  assign n6952 = ~n2569 & ~n6937;
  assign n6953 = ~n6948 & ~n6952;
  assign n6954 = pi0054 & ~n6953;
  assign n6955 = ~pi0075 & n6947;
  assign n6956 = pi0075 & ~n6937;
  assign n6957 = pi0092 & ~n6956;
  assign n6958 = ~n6955 & n6957;
  assign n6959 = pi0075 & n6947;
  assign n6960 = pi0087 & n6937;
  assign n6961 = ~n2530 & n6937;
  assign n6962 = pi0960 & n6745;
  assign n6963 = n6940 & ~n6962;
  assign n6964 = pi0977 & n6752;
  assign n6965 = ~pi0299 & ~n6964;
  assign n6966 = n2530 & ~n6963;
  assign n6967 = ~n6965 & n6966;
  assign n6968 = pi0100 & ~n6961;
  assign n6969 = ~n6967 & n6968;
  assign n6970 = ~n6764 & n6934;
  assign n6971 = ~n6761 & n6935;
  assign n6972 = ~n6970 & ~n6971;
  assign n6973 = n6767 & ~n6972;
  assign n6974 = pi0977 & n6775;
  assign n6975 = ~pi0299 & ~n6974;
  assign n6976 = n6778 & n6922;
  assign n6977 = n6940 & ~n6976;
  assign n6978 = ~n6781 & ~n6977;
  assign n6979 = n6786 & n6922;
  assign n6980 = ~n6921 & ~n6979;
  assign n6981 = n6416 & ~n6980;
  assign n6982 = ~n6978 & ~n6981;
  assign n6983 = pi0232 & ~n6975;
  assign n6984 = ~n6982 & n6983;
  assign n6985 = pi0977 & n6769;
  assign n6986 = ~pi0299 & ~n6985;
  assign n6987 = ~pi0232 & ~n6977;
  assign n6988 = ~n6986 & n6987;
  assign n6989 = ~n6984 & ~n6988;
  assign n6990 = ~pi0039 & ~n6989;
  assign n6991 = ~pi0038 & ~n6973;
  assign n6992 = ~n6990 & n6991;
  assign n6993 = pi0039 & n6937;
  assign n6994 = pi0038 & ~n6993;
  assign n6995 = ~n6945 & n6994;
  assign n6996 = ~n6992 & ~n6995;
  assign n6997 = ~pi0100 & ~n6996;
  assign n6998 = ~pi0087 & ~n6969;
  assign n6999 = ~n6997 & n6998;
  assign n7000 = ~pi0075 & ~n6960;
  assign n7001 = ~n6999 & n7000;
  assign n7002 = ~pi0092 & ~n6959;
  assign n7003 = ~n7001 & n7002;
  assign n7004 = ~pi0054 & ~n6958;
  assign n7005 = ~n7003 & n7004;
  assign n7006 = ~pi0074 & ~n6954;
  assign n7007 = ~n7005 & n7006;
  assign n7008 = ~pi0055 & ~n6951;
  assign n7009 = ~n7007 & n7008;
  assign n7010 = n2529 & ~n6933;
  assign n7011 = ~n7009 & n7010;
  assign n7012 = ~pi0059 & ~n6931;
  assign n7013 = ~n7011 & n7012;
  assign n7014 = ~pi0057 & ~n6930;
  assign n7015 = ~n7013 & n7014;
  assign po0175 = ~n6927 & ~n7015;
  assign n7017 = pi0963 & n6696;
  assign n7018 = ~pi0228 & pi0963;
  assign n7019 = n6222 & n7018;
  assign n7020 = n2572 & n7019;
  assign n7021 = n6305 & n7020;
  assign n7022 = ~n7017 & ~n7021;
  assign n7023 = pi0057 & ~n7022;
  assign n7024 = n6304 & n7020;
  assign n7025 = pi0059 & ~n7017;
  assign n7026 = ~n7024 & n7025;
  assign n7027 = ~n2529 & n7017;
  assign n7028 = pi0055 & ~n7017;
  assign n7029 = ~n7020 & n7028;
  assign n7030 = ~pi0299 & pi0969;
  assign n7031 = pi0299 & pi0963;
  assign n7032 = ~n7030 & ~n7031;
  assign n7033 = n6696 & ~n7032;
  assign n7034 = ~n6323 & ~n7033;
  assign n7035 = ~n2610 & n7033;
  assign n7036 = pi0299 & ~n7017;
  assign n7037 = ~n7019 & n7036;
  assign n7038 = pi0969 & n6720;
  assign n7039 = ~pi0299 & ~n7038;
  assign n7040 = ~pi0039 & ~n7037;
  assign n7041 = ~n7039 & n7040;
  assign n7042 = n2620 & n7041;
  assign n7043 = ~n7035 & ~n7042;
  assign n7044 = n2569 & n7043;
  assign n7045 = ~pi0054 & n7044;
  assign n7046 = pi0074 & ~n7034;
  assign n7047 = ~n7045 & n7046;
  assign n7048 = ~n2569 & ~n7033;
  assign n7049 = ~n7044 & ~n7048;
  assign n7050 = pi0054 & ~n7049;
  assign n7051 = ~pi0075 & n7043;
  assign n7052 = pi0075 & ~n7033;
  assign n7053 = pi0092 & ~n7052;
  assign n7054 = ~n7051 & n7053;
  assign n7055 = pi0075 & n7043;
  assign n7056 = pi0087 & n7033;
  assign n7057 = ~n2530 & n7033;
  assign n7058 = pi0963 & n6745;
  assign n7059 = n7036 & ~n7058;
  assign n7060 = pi0969 & n6752;
  assign n7061 = ~pi0299 & ~n7060;
  assign n7062 = n2530 & ~n7059;
  assign n7063 = ~n7061 & n7062;
  assign n7064 = pi0100 & ~n7057;
  assign n7065 = ~n7063 & n7064;
  assign n7066 = ~n6764 & n7030;
  assign n7067 = ~n6761 & n7031;
  assign n7068 = ~n7066 & ~n7067;
  assign n7069 = n6767 & ~n7068;
  assign n7070 = pi0969 & n6775;
  assign n7071 = ~pi0299 & ~n7070;
  assign n7072 = n6778 & n7018;
  assign n7073 = n7036 & ~n7072;
  assign n7074 = ~n6781 & ~n7073;
  assign n7075 = n6786 & n7018;
  assign n7076 = ~n7017 & ~n7075;
  assign n7077 = n6416 & ~n7076;
  assign n7078 = ~n7074 & ~n7077;
  assign n7079 = pi0232 & ~n7071;
  assign n7080 = ~n7078 & n7079;
  assign n7081 = pi0969 & n6769;
  assign n7082 = ~pi0299 & ~n7081;
  assign n7083 = ~pi0232 & ~n7073;
  assign n7084 = ~n7082 & n7083;
  assign n7085 = ~n7080 & ~n7084;
  assign n7086 = ~pi0039 & ~n7085;
  assign n7087 = ~pi0038 & ~n7069;
  assign n7088 = ~n7086 & n7087;
  assign n7089 = pi0039 & n7033;
  assign n7090 = pi0038 & ~n7089;
  assign n7091 = ~n7041 & n7090;
  assign n7092 = ~n7088 & ~n7091;
  assign n7093 = ~pi0100 & ~n7092;
  assign n7094 = ~pi0087 & ~n7065;
  assign n7095 = ~n7093 & n7094;
  assign n7096 = ~pi0075 & ~n7056;
  assign n7097 = ~n7095 & n7096;
  assign n7098 = ~pi0092 & ~n7055;
  assign n7099 = ~n7097 & n7098;
  assign n7100 = ~pi0054 & ~n7054;
  assign n7101 = ~n7099 & n7100;
  assign n7102 = ~pi0074 & ~n7050;
  assign n7103 = ~n7101 & n7102;
  assign n7104 = ~pi0055 & ~n7047;
  assign n7105 = ~n7103 & n7104;
  assign n7106 = n2529 & ~n7029;
  assign n7107 = ~n7105 & n7106;
  assign n7108 = ~pi0059 & ~n7027;
  assign n7109 = ~n7107 & n7108;
  assign n7110 = ~pi0057 & ~n7026;
  assign n7111 = ~n7109 & n7110;
  assign po0176 = ~n7023 & ~n7111;
  assign n7113 = pi0975 & n6696;
  assign n7114 = ~pi0228 & pi0975;
  assign n7115 = n6222 & n7114;
  assign n7116 = n2572 & n7115;
  assign n7117 = n6305 & n7116;
  assign n7118 = ~n7113 & ~n7117;
  assign n7119 = pi0057 & ~n7118;
  assign n7120 = n6304 & n7116;
  assign n7121 = pi0059 & ~n7113;
  assign n7122 = ~n7120 & n7121;
  assign n7123 = ~n2529 & n7113;
  assign n7124 = pi0055 & ~n7113;
  assign n7125 = ~n7116 & n7124;
  assign n7126 = ~pi0299 & pi0971;
  assign n7127 = pi0299 & pi0975;
  assign n7128 = ~n7126 & ~n7127;
  assign n7129 = n6696 & ~n7128;
  assign n7130 = ~n6323 & ~n7129;
  assign n7131 = ~n2610 & n7129;
  assign n7132 = pi0299 & ~n7113;
  assign n7133 = ~n7115 & n7132;
  assign n7134 = pi0971 & n6720;
  assign n7135 = ~pi0299 & ~n7134;
  assign n7136 = ~pi0039 & ~n7133;
  assign n7137 = ~n7135 & n7136;
  assign n7138 = n2620 & n7137;
  assign n7139 = ~n7131 & ~n7138;
  assign n7140 = n2569 & n7139;
  assign n7141 = ~pi0054 & n7140;
  assign n7142 = pi0074 & ~n7130;
  assign n7143 = ~n7141 & n7142;
  assign n7144 = ~n2569 & ~n7129;
  assign n7145 = ~n7140 & ~n7144;
  assign n7146 = pi0054 & ~n7145;
  assign n7147 = ~pi0075 & n7139;
  assign n7148 = pi0075 & ~n7129;
  assign n7149 = pi0092 & ~n7148;
  assign n7150 = ~n7147 & n7149;
  assign n7151 = pi0075 & n7139;
  assign n7152 = pi0087 & n7129;
  assign n7153 = ~n2530 & n7129;
  assign n7154 = pi0975 & n6745;
  assign n7155 = n7132 & ~n7154;
  assign n7156 = pi0971 & n6752;
  assign n7157 = ~pi0299 & ~n7156;
  assign n7158 = n2530 & ~n7155;
  assign n7159 = ~n7157 & n7158;
  assign n7160 = pi0100 & ~n7153;
  assign n7161 = ~n7159 & n7160;
  assign n7162 = ~n6764 & n7126;
  assign n7163 = ~n6761 & n7127;
  assign n7164 = ~n7162 & ~n7163;
  assign n7165 = n6767 & ~n7164;
  assign n7166 = pi0971 & n6775;
  assign n7167 = ~pi0299 & ~n7166;
  assign n7168 = n6778 & n7114;
  assign n7169 = n7132 & ~n7168;
  assign n7170 = ~n6781 & ~n7169;
  assign n7171 = n6786 & n7114;
  assign n7172 = ~n7113 & ~n7171;
  assign n7173 = n6416 & ~n7172;
  assign n7174 = ~n7170 & ~n7173;
  assign n7175 = pi0232 & ~n7167;
  assign n7176 = ~n7174 & n7175;
  assign n7177 = pi0971 & n6769;
  assign n7178 = ~pi0299 & ~n7177;
  assign n7179 = ~pi0232 & ~n7169;
  assign n7180 = ~n7178 & n7179;
  assign n7181 = ~n7176 & ~n7180;
  assign n7182 = ~pi0039 & ~n7181;
  assign n7183 = ~pi0038 & ~n7165;
  assign n7184 = ~n7182 & n7183;
  assign n7185 = pi0039 & n7129;
  assign n7186 = pi0038 & ~n7185;
  assign n7187 = ~n7137 & n7186;
  assign n7188 = ~n7184 & ~n7187;
  assign n7189 = ~pi0100 & ~n7188;
  assign n7190 = ~pi0087 & ~n7161;
  assign n7191 = ~n7189 & n7190;
  assign n7192 = ~pi0075 & ~n7152;
  assign n7193 = ~n7191 & n7192;
  assign n7194 = ~pi0092 & ~n7151;
  assign n7195 = ~n7193 & n7194;
  assign n7196 = ~pi0054 & ~n7150;
  assign n7197 = ~n7195 & n7196;
  assign n7198 = ~pi0074 & ~n7146;
  assign n7199 = ~n7197 & n7198;
  assign n7200 = ~pi0055 & ~n7143;
  assign n7201 = ~n7199 & n7200;
  assign n7202 = n2529 & ~n7125;
  assign n7203 = ~n7201 & n7202;
  assign n7204 = ~pi0059 & ~n7123;
  assign n7205 = ~n7203 & n7204;
  assign n7206 = ~pi0057 & ~n7122;
  assign n7207 = ~n7205 & n7206;
  assign po0177 = ~n7119 & ~n7207;
  assign n7209 = pi0978 & n6696;
  assign n7210 = ~pi0228 & pi0978;
  assign n7211 = n2572 & n7210;
  assign n7212 = n6222 & n7211;
  assign n7213 = n6305 & n7212;
  assign n7214 = ~n7209 & ~n7213;
  assign n7215 = pi0057 & ~n7214;
  assign n7216 = n6304 & n7212;
  assign n7217 = pi0059 & ~n7209;
  assign n7218 = ~n7216 & n7217;
  assign n7219 = ~n2529 & n7209;
  assign n7220 = pi0055 & ~n7209;
  assign n7221 = ~n7212 & n7220;
  assign n7222 = ~pi0299 & pi0974;
  assign n7223 = pi0299 & pi0978;
  assign n7224 = ~n7222 & ~n7223;
  assign n7225 = n6696 & ~n7224;
  assign n7226 = ~n6323 & ~n7225;
  assign n7227 = n6720 & ~n7224;
  assign n7228 = ~pi0228 & ~n2610;
  assign n7229 = n7227 & ~n7228;
  assign n7230 = n2569 & ~n7229;
  assign n7231 = ~pi0054 & n7230;
  assign n7232 = pi0074 & ~n7226;
  assign n7233 = ~n7231 & n7232;
  assign n7234 = ~n2569 & ~n7225;
  assign n7235 = ~n7230 & ~n7234;
  assign n7236 = pi0054 & ~n7235;
  assign n7237 = ~pi0075 & ~n7229;
  assign n7238 = pi0075 & ~n7225;
  assign n7239 = pi0092 & ~n7238;
  assign n7240 = ~n7237 & n7239;
  assign n7241 = pi0075 & ~n7229;
  assign n7242 = pi0087 & n7225;
  assign n7243 = ~n2530 & n7225;
  assign n7244 = pi0299 & ~n7209;
  assign n7245 = pi0978 & n6745;
  assign n7246 = n7244 & ~n7245;
  assign n7247 = pi0974 & n6752;
  assign n7248 = ~pi0299 & ~n7247;
  assign n7249 = n2530 & ~n7246;
  assign n7250 = ~n7248 & n7249;
  assign n7251 = pi0100 & ~n7243;
  assign n7252 = ~n7250 & n7251;
  assign n7253 = pi0039 & n7225;
  assign n7254 = ~pi0039 & n7227;
  assign n7255 = pi0038 & ~n7253;
  assign n7256 = ~n7254 & n7255;
  assign n7257 = ~n6764 & n7222;
  assign n7258 = ~n6761 & n7223;
  assign n7259 = ~n7257 & ~n7258;
  assign n7260 = n6767 & ~n7259;
  assign n7261 = pi0974 & n6775;
  assign n7262 = ~pi0299 & ~n7261;
  assign n7263 = n6778 & n7210;
  assign n7264 = n7244 & ~n7263;
  assign n7265 = ~n6781 & ~n7264;
  assign n7266 = n6786 & n7210;
  assign n7267 = ~n7209 & ~n7266;
  assign n7268 = n6416 & ~n7267;
  assign n7269 = ~n7265 & ~n7268;
  assign n7270 = pi0232 & ~n7262;
  assign n7271 = ~n7269 & n7270;
  assign n7272 = pi0974 & n6769;
  assign n7273 = ~pi0299 & ~n7272;
  assign n7274 = ~pi0232 & ~n7264;
  assign n7275 = ~n7273 & n7274;
  assign n7276 = ~n7271 & ~n7275;
  assign n7277 = ~pi0039 & ~n7276;
  assign n7278 = ~pi0038 & ~n7260;
  assign n7279 = ~n7277 & n7278;
  assign n7280 = ~n7256 & ~n7279;
  assign n7281 = ~pi0100 & ~n7280;
  assign n7282 = ~pi0087 & ~n7252;
  assign n7283 = ~n7281 & n7282;
  assign n7284 = ~pi0075 & ~n7242;
  assign n7285 = ~n7283 & n7284;
  assign n7286 = ~pi0092 & ~n7241;
  assign n7287 = ~n7285 & n7286;
  assign n7288 = ~pi0054 & ~n7240;
  assign n7289 = ~n7287 & n7288;
  assign n7290 = ~pi0074 & ~n7236;
  assign n7291 = ~n7289 & n7290;
  assign n7292 = ~pi0055 & ~n7233;
  assign n7293 = ~n7291 & n7292;
  assign n7294 = n2529 & ~n7221;
  assign n7295 = ~n7293 & n7294;
  assign n7296 = ~pi0059 & ~n7219;
  assign n7297 = ~n7295 & n7296;
  assign n7298 = ~pi0057 & ~n7218;
  assign n7299 = ~n7297 & n7298;
  assign po0178 = ~n7215 & ~n7299;
  assign n7301 = n2620 & n6284;
  assign n7302 = pi0075 & ~n7301;
  assign n7303 = n2533 & n2608;
  assign n7304 = n6284 & n7303;
  assign n7305 = pi0092 & ~n7304;
  assign n7306 = ~n7302 & ~n7305;
  assign n7307 = pi0299 & ~n6244;
  assign n7308 = n6759 & n7307;
  assign n7309 = ~pi0299 & ~n6207;
  assign n7310 = n6409 & n7309;
  assign n7311 = pi0039 & ~n7310;
  assign n7312 = ~n7308 & n7311;
  assign n7313 = pi0299 & n6489;
  assign n7314 = ~pi0299 & n6520;
  assign n7315 = ~pi0232 & ~n7313;
  assign n7316 = ~n7314 & n7315;
  assign n7317 = n6527 & n6532;
  assign n7318 = ~pi0299 & ~n6530;
  assign n7319 = ~n6771 & n7318;
  assign n7320 = ~n7317 & n7319;
  assign n7321 = ~n6416 & n7313;
  assign n7322 = ~n6490 & n6781;
  assign n7323 = ~n6785 & n7322;
  assign n7324 = pi0232 & ~n7321;
  assign n7325 = ~n7320 & n7324;
  assign n7326 = ~n7323 & n7325;
  assign n7327 = ~pi0039 & ~n7316;
  assign n7328 = ~n7326 & n7327;
  assign n7329 = ~n7312 & ~n7328;
  assign n7330 = ~pi0038 & ~n7329;
  assign n7331 = ~n6136 & ~n7330;
  assign n7332 = ~pi0100 & ~n7331;
  assign n7333 = ~pi0038 & n6284;
  assign n7334 = pi0100 & ~n7333;
  assign n7335 = n6289 & ~n7334;
  assign n7336 = ~n7332 & n7335;
  assign n7337 = n2569 & ~n7336;
  assign n7338 = n7306 & ~n7337;
  assign n7339 = ~pi0054 & ~n7338;
  assign n7340 = ~pi0092 & n7304;
  assign n7341 = pi0054 & ~n7340;
  assign n7342 = ~n7339 & ~n7341;
  assign n7343 = ~pi0074 & ~n7342;
  assign n7344 = ~n6130 & ~n7343;
  assign n7345 = ~pi0055 & ~n7344;
  assign n7346 = n2535 & n6125;
  assign n7347 = pi0055 & ~n7346;
  assign n7348 = ~pi0056 & ~n7347;
  assign n7349 = ~pi0062 & n7348;
  assign n7350 = ~n7345 & n7349;
  assign n7351 = n3328 & ~n7350;
  assign po0195 = n6123 & ~n7351;
  assign n7353 = ~pi0954 & ~po0195;
  assign n7354 = pi0024 & pi0954;
  assign po0182 = ~n7353 & ~n7354;
  assign n7356 = n2531 & n3335;
  assign n7357 = n3330 & n7356;
  assign n7358 = ~n2441 & ~n7357;
  assign n7359 = pi0062 & ~n7358;
  assign n7360 = n2537 & n3335;
  assign n7361 = pi0056 & ~n2441;
  assign n7362 = ~n7360 & n7361;
  assign n7363 = n2531 & n6128;
  assign n7364 = n3335 & n7363;
  assign n7365 = ~pi0074 & n7364;
  assign n7366 = ~n2441 & ~n7365;
  assign n7367 = pi0055 & ~n7366;
  assign n7368 = ~n2441 & ~n2532;
  assign n7369 = n3335 & n3373;
  assign n7370 = ~n2441 & ~n7369;
  assign n7371 = pi0092 & ~n7370;
  assign n7372 = pi0075 & ~n2441;
  assign n7373 = ~n2441 & ~n7356;
  assign n7374 = pi0087 & ~n7373;
  assign n7375 = ~pi0100 & n4730;
  assign n7376 = n2521 & ~n6356;
  assign n7377 = ~pi0299 & ~n7376;
  assign n7378 = pi0299 & ~n3394;
  assign n7379 = ~n7377 & ~n7378;
  assign n7380 = pi0100 & n3335;
  assign n7381 = n7379 & n7380;
  assign n7382 = ~pi0039 & ~n7381;
  assign n7383 = ~n7375 & n7382;
  assign n7384 = ~pi0100 & n3335;
  assign n7385 = pi0039 & ~n7384;
  assign n7386 = ~pi0038 & ~n7385;
  assign n7387 = ~n7383 & n7386;
  assign n7388 = ~n2441 & ~n7387;
  assign n7389 = ~pi0087 & ~n7388;
  assign n7390 = ~pi0075 & ~n7374;
  assign n7391 = ~n7389 & n7390;
  assign n7392 = ~pi0092 & ~n7372;
  assign n7393 = ~n7391 & n7392;
  assign n7394 = n2532 & ~n7371;
  assign n7395 = ~n7393 & n7394;
  assign n7396 = ~pi0055 & ~n7368;
  assign n7397 = ~n7395 & n7396;
  assign n7398 = ~pi0056 & ~n7367;
  assign n7399 = ~n7397 & n7398;
  assign n7400 = ~pi0062 & ~n7362;
  assign n7401 = ~n7399 & n7400;
  assign n7402 = ~n7359 & ~n7401;
  assign n7403 = n3328 & ~n7402;
  assign n7404 = n2441 & ~n3328;
  assign po0183 = n7403 | n7404;
  assign n7406 = pi0119 & pi1056;
  assign n7407 = ~pi0228 & pi0252;
  assign n7408 = ~pi0119 & ~n7407;
  assign n7409 = ~pi0468 & ~n7408;
  assign po0184 = n7406 | ~n7409;
  assign n7411 = pi0119 & pi1077;
  assign po0185 = ~n7409 | n7411;
  assign n7413 = pi0119 & pi1073;
  assign po0186 = ~n7409 | n7413;
  assign n7415 = pi0119 & pi1041;
  assign po0187 = ~n7409 | n7415;
  assign n7417 = pi0824 & n2932;
  assign n7418 = ~pi0122 & pi1093;
  assign n7419 = n7417 & n7418;
  assign n7420 = ~pi1091 & n7419;
  assign n7421 = ~pi0098 & n7420;
  assign n7422 = pi0567 & n7421;
  assign n7423 = ~pi0285 & ~pi0286;
  assign n7424 = ~pi0289 & n7423;
  assign n7425 = ~pi0288 & n7424;
  assign po1038 = pi0057 | ~n6305;
  assign n7427 = ~n7425 & po1038;
  assign n7428 = n7422 & n7427;
  assign n7429 = ~pi0074 & n6134;
  assign n7430 = ~pi0122 & pi0829;
  assign n7431 = n2961 & ~n6157;
  assign n7432 = ~pi0841 & n2703;
  assign n7433 = pi0090 & n7432;
  assign n7434 = ~pi0093 & ~n7433;
  assign n7435 = n7431 & ~n7434;
  assign n7436 = ~pi0051 & ~n7435;
  assign n7437 = ~pi0088 & pi0098;
  assign n7438 = ~pi0050 & ~pi0077;
  assign n7439 = ~pi0094 & n7438;
  assign n7440 = n2767 & n7439;
  assign n7441 = n2495 & n7437;
  assign n7442 = n7440 & n7441;
  assign n7443 = ~pi0097 & ~n7442;
  assign n7444 = n2717 & ~n7443;
  assign n7445 = ~pi0035 & n2704;
  assign n7446 = ~pi0070 & n7445;
  assign n7447 = n7444 & n7446;
  assign n7448 = n7436 & ~n7447;
  assign n7449 = ~n2747 & ~n7448;
  assign n7450 = ~pi0096 & n2519;
  assign n7451 = n7449 & n7450;
  assign n7452 = n6277 & n7451;
  assign n7453 = ~n7430 & n7452;
  assign n7454 = ~pi0096 & ~n7449;
  assign n7455 = pi0096 & ~n6484;
  assign n7456 = n2519 & ~n7455;
  assign n7457 = n2932 & n7430;
  assign n7458 = n7456 & n7457;
  assign n7459 = ~n7454 & n7458;
  assign n7460 = ~n7453 & ~n7459;
  assign n7461 = ~pi1093 & ~n7460;
  assign n7462 = ~pi0087 & ~n7461;
  assign n7463 = n2521 & po0740;
  assign n7464 = pi0087 & ~n7463;
  assign n7465 = ~pi0075 & n2531;
  assign n7466 = ~n7464 & n7465;
  assign n7467 = ~n7462 & n7466;
  assign n7468 = ~pi0567 & ~n7467;
  assign n7469 = n7429 & ~n7468;
  assign n7470 = ~pi0299 & ~n2669;
  assign n7471 = pi0299 & ~n2639;
  assign n7472 = ~n7470 & ~n7471;
  assign n7473 = pi0232 & n6197;
  assign n7474 = n7472 & n7473;
  assign n7475 = n2610 & ~n7474;
  assign n7476 = n7421 & ~n7475;
  assign n7477 = ~pi0024 & n6359;
  assign n7478 = ~n2923 & po1057;
  assign n7479 = pi1093 & n7457;
  assign n7480 = n7478 & n7479;
  assign n7481 = n7477 & n7480;
  assign n7482 = pi1091 & ~n7481;
  assign n7483 = n7475 & ~n7482;
  assign n7484 = ~pi0098 & n7417;
  assign n7485 = n7418 & n7484;
  assign n7486 = ~pi1091 & ~n7485;
  assign n7487 = n7483 & ~n7486;
  assign n7488 = pi0075 & ~n7476;
  assign n7489 = ~n7487 & n7488;
  assign n7490 = pi1093 & n2923;
  assign n7491 = n6277 & ~n7490;
  assign n7492 = n2521 & n7491;
  assign n7493 = pi1091 & ~n7492;
  assign n7494 = ~pi1091 & ~n7463;
  assign n7495 = n2521 & n7417;
  assign n7496 = pi0122 & n7495;
  assign n7497 = ~pi0122 & n7484;
  assign n7498 = ~n7496 & ~n7497;
  assign n7499 = pi1093 & ~n7498;
  assign n7500 = n7494 & ~n7499;
  assign n7501 = n2625 & ~n7493;
  assign n7502 = ~n7500 & n7501;
  assign n7503 = ~n7421 & ~n7502;
  assign n7504 = pi0087 & ~n7503;
  assign n7505 = ~n2530 & n7421;
  assign n7506 = pi0228 & ~n7474;
  assign n7507 = ~n7421 & ~n7506;
  assign n7508 = n2521 & n7480;
  assign n7509 = pi1091 & ~n7508;
  assign n7510 = ~n7486 & ~n7509;
  assign n7511 = n7506 & ~n7510;
  assign n7512 = n2530 & ~n7507;
  assign n7513 = ~n7511 & n7512;
  assign n7514 = pi0100 & ~n7505;
  assign n7515 = ~n7513 & n7514;
  assign n7516 = pi0038 & n7421;
  assign n7517 = pi1093 & ~n2923;
  assign n7518 = ~n2747 & n7450;
  assign n7519 = ~n7436 & n7518;
  assign n7520 = n7417 & n7519;
  assign n7521 = ~pi0829 & n7520;
  assign n7522 = ~pi0024 & n2756;
  assign n7523 = ~pi0046 & pi0097;
  assign n7524 = ~pi0108 & n7523;
  assign n7525 = n6491 & n7524;
  assign n7526 = n2772 & n7525;
  assign n7527 = ~pi0091 & n7526;
  assign n7528 = ~n7522 & ~n7527;
  assign n7529 = n2461 & n7431;
  assign n7530 = ~n7528 & n7529;
  assign n7531 = n7436 & ~n7530;
  assign n7532 = ~n2747 & ~n7531;
  assign n7533 = ~pi0096 & ~n7532;
  assign n7534 = n2933 & n7456;
  assign n7535 = ~n7533 & n7534;
  assign n7536 = ~n7521 & ~n7535;
  assign n7537 = ~pi0122 & ~n7536;
  assign n7538 = pi0122 & n6277;
  assign n7539 = n7519 & n7538;
  assign n7540 = ~n7537 & ~n7539;
  assign n7541 = n7517 & ~n7540;
  assign n7542 = pi1091 & ~n7541;
  assign n7543 = ~n7461 & n7542;
  assign n7544 = ~pi0039 & ~n7543;
  assign n7545 = ~pi1091 & ~n7461;
  assign n7546 = pi0122 & n7520;
  assign n7547 = ~n7497 & ~n7546;
  assign n7548 = pi1093 & ~n7547;
  assign n7549 = n7545 & ~n7548;
  assign n7550 = n7544 & ~n7549;
  assign n7551 = ~pi0223 & n5810;
  assign n7552 = n7421 & ~n7551;
  assign n7553 = ~n2923 & n2925;
  assign n7554 = n6382 & n7553;
  assign n7555 = n2926 & n7554;
  assign n7556 = pi1091 & ~n7555;
  assign n7557 = ~n7486 & ~n7556;
  assign n7558 = n6198 & n7557;
  assign n7559 = ~n6198 & n7421;
  assign n7560 = ~n7558 & ~n7559;
  assign n7561 = n6205 & n7560;
  assign n7562 = ~n6227 & n7557;
  assign n7563 = n6227 & n7421;
  assign n7564 = ~n7562 & ~n7563;
  assign n7565 = ~n6205 & n7564;
  assign n7566 = n7551 & ~n7561;
  assign n7567 = ~n7565 & n7566;
  assign n7568 = ~pi0299 & ~n7552;
  assign n7569 = ~n7567 & n7568;
  assign n7570 = ~pi0216 & n6379;
  assign n7571 = n7421 & ~n7570;
  assign n7572 = n6242 & n7560;
  assign n7573 = ~n6242 & n7564;
  assign n7574 = n7570 & ~n7572;
  assign n7575 = ~n7573 & n7574;
  assign n7576 = pi0299 & ~n7571;
  assign n7577 = ~n7575 & n7576;
  assign n7578 = pi0039 & ~n7569;
  assign n7579 = ~n7577 & n7578;
  assign n7580 = ~n7550 & ~n7579;
  assign n7581 = ~pi0038 & ~n7580;
  assign n7582 = ~pi0100 & ~n7516;
  assign n7583 = ~n7581 & n7582;
  assign n7584 = ~pi0087 & ~n7515;
  assign n7585 = ~n7583 & n7584;
  assign n7586 = ~pi0075 & ~n7504;
  assign n7587 = ~n7585 & n7586;
  assign n7588 = ~n7489 & ~n7587;
  assign n7589 = pi0567 & ~n7588;
  assign n7590 = n7469 & ~n7589;
  assign n7591 = n7422 & ~n7429;
  assign n7592 = ~n7590 & ~n7591;
  assign n7593 = ~n7425 & n7592;
  assign n7594 = pi1091 & n7478;
  assign n7595 = n7457 & n7594;
  assign n7596 = n7477 & n7595;
  assign n7597 = pi1093 & n7596;
  assign n7598 = n7475 & n7597;
  assign n7599 = pi0075 & ~n7598;
  assign n7600 = ~n7543 & ~n7545;
  assign n7601 = ~pi0039 & ~n7600;
  assign n7602 = pi1091 & n7555;
  assign n7603 = ~n6244 & n7602;
  assign n7604 = ~pi0216 & n6640;
  assign n7605 = n7603 & n7604;
  assign n7606 = ~n6207 & n7602;
  assign n7607 = ~pi0299 & n6405;
  assign n7608 = ~pi0224 & n7607;
  assign n7609 = n7606 & n7608;
  assign n7610 = pi0039 & ~n7605;
  assign n7611 = ~n7609 & n7610;
  assign n7612 = ~pi0038 & ~n7611;
  assign n7613 = ~n7601 & n7612;
  assign n7614 = ~pi0100 & ~n7613;
  assign n7615 = n6384 & n7519;
  assign n7616 = n7612 & n7615;
  assign n7617 = ~n7542 & n7616;
  assign n7618 = n7614 & ~n7617;
  assign n7619 = pi1091 & n7508;
  assign n7620 = pi0228 & n7619;
  assign n7621 = n2530 & ~n7474;
  assign n7622 = n7620 & n7621;
  assign n7623 = pi0100 & ~n7622;
  assign n7624 = ~n7618 & ~n7623;
  assign n7625 = ~pi0087 & ~n7624;
  assign n7626 = ~pi1091 & pi1093;
  assign n7627 = ~n7495 & n7626;
  assign n7628 = ~n7492 & ~n7626;
  assign n7629 = n2625 & ~n7628;
  assign n7630 = ~n7627 & n7629;
  assign n7631 = pi0087 & ~n7630;
  assign n7632 = ~n7625 & ~n7631;
  assign n7633 = ~pi0075 & ~n7632;
  assign n7634 = ~n7599 & ~n7633;
  assign n7635 = pi0567 & ~n7634;
  assign n7636 = n7469 & ~n7635;
  assign n7637 = n7425 & ~n7636;
  assign n7638 = ~po1038 & ~n7593;
  assign n7639 = ~n7637 & n7638;
  assign n7640 = pi0217 & ~n7428;
  assign n7641 = ~n7639 & n7640;
  assign n7642 = ~pi1161 & ~pi1162;
  assign n7643 = ~pi1163 & n7642;
  assign n7644 = ~pi0592 & n7422;
  assign n7645 = pi0592 & n7422;
  assign n7646 = ~pi0363 & ~pi0372;
  assign n7647 = pi0363 & pi0372;
  assign n7648 = ~n7646 & ~n7647;
  assign n7649 = pi0386 & ~n7648;
  assign n7650 = ~pi0386 & n7648;
  assign n7651 = ~n7649 & ~n7650;
  assign n7652 = pi0338 & ~pi0388;
  assign n7653 = ~pi0338 & pi0388;
  assign n7654 = ~n7652 & ~n7653;
  assign n7655 = pi0337 & ~pi0339;
  assign n7656 = ~pi0337 & pi0339;
  assign n7657 = ~n7655 & ~n7656;
  assign n7658 = pi0387 & n7657;
  assign n7659 = ~pi0387 & ~n7657;
  assign n7660 = ~n7658 & ~n7659;
  assign n7661 = pi0380 & ~n7660;
  assign n7662 = ~pi0380 & n7660;
  assign n7663 = ~n7661 & ~n7662;
  assign n7664 = n7654 & ~n7663;
  assign n7665 = ~n7654 & n7663;
  assign n7666 = ~n7664 & ~n7665;
  assign n7667 = n7651 & n7666;
  assign n7668 = ~n7651 & ~n7666;
  assign n7669 = ~n7667 & ~n7668;
  assign n7670 = pi1196 & ~n7669;
  assign n7671 = ~pi0368 & ~pi0389;
  assign n7672 = pi0368 & pi0389;
  assign n7673 = ~n7671 & ~n7672;
  assign n7674 = pi0365 & ~pi0447;
  assign n7675 = ~pi0365 & pi0447;
  assign n7676 = ~n7674 & ~n7675;
  assign n7677 = pi0336 & ~pi0383;
  assign n7678 = ~pi0336 & pi0383;
  assign n7679 = ~n7677 & ~n7678;
  assign n7680 = pi0364 & ~pi0366;
  assign n7681 = ~pi0364 & pi0366;
  assign n7682 = ~n7680 & ~n7681;
  assign n7683 = n7679 & n7682;
  assign n7684 = ~n7679 & ~n7682;
  assign n7685 = ~n7683 & ~n7684;
  assign n7686 = n7676 & n7685;
  assign n7687 = ~n7676 & ~n7685;
  assign n7688 = ~n7686 & ~n7687;
  assign n7689 = pi0367 & ~n7688;
  assign n7690 = ~pi0367 & n7688;
  assign n7691 = ~n7689 & ~n7690;
  assign n7692 = n7673 & n7691;
  assign n7693 = ~n7673 & ~n7691;
  assign n7694 = pi1197 & ~n7692;
  assign n7695 = ~n7693 & n7694;
  assign n7696 = ~n7670 & ~n7695;
  assign n7697 = pi0592 & ~n7696;
  assign n7698 = pi0379 & ~pi0382;
  assign n7699 = ~pi0379 & pi0382;
  assign n7700 = ~n7698 & ~n7699;
  assign n7701 = pi0376 & ~pi0439;
  assign n7702 = ~pi0376 & pi0439;
  assign n7703 = ~n7701 & ~n7702;
  assign n7704 = pi0381 & n7703;
  assign n7705 = ~pi0381 & ~n7703;
  assign n7706 = ~n7704 & ~n7705;
  assign n7707 = pi0317 & ~pi0385;
  assign n7708 = ~pi0317 & pi0385;
  assign n7709 = ~n7707 & ~n7708;
  assign n7710 = pi0378 & n7709;
  assign n7711 = ~pi0378 & ~n7709;
  assign n7712 = ~n7710 & ~n7711;
  assign n7713 = n7706 & ~n7712;
  assign n7714 = ~n7706 & n7712;
  assign n7715 = ~n7713 & ~n7714;
  assign n7716 = n7700 & n7715;
  assign n7717 = ~n7700 & ~n7715;
  assign n7718 = ~n7716 & ~n7717;
  assign n7719 = ~pi0377 & ~n7718;
  assign n7720 = pi0377 & n7718;
  assign n7721 = ~n7719 & ~n7720;
  assign n7722 = n7696 & ~n7721;
  assign n7723 = pi0592 & ~n7722;
  assign n7724 = n7422 & ~n7723;
  assign n7725 = pi1199 & ~n7724;
  assign n7726 = ~n7697 & ~n7725;
  assign n7727 = n7645 & n7726;
  assign n7728 = ~pi1198 & n7727;
  assign n7729 = pi0384 & ~pi0442;
  assign n7730 = ~pi0384 & pi0442;
  assign n7731 = ~n7729 & ~n7730;
  assign n7732 = pi0440 & ~n7731;
  assign n7733 = ~pi0440 & n7731;
  assign n7734 = ~n7732 & ~n7733;
  assign n7735 = ~pi0369 & ~pi0374;
  assign n7736 = pi0369 & pi0374;
  assign n7737 = ~n7735 & ~n7736;
  assign n7738 = ~pi0370 & ~n7737;
  assign n7739 = pi0370 & n7737;
  assign n7740 = ~n7738 & ~n7739;
  assign n7741 = ~pi0371 & ~n7740;
  assign n7742 = pi0371 & n7740;
  assign n7743 = ~n7741 & ~n7742;
  assign n7744 = ~pi0373 & ~n7743;
  assign n7745 = pi0373 & n7743;
  assign n7746 = ~n7744 & ~n7745;
  assign n7747 = pi0375 & ~n7746;
  assign n7748 = ~pi0375 & n7746;
  assign n7749 = ~n7747 & ~n7748;
  assign n7750 = ~n7734 & ~n7749;
  assign n7751 = n7734 & n7749;
  assign n7752 = ~n7750 & ~n7751;
  assign n7753 = n7727 & n7752;
  assign n7754 = ~n7644 & ~n7728;
  assign n7755 = ~n7753 & n7754;
  assign n7756 = ~pi0590 & ~n7755;
  assign n7757 = pi0351 & pi1199;
  assign n7758 = pi0345 & ~pi0346;
  assign n7759 = ~pi0345 & pi0346;
  assign n7760 = ~n7758 & ~n7759;
  assign n7761 = pi0323 & ~n7760;
  assign n7762 = ~pi0323 & n7760;
  assign n7763 = ~n7761 & ~n7762;
  assign n7764 = pi0358 & ~pi0450;
  assign n7765 = ~pi0358 & pi0450;
  assign n7766 = ~n7764 & ~n7765;
  assign n7767 = n7763 & ~n7766;
  assign n7768 = ~n7763 & n7766;
  assign n7769 = ~n7767 & ~n7768;
  assign n7770 = ~pi0327 & ~pi0362;
  assign n7771 = pi0327 & pi0362;
  assign n7772 = ~n7770 & ~n7771;
  assign n7773 = pi0343 & ~pi0344;
  assign n7774 = ~pi0343 & pi0344;
  assign n7775 = ~n7773 & ~n7774;
  assign n7776 = n7772 & ~n7775;
  assign n7777 = ~n7772 & n7775;
  assign n7778 = ~n7776 & ~n7777;
  assign n7779 = n7769 & n7778;
  assign n7780 = ~n7769 & ~n7778;
  assign n7781 = pi1197 & ~n7779;
  assign n7782 = ~n7780 & n7781;
  assign n7783 = pi0320 & ~pi0460;
  assign n7784 = ~pi0320 & pi0460;
  assign n7785 = ~n7783 & ~n7784;
  assign n7786 = pi0342 & ~n7785;
  assign n7787 = ~pi0342 & n7785;
  assign n7788 = ~n7786 & ~n7787;
  assign n7789 = pi0452 & ~pi0455;
  assign n7790 = ~pi0452 & pi0455;
  assign n7791 = ~n7789 & ~n7790;
  assign n7792 = pi0355 & n7791;
  assign n7793 = ~pi0355 & ~n7791;
  assign n7794 = ~n7792 & ~n7793;
  assign n7795 = pi0361 & ~pi0458;
  assign n7796 = ~pi0361 & pi0458;
  assign n7797 = ~n7795 & ~n7796;
  assign n7798 = n7794 & n7797;
  assign n7799 = ~n7794 & ~n7797;
  assign n7800 = ~n7798 & ~n7799;
  assign n7801 = ~pi0441 & n7800;
  assign n7802 = pi0441 & ~n7800;
  assign n7803 = ~pi0592 & ~n7801;
  assign n7804 = ~n7802 & n7803;
  assign n7805 = n7422 & n7788;
  assign n7806 = ~n7804 & n7805;
  assign n7807 = pi0361 & ~pi0441;
  assign n7808 = ~pi0361 & pi0441;
  assign n7809 = ~n7807 & ~n7808;
  assign n7810 = n7788 & n7809;
  assign n7811 = ~n7788 & ~n7809;
  assign n7812 = ~n7810 & ~n7811;
  assign n7813 = pi0458 & n7812;
  assign n7814 = ~pi0458 & ~n7812;
  assign n7815 = ~n7813 & ~n7814;
  assign n7816 = n7794 & n7815;
  assign n7817 = ~n7794 & ~n7815;
  assign n7818 = ~n7816 & ~n7817;
  assign n7819 = ~pi0592 & n7818;
  assign n7820 = n7422 & ~n7788;
  assign n7821 = ~n7819 & n7820;
  assign n7822 = pi1196 & ~n7806;
  assign n7823 = ~n7821 & n7822;
  assign n7824 = ~pi1198 & ~n7823;
  assign n7825 = pi1196 & n7818;
  assign n7826 = pi0321 & ~pi0347;
  assign n7827 = ~pi0321 & pi0347;
  assign n7828 = ~n7826 & ~n7827;
  assign n7829 = pi0316 & ~pi0349;
  assign n7830 = ~pi0316 & pi0349;
  assign n7831 = ~n7829 & ~n7830;
  assign n7832 = pi0348 & n7831;
  assign n7833 = ~pi0348 & ~n7831;
  assign n7834 = ~n7832 & ~n7833;
  assign n7835 = pi0315 & ~pi0359;
  assign n7836 = ~pi0315 & pi0359;
  assign n7837 = ~n7835 & ~n7836;
  assign n7838 = pi0322 & n7837;
  assign n7839 = ~pi0322 & ~n7837;
  assign n7840 = ~n7838 & ~n7839;
  assign n7841 = n7834 & ~n7840;
  assign n7842 = ~n7834 & n7840;
  assign n7843 = ~n7841 & ~n7842;
  assign n7844 = n7828 & n7843;
  assign n7845 = ~n7828 & ~n7843;
  assign n7846 = ~n7844 & ~n7845;
  assign n7847 = pi0350 & ~n7846;
  assign n7848 = ~pi0350 & n7846;
  assign n7849 = ~n7847 & ~n7848;
  assign n7850 = ~n7825 & n7849;
  assign n7851 = pi1198 & n7644;
  assign n7852 = n7850 & n7851;
  assign n7853 = ~n7824 & ~n7852;
  assign n7854 = ~n7782 & ~n7853;
  assign n7855 = ~pi0592 & ~n7854;
  assign n7856 = n7422 & ~n7855;
  assign n7857 = ~n7757 & ~n7856;
  assign n7858 = pi1199 & ~n7645;
  assign n7859 = pi0351 & n7858;
  assign n7860 = ~n7857 & ~n7859;
  assign n7861 = ~pi0461 & ~n7860;
  assign n7862 = ~pi0351 & pi1199;
  assign n7863 = ~n7856 & ~n7862;
  assign n7864 = ~pi0351 & n7858;
  assign n7865 = ~n7863 & ~n7864;
  assign n7866 = pi0461 & ~n7865;
  assign n7867 = ~n7861 & ~n7866;
  assign n7868 = ~pi0357 & ~n7867;
  assign n7869 = ~pi0461 & ~n7865;
  assign n7870 = pi0461 & ~n7860;
  assign n7871 = ~n7869 & ~n7870;
  assign n7872 = pi0357 & ~n7871;
  assign n7873 = ~n7868 & ~n7872;
  assign n7874 = ~pi0356 & ~n7873;
  assign n7875 = ~pi0357 & ~n7871;
  assign n7876 = pi0357 & ~n7867;
  assign n7877 = ~n7875 & ~n7876;
  assign n7878 = pi0356 & ~n7877;
  assign n7879 = pi0360 & ~pi0462;
  assign n7880 = ~pi0360 & pi0462;
  assign n7881 = ~n7879 & ~n7880;
  assign n7882 = pi0352 & ~pi0353;
  assign n7883 = ~pi0352 & pi0353;
  assign n7884 = ~n7882 & ~n7883;
  assign n7885 = n7881 & n7884;
  assign n7886 = ~n7881 & ~n7884;
  assign n7887 = ~n7885 & ~n7886;
  assign n7888 = pi0354 & ~n7887;
  assign n7889 = ~pi0354 & n7887;
  assign n7890 = ~n7888 & ~n7889;
  assign n7891 = ~n7874 & n7890;
  assign n7892 = ~n7878 & n7891;
  assign n7893 = ~pi0356 & ~n7877;
  assign n7894 = pi0356 & ~n7873;
  assign n7895 = ~n7890 & ~n7893;
  assign n7896 = ~n7894 & n7895;
  assign n7897 = ~n7892 & ~n7896;
  assign n7898 = pi0590 & ~n7897;
  assign n7899 = ~pi0591 & ~n7756;
  assign n7900 = ~n7898 & n7899;
  assign n7901 = pi0590 & n7422;
  assign n7902 = pi1197 & ~n7645;
  assign n7903 = pi0318 & ~pi0409;
  assign n7904 = ~pi0318 & pi0409;
  assign n7905 = ~n7903 & ~n7904;
  assign n7906 = pi0401 & ~pi0402;
  assign n7907 = ~pi0401 & pi0402;
  assign n7908 = ~n7906 & ~n7907;
  assign n7909 = pi0406 & n7908;
  assign n7910 = ~pi0406 & ~n7908;
  assign n7911 = ~n7909 & ~n7910;
  assign n7912 = ~pi0403 & ~pi0405;
  assign n7913 = pi0403 & pi0405;
  assign n7914 = ~n7912 & ~n7913;
  assign n7915 = pi0325 & ~pi0326;
  assign n7916 = ~pi0325 & pi0326;
  assign n7917 = ~n7915 & ~n7916;
  assign n7918 = n7914 & n7917;
  assign n7919 = ~n7914 & ~n7917;
  assign n7920 = ~n7918 & ~n7919;
  assign n7921 = n7911 & ~n7920;
  assign n7922 = ~n7911 & n7920;
  assign n7923 = ~n7921 & ~n7922;
  assign n7924 = n7905 & n7923;
  assign n7925 = ~n7905 & ~n7923;
  assign n7926 = ~n7924 & ~n7925;
  assign n7927 = n7485 & ~n7926;
  assign n7928 = ~pi1091 & n7927;
  assign n7929 = pi0567 & n7928;
  assign n7930 = pi0390 & ~pi0410;
  assign n7931 = ~pi0390 & pi0410;
  assign n7932 = ~n7930 & ~n7931;
  assign n7933 = pi0397 & ~pi0412;
  assign n7934 = ~pi0397 & pi0412;
  assign n7935 = ~n7933 & ~n7934;
  assign n7936 = pi0404 & n7935;
  assign n7937 = ~pi0404 & ~n7935;
  assign n7938 = ~n7936 & ~n7937;
  assign n7939 = pi0319 & ~pi0324;
  assign n7940 = ~pi0319 & pi0324;
  assign n7941 = ~n7939 & ~n7940;
  assign n7942 = pi0456 & ~n7941;
  assign n7943 = ~pi0456 & n7941;
  assign n7944 = ~n7942 & ~n7943;
  assign n7945 = n7938 & ~n7944;
  assign n7946 = ~n7938 & n7944;
  assign n7947 = ~n7945 & ~n7946;
  assign n7948 = n7932 & n7947;
  assign n7949 = ~n7932 & ~n7947;
  assign n7950 = ~n7948 & ~n7949;
  assign n7951 = pi0411 & n7950;
  assign n7952 = ~pi0411 & ~n7950;
  assign n7953 = ~n7951 & ~n7952;
  assign n7954 = pi1196 & ~n7953;
  assign n7955 = ~pi0592 & n7929;
  assign n7956 = ~n7954 & n7955;
  assign n7957 = n7858 & ~n7956;
  assign n7958 = ~pi0592 & pi1196;
  assign n7959 = n7422 & ~n7958;
  assign n7960 = n7485 & n7953;
  assign n7961 = ~pi1091 & n7960;
  assign n7962 = pi0567 & n7961;
  assign n7963 = n7958 & n7962;
  assign n7964 = ~pi1199 & ~n7959;
  assign n7965 = ~n7963 & n7964;
  assign n7966 = ~n7957 & ~n7965;
  assign n7967 = ~pi1197 & ~n7966;
  assign n7968 = ~n7902 & ~n7967;
  assign n7969 = pi0333 & ~n7968;
  assign n7970 = pi1198 & ~n7645;
  assign n7971 = n7966 & ~n7970;
  assign n7972 = pi0328 & ~pi0408;
  assign n7973 = ~pi0328 & pi0408;
  assign n7974 = ~n7972 & ~n7973;
  assign n7975 = ~pi0394 & ~pi0396;
  assign n7976 = pi0394 & pi0396;
  assign n7977 = ~n7975 & ~n7976;
  assign n7978 = n7974 & ~n7977;
  assign n7979 = ~n7974 & n7977;
  assign n7980 = ~n7978 & ~n7979;
  assign n7981 = pi0398 & ~pi0399;
  assign n7982 = ~pi0398 & pi0399;
  assign n7983 = ~n7981 & ~n7982;
  assign n7984 = pi0395 & n7983;
  assign n7985 = ~pi0395 & ~n7983;
  assign n7986 = ~n7984 & ~n7985;
  assign n7987 = pi0329 & ~n7986;
  assign n7988 = ~pi0329 & n7986;
  assign n7989 = ~n7987 & ~n7988;
  assign n7990 = pi0400 & ~n7989;
  assign n7991 = ~pi0400 & n7989;
  assign n7992 = ~n7990 & ~n7991;
  assign n7993 = n7980 & n7992;
  assign n7994 = ~n7980 & ~n7992;
  assign n7995 = ~n7993 & ~n7994;
  assign n7996 = ~n7971 & ~n7995;
  assign n7997 = ~pi0333 & ~n7966;
  assign n7998 = ~n7996 & ~n7997;
  assign n7999 = ~n7969 & n7998;
  assign n8000 = ~pi0391 & ~n7999;
  assign n8001 = ~pi0333 & ~n7968;
  assign n8002 = n7966 & ~n7996;
  assign n8003 = ~n8001 & n8002;
  assign n8004 = pi0391 & ~n8003;
  assign n8005 = ~n8000 & ~n8004;
  assign n8006 = ~pi0392 & ~n8005;
  assign n8007 = ~pi0391 & ~n8003;
  assign n8008 = pi0391 & ~n7999;
  assign n8009 = ~n8007 & ~n8008;
  assign n8010 = pi0392 & ~n8009;
  assign n8011 = ~n8006 & ~n8010;
  assign n8012 = ~pi0393 & ~n8011;
  assign n8013 = ~pi0392 & ~n8009;
  assign n8014 = pi0392 & ~n8005;
  assign n8015 = ~n8013 & ~n8014;
  assign n8016 = pi0393 & ~n8015;
  assign n8017 = pi0407 & ~pi0463;
  assign n8018 = ~pi0407 & pi0463;
  assign n8019 = ~n8017 & ~n8018;
  assign n8020 = pi0335 & ~pi0413;
  assign n8021 = ~pi0335 & pi0413;
  assign n8022 = ~n8020 & ~n8021;
  assign n8023 = n8019 & n8022;
  assign n8024 = ~n8019 & ~n8022;
  assign n8025 = ~n8023 & ~n8024;
  assign n8026 = pi0334 & ~n8025;
  assign n8027 = ~pi0334 & n8025;
  assign n8028 = ~n8026 & ~n8027;
  assign n8029 = ~n8012 & n8028;
  assign n8030 = ~n8016 & n8029;
  assign n8031 = ~pi0393 & ~n8015;
  assign n8032 = pi0393 & ~n8011;
  assign n8033 = ~n8028 & ~n8031;
  assign n8034 = ~n8032 & n8033;
  assign n8035 = ~n8030 & ~n8034;
  assign n8036 = ~pi0590 & ~n8035;
  assign n8037 = pi0591 & ~n7901;
  assign n8038 = ~n8036 & n8037;
  assign n8039 = ~n7900 & ~n8038;
  assign n8040 = ~pi0588 & ~n8039;
  assign n8041 = ~pi0590 & ~pi0591;
  assign n8042 = n7422 & ~n8041;
  assign n8043 = ~pi0417 & ~pi0418;
  assign n8044 = pi0417 & pi0418;
  assign n8045 = ~n8043 & ~n8044;
  assign n8046 = pi0437 & n8045;
  assign n8047 = ~pi0437 & ~n8045;
  assign n8048 = ~n8046 & ~n8047;
  assign n8049 = pi0453 & ~pi0464;
  assign n8050 = ~pi0453 & pi0464;
  assign n8051 = ~n8049 & ~n8050;
  assign n8052 = n8048 & n8051;
  assign n8053 = ~n8048 & ~n8051;
  assign n8054 = ~n8052 & ~n8053;
  assign n8055 = pi0415 & ~pi0431;
  assign n8056 = ~pi0415 & pi0431;
  assign n8057 = ~n8055 & ~n8056;
  assign n8058 = pi0416 & ~pi0438;
  assign n8059 = ~pi0416 & pi0438;
  assign n8060 = ~n8058 & ~n8059;
  assign n8061 = n8057 & n8060;
  assign n8062 = ~n8057 & ~n8060;
  assign n8063 = ~n8061 & ~n8062;
  assign n8064 = n8054 & ~n8063;
  assign n8065 = ~n8054 & n8063;
  assign n8066 = pi1197 & ~n8064;
  assign n8067 = ~n8065 & n8066;
  assign n8068 = pi0421 & ~pi0454;
  assign n8069 = ~pi0421 & pi0454;
  assign n8070 = ~n8068 & ~n8069;
  assign n8071 = pi0432 & ~pi0459;
  assign n8072 = ~pi0432 & pi0459;
  assign n8073 = ~n8071 & ~n8072;
  assign n8074 = n8070 & ~n8073;
  assign n8075 = ~n8070 & n8073;
  assign n8076 = ~n8074 & ~n8075;
  assign n8077 = ~pi0419 & ~pi0420;
  assign n8078 = pi0419 & pi0420;
  assign n8079 = ~n8077 & ~n8078;
  assign n8080 = pi0423 & ~pi0424;
  assign n8081 = ~pi0423 & pi0424;
  assign n8082 = ~n8080 & ~n8081;
  assign n8083 = n8079 & ~n8082;
  assign n8084 = ~n8079 & n8082;
  assign n8085 = ~n8083 & ~n8084;
  assign n8086 = n8076 & n8085;
  assign n8087 = ~n8076 & ~n8085;
  assign n8088 = ~n8086 & ~n8087;
  assign n8089 = pi0425 & ~n8088;
  assign n8090 = ~pi0425 & n8088;
  assign n8091 = pi1198 & ~n8089;
  assign n8092 = ~n8090 & n8091;
  assign n8093 = ~n8067 & ~n8092;
  assign n8094 = ~pi0429 & ~pi0435;
  assign n8095 = pi0429 & pi0435;
  assign n8096 = ~n8094 & ~n8095;
  assign n8097 = pi0434 & ~pi0446;
  assign n8098 = ~pi0434 & pi0446;
  assign n8099 = ~n8097 & ~n8098;
  assign n8100 = pi0414 & ~pi0422;
  assign n8101 = ~pi0414 & pi0422;
  assign n8102 = ~n8100 & ~n8101;
  assign n8103 = n8099 & n8102;
  assign n8104 = ~n8099 & ~n8102;
  assign n8105 = ~n8103 & ~n8104;
  assign n8106 = n8096 & n8105;
  assign n8107 = ~n8096 & ~n8105;
  assign n8108 = ~n8106 & ~n8107;
  assign n8109 = pi0436 & ~pi0443;
  assign n8110 = ~pi0436 & pi0443;
  assign n8111 = ~n8109 & ~n8110;
  assign n8112 = ~pi0444 & n8111;
  assign n8113 = pi0444 & ~n8111;
  assign n8114 = ~n8112 & ~n8113;
  assign n8115 = ~n8108 & ~n8114;
  assign n8116 = n8108 & n8114;
  assign n8117 = n7958 & ~n8115;
  assign n8118 = ~n8116 & n8117;
  assign n8119 = n8093 & ~n8118;
  assign n8120 = n7644 & n8119;
  assign n8121 = ~pi1199 & ~n7645;
  assign n8122 = ~n8120 & n8121;
  assign n8123 = pi0433 & ~pi0451;
  assign n8124 = ~pi0433 & pi0451;
  assign n8125 = ~n8123 & ~n8124;
  assign n8126 = pi0449 & n8125;
  assign n8127 = ~pi0449 & ~n8125;
  assign n8128 = ~n8126 & ~n8127;
  assign n8129 = ~pi0427 & pi0428;
  assign n8130 = pi0427 & ~pi0428;
  assign n8131 = ~n8129 & ~n8130;
  assign n8132 = pi0430 & ~n8131;
  assign n8133 = ~pi0430 & n8131;
  assign n8134 = ~n8132 & ~n8133;
  assign n8135 = ~pi0426 & ~n8134;
  assign n8136 = pi0426 & n8134;
  assign n8137 = ~n8135 & ~n8136;
  assign n8138 = ~pi0445 & ~n8137;
  assign n8139 = pi0445 & n8137;
  assign n8140 = ~n8138 & ~n8139;
  assign n8141 = ~pi0448 & ~n8140;
  assign n8142 = pi0448 & n8140;
  assign n8143 = ~n8141 & ~n8142;
  assign n8144 = n8120 & ~n8143;
  assign n8145 = ~n7645 & ~n8144;
  assign n8146 = n8128 & ~n8145;
  assign n8147 = n8120 & n8143;
  assign n8148 = ~n7645 & ~n8147;
  assign n8149 = ~n8128 & ~n8148;
  assign n8150 = pi1199 & ~n8146;
  assign n8151 = ~n8149 & n8150;
  assign n8152 = n8041 & ~n8122;
  assign n8153 = ~n8151 & n8152;
  assign n8154 = pi0588 & ~n8042;
  assign n8155 = ~n8153 & n8154;
  assign n8156 = n7427 & ~n8155;
  assign n8157 = ~n8040 & n8156;
  assign n8158 = n7636 & ~n8041;
  assign n8159 = ~pi0087 & ~n7623;
  assign n8160 = ~n7614 & n8159;
  assign n8161 = pi0087 & ~pi0100;
  assign n8162 = n2530 & n8161;
  assign n8163 = ~n7493 & n8162;
  assign n8164 = ~n7494 & n8163;
  assign n8165 = ~pi0075 & ~n8164;
  assign n8166 = ~n8160 & n8165;
  assign n8167 = ~n7599 & ~n8166;
  assign n8168 = pi0567 & ~n8167;
  assign n8169 = n7469 & ~n8168;
  assign n8170 = ~pi0592 & ~n8169;
  assign n8171 = pi0592 & ~n7636;
  assign n8172 = ~n8170 & ~n8171;
  assign n8173 = ~n8093 & n8172;
  assign n8174 = ~pi1196 & ~n7636;
  assign n8175 = ~pi0443 & ~pi0592;
  assign n8176 = ~n7636 & ~n8175;
  assign n8177 = ~n8169 & n8175;
  assign n8178 = ~n8176 & ~n8177;
  assign n8179 = ~pi0444 & ~n8178;
  assign n8180 = pi0443 & ~pi0592;
  assign n8181 = ~n7636 & ~n8180;
  assign n8182 = ~n8169 & n8180;
  assign n8183 = ~n8181 & ~n8182;
  assign n8184 = pi0444 & ~n8183;
  assign n8185 = ~n8179 & ~n8184;
  assign n8186 = ~pi0436 & ~n8185;
  assign n8187 = ~pi0444 & ~n8183;
  assign n8188 = pi0444 & ~n8178;
  assign n8189 = ~n8187 & ~n8188;
  assign n8190 = pi0436 & ~n8189;
  assign n8191 = n8108 & ~n8186;
  assign n8192 = ~n8190 & n8191;
  assign n8193 = ~pi0436 & ~n8189;
  assign n8194 = pi0436 & ~n8185;
  assign n8195 = ~n8108 & ~n8193;
  assign n8196 = ~n8194 & n8195;
  assign n8197 = pi1196 & ~n8192;
  assign n8198 = ~n8196 & n8197;
  assign n8199 = n8093 & ~n8174;
  assign n8200 = ~n8198 & n8199;
  assign n8201 = ~n8173 & ~n8200;
  assign n8202 = ~pi1199 & n8201;
  assign n8203 = pi0428 & ~n8201;
  assign n8204 = ~pi0428 & n8172;
  assign n8205 = ~n8203 & ~n8204;
  assign n8206 = ~pi0427 & ~n8205;
  assign n8207 = ~pi0428 & ~n8201;
  assign n8208 = pi0428 & n8172;
  assign n8209 = ~n8207 & ~n8208;
  assign n8210 = pi0427 & ~n8209;
  assign n8211 = ~n8206 & ~n8210;
  assign n8212 = pi0430 & ~n8211;
  assign n8213 = ~pi0427 & ~n8209;
  assign n8214 = pi0427 & ~n8205;
  assign n8215 = ~n8213 & ~n8214;
  assign n8216 = ~pi0430 & ~n8215;
  assign n8217 = ~n8212 & ~n8216;
  assign n8218 = pi0426 & ~n8217;
  assign n8219 = pi0430 & ~n8215;
  assign n8220 = ~pi0430 & ~n8211;
  assign n8221 = ~n8219 & ~n8220;
  assign n8222 = ~pi0426 & ~n8221;
  assign n8223 = ~n8218 & ~n8222;
  assign n8224 = pi0445 & ~n8223;
  assign n8225 = pi0426 & ~n8221;
  assign n8226 = ~pi0426 & ~n8217;
  assign n8227 = ~n8225 & ~n8226;
  assign n8228 = ~pi0445 & ~n8227;
  assign n8229 = ~n8224 & ~n8228;
  assign n8230 = pi0448 & ~n8128;
  assign n8231 = ~pi0448 & n8128;
  assign n8232 = ~n8230 & ~n8231;
  assign n8233 = ~n8229 & ~n8232;
  assign n8234 = pi0445 & ~n8227;
  assign n8235 = ~pi0445 & ~n8223;
  assign n8236 = ~n8234 & ~n8235;
  assign n8237 = n8232 & ~n8236;
  assign n8238 = pi1199 & ~n8233;
  assign n8239 = ~n8237 & n8238;
  assign n8240 = n8041 & ~n8202;
  assign n8241 = ~n8239 & n8240;
  assign n8242 = n7425 & ~n8158;
  assign n8243 = ~n8241 & n8242;
  assign n8244 = ~n7592 & ~n8041;
  assign n8245 = ~pi1196 & n7592;
  assign n8246 = n7592 & ~n8175;
  assign n8247 = ~pi0436 & pi0444;
  assign n8248 = pi0436 & ~pi0444;
  assign n8249 = ~n8247 & ~n8248;
  assign n8250 = n8108 & ~n8249;
  assign n8251 = ~n8108 & n8249;
  assign n8252 = ~n8250 & ~n8251;
  assign n8253 = ~n8177 & n8252;
  assign n8254 = ~n8246 & n8253;
  assign n8255 = n7592 & ~n8180;
  assign n8256 = ~n8182 & ~n8252;
  assign n8257 = ~n8255 & n8256;
  assign n8258 = pi1196 & ~n8254;
  assign n8259 = ~n8257 & n8258;
  assign n8260 = ~n8245 & ~n8259;
  assign n8261 = n8093 & ~n8260;
  assign n8262 = pi0592 & n7592;
  assign n8263 = ~n8170 & ~n8262;
  assign n8264 = ~n8093 & ~n8263;
  assign n8265 = ~n8261 & ~n8264;
  assign n8266 = ~pi1199 & ~n8265;
  assign n8267 = ~pi0428 & n8263;
  assign n8268 = pi0428 & n8265;
  assign n8269 = pi0427 & ~n8267;
  assign n8270 = ~n8268 & n8269;
  assign n8271 = ~pi0428 & n8265;
  assign n8272 = pi0428 & n8263;
  assign n8273 = ~pi0427 & ~n8272;
  assign n8274 = ~n8271 & n8273;
  assign n8275 = ~n8270 & ~n8274;
  assign n8276 = ~pi0430 & ~n8275;
  assign n8277 = n8131 & n8263;
  assign n8278 = ~n8131 & n8265;
  assign n8279 = ~n8277 & ~n8278;
  assign n8280 = pi0430 & n8279;
  assign n8281 = ~n8276 & ~n8280;
  assign n8282 = ~pi0426 & ~n8281;
  assign n8283 = pi0430 & ~n8275;
  assign n8284 = ~pi0430 & n8279;
  assign n8285 = ~n8283 & ~n8284;
  assign n8286 = pi0426 & ~n8285;
  assign n8287 = ~n8282 & ~n8286;
  assign n8288 = ~pi0445 & ~n8287;
  assign n8289 = ~pi0426 & ~n8285;
  assign n8290 = pi0426 & ~n8281;
  assign n8291 = ~n8289 & ~n8290;
  assign n8292 = pi0445 & ~n8291;
  assign n8293 = ~n8288 & ~n8292;
  assign n8294 = pi0448 & n8293;
  assign n8295 = ~pi0445 & ~n8291;
  assign n8296 = pi0445 & ~n8287;
  assign n8297 = ~n8295 & ~n8296;
  assign n8298 = ~pi0448 & n8297;
  assign n8299 = ~n8128 & ~n8294;
  assign n8300 = ~n8298 & n8299;
  assign n8301 = ~pi0448 & n8293;
  assign n8302 = pi0448 & n8297;
  assign n8303 = n8128 & ~n8301;
  assign n8304 = ~n8302 & n8303;
  assign n8305 = ~n8300 & ~n8304;
  assign n8306 = pi1199 & ~n8305;
  assign n8307 = n8041 & ~n8266;
  assign n8308 = ~n8306 & n8307;
  assign n8309 = ~n7425 & ~n8244;
  assign n8310 = ~n8308 & n8309;
  assign n8311 = ~n8243 & ~n8310;
  assign n8312 = pi0588 & ~n8311;
  assign n8313 = pi0591 & n7636;
  assign n8314 = n7825 & ~n8172;
  assign n8315 = ~pi0350 & ~pi0592;
  assign n8316 = ~n7636 & ~n8315;
  assign n8317 = ~n8169 & n8315;
  assign n8318 = n7846 & ~n8317;
  assign n8319 = ~n8316 & n8318;
  assign n8320 = pi0350 & ~pi0592;
  assign n8321 = ~n7636 & ~n8320;
  assign n8322 = ~n8169 & n8320;
  assign n8323 = ~n7846 & ~n8322;
  assign n8324 = ~n8321 & n8323;
  assign n8325 = ~n7825 & ~n8319;
  assign n8326 = ~n8324 & n8325;
  assign n8327 = pi1198 & ~n8314;
  assign n8328 = ~n8326 & n8327;
  assign n8329 = ~pi0455 & ~n8172;
  assign n8330 = pi0455 & ~n7636;
  assign n8331 = ~n8329 & ~n8330;
  assign n8332 = ~pi0452 & ~n8331;
  assign n8333 = pi0455 & ~n8172;
  assign n8334 = ~pi0455 & ~n7636;
  assign n8335 = ~n8333 & ~n8334;
  assign n8336 = pi0452 & ~n8335;
  assign n8337 = ~n8332 & ~n8336;
  assign n8338 = ~pi0355 & ~n8337;
  assign n8339 = ~pi0452 & ~n8335;
  assign n8340 = pi0452 & ~n8331;
  assign n8341 = ~n8339 & ~n8340;
  assign n8342 = pi0355 & ~n8341;
  assign n8343 = ~n8338 & ~n8342;
  assign n8344 = pi0458 & ~n8343;
  assign n8345 = ~pi0355 & ~n8341;
  assign n8346 = pi0355 & ~n8337;
  assign n8347 = ~n8345 & ~n8346;
  assign n8348 = ~pi0458 & ~n8347;
  assign n8349 = n7812 & ~n8344;
  assign n8350 = ~n8348 & n8349;
  assign n8351 = pi0458 & ~n8347;
  assign n8352 = ~pi0458 & ~n8343;
  assign n8353 = ~n7812 & ~n8351;
  assign n8354 = ~n8352 & n8353;
  assign n8355 = pi1196 & ~n8350;
  assign n8356 = ~n8354 & n8355;
  assign n8357 = ~pi1198 & ~n8174;
  assign n8358 = ~n8356 & n8357;
  assign n8359 = ~n8328 & ~n8358;
  assign n8360 = ~n7782 & ~n8359;
  assign n8361 = n7782 & n8172;
  assign n8362 = ~n8360 & ~n8361;
  assign n8363 = ~n7862 & n8362;
  assign n8364 = pi1199 & ~n8172;
  assign n8365 = ~pi0351 & n8364;
  assign n8366 = ~n8363 & ~n8365;
  assign n8367 = ~pi0461 & ~n8366;
  assign n8368 = ~n7757 & n8362;
  assign n8369 = pi0351 & n8364;
  assign n8370 = ~n8368 & ~n8369;
  assign n8371 = pi0461 & ~n8370;
  assign n8372 = ~n8367 & ~n8371;
  assign n8373 = ~pi0357 & ~n8372;
  assign n8374 = ~pi0461 & ~n8370;
  assign n8375 = pi0461 & ~n8366;
  assign n8376 = ~n8374 & ~n8375;
  assign n8377 = pi0357 & ~n8376;
  assign n8378 = ~n8373 & ~n8377;
  assign n8379 = ~pi0356 & ~n8378;
  assign n8380 = ~pi0357 & ~n8376;
  assign n8381 = pi0357 & ~n8372;
  assign n8382 = ~n8380 & ~n8381;
  assign n8383 = pi0356 & ~n8382;
  assign n8384 = ~n8379 & ~n8383;
  assign n8385 = ~n7890 & ~n8384;
  assign n8386 = ~pi0356 & ~n8382;
  assign n8387 = pi0356 & ~n8378;
  assign n8388 = ~n8386 & ~n8387;
  assign n8389 = n7890 & ~n8388;
  assign n8390 = ~pi0591 & ~n8385;
  assign n8391 = ~n8389 & n8390;
  assign n8392 = pi0590 & ~n8313;
  assign n8393 = ~n8391 & n8392;
  assign n8394 = pi1197 & ~n8172;
  assign n8395 = pi1198 & ~n7995;
  assign n8396 = n8172 & n8395;
  assign n8397 = ~pi0075 & n7954;
  assign n8398 = ~n7926 & ~n8397;
  assign n8399 = n7617 & n8398;
  assign n8400 = n7614 & ~n8399;
  assign n8401 = n8159 & ~n8400;
  assign n8402 = ~n7628 & n8162;
  assign n8403 = n7495 & ~n7926;
  assign n8404 = n7626 & ~n8403;
  assign n8405 = n8402 & ~n8404;
  assign n8406 = ~pi1196 & n8405;
  assign n8407 = n7495 & n7953;
  assign n8408 = n7626 & ~n8407;
  assign n8409 = n8405 & ~n8408;
  assign n8410 = ~pi0075 & ~pi0592;
  assign n8411 = pi1199 & n8410;
  assign n8412 = ~n8406 & n8411;
  assign n8413 = ~n8409 & n8412;
  assign n8414 = ~n8401 & n8413;
  assign n8415 = ~n7634 & ~n8410;
  assign n8416 = n8402 & ~n8408;
  assign n8417 = n7617 & n7953;
  assign n8418 = n7614 & ~n8417;
  assign n8419 = n8159 & ~n8418;
  assign n8420 = pi1196 & n8410;
  assign n8421 = ~n8416 & n8420;
  assign n8422 = ~n8419 & n8421;
  assign n8423 = ~pi1196 & n7633;
  assign n8424 = ~n8422 & ~n8423;
  assign n8425 = ~pi1199 & ~n8424;
  assign n8426 = ~n8414 & ~n8415;
  assign n8427 = ~n8425 & n8426;
  assign n8428 = pi0567 & ~n8427;
  assign n8429 = n7469 & ~n8395;
  assign n8430 = ~n8428 & n8429;
  assign n8431 = ~n8396 & ~n8430;
  assign n8432 = ~pi1197 & n8431;
  assign n8433 = ~n8394 & ~n8432;
  assign n8434 = pi0333 & ~n8433;
  assign n8435 = ~pi0333 & n8431;
  assign n8436 = ~n8434 & ~n8435;
  assign n8437 = pi0391 & ~n8436;
  assign n8438 = pi0333 & ~n8431;
  assign n8439 = ~pi0333 & n8433;
  assign n8440 = ~n8438 & ~n8439;
  assign n8441 = ~pi0391 & n8440;
  assign n8442 = ~n8437 & ~n8441;
  assign n8443 = ~pi0392 & ~n8442;
  assign n8444 = ~pi0391 & ~n8436;
  assign n8445 = pi0391 & n8440;
  assign n8446 = ~n8444 & ~n8445;
  assign n8447 = pi0392 & ~n8446;
  assign n8448 = ~n8443 & ~n8447;
  assign n8449 = ~pi0393 & ~n8448;
  assign n8450 = ~pi0392 & ~n8446;
  assign n8451 = pi0392 & ~n8442;
  assign n8452 = ~n8450 & ~n8451;
  assign n8453 = pi0393 & ~n8452;
  assign n8454 = ~n8449 & ~n8453;
  assign n8455 = ~pi0334 & n8454;
  assign n8456 = ~pi0393 & ~n8452;
  assign n8457 = pi0393 & ~n8448;
  assign n8458 = ~n8456 & ~n8457;
  assign n8459 = pi0334 & n8458;
  assign n8460 = n8025 & ~n8455;
  assign n8461 = ~n8459 & n8460;
  assign n8462 = ~pi0334 & n8458;
  assign n8463 = pi0334 & n8454;
  assign n8464 = ~n8025 & ~n8462;
  assign n8465 = ~n8463 & n8464;
  assign n8466 = pi0591 & ~n8461;
  assign n8467 = ~n8465 & n8466;
  assign n8468 = pi0377 & pi0592;
  assign n8469 = ~n7636 & ~n8468;
  assign n8470 = ~n8169 & n8468;
  assign n8471 = ~n7718 & ~n8470;
  assign n8472 = ~n8469 & n8471;
  assign n8473 = ~pi0377 & pi0592;
  assign n8474 = ~n7636 & ~n8473;
  assign n8475 = ~n8169 & n8473;
  assign n8476 = n7718 & ~n8475;
  assign n8477 = ~n8474 & n8476;
  assign n8478 = ~n8472 & ~n8477;
  assign n8479 = n7696 & ~n8478;
  assign n8480 = pi0592 & ~n8169;
  assign n8481 = ~pi0592 & ~n7636;
  assign n8482 = ~n8480 & ~n8481;
  assign n8483 = ~n7696 & n8482;
  assign n8484 = ~n8479 & ~n8483;
  assign n8485 = pi1199 & n8484;
  assign n8486 = n7636 & ~n7695;
  assign n8487 = n7695 & n8482;
  assign n8488 = ~n8486 & ~n8487;
  assign n8489 = n7669 & ~n8488;
  assign n8490 = ~pi1196 & ~n7695;
  assign n8491 = n8482 & ~n8490;
  assign n8492 = ~pi1196 & n8486;
  assign n8493 = ~n8491 & ~n8492;
  assign n8494 = ~n7669 & ~n8493;
  assign n8495 = ~pi1199 & ~n8489;
  assign n8496 = ~n8494 & n8495;
  assign n8497 = ~n8485 & ~n8496;
  assign n8498 = ~pi0374 & ~n8497;
  assign n8499 = ~pi1198 & pi1199;
  assign n8500 = n8484 & n8499;
  assign n8501 = ~pi1198 & n8496;
  assign n8502 = pi1198 & ~n8482;
  assign n8503 = ~n8500 & ~n8502;
  assign n8504 = ~n8501 & n8503;
  assign n8505 = pi0374 & ~n8504;
  assign n8506 = ~n8498 & ~n8505;
  assign n8507 = pi0369 & ~n8506;
  assign n8508 = ~pi0374 & ~n8504;
  assign n8509 = pi0374 & ~n8497;
  assign n8510 = ~n8508 & ~n8509;
  assign n8511 = ~pi0369 & ~n8510;
  assign n8512 = ~n8507 & ~n8511;
  assign n8513 = ~pi0370 & ~n8512;
  assign n8514 = ~pi0369 & ~n8506;
  assign n8515 = pi0369 & ~n8510;
  assign n8516 = ~n8514 & ~n8515;
  assign n8517 = pi0370 & ~n8516;
  assign n8518 = ~n8513 & ~n8517;
  assign n8519 = ~pi0371 & ~n8518;
  assign n8520 = ~pi0370 & ~n8516;
  assign n8521 = pi0370 & ~n8512;
  assign n8522 = ~n8520 & ~n8521;
  assign n8523 = pi0371 & ~n8522;
  assign n8524 = ~n8519 & ~n8523;
  assign n8525 = ~pi0373 & ~n8524;
  assign n8526 = ~pi0371 & ~n8522;
  assign n8527 = pi0371 & ~n8518;
  assign n8528 = ~n8526 & ~n8527;
  assign n8529 = pi0373 & ~n8528;
  assign n8530 = ~n8525 & ~n8529;
  assign n8531 = ~pi0375 & n8530;
  assign n8532 = ~pi0373 & ~n8528;
  assign n8533 = pi0373 & ~n8524;
  assign n8534 = ~n8532 & ~n8533;
  assign n8535 = pi0375 & n8534;
  assign n8536 = n7734 & ~n8531;
  assign n8537 = ~n8535 & n8536;
  assign n8538 = pi0375 & n8530;
  assign n8539 = ~pi0375 & n8534;
  assign n8540 = ~n7734 & ~n8538;
  assign n8541 = ~n8539 & n8540;
  assign n8542 = ~pi0591 & ~n8537;
  assign n8543 = ~n8541 & n8542;
  assign n8544 = ~pi0590 & ~n8467;
  assign n8545 = ~n8543 & n8544;
  assign n8546 = n7425 & ~n8545;
  assign n8547 = ~n8393 & n8546;
  assign n8548 = pi0591 & ~n7592;
  assign n8549 = n7782 & ~n8263;
  assign n8550 = n7825 & ~n8263;
  assign n8551 = n7592 & ~n8320;
  assign n8552 = n8323 & ~n8551;
  assign n8553 = n7592 & ~n8315;
  assign n8554 = n8318 & ~n8553;
  assign n8555 = ~n7825 & ~n8552;
  assign n8556 = ~n8554 & n8555;
  assign n8557 = pi1198 & ~n8550;
  assign n8558 = ~n8556 & n8557;
  assign n8559 = pi0455 & ~n8263;
  assign n8560 = ~pi0455 & n7592;
  assign n8561 = ~n8559 & ~n8560;
  assign n8562 = ~pi0452 & ~n8561;
  assign n8563 = ~pi0455 & ~n8263;
  assign n8564 = pi0455 & n7592;
  assign n8565 = ~n8563 & ~n8564;
  assign n8566 = pi0452 & ~n8565;
  assign n8567 = pi0355 & ~n7815;
  assign n8568 = ~pi0355 & n7815;
  assign n8569 = ~n8567 & ~n8568;
  assign n8570 = ~n8562 & ~n8569;
  assign n8571 = ~n8566 & n8570;
  assign n8572 = ~pi0452 & ~n8565;
  assign n8573 = pi0452 & ~n8561;
  assign n8574 = n8569 & ~n8572;
  assign n8575 = ~n8573 & n8574;
  assign n8576 = pi1196 & ~n8571;
  assign n8577 = ~n8575 & n8576;
  assign n8578 = ~pi1198 & ~n8245;
  assign n8579 = ~n8577 & n8578;
  assign n8580 = ~n7782 & ~n8558;
  assign n8581 = ~n8579 & n8580;
  assign n8582 = ~n8549 & ~n8581;
  assign n8583 = ~n7862 & ~n8582;
  assign n8584 = pi1199 & ~n8263;
  assign n8585 = ~pi0351 & n8584;
  assign n8586 = ~n8583 & ~n8585;
  assign n8587 = ~pi0461 & ~n8586;
  assign n8588 = ~n7757 & ~n8582;
  assign n8589 = pi0351 & n8584;
  assign n8590 = ~n8588 & ~n8589;
  assign n8591 = pi0461 & ~n8590;
  assign n8592 = ~n8587 & ~n8591;
  assign n8593 = ~pi0357 & ~n8592;
  assign n8594 = ~pi0461 & ~n8590;
  assign n8595 = pi0461 & ~n8586;
  assign n8596 = ~n8594 & ~n8595;
  assign n8597 = pi0357 & ~n8596;
  assign n8598 = ~n8593 & ~n8597;
  assign n8599 = ~pi0356 & ~n8598;
  assign n8600 = ~pi0357 & ~n8596;
  assign n8601 = pi0357 & ~n8592;
  assign n8602 = ~n8600 & ~n8601;
  assign n8603 = pi0356 & ~n8602;
  assign n8604 = ~n8599 & ~n8603;
  assign n8605 = ~n7890 & ~n8604;
  assign n8606 = ~pi0356 & ~n8602;
  assign n8607 = pi0356 & ~n8598;
  assign n8608 = ~n8606 & ~n8607;
  assign n8609 = n7890 & ~n8608;
  assign n8610 = ~pi0591 & ~n8605;
  assign n8611 = ~n8609 & n8610;
  assign n8612 = pi0590 & ~n8548;
  assign n8613 = ~n8611 & n8612;
  assign n8614 = ~n7429 & n7962;
  assign n8615 = pi0038 & n7961;
  assign n8616 = ~pi0100 & ~n8615;
  assign n8617 = n7545 & ~n7953;
  assign n8618 = n7550 & ~n8617;
  assign n8619 = ~n7570 & n7961;
  assign n8620 = pi0299 & ~n8619;
  assign n8621 = ~n6227 & n7602;
  assign n8622 = ~n7961 & ~n8621;
  assign n8623 = ~n6242 & n8622;
  assign n8624 = n6198 & n7602;
  assign n8625 = ~n7961 & ~n8624;
  assign n8626 = n6242 & n8625;
  assign n8627 = n7570 & ~n8623;
  assign n8628 = ~n8626 & n8627;
  assign n8629 = n8620 & ~n8628;
  assign n8630 = ~n7551 & n7961;
  assign n8631 = ~pi0299 & ~n8630;
  assign n8632 = ~n6205 & n8622;
  assign n8633 = n6205 & n8625;
  assign n8634 = n7551 & ~n8632;
  assign n8635 = ~n8633 & n8634;
  assign n8636 = n8631 & ~n8635;
  assign n8637 = pi0039 & ~n8629;
  assign n8638 = ~n8636 & n8637;
  assign n8639 = ~n8618 & ~n8638;
  assign n8640 = ~pi0038 & ~n8639;
  assign n8641 = n8616 & ~n8640;
  assign n8642 = n7623 & ~n7961;
  assign n8643 = ~n8641 & ~n8642;
  assign n8644 = ~pi0087 & ~n8643;
  assign n8645 = ~n2625 & n7961;
  assign n8646 = pi0087 & ~n8645;
  assign n8647 = n7494 & ~n7953;
  assign n8648 = n7502 & ~n8647;
  assign n8649 = n8646 & ~n8648;
  assign n8650 = ~n8644 & ~n8649;
  assign n8651 = ~pi0075 & ~n8650;
  assign n8652 = ~n7475 & n7961;
  assign n8653 = pi0075 & ~n8652;
  assign n8654 = ~pi1091 & ~n7960;
  assign n8655 = n7483 & ~n8654;
  assign n8656 = n8653 & ~n8655;
  assign n8657 = ~n8651 & ~n8656;
  assign n8658 = pi0567 & ~n8657;
  assign n8659 = n7469 & ~n8658;
  assign n8660 = n7958 & ~n8614;
  assign n8661 = ~n8659 & n8660;
  assign n8662 = ~pi1199 & ~n8245;
  assign n8663 = ~n8661 & n8662;
  assign n8664 = n7484 & ~n7926;
  assign n8665 = n8614 & n8664;
  assign n8666 = n7958 & ~n8665;
  assign n8667 = ~n7429 & n7929;
  assign n8668 = ~pi0592 & ~pi1196;
  assign n8669 = ~n8667 & n8668;
  assign n8670 = ~n8666 & ~n8669;
  assign n8671 = ~n7469 & ~n8670;
  assign n8672 = ~n7570 & n7928;
  assign n8673 = pi0299 & ~n8672;
  assign n8674 = ~n8620 & ~n8673;
  assign n8675 = ~n7926 & n7961;
  assign n8676 = ~n8624 & ~n8675;
  assign n8677 = n6242 & n8676;
  assign n8678 = ~n8621 & ~n8675;
  assign n8679 = ~n6242 & n8678;
  assign n8680 = n7570 & ~n8677;
  assign n8681 = ~n8679 & n8680;
  assign n8682 = ~n8674 & ~n8681;
  assign n8683 = ~n7551 & n7928;
  assign n8684 = ~pi0299 & ~n8683;
  assign n8685 = ~n8631 & ~n8684;
  assign n8686 = n6205 & n8676;
  assign n8687 = ~n6205 & n8678;
  assign n8688 = n7551 & ~n8686;
  assign n8689 = ~n8687 & n8688;
  assign n8690 = ~n8685 & ~n8689;
  assign n8691 = pi0039 & ~n8682;
  assign n8692 = ~n8690 & n8691;
  assign n8693 = n7520 & ~n7926;
  assign n8694 = pi0122 & ~n8693;
  assign n8695 = ~pi0122 & ~n8664;
  assign n8696 = pi1093 & ~n8695;
  assign n8697 = ~n8694 & n8696;
  assign n8698 = n7545 & ~n8697;
  assign n8699 = n8618 & ~n8698;
  assign n8700 = ~n8692 & ~n8699;
  assign n8701 = ~pi0038 & ~n8700;
  assign n8702 = pi0038 & n7928;
  assign n8703 = ~pi0100 & ~n8702;
  assign n8704 = ~n8616 & ~n8703;
  assign n8705 = ~n8701 & ~n8704;
  assign n8706 = ~n2530 & n8675;
  assign n8707 = ~pi0232 & ~n8675;
  assign n8708 = ~n7620 & n8707;
  assign n8709 = n6197 & ~n7471;
  assign n8710 = ~n7470 & ~n8709;
  assign n8711 = pi0228 & n8710;
  assign n8712 = n8675 & ~n8711;
  assign n8713 = n7470 & n7619;
  assign n8714 = ~pi1091 & ~n8675;
  assign n8715 = n8710 & ~n8714;
  assign n8716 = ~n7509 & n8715;
  assign n8717 = ~n8713 & ~n8716;
  assign n8718 = pi0228 & ~n8717;
  assign n8719 = pi0232 & ~n8712;
  assign n8720 = ~n8718 & n8719;
  assign n8721 = n2530 & ~n8708;
  assign n8722 = ~n8720 & n8721;
  assign n8723 = pi0100 & ~n8706;
  assign n8724 = ~n8722 & n8723;
  assign n8725 = ~n8705 & ~n8724;
  assign n8726 = ~pi0087 & ~n8725;
  assign n8727 = ~n2625 & n7928;
  assign n8728 = pi0087 & ~n8727;
  assign n8729 = ~n8646 & ~n8728;
  assign n8730 = n7494 & n7926;
  assign n8731 = n7502 & ~n8730;
  assign n8732 = ~n8647 & n8731;
  assign n8733 = ~n8729 & ~n8732;
  assign n8734 = ~n8726 & ~n8733;
  assign n8735 = ~pi0075 & ~n8734;
  assign n8736 = ~n7475 & n7928;
  assign n8737 = pi0075 & ~n8736;
  assign n8738 = ~n8653 & ~n8737;
  assign n8739 = n7483 & ~n8714;
  assign n8740 = ~n8738 & ~n8739;
  assign n8741 = ~n8735 & ~n8740;
  assign n8742 = n8666 & ~n8741;
  assign n8743 = n8728 & ~n8731;
  assign n8744 = n7623 & ~n7928;
  assign n8745 = n7544 & ~n8698;
  assign n8746 = ~n7928 & ~n8621;
  assign n8747 = ~n6242 & n8746;
  assign n8748 = ~n7928 & ~n8624;
  assign n8749 = n6242 & n8748;
  assign n8750 = n7570 & ~n8747;
  assign n8751 = ~n8749 & n8750;
  assign n8752 = n8673 & ~n8751;
  assign n8753 = ~n6205 & n8746;
  assign n8754 = n6205 & n8748;
  assign n8755 = n7551 & ~n8753;
  assign n8756 = ~n8754 & n8755;
  assign n8757 = n8684 & ~n8756;
  assign n8758 = pi0039 & ~n8752;
  assign n8759 = ~n8757 & n8758;
  assign n8760 = ~n8745 & ~n8759;
  assign n8761 = ~pi0038 & ~n8760;
  assign n8762 = n8703 & ~n8761;
  assign n8763 = ~n8744 & ~n8762;
  assign n8764 = ~pi0087 & ~n8763;
  assign n8765 = ~n8743 & ~n8764;
  assign n8766 = ~pi0075 & ~n8765;
  assign n8767 = ~pi1091 & ~n7927;
  assign n8768 = n7483 & ~n8767;
  assign n8769 = n8737 & ~n8768;
  assign n8770 = ~n8766 & ~n8769;
  assign n8771 = n8669 & ~n8770;
  assign n8772 = ~n8742 & ~n8771;
  assign n8773 = pi0567 & ~n8772;
  assign n8774 = pi1199 & ~n8671;
  assign n8775 = ~n8773 & n8774;
  assign n8776 = ~n8395 & ~n8663;
  assign n8777 = ~n8775 & n8776;
  assign n8778 = n8170 & n8395;
  assign n8779 = ~n8262 & ~n8778;
  assign n8780 = ~n8777 & n8779;
  assign n8781 = ~pi1197 & ~n8780;
  assign n8782 = pi1197 & ~n8263;
  assign n8783 = ~n8781 & ~n8782;
  assign n8784 = ~pi0333 & ~n8783;
  assign n8785 = pi0333 & ~n8780;
  assign n8786 = ~n8784 & ~n8785;
  assign n8787 = ~pi0391 & ~n8786;
  assign n8788 = ~pi0333 & ~n8780;
  assign n8789 = pi0333 & ~n8783;
  assign n8790 = ~n8788 & ~n8789;
  assign n8791 = pi0391 & ~n8790;
  assign n8792 = ~n8787 & ~n8791;
  assign n8793 = ~pi0392 & ~n8792;
  assign n8794 = ~pi0391 & ~n8790;
  assign n8795 = pi0391 & ~n8786;
  assign n8796 = ~n8794 & ~n8795;
  assign n8797 = pi0392 & ~n8796;
  assign n8798 = ~n8793 & ~n8797;
  assign n8799 = pi0393 & n8028;
  assign n8800 = ~pi0393 & ~n8028;
  assign n8801 = ~n8799 & ~n8800;
  assign n8802 = ~n8798 & ~n8801;
  assign n8803 = ~pi0392 & ~n8796;
  assign n8804 = pi0392 & ~n8792;
  assign n8805 = ~n8803 & ~n8804;
  assign n8806 = n8801 & ~n8805;
  assign n8807 = pi0591 & ~n8802;
  assign n8808 = ~n8806 & n8807;
  assign n8809 = ~pi0592 & n7592;
  assign n8810 = ~n8480 & ~n8809;
  assign n8811 = ~n7696 & n8810;
  assign n8812 = ~n7592 & n7696;
  assign n8813 = ~pi1199 & ~n8812;
  assign n8814 = ~n8811 & n8813;
  assign n8815 = n7592 & ~n8473;
  assign n8816 = n8476 & ~n8815;
  assign n8817 = n7592 & ~n8468;
  assign n8818 = n8471 & ~n8817;
  assign n8819 = ~n8816 & ~n8818;
  assign n8820 = n7696 & ~n8819;
  assign n8821 = pi1199 & ~n8811;
  assign n8822 = ~n8820 & n8821;
  assign n8823 = ~n8814 & ~n8822;
  assign n8824 = ~pi0374 & ~n8823;
  assign n8825 = ~pi1198 & ~n8823;
  assign n8826 = pi1198 & ~n8810;
  assign n8827 = ~n8825 & ~n8826;
  assign n8828 = pi0374 & ~n8827;
  assign n8829 = ~n8824 & ~n8828;
  assign n8830 = pi0369 & ~n8829;
  assign n8831 = ~pi0374 & ~n8827;
  assign n8832 = pi0374 & ~n8823;
  assign n8833 = ~n8831 & ~n8832;
  assign n8834 = ~pi0369 & ~n8833;
  assign n8835 = ~n8830 & ~n8834;
  assign n8836 = ~pi0370 & ~n8835;
  assign n8837 = ~pi0369 & ~n8829;
  assign n8838 = pi0369 & ~n8833;
  assign n8839 = ~n8837 & ~n8838;
  assign n8840 = pi0370 & ~n8839;
  assign n8841 = ~n8836 & ~n8840;
  assign n8842 = ~pi0371 & ~n8841;
  assign n8843 = ~pi0370 & ~n8839;
  assign n8844 = pi0370 & ~n8835;
  assign n8845 = ~n8843 & ~n8844;
  assign n8846 = pi0371 & ~n8845;
  assign n8847 = ~n8842 & ~n8846;
  assign n8848 = pi0375 & n7734;
  assign n8849 = ~pi0375 & ~n7734;
  assign n8850 = ~n8848 & ~n8849;
  assign n8851 = pi0373 & ~n8850;
  assign n8852 = ~pi0373 & n8850;
  assign n8853 = ~n8851 & ~n8852;
  assign n8854 = ~n8847 & ~n8853;
  assign n8855 = ~pi0371 & ~n8845;
  assign n8856 = pi0371 & ~n8841;
  assign n8857 = ~n8855 & ~n8856;
  assign n8858 = n8853 & ~n8857;
  assign n8859 = ~pi0591 & ~n8854;
  assign n8860 = ~n8858 & n8859;
  assign n8861 = ~pi0590 & ~n8808;
  assign n8862 = ~n8860 & n8861;
  assign n8863 = ~n7425 & ~n8862;
  assign n8864 = ~n8613 & n8863;
  assign n8865 = ~pi0588 & ~n8864;
  assign n8866 = ~n8547 & n8865;
  assign n8867 = ~po1038 & ~n8312;
  assign n8868 = ~n8866 & n8867;
  assign n8869 = ~pi0217 & ~n8157;
  assign n8870 = ~n8868 & n8869;
  assign n8871 = ~n7641 & n7643;
  assign n8872 = ~n8870 & n8871;
  assign n8873 = pi1161 & ~pi1163;
  assign n8874 = n2926 & n8873;
  assign n8875 = ~pi0031 & pi1162;
  assign n8876 = n8874 & n8875;
  assign po0189 = n8872 | n8876;
  assign n8878 = n2529 & n3328;
  assign n8879 = ~pi0055 & ~pi0074;
  assign n8880 = n8878 & n8879;
  assign n8881 = n6134 & n8880;
  assign n8882 = pi0100 & n2530;
  assign n8883 = ~n6263 & ~po1057;
  assign n8884 = n6351 & n8883;
  assign n8885 = ~pi0137 & n8884;
  assign n8886 = ~pi0137 & pi0252;
  assign n8887 = pi0129 & n2521;
  assign n8888 = po1057 & ~n7474;
  assign n8889 = n6263 & ~n8888;
  assign n8890 = n8886 & n8889;
  assign n8891 = n8887 & n8890;
  assign n8892 = ~n8885 & ~n8891;
  assign n8893 = n8882 & ~n8892;
  assign n8894 = ~pi0024 & ~pi0090;
  assign n8895 = n6171 & n8894;
  assign n8896 = n2497 & n2714;
  assign n8897 = n2701 & n8896;
  assign n8898 = pi0050 & n2777;
  assign n8899 = n2495 & n8898;
  assign n8900 = ~pi0093 & n8897;
  assign n8901 = n8899 & n8900;
  assign n8902 = n8895 & n8901;
  assign n8903 = pi0829 & ~pi1093;
  assign n8904 = n2932 & n8903;
  assign po0840 = n2928 | n8904;
  assign n8906 = ~n7425 & ~po0840;
  assign n8907 = ~pi0137 & ~n8906;
  assign n8908 = n8902 & ~n8907;
  assign n8909 = ~pi0068 & ~pi0073;
  assign n8910 = n2462 & n2804;
  assign n8911 = ~pi0103 & n2471;
  assign n8912 = n8910 & n8911;
  assign n8913 = ~pi0089 & ~pi0102;
  assign n8914 = n7438 & n8913;
  assign n8915 = ~pi0045 & ~pi0048;
  assign n8916 = n2466 & n2797;
  assign n8917 = ~pi0061 & ~pi0104;
  assign n8918 = n8915 & n8917;
  assign n8919 = n8916 & n8918;
  assign n8920 = ~pi0049 & ~pi0066;
  assign n8921 = ~pi0064 & ~pi0081;
  assign n8922 = n2487 & n8921;
  assign n8923 = pi0076 & ~pi0084;
  assign n8924 = n2479 & n8923;
  assign n8925 = n8909 & n8920;
  assign n8926 = n8924 & n8925;
  assign n8927 = n8914 & n8922;
  assign n8928 = n8926 & n8927;
  assign n8929 = n8912 & n8919;
  assign n8930 = n8928 & n8929;
  assign n8931 = n2495 & n8930;
  assign n8932 = n8897 & n8931;
  assign n8933 = pi0024 & ~n8932;
  assign n8934 = ~n8898 & ~n8930;
  assign n8935 = n2499 & n2702;
  assign n8936 = ~n8934 & n8935;
  assign n8937 = ~pi0024 & ~n8936;
  assign n8938 = n2507 & n2736;
  assign n8939 = ~pi0137 & n7445;
  assign n8940 = n8938 & n8939;
  assign n8941 = ~n8906 & n8940;
  assign n8942 = ~n8933 & n8941;
  assign n8943 = ~n8937 & n8942;
  assign n8944 = ~n8908 & ~n8943;
  assign n8945 = ~pi0032 & ~n8944;
  assign n8946 = ~pi0024 & ~pi0841;
  assign n8947 = pi0032 & ~n8946;
  assign n8948 = n2710 & n8947;
  assign n8949 = ~n8945 & ~n8948;
  assign n8950 = ~n6169 & ~n8949;
  assign n8951 = ~pi0032 & ~n8902;
  assign n8952 = n6169 & ~n6173;
  assign n8953 = ~n8951 & n8952;
  assign n8954 = ~n8950 & ~n8953;
  assign n8955 = ~pi0095 & n2531;
  assign n8956 = ~n8954 & n8955;
  assign n8957 = ~n8893 & ~n8956;
  assign n8958 = n2533 & ~n8957;
  assign n8959 = ~pi0024 & n2505;
  assign n8960 = n2519 & n2705;
  assign n8961 = ~pi0051 & n8960;
  assign n8962 = n8959 & n8961;
  assign n8963 = ~po0840 & n8962;
  assign n8964 = pi0252 & ~n8888;
  assign n8965 = ~pi0087 & n2530;
  assign n8966 = pi0075 & ~pi0100;
  assign n8967 = n8965 & n8966;
  assign n8968 = ~pi0137 & n8967;
  assign n8969 = ~n6282 & n8968;
  assign n8970 = ~n8964 & n8969;
  assign n8971 = n8963 & n8970;
  assign n8972 = ~n8958 & ~n8971;
  assign po0190 = n8881 & ~n8972;
  assign n8974 = ~pi0195 & ~pi0196;
  assign n8975 = ~pi0138 & n8974;
  assign n8976 = ~pi0139 & n8975;
  assign n8977 = ~pi0118 & n8976;
  assign n8978 = ~pi0079 & n8977;
  assign n8979 = ~pi0034 & n8978;
  assign n8980 = ~pi0033 & ~n8979;
  assign n8981 = pi0149 & pi0157;
  assign n8982 = ~pi0149 & ~pi0157;
  assign n8983 = n6197 & ~n8982;
  assign n8984 = ~n8981 & n8983;
  assign n8985 = pi0232 & n8984;
  assign n8986 = pi0075 & ~n8985;
  assign n8987 = pi0100 & ~n8985;
  assign n8988 = ~n8986 & ~n8987;
  assign n8989 = ~pi0075 & ~pi0100;
  assign n8990 = n7473 & n8989;
  assign n8991 = pi0164 & n8990;
  assign n8992 = n8988 & ~n8991;
  assign n8993 = ~pi0074 & ~n8992;
  assign n8994 = pi0169 & n8990;
  assign n8995 = n8988 & ~n8994;
  assign n8996 = pi0074 & ~n8995;
  assign n8997 = ~n3328 & ~n8993;
  assign n8998 = ~n8996 & n8997;
  assign n8999 = pi0054 & ~n8992;
  assign n9000 = pi0164 & n7473;
  assign n9001 = pi0038 & n9000;
  assign n9002 = n8989 & n9001;
  assign n9003 = n8988 & ~n9002;
  assign n9004 = ~n8999 & n9003;
  assign n9005 = ~pi0074 & ~n9004;
  assign n9006 = ~n8996 & ~n9005;
  assign n9007 = ~n2529 & ~n9006;
  assign n9008 = n3328 & ~n9007;
  assign n9009 = pi0299 & ~n8984;
  assign n9010 = pi0178 & pi0183;
  assign n9011 = ~pi0178 & ~pi0183;
  assign n9012 = n6197 & ~n9011;
  assign n9013 = ~n9010 & n9012;
  assign n9014 = ~pi0299 & ~n9013;
  assign n9015 = pi0232 & ~n9009;
  assign n9016 = ~n9014 & n9015;
  assign n9017 = pi0100 & ~n9016;
  assign n9018 = pi0075 & ~n9016;
  assign n9019 = ~n9017 & ~n9018;
  assign n9020 = pi0191 & ~pi0299;
  assign n9021 = pi0169 & pi0299;
  assign n9022 = ~n9020 & ~n9021;
  assign n9023 = n8990 & ~n9022;
  assign n9024 = n9019 & ~n9023;
  assign n9025 = pi0074 & ~n9024;
  assign n9026 = ~pi0055 & ~n9025;
  assign n9027 = ~pi0186 & ~pi0299;
  assign n9028 = ~pi0164 & pi0299;
  assign n9029 = ~n9027 & ~n9028;
  assign n9030 = n7473 & n9029;
  assign n9031 = n8989 & n9030;
  assign n9032 = n9019 & ~n9031;
  assign n9033 = pi0054 & ~n9032;
  assign n9034 = pi0038 & n9030;
  assign n9035 = pi0087 & ~n9034;
  assign n9036 = pi0216 & n6379;
  assign n9037 = n6243 & ~n6392;
  assign n9038 = pi0154 & ~n9037;
  assign n9039 = n6243 & n6396;
  assign n9040 = ~pi0154 & ~n9039;
  assign n9041 = ~pi0152 & ~n9040;
  assign n9042 = ~n9038 & n9041;
  assign n9043 = n6197 & n7602;
  assign n9044 = ~n6242 & n9043;
  assign n9045 = pi0152 & pi0154;
  assign n9046 = n9044 & n9045;
  assign n9047 = ~n9042 & ~n9046;
  assign n9048 = n9036 & ~n9047;
  assign n9049 = pi0299 & ~n9048;
  assign n9050 = ~pi0176 & pi0232;
  assign n9051 = pi0224 & n6405;
  assign n9052 = n6206 & n6396;
  assign n9053 = n9051 & n9052;
  assign n9054 = ~pi0174 & n9053;
  assign n9055 = ~pi0299 & ~n9054;
  assign n9056 = n9050 & ~n9055;
  assign n9057 = pi0176 & pi0232;
  assign n9058 = n6206 & n9051;
  assign n9059 = n7602 & n9058;
  assign n9060 = pi0174 & n9059;
  assign n9061 = ~n6392 & n9051;
  assign n9062 = n6206 & n9061;
  assign n9063 = ~pi0174 & n9062;
  assign n9064 = ~pi0299 & ~n9060;
  assign n9065 = ~n9063 & n9064;
  assign n9066 = n9057 & ~n9065;
  assign n9067 = ~n9056 & ~n9066;
  assign n9068 = pi0039 & ~n9049;
  assign n9069 = ~n9067 & n9068;
  assign n9070 = n3181 & n6197;
  assign n9071 = pi0180 & n9070;
  assign n9072 = pi0090 & ~n7432;
  assign n9073 = ~pi0072 & ~pi0093;
  assign n9074 = n2707 & n9073;
  assign n9075 = ~n9072 & n9074;
  assign n9076 = ~pi0066 & ~pi0084;
  assign n9077 = ~pi0068 & n2468;
  assign n9078 = ~pi0111 & n2467;
  assign n9079 = ~pi0036 & n9077;
  assign n9080 = n9078 & n9079;
  assign n9081 = ~pi0102 & n8921;
  assign n9082 = n2466 & n9081;
  assign n9083 = n2464 & n9082;
  assign n9084 = pi0073 & ~pi0082;
  assign n9085 = n9076 & n9084;
  assign n9086 = n9080 & n9085;
  assign n9087 = n9083 & n9086;
  assign n9088 = n2477 & n9087;
  assign n9089 = n8935 & n9088;
  assign n9090 = n2487 & n9089;
  assign n9091 = n6139 & ~n9090;
  assign n9092 = n9075 & ~n9091;
  assign n9093 = n2518 & n6197;
  assign n9094 = ~pi0040 & n9093;
  assign n9095 = n9092 & n9094;
  assign n9096 = ~pi0183 & n9095;
  assign n9097 = pi0183 & n6197;
  assign n9098 = n2504 & ~n6139;
  assign n9099 = ~n9072 & n9098;
  assign n9100 = n2485 & n9083;
  assign n9101 = ~pi0060 & n9100;
  assign n9102 = pi0053 & ~n9101;
  assign n9103 = ~pi0060 & n8898;
  assign n9104 = n2719 & ~n9103;
  assign n9105 = ~n9102 & ~n9104;
  assign n9106 = n2494 & n9088;
  assign n9107 = n2487 & ~n9106;
  assign n9108 = ~n9105 & n9107;
  assign n9109 = n2720 & ~n9108;
  assign n9110 = ~pi0090 & n2717;
  assign n9111 = n2504 & n9110;
  assign n9112 = n2723 & n9111;
  assign n9113 = n2487 & n9112;
  assign n9114 = n9109 & n9113;
  assign n9115 = ~pi0070 & ~n9114;
  assign n9116 = ~n9099 & n9115;
  assign n9117 = n2519 & n3100;
  assign n9118 = ~n9116 & n9117;
  assign n9119 = ~n9115 & n9117;
  assign n9120 = ~n6487 & ~n9119;
  assign n9121 = ~pi0198 & ~n9120;
  assign n9122 = ~n9118 & ~n9121;
  assign n9123 = n9097 & ~n9122;
  assign n9124 = ~pi0174 & ~n9096;
  assign n9125 = ~n9123 & n9124;
  assign n9126 = ~n9104 & n9112;
  assign n9127 = ~pi0070 & ~n9126;
  assign n9128 = ~n9099 & n9127;
  assign n9129 = n9117 & ~n9128;
  assign n9130 = ~n6519 & ~n9129;
  assign n9131 = n6197 & ~n9130;
  assign n9132 = pi0183 & n9131;
  assign n9133 = ~n6139 & n9075;
  assign n9134 = n9094 & n9133;
  assign n9135 = ~pi0183 & n9134;
  assign n9136 = pi0174 & ~n9135;
  assign n9137 = ~n9132 & n9136;
  assign n9138 = ~n9125 & ~n9137;
  assign n9139 = pi0193 & ~n9138;
  assign n9140 = ~pi0040 & n6197;
  assign n9141 = ~pi0090 & n9074;
  assign n9142 = n9090 & n9141;
  assign n9143 = n2518 & n9142;
  assign n9144 = n9140 & n9143;
  assign n9145 = ~pi0174 & ~pi0183;
  assign n9146 = n9144 & n9145;
  assign n9147 = ~n6519 & ~n9119;
  assign n9148 = ~pi0174 & n9147;
  assign n9149 = n9117 & ~n9127;
  assign n9150 = ~n6519 & ~n9149;
  assign n9151 = pi0174 & n9150;
  assign n9152 = n9097 & ~n9151;
  assign n9153 = ~n9148 & n9152;
  assign n9154 = ~pi0193 & ~n9146;
  assign n9155 = ~n9153 & n9154;
  assign n9156 = ~n9139 & ~n9155;
  assign n9157 = ~pi0299 & ~n9071;
  assign n9158 = ~n9156 & n9157;
  assign n9159 = ~pi0039 & pi0232;
  assign n9160 = pi0158 & n9070;
  assign n9161 = pi0172 & n9118;
  assign n9162 = ~n6488 & ~n9119;
  assign n9163 = ~pi0152 & n9162;
  assign n9164 = ~n9161 & n9163;
  assign n9165 = pi0172 & n9129;
  assign n9166 = ~n6488 & ~n9149;
  assign n9167 = pi0152 & ~n9165;
  assign n9168 = n9166 & n9167;
  assign n9169 = pi0149 & n6197;
  assign n9170 = ~n9168 & n9169;
  assign n9171 = ~n9164 & n9170;
  assign n9172 = ~pi0152 & n9095;
  assign n9173 = ~n9134 & ~n9172;
  assign n9174 = pi0172 & ~n9173;
  assign n9175 = ~pi0152 & ~pi0172;
  assign n9176 = n9144 & n9175;
  assign n9177 = ~n9174 & ~n9176;
  assign n9178 = ~pi0149 & ~n9177;
  assign n9179 = pi0299 & ~n9160;
  assign n9180 = ~n9178 & n9179;
  assign n9181 = ~n9171 & n9180;
  assign n9182 = n9159 & ~n9181;
  assign n9183 = ~n9158 & n9182;
  assign n9184 = ~n9069 & ~n9183;
  assign n9185 = ~pi0038 & ~n9184;
  assign n9186 = pi0299 & n7473;
  assign n9187 = ~n6135 & n9186;
  assign n9188 = ~pi0186 & ~n9187;
  assign n9189 = ~n6284 & n7473;
  assign n9190 = pi0186 & ~n9189;
  assign n9191 = pi0164 & ~n9190;
  assign n9192 = ~n9188 & n9191;
  assign n9193 = ~pi0299 & n7473;
  assign n9194 = ~n6135 & n9193;
  assign n9195 = ~pi0164 & pi0186;
  assign n9196 = n9194 & n9195;
  assign n9197 = ~n9192 & ~n9196;
  assign n9198 = pi0038 & ~n9197;
  assign n9199 = ~pi0087 & ~n9198;
  assign n9200 = ~n9185 & n9199;
  assign n9201 = ~pi0100 & ~n9035;
  assign n9202 = ~n9200 & n9201;
  assign n9203 = ~n9017 & ~n9202;
  assign n9204 = n2569 & ~n9203;
  assign n9205 = ~pi0075 & pi0092;
  assign n9206 = ~pi0100 & n9034;
  assign n9207 = ~n9017 & ~n9206;
  assign n9208 = ~pi0038 & ~pi0087;
  assign n9209 = pi0232 & ~n3383;
  assign n9210 = ~pi0176 & ~pi0299;
  assign n9211 = n6197 & ~n9210;
  assign n9212 = n9209 & n9211;
  assign n9213 = ~pi0100 & n9208;
  assign n9214 = n9212 & n9213;
  assign n9215 = n6135 & n9214;
  assign n9216 = n9207 & ~n9215;
  assign n9217 = n9205 & ~n9216;
  assign n9218 = ~n9018 & ~n9217;
  assign n9219 = ~n9204 & n9218;
  assign n9220 = ~pi0054 & ~n9219;
  assign n9221 = ~n9033 & ~n9220;
  assign n9222 = ~pi0074 & ~n9221;
  assign n9223 = n9026 & ~n9222;
  assign n9224 = pi0055 & ~n8996;
  assign n9225 = ~pi0092 & ~n8986;
  assign n9226 = pi0038 & ~n9000;
  assign n9227 = n2568 & ~n9226;
  assign n9228 = pi0149 & n7473;
  assign n9229 = n6135 & n9228;
  assign n9230 = ~pi0038 & ~n9229;
  assign n9231 = n9227 & ~n9230;
  assign n9232 = n8161 & n9001;
  assign n9233 = ~n8987 & ~n9232;
  assign n9234 = ~n9231 & n9233;
  assign n9235 = ~pi0075 & ~n9234;
  assign n9236 = n9225 & ~n9235;
  assign n9237 = pi0092 & n9003;
  assign n9238 = ~pi0054 & ~n9237;
  assign n9239 = ~n9236 & n9238;
  assign n9240 = ~n8999 & ~n9239;
  assign n9241 = ~pi0074 & ~n9240;
  assign n9242 = n9224 & ~n9241;
  assign n9243 = n2529 & ~n9242;
  assign n9244 = ~n9223 & n9243;
  assign n9245 = n9008 & ~n9244;
  assign n9246 = ~n8998 & ~n9245;
  assign n9247 = n8980 & ~n9246;
  assign n9248 = ~pi0040 & n2487;
  assign n9249 = ~pi0038 & n9248;
  assign n9250 = n8989 & n9249;
  assign n9251 = n2532 & n9250;
  assign n9252 = ~n2529 & n9251;
  assign n9253 = n2716 & n2720;
  assign n9254 = ~pi0053 & n9253;
  assign n9255 = n9101 & n9254;
  assign n9256 = ~pi0058 & n9255;
  assign n9257 = n7445 & n9256;
  assign n9258 = ~pi0032 & n2508;
  assign n9259 = n9257 & n9258;
  assign n9260 = ~pi0095 & n9259;
  assign n9261 = ~pi0039 & ~n9228;
  assign n9262 = n9260 & n9261;
  assign n9263 = n9248 & ~n9262;
  assign n9264 = ~pi0038 & ~n9263;
  assign n9265 = n9227 & ~n9264;
  assign n9266 = ~pi0038 & ~n9248;
  assign n9267 = ~pi0100 & ~n9266;
  assign n9268 = ~n9226 & n9267;
  assign n9269 = pi0087 & n9268;
  assign n9270 = ~n8987 & ~n9269;
  assign n9271 = ~n9265 & n9270;
  assign n9272 = ~pi0075 & ~n9271;
  assign n9273 = n9225 & ~n9272;
  assign n9274 = ~pi0075 & n9268;
  assign n9275 = pi0092 & n8988;
  assign n9276 = ~n9274 & n9275;
  assign n9277 = ~pi0054 & ~n9276;
  assign n9278 = ~n9273 & n9277;
  assign n9279 = ~n8999 & ~n9278;
  assign n9280 = ~pi0074 & ~n9279;
  assign n9281 = n9224 & ~n9280;
  assign n9282 = n2609 & n9260;
  assign n9283 = ~n9212 & n9282;
  assign n9284 = n2608 & n9248;
  assign n9285 = ~n9283 & n9284;
  assign n9286 = n9207 & ~n9285;
  assign n9287 = n9205 & ~n9286;
  assign n9288 = pi0087 & ~n9284;
  assign n9289 = n9207 & n9288;
  assign n9290 = ~n9036 & n9248;
  assign n9291 = pi0299 & ~n9290;
  assign n9292 = n6383 & ~n6395;
  assign n9293 = n6212 & n9292;
  assign n9294 = ~n6188 & ~n9293;
  assign n9295 = n9260 & ~n9294;
  assign n9296 = n6198 & n9295;
  assign n9297 = n9248 & ~n9296;
  assign n9298 = n6197 & n9295;
  assign n9299 = n9248 & ~n9298;
  assign n9300 = ~n6242 & ~n9299;
  assign n9301 = n9297 & ~n9300;
  assign n9302 = n9291 & ~n9301;
  assign n9303 = ~n9051 & n9248;
  assign n9304 = ~n9297 & ~n9303;
  assign n9305 = ~n6205 & ~n9299;
  assign n9306 = ~n9303 & n9305;
  assign n9307 = ~n9304 & ~n9306;
  assign n9308 = ~pi0299 & ~n9307;
  assign n9309 = ~n9302 & ~n9308;
  assign n9310 = ~pi0232 & ~n9309;
  assign n9311 = n9260 & n9293;
  assign n9312 = n6197 & n9311;
  assign n9313 = n9248 & ~n9312;
  assign n9314 = ~n6205 & ~n9313;
  assign n9315 = ~n9303 & n9314;
  assign n9316 = pi0174 & n9315;
  assign n9317 = ~n9304 & ~n9316;
  assign n9318 = ~pi0299 & ~n9317;
  assign n9319 = n9248 & ~n9311;
  assign n9320 = n6243 & ~n9319;
  assign n9321 = pi0152 & n9320;
  assign n9322 = n9297 & ~n9321;
  assign n9323 = pi0154 & ~n9322;
  assign n9324 = n6188 & n9260;
  assign n9325 = ~n6227 & n9324;
  assign n9326 = n9248 & ~n9325;
  assign n9327 = n6197 & n9326;
  assign n9328 = ~pi0152 & n9327;
  assign n9329 = ~pi0154 & ~n9301;
  assign n9330 = ~n9328 & n9329;
  assign n9331 = n9036 & ~n9323;
  assign n9332 = ~n9330 & n9331;
  assign n9333 = n9291 & ~n9332;
  assign n9334 = ~n9318 & ~n9333;
  assign n9335 = n6206 & n9324;
  assign n9336 = n9051 & n9248;
  assign n9337 = ~n9335 & n9336;
  assign n9338 = ~n9303 & ~n9337;
  assign n9339 = ~pi0299 & n9338;
  assign n9340 = n9334 & ~n9339;
  assign n9341 = n9050 & ~n9340;
  assign n9342 = n9057 & ~n9334;
  assign n9343 = pi0039 & ~n9310;
  assign n9344 = ~n9342 & n9343;
  assign n9345 = ~n9341 & n9344;
  assign n9346 = pi0095 & ~n9248;
  assign n9347 = ~n2442 & ~n9346;
  assign n9348 = ~pi0040 & ~pi0479;
  assign n9349 = n2487 & ~n9259;
  assign n9350 = n9348 & n9349;
  assign n9351 = ~n9347 & ~n9350;
  assign n9352 = pi0032 & ~n9248;
  assign n9353 = n2487 & ~n2506;
  assign n9354 = n2487 & ~n9257;
  assign n9355 = pi0070 & ~n9354;
  assign n9356 = n2487 & ~n9255;
  assign n9357 = pi0058 & ~n9356;
  assign n9358 = n2487 & ~n2716;
  assign n9359 = ~n2487 & ~n2720;
  assign n9360 = n2716 & ~n9359;
  assign n9361 = ~n9109 & n9360;
  assign n9362 = ~pi0058 & ~n9358;
  assign n9363 = ~n9361 & n9362;
  assign n9364 = ~n9357 & ~n9363;
  assign n9365 = ~pi0090 & ~n9364;
  assign n9366 = ~pi0841 & n9256;
  assign n9367 = n2487 & ~n9366;
  assign n9368 = pi0090 & ~n9367;
  assign n9369 = n2504 & ~n9368;
  assign n9370 = ~n9365 & n9369;
  assign n9371 = n2487 & ~n2504;
  assign n9372 = ~pi0070 & ~n9371;
  assign n9373 = ~n9370 & n9372;
  assign n9374 = ~n9355 & ~n9373;
  assign n9375 = ~pi0051 & ~n9374;
  assign n9376 = pi0051 & ~n2487;
  assign n9377 = n2506 & ~n9376;
  assign n9378 = ~n9375 & n9377;
  assign n9379 = ~n9353 & ~n9378;
  assign n9380 = ~pi0040 & ~n9379;
  assign n9381 = ~pi0032 & ~n9380;
  assign n9382 = ~n9352 & ~n9381;
  assign n9383 = ~pi0095 & ~n9382;
  assign n9384 = ~n9351 & ~n9383;
  assign n9385 = n9141 & n9366;
  assign n9386 = n9248 & ~n9385;
  assign n9387 = pi0032 & ~n9386;
  assign n9388 = ~n9381 & ~n9387;
  assign n9389 = ~pi0095 & ~n9388;
  assign n9390 = ~pi0198 & n9389;
  assign n9391 = n9384 & ~n9390;
  assign n9392 = ~n6197 & n9391;
  assign n9393 = n9105 & n9253;
  assign n9394 = n2487 & ~n9393;
  assign n9395 = ~pi0058 & ~n9394;
  assign n9396 = ~n9357 & ~n9395;
  assign n9397 = ~pi0090 & ~n9396;
  assign n9398 = n9369 & ~n9397;
  assign n9399 = n9372 & ~n9398;
  assign n9400 = ~n9355 & ~n9399;
  assign n9401 = ~pi0051 & ~n9400;
  assign n9402 = n9377 & ~n9401;
  assign n9403 = ~n9353 & ~n9402;
  assign n9404 = ~pi0040 & ~n9403;
  assign n9405 = ~pi0032 & ~n9404;
  assign n9406 = ~n9387 & ~n9405;
  assign n9407 = ~pi0095 & ~n9406;
  assign n9408 = ~pi0198 & n9407;
  assign n9409 = n6197 & ~n9346;
  assign n9410 = ~n9352 & ~n9405;
  assign n9411 = ~pi0095 & ~n9410;
  assign n9412 = n9409 & ~n9411;
  assign n9413 = ~n9408 & n9412;
  assign n9414 = ~n9392 & ~n9413;
  assign n9415 = ~pi0183 & ~n9414;
  assign n9416 = ~pi0040 & ~n9352;
  assign n9417 = n2487 & ~n6170;
  assign n9418 = ~pi0032 & ~n9417;
  assign n9419 = pi0093 & ~n2487;
  assign n9420 = n6170 & ~n9419;
  assign n9421 = n2487 & ~n9357;
  assign n9422 = ~pi0090 & ~n9421;
  assign n9423 = ~n9368 & ~n9422;
  assign n9424 = ~pi0093 & ~n9423;
  assign n9425 = n9420 & ~n9424;
  assign n9426 = n9418 & ~n9425;
  assign n9427 = n9416 & ~n9426;
  assign n9428 = ~pi0095 & ~n9427;
  assign n9429 = n9409 & ~n9428;
  assign n9430 = ~n9392 & ~n9429;
  assign n9431 = pi0183 & ~n9430;
  assign n9432 = ~n9415 & ~n9431;
  assign n9433 = ~pi0095 & n9432;
  assign n9434 = ~pi0174 & ~n9351;
  assign n9435 = ~n9433 & n9434;
  assign n9436 = ~n9097 & ~n9391;
  assign n9437 = ~pi0090 & n9089;
  assign n9438 = n9423 & ~n9437;
  assign n9439 = ~pi0093 & ~n9438;
  assign n9440 = n9420 & ~n9439;
  assign n9441 = n9418 & ~n9440;
  assign n9442 = n9416 & ~n9441;
  assign n9443 = ~pi0095 & ~n9442;
  assign n9444 = ~n9351 & ~n9443;
  assign n9445 = n6197 & ~n9444;
  assign n9446 = pi0183 & n9445;
  assign n9447 = pi0174 & ~n9446;
  assign n9448 = ~n9436 & n9447;
  assign n9449 = ~pi0180 & ~n9448;
  assign n9450 = ~n9435 & n9449;
  assign n9451 = ~pi0174 & ~n9432;
  assign n9452 = n9409 & ~n9443;
  assign n9453 = ~n9392 & ~n9452;
  assign n9454 = pi0183 & ~n9453;
  assign n9455 = ~n9346 & ~n9383;
  assign n9456 = ~n9390 & n9455;
  assign n9457 = n9140 & n9456;
  assign n9458 = ~n9392 & ~n9457;
  assign n9459 = ~pi0183 & ~n9458;
  assign n9460 = ~n9454 & ~n9459;
  assign n9461 = pi0174 & ~n9460;
  assign n9462 = pi0180 & ~n9451;
  assign n9463 = ~n9461 & n9462;
  assign n9464 = ~n9450 & ~n9463;
  assign n9465 = ~pi0193 & ~n9464;
  assign n9466 = ~pi0040 & ~n2487;
  assign n9467 = pi0032 & ~n9466;
  assign n9468 = n2461 & n2504;
  assign n9469 = ~n2487 & ~n9468;
  assign n9470 = n7445 & n9363;
  assign n9471 = ~n9469 & ~n9470;
  assign n9472 = ~pi0070 & ~n9471;
  assign n9473 = ~n9355 & ~n9472;
  assign n9474 = ~pi0051 & ~n9473;
  assign n9475 = n9377 & ~n9474;
  assign n9476 = ~pi0040 & ~n9353;
  assign n9477 = ~n9475 & n9476;
  assign n9478 = ~pi0032 & ~n9477;
  assign n9479 = ~n9467 & ~n9478;
  assign n9480 = ~n2736 & ~n9248;
  assign n9481 = ~n9479 & ~n9480;
  assign n9482 = ~pi0095 & ~n9481;
  assign n9483 = ~n9351 & ~n9482;
  assign n9484 = ~n9346 & ~n9482;
  assign n9485 = pi0095 & ~n9466;
  assign n9486 = ~pi0040 & ~n9386;
  assign n9487 = pi0032 & ~n9486;
  assign n9488 = ~n9478 & ~n9487;
  assign n9489 = ~pi0095 & ~n9488;
  assign n9490 = ~n9485 & ~n9489;
  assign n9491 = n9484 & ~n9490;
  assign n9492 = ~pi0198 & ~n9491;
  assign n9493 = n6197 & ~n9492;
  assign n9494 = n6197 & ~n9248;
  assign n9495 = ~n9493 & ~n9494;
  assign n9496 = n9483 & ~n9495;
  assign n9497 = ~n9392 & ~n9496;
  assign n9498 = ~pi0183 & ~n9497;
  assign n9499 = n2704 & n6170;
  assign n9500 = n8935 & n9499;
  assign n9501 = ~pi0032 & n9500;
  assign n9502 = n9088 & n9501;
  assign n9503 = n9248 & ~n9502;
  assign n9504 = ~pi0095 & ~n9503;
  assign n9505 = n6197 & ~n9504;
  assign n9506 = ~n9351 & n9505;
  assign n9507 = ~n9392 & ~n9506;
  assign n9508 = pi0183 & ~n9507;
  assign n9509 = pi0174 & ~n9508;
  assign n9510 = ~n9498 & n9509;
  assign n9511 = ~n6197 & ~n9391;
  assign n9512 = n7445 & n9395;
  assign n9513 = ~n9469 & ~n9512;
  assign n9514 = ~pi0070 & ~n9513;
  assign n9515 = ~n9355 & ~n9514;
  assign n9516 = ~pi0051 & ~n9515;
  assign n9517 = n9377 & ~n9516;
  assign n9518 = ~n9353 & ~n9517;
  assign n9519 = ~pi0040 & ~n9518;
  assign n9520 = ~pi0032 & ~n9519;
  assign n9521 = ~n9352 & ~n9520;
  assign n9522 = ~pi0095 & ~n9521;
  assign n9523 = ~n9351 & ~n9522;
  assign n9524 = ~n9387 & ~n9520;
  assign n9525 = ~pi0095 & ~n9524;
  assign n9526 = ~pi0198 & n9525;
  assign n9527 = n9523 & ~n9526;
  assign n9528 = n6197 & ~n9527;
  assign n9529 = ~n9511 & ~n9528;
  assign n9530 = ~pi0183 & n9529;
  assign n9531 = ~pi0095 & ~n9248;
  assign n9532 = ~n9351 & ~n9531;
  assign n9533 = n6197 & n9532;
  assign n9534 = ~n9392 & ~n9533;
  assign n9535 = pi0183 & ~n9534;
  assign n9536 = ~pi0174 & ~n9530;
  assign n9537 = ~n9535 & n9536;
  assign n9538 = ~pi0180 & ~n9537;
  assign n9539 = ~n9510 & n9538;
  assign n9540 = n9409 & ~n9504;
  assign n9541 = ~n9392 & ~n9540;
  assign n9542 = pi0183 & ~n9541;
  assign n9543 = n9484 & n9493;
  assign n9544 = ~n9392 & ~n9543;
  assign n9545 = ~pi0183 & ~n9544;
  assign n9546 = pi0174 & ~n9542;
  assign n9547 = ~n9545 & n9546;
  assign n9548 = ~n9494 & ~n9511;
  assign n9549 = pi0183 & n9548;
  assign n9550 = ~pi0040 & n9518;
  assign n9551 = ~pi0032 & ~n9550;
  assign n9552 = ~n9467 & ~n9551;
  assign n9553 = ~pi0095 & ~n9552;
  assign n9554 = ~n9485 & ~n9553;
  assign n9555 = pi0198 & ~n9554;
  assign n9556 = ~n9487 & ~n9551;
  assign n9557 = ~pi0095 & ~n9556;
  assign n9558 = ~n9485 & ~n9557;
  assign n9559 = ~pi0198 & ~n9558;
  assign n9560 = ~n9555 & ~n9559;
  assign n9561 = n9140 & ~n9560;
  assign n9562 = ~n9392 & ~n9561;
  assign n9563 = ~pi0183 & ~n9562;
  assign n9564 = ~pi0174 & ~n9549;
  assign n9565 = ~n9563 & n9564;
  assign n9566 = pi0180 & ~n9547;
  assign n9567 = ~n9565 & n9566;
  assign n9568 = pi0193 & ~n9539;
  assign n9569 = ~n9567 & n9568;
  assign n9570 = ~n9465 & ~n9569;
  assign n9571 = ~pi0299 & ~n9570;
  assign n9572 = pi0158 & pi0299;
  assign n9573 = ~pi0210 & n9389;
  assign n9574 = n9384 & ~n9573;
  assign n9575 = ~n6197 & n9574;
  assign n9576 = ~pi0210 & n9407;
  assign n9577 = n9412 & ~n9576;
  assign n9578 = ~n9575 & ~n9577;
  assign n9579 = ~pi0152 & ~n9578;
  assign n9580 = ~n6197 & ~n9574;
  assign n9581 = n9455 & ~n9573;
  assign n9582 = n6197 & ~n9581;
  assign n9583 = ~n9580 & ~n9582;
  assign n9584 = pi0152 & n9583;
  assign n9585 = ~pi0172 & ~n9579;
  assign n9586 = ~n9584 & n9585;
  assign n9587 = ~n9346 & ~n9525;
  assign n9588 = ~pi0210 & ~n9587;
  assign n9589 = n6197 & ~n9588;
  assign n9590 = ~n9346 & ~n9522;
  assign n9591 = n9589 & n9590;
  assign n9592 = ~n9575 & ~n9591;
  assign n9593 = ~pi0152 & ~n9592;
  assign n9594 = ~pi0210 & ~n9491;
  assign n9595 = n6197 & ~n9594;
  assign n9596 = n9484 & n9595;
  assign n9597 = ~n9575 & ~n9596;
  assign n9598 = pi0152 & ~n9597;
  assign n9599 = pi0172 & ~n9593;
  assign n9600 = ~n9598 & n9599;
  assign n9601 = ~n9586 & ~n9600;
  assign n9602 = n9572 & ~n9601;
  assign n9603 = ~pi0158 & pi0299;
  assign n9604 = ~n9351 & ~n9411;
  assign n9605 = ~n9576 & n9604;
  assign n9606 = n6197 & n9605;
  assign n9607 = ~pi0152 & ~n9606;
  assign n9608 = pi0152 & ~n9574;
  assign n9609 = ~pi0172 & ~n9607;
  assign n9610 = ~n9608 & n9609;
  assign n9611 = ~n9494 & ~n9595;
  assign n9612 = n9483 & ~n9611;
  assign n9613 = pi0152 & ~n9612;
  assign n9614 = ~n9494 & ~n9589;
  assign n9615 = n9523 & ~n9614;
  assign n9616 = ~pi0152 & ~n9615;
  assign n9617 = pi0172 & ~n9616;
  assign n9618 = ~n9613 & n9617;
  assign n9619 = ~n9575 & n9603;
  assign n9620 = ~n9610 & n9619;
  assign n9621 = ~n9618 & n9620;
  assign n9622 = ~pi0149 & ~n9621;
  assign n9623 = ~n9602 & n9622;
  assign n9624 = ~n9452 & ~n9575;
  assign n9625 = pi0152 & ~n9624;
  assign n9626 = ~n9429 & ~n9575;
  assign n9627 = ~pi0152 & ~n9626;
  assign n9628 = ~pi0172 & ~n9625;
  assign n9629 = ~n9627 & n9628;
  assign n9630 = ~n9540 & ~n9575;
  assign n9631 = pi0152 & ~n9630;
  assign n9632 = ~n9494 & ~n9580;
  assign n9633 = ~pi0152 & n9632;
  assign n9634 = pi0172 & ~n9631;
  assign n9635 = ~n9633 & n9634;
  assign n9636 = ~n9629 & ~n9635;
  assign n9637 = n9572 & ~n9636;
  assign n9638 = ~n9506 & ~n9575;
  assign n9639 = pi0152 & ~n9638;
  assign n9640 = ~n9533 & ~n9575;
  assign n9641 = ~pi0152 & ~n9640;
  assign n9642 = pi0172 & ~n9639;
  assign n9643 = ~n9641 & n9642;
  assign n9644 = ~n9351 & ~n9428;
  assign n9645 = n6197 & ~n9644;
  assign n9646 = ~n9580 & ~n9645;
  assign n9647 = ~pi0152 & n9646;
  assign n9648 = ~n9445 & ~n9580;
  assign n9649 = pi0152 & n9648;
  assign n9650 = ~pi0172 & ~n9647;
  assign n9651 = ~n9649 & n9650;
  assign n9652 = ~n9643 & ~n9651;
  assign n9653 = n9603 & ~n9652;
  assign n9654 = pi0149 & ~n9637;
  assign n9655 = ~n9653 & n9654;
  assign n9656 = ~n9623 & ~n9655;
  assign n9657 = ~n9571 & ~n9656;
  assign n9658 = pi0232 & ~n9657;
  assign n9659 = ~n6169 & n9389;
  assign n9660 = n9384 & ~n9659;
  assign n9661 = ~pi0232 & ~n9660;
  assign n9662 = ~pi0039 & ~n9661;
  assign n9663 = ~n9658 & n9662;
  assign n9664 = ~n9345 & ~n9663;
  assign n9665 = ~pi0038 & ~n9664;
  assign n9666 = ~n9198 & ~n9665;
  assign n9667 = ~pi0100 & ~n9666;
  assign n9668 = ~pi0087 & ~n9017;
  assign n9669 = ~n9667 & n9668;
  assign n9670 = n2569 & ~n9289;
  assign n9671 = ~n9669 & n9670;
  assign n9672 = ~n9018 & ~n9287;
  assign n9673 = ~n9671 & n9672;
  assign n9674 = ~pi0054 & ~n9673;
  assign n9675 = ~n9033 & ~n9674;
  assign n9676 = ~pi0074 & ~n9675;
  assign n9677 = n9026 & ~n9676;
  assign n9678 = n2529 & ~n9281;
  assign n9679 = ~n9677 & n9678;
  assign n9680 = n9008 & ~n9252;
  assign n9681 = ~n9679 & n9680;
  assign n9682 = ~n8998 & ~n9681;
  assign n9683 = ~n8980 & ~n9682;
  assign n9684 = ~pi0954 & ~n9247;
  assign n9685 = ~n9683 & n9684;
  assign n9686 = pi0033 & ~n9246;
  assign n9687 = ~pi0033 & ~n9682;
  assign n9688 = pi0954 & ~n9686;
  assign n9689 = ~n9687 & n9688;
  assign po0191 = ~n9685 & ~n9689;
  assign n9691 = pi0197 & n8982;
  assign n9692 = ~pi0197 & ~n8982;
  assign n9693 = ~n9691 & ~n9692;
  assign n9694 = pi0162 & n6197;
  assign n9695 = n9693 & ~n9694;
  assign n9696 = n9691 & n9694;
  assign n9697 = ~pi0162 & ~pi0197;
  assign n9698 = n8983 & ~n9697;
  assign n9699 = n6197 & ~n9698;
  assign n9700 = ~n9696 & n9699;
  assign n9701 = ~n9693 & ~n9700;
  assign n9702 = ~n9695 & ~n9701;
  assign n9703 = pi0232 & n9702;
  assign n9704 = ~n8989 & n9703;
  assign n9705 = pi0167 & n7473;
  assign n9706 = n8989 & n9705;
  assign n9707 = ~n9704 & ~n9706;
  assign n9708 = ~pi0074 & n9707;
  assign n9709 = pi0148 & n8990;
  assign n9710 = pi0074 & ~n9709;
  assign n9711 = ~n9704 & n9710;
  assign n9712 = ~n9708 & ~n9711;
  assign n9713 = ~n3328 & n9712;
  assign n9714 = ~pi0054 & ~n9704;
  assign n9715 = pi0038 & n9706;
  assign n9716 = n9714 & ~n9715;
  assign n9717 = ~pi0074 & n9716;
  assign n9718 = n9712 & ~n9717;
  assign n9719 = ~n2529 & ~n9718;
  assign n9720 = n3328 & ~n9719;
  assign n9721 = pi0140 & pi0145;
  assign n9722 = n9011 & ~n9721;
  assign n9723 = ~pi0140 & ~pi0145;
  assign n9724 = n6197 & ~n9723;
  assign n9725 = n9722 & n9724;
  assign n9726 = ~n9721 & ~n9723;
  assign n9727 = n9012 & ~n9726;
  assign n9728 = ~pi0299 & ~n9725;
  assign n9729 = ~n9727 & n9728;
  assign n9730 = pi0299 & ~n9702;
  assign n9731 = pi0232 & ~n9729;
  assign n9732 = ~n9730 & n9731;
  assign n9733 = pi0100 & ~n9732;
  assign n9734 = pi0075 & ~n9732;
  assign n9735 = ~n9733 & ~n9734;
  assign n9736 = pi0141 & ~pi0299;
  assign n9737 = pi0148 & pi0299;
  assign n9738 = ~n9736 & ~n9737;
  assign n9739 = n7473 & ~n9738;
  assign n9740 = n8989 & ~n9739;
  assign n9741 = n9735 & ~n9740;
  assign n9742 = pi0074 & ~n9741;
  assign n9743 = ~pi0055 & ~n9742;
  assign n9744 = pi0188 & ~pi0299;
  assign n9745 = pi0167 & pi0299;
  assign n9746 = ~n9744 & ~n9745;
  assign n9747 = n7473 & ~n9746;
  assign n9748 = ~pi0100 & ~n9747;
  assign n9749 = ~pi0075 & n9748;
  assign n9750 = n9735 & ~n9749;
  assign n9751 = pi0054 & ~n9750;
  assign n9752 = ~pi0188 & ~n9187;
  assign n9753 = pi0188 & n9194;
  assign n9754 = ~pi0167 & ~n9753;
  assign n9755 = pi0167 & pi0188;
  assign n9756 = ~n9189 & n9755;
  assign n9757 = ~n9752 & ~n9756;
  assign n9758 = ~n9754 & n9757;
  assign n9759 = pi0038 & ~n9758;
  assign n9760 = ~pi0038 & pi0155;
  assign n9761 = pi0161 & ~n9044;
  assign n9762 = ~pi0161 & ~n9037;
  assign n9763 = n9036 & ~n9762;
  assign n9764 = ~n9761 & n9763;
  assign n9765 = n9760 & ~n9764;
  assign n9766 = ~pi0038 & ~pi0155;
  assign n9767 = ~pi0161 & n9036;
  assign n9768 = n9039 & n9767;
  assign n9769 = n9766 & ~n9768;
  assign n9770 = ~n9765 & ~n9769;
  assign n9771 = pi0299 & ~n9770;
  assign n9772 = ~pi0177 & ~pi0299;
  assign n9773 = ~pi0144 & n9053;
  assign n9774 = n9772 & ~n9773;
  assign n9775 = ~pi0144 & n9062;
  assign n9776 = pi0177 & ~pi0299;
  assign n9777 = pi0144 & n9059;
  assign n9778 = n9776 & ~n9777;
  assign n9779 = ~n9775 & n9778;
  assign n9780 = pi0232 & ~n9774;
  assign n9781 = ~n9779 & n9780;
  assign n9782 = ~pi0038 & ~n9781;
  assign n9783 = ~n9771 & ~n9782;
  assign n9784 = pi0039 & ~n9783;
  assign n9785 = ~pi0146 & ~n9095;
  assign n9786 = pi0146 & ~n9144;
  assign n9787 = ~pi0161 & ~n9786;
  assign n9788 = ~n9785 & n9787;
  assign n9789 = ~pi0146 & pi0161;
  assign n9790 = n9134 & n9789;
  assign n9791 = ~n9788 & ~n9790;
  assign n9792 = ~pi0162 & ~n9791;
  assign n9793 = ~pi0159 & pi0299;
  assign n9794 = pi0159 & pi0299;
  assign n9795 = ~pi0162 & n9070;
  assign n9796 = n9794 & ~n9795;
  assign n9797 = ~n9793 & ~n9796;
  assign n9798 = ~n9694 & ~n9797;
  assign n9799 = pi0159 & n3181;
  assign n9800 = ~pi0146 & n9129;
  assign n9801 = n9166 & ~n9800;
  assign n9802 = pi0161 & ~n9801;
  assign n9803 = ~pi0146 & n9118;
  assign n9804 = n9162 & ~n9803;
  assign n9805 = ~pi0161 & ~n9804;
  assign n9806 = pi0299 & ~n9799;
  assign n9807 = ~n9802 & n9806;
  assign n9808 = ~n9805 & n9807;
  assign n9809 = ~n9798 & ~n9808;
  assign n9810 = ~n9792 & ~n9809;
  assign n9811 = pi0181 & n9070;
  assign n9812 = pi0140 & ~n6197;
  assign n9813 = ~pi0142 & n9134;
  assign n9814 = ~pi0140 & ~n9813;
  assign n9815 = ~pi0142 & n9129;
  assign n9816 = pi0140 & ~n9815;
  assign n9817 = n9150 & n9816;
  assign n9818 = ~n9814 & ~n9817;
  assign n9819 = pi0144 & ~n9818;
  assign n9820 = ~pi0142 & n9095;
  assign n9821 = pi0142 & n9144;
  assign n9822 = ~pi0140 & ~n9821;
  assign n9823 = ~n9820 & n9822;
  assign n9824 = ~pi0142 & n9118;
  assign n9825 = pi0140 & n9147;
  assign n9826 = ~n9824 & n9825;
  assign n9827 = ~n9823 & ~n9826;
  assign n9828 = ~pi0144 & ~n9827;
  assign n9829 = ~n9812 & ~n9819;
  assign n9830 = ~n9828 & n9829;
  assign n9831 = ~pi0299 & ~n9811;
  assign n9832 = ~n9830 & n9831;
  assign n9833 = pi0232 & ~n9810;
  assign n9834 = ~n9832 & n9833;
  assign n9835 = n2530 & ~n9834;
  assign n9836 = ~n9759 & ~n9784;
  assign n9837 = ~n9835 & n9836;
  assign n9838 = ~pi0100 & ~n9837;
  assign n9839 = ~n9733 & ~n9838;
  assign n9840 = ~pi0087 & ~n9839;
  assign n9841 = ~n2608 & ~n9748;
  assign n9842 = ~n9733 & n9841;
  assign n9843 = pi0087 & ~n9842;
  assign n9844 = ~n9840 & ~n9843;
  assign n9845 = n2569 & ~n9844;
  assign n9846 = pi0038 & ~n9746;
  assign n9847 = pi0155 & pi0299;
  assign n9848 = ~n9776 & ~n9847;
  assign n9849 = n2530 & ~n9848;
  assign n9850 = n2512 & n9849;
  assign n9851 = ~n9846 & ~n9850;
  assign n9852 = n7473 & ~n9851;
  assign n9853 = ~pi0100 & ~n9852;
  assign n9854 = ~n9733 & ~n9853;
  assign n9855 = ~pi0087 & ~n9854;
  assign n9856 = ~n9843 & ~n9855;
  assign n9857 = n9205 & ~n9856;
  assign n9858 = ~n9734 & ~n9857;
  assign n9859 = ~n9845 & n9858;
  assign n9860 = ~pi0054 & ~n9859;
  assign n9861 = ~n9751 & ~n9860;
  assign n9862 = ~pi0074 & ~n9861;
  assign n9863 = n9743 & ~n9862;
  assign n9864 = pi0055 & ~n9711;
  assign n9865 = pi0054 & n9707;
  assign n9866 = pi0038 & n9705;
  assign n9867 = ~pi0092 & pi0162;
  assign n9868 = n9159 & n9867;
  assign n9869 = n9208 & n9868;
  assign n9870 = n6222 & n9869;
  assign n9871 = ~n9866 & ~n9870;
  assign n9872 = n8989 & ~n9871;
  assign n9873 = n9714 & ~n9872;
  assign n9874 = ~n9865 & ~n9873;
  assign n9875 = ~pi0074 & ~n9874;
  assign n9876 = n9864 & ~n9875;
  assign n9877 = n2529 & ~n9876;
  assign n9878 = ~n9863 & n9877;
  assign n9879 = n9720 & ~n9878;
  assign n9880 = ~n9713 & ~n9879;
  assign n9881 = pi0034 & n9880;
  assign n9882 = ~n2529 & ~n9251;
  assign n9883 = n3328 & ~n9882;
  assign n9884 = ~n9720 & ~n9883;
  assign n9885 = ~n9250 & n9716;
  assign n9886 = ~n6134 & ~n9885;
  assign n9887 = pi0075 & ~n9703;
  assign n9888 = pi0100 & ~n9703;
  assign n9889 = n9282 & ~n9694;
  assign n9890 = n9249 & ~n9889;
  assign n9891 = ~pi0100 & ~n9890;
  assign n9892 = ~pi0232 & n9282;
  assign n9893 = ~n9891 & ~n9892;
  assign n9894 = ~n9866 & ~n9893;
  assign n9895 = ~n9888 & ~n9894;
  assign n9896 = ~pi0075 & ~n9895;
  assign n9897 = ~pi0092 & ~n9887;
  assign n9898 = ~n9896 & n9897;
  assign n9899 = ~n9886 & ~n9898;
  assign n9900 = ~n9865 & ~n9899;
  assign n9901 = ~pi0074 & ~n9900;
  assign n9902 = n9864 & ~n9901;
  assign n9903 = pi0146 & n9646;
  assign n9904 = ~pi0146 & ~n9640;
  assign n9905 = ~pi0161 & ~n9903;
  assign n9906 = ~n9904 & n9905;
  assign n9907 = pi0146 & n9648;
  assign n9908 = ~pi0146 & ~n9638;
  assign n9909 = pi0161 & ~n9907;
  assign n9910 = ~n9908 & n9909;
  assign n9911 = ~n9906 & ~n9910;
  assign n9912 = pi0162 & ~n9911;
  assign n9913 = ~pi0161 & ~n9606;
  assign n9914 = pi0161 & ~n9574;
  assign n9915 = pi0146 & ~n9913;
  assign n9916 = ~n9914 & n9915;
  assign n9917 = ~pi0161 & ~n9615;
  assign n9918 = pi0161 & ~n9612;
  assign n9919 = ~pi0146 & ~n9917;
  assign n9920 = ~n9918 & n9919;
  assign n9921 = ~pi0162 & ~n9575;
  assign n9922 = ~n9916 & n9921;
  assign n9923 = ~n9920 & n9922;
  assign n9924 = ~n9912 & ~n9923;
  assign n9925 = n9793 & ~n9924;
  assign n9926 = pi0142 & n9391;
  assign n9927 = ~pi0142 & ~n9497;
  assign n9928 = ~pi0140 & ~n9926;
  assign n9929 = ~n9927 & n9928;
  assign n9930 = pi0142 & ~n9445;
  assign n9931 = ~n9511 & n9930;
  assign n9932 = ~pi0142 & ~n9507;
  assign n9933 = pi0140 & ~n9931;
  assign n9934 = ~n9932 & n9933;
  assign n9935 = ~n9929 & ~n9934;
  assign n9936 = ~pi0181 & ~n9935;
  assign n9937 = ~pi0142 & ~n9544;
  assign n9938 = pi0142 & ~n9458;
  assign n9939 = ~pi0140 & ~n9938;
  assign n9940 = ~n9937 & n9939;
  assign n9941 = pi0142 & ~n9453;
  assign n9942 = ~pi0142 & ~n9541;
  assign n9943 = pi0140 & ~n9941;
  assign n9944 = ~n9942 & n9943;
  assign n9945 = ~n9940 & ~n9944;
  assign n9946 = pi0181 & ~n9945;
  assign n9947 = pi0144 & ~n9946;
  assign n9948 = ~n9936 & n9947;
  assign n9949 = ~n9408 & n9604;
  assign n9950 = n6197 & ~n9949;
  assign n9951 = pi0142 & ~n9950;
  assign n9952 = ~n9511 & n9951;
  assign n9953 = ~pi0142 & n9529;
  assign n9954 = ~pi0140 & ~n9952;
  assign n9955 = ~n9953 & n9954;
  assign n9956 = pi0142 & ~n9645;
  assign n9957 = ~n9511 & n9956;
  assign n9958 = ~pi0142 & ~n9534;
  assign n9959 = pi0140 & ~n9957;
  assign n9960 = ~n9958 & n9959;
  assign n9961 = ~n9955 & ~n9960;
  assign n9962 = ~pi0181 & ~n9961;
  assign n9963 = pi0142 & ~n9414;
  assign n9964 = ~pi0142 & ~n9562;
  assign n9965 = ~pi0140 & ~n9963;
  assign n9966 = ~n9964 & n9965;
  assign n9967 = ~pi0142 & n9548;
  assign n9968 = pi0142 & ~n9430;
  assign n9969 = pi0140 & ~n9967;
  assign n9970 = ~n9968 & n9969;
  assign n9971 = ~n9966 & ~n9970;
  assign n9972 = pi0181 & ~n9971;
  assign n9973 = ~pi0144 & ~n9962;
  assign n9974 = ~n9972 & n9973;
  assign n9975 = ~pi0299 & ~n9974;
  assign n9976 = ~n9948 & n9975;
  assign n9977 = pi0146 & n9583;
  assign n9978 = ~pi0146 & ~n9597;
  assign n9979 = pi0161 & ~n9977;
  assign n9980 = ~n9978 & n9979;
  assign n9981 = pi0146 & ~n9578;
  assign n9982 = ~pi0146 & ~n9592;
  assign n9983 = ~pi0161 & ~n9981;
  assign n9984 = ~n9982 & n9983;
  assign n9985 = ~pi0162 & ~n9980;
  assign n9986 = ~n9984 & n9985;
  assign n9987 = ~pi0146 & n9632;
  assign n9988 = pi0146 & ~n9626;
  assign n9989 = ~pi0161 & ~n9987;
  assign n9990 = ~n9988 & n9989;
  assign n9991 = pi0146 & ~n9624;
  assign n9992 = ~pi0146 & ~n9630;
  assign n9993 = pi0161 & ~n9991;
  assign n9994 = ~n9992 & n9993;
  assign n9995 = pi0162 & ~n9990;
  assign n9996 = ~n9994 & n9995;
  assign n9997 = n9794 & ~n9986;
  assign n9998 = ~n9996 & n9997;
  assign n9999 = ~n9925 & ~n9998;
  assign n10000 = ~n9976 & n9999;
  assign n10001 = pi0232 & ~n10000;
  assign n10002 = ~n9661 & ~n10001;
  assign n10003 = n2530 & ~n10002;
  assign n10004 = pi0144 & n9307;
  assign n10005 = ~pi0144 & ~n9304;
  assign n10006 = ~n9338 & n10005;
  assign n10007 = n9772 & ~n10006;
  assign n10008 = ~n10004 & n10007;
  assign n10009 = ~n9304 & ~n9315;
  assign n10010 = n9776 & ~n10005;
  assign n10011 = ~n10009 & n10010;
  assign n10012 = ~n10008 & ~n10011;
  assign n10013 = pi0232 & ~n10012;
  assign n10014 = ~n9310 & ~n10013;
  assign n10015 = ~pi0038 & ~n10014;
  assign n10016 = ~pi0161 & n9327;
  assign n10017 = ~n9301 & ~n10016;
  assign n10018 = n9036 & ~n10017;
  assign n10019 = n9291 & n9766;
  assign n10020 = ~n10018 & n10019;
  assign n10021 = pi0161 & n9320;
  assign n10022 = n9036 & n9297;
  assign n10023 = ~n10021 & n10022;
  assign n10024 = n9291 & n9760;
  assign n10025 = ~n10023 & n10024;
  assign n10026 = ~n10020 & ~n10025;
  assign n10027 = pi0232 & ~n10026;
  assign n10028 = ~n10015 & ~n10027;
  assign n10029 = pi0039 & ~n10028;
  assign n10030 = ~pi0087 & ~n9759;
  assign n10031 = ~n10029 & n10030;
  assign n10032 = ~n10003 & n10031;
  assign n10033 = pi0038 & ~n9747;
  assign n10034 = ~n9266 & ~n10033;
  assign n10035 = pi0087 & n10034;
  assign n10036 = ~pi0100 & ~n10035;
  assign n10037 = ~n10032 & n10036;
  assign n10038 = ~n9733 & ~n10037;
  assign n10039 = n2569 & ~n10038;
  assign n10040 = ~pi0038 & n9848;
  assign n10041 = n7473 & ~n10040;
  assign n10042 = n9282 & ~n10041;
  assign n10043 = n10034 & ~n10042;
  assign n10044 = ~pi0100 & ~n10043;
  assign n10045 = ~n9733 & ~n10044;
  assign n10046 = n9205 & ~n10045;
  assign n10047 = ~n9734 & ~n10046;
  assign n10048 = ~n10039 & n10047;
  assign n10049 = ~pi0054 & ~n10048;
  assign n10050 = ~n9751 & ~n10049;
  assign n10051 = ~pi0074 & ~n10050;
  assign n10052 = n9743 & ~n10051;
  assign n10053 = n2529 & ~n9902;
  assign n10054 = ~n10052 & n10053;
  assign n10055 = ~n9884 & ~n10054;
  assign n10056 = ~n9713 & ~n10055;
  assign n10057 = ~pi0034 & n10056;
  assign n10058 = ~pi0033 & ~pi0954;
  assign n10059 = ~n9881 & ~n10058;
  assign n10060 = ~n10057 & n10059;
  assign n10061 = ~pi0034 & ~n8978;
  assign n10062 = n9880 & n10061;
  assign n10063 = n10056 & ~n10061;
  assign n10064 = n10058 & ~n10062;
  assign n10065 = ~n10063 & n10064;
  assign po0192 = ~n10060 & ~n10065;
  assign n10067 = n2529 & n2572;
  assign n10068 = n8962 & n10067;
  assign n10069 = ~pi0055 & n10068;
  assign n10070 = pi0059 & ~n10069;
  assign n10071 = ~pi0024 & n7340;
  assign n10072 = pi0054 & ~n10071;
  assign n10073 = pi0137 & n8884;
  assign n10074 = n2923 & n2930;
  assign n10075 = n7417 & ~n10074;
  assign n10076 = pi0683 & n10075;
  assign n10077 = pi0252 & po1057;
  assign n10078 = ~n10076 & n10077;
  assign n10079 = pi0146 & n7471;
  assign n10080 = pi0142 & n7470;
  assign n10081 = ~n10079 & ~n10080;
  assign n10082 = ~n7472 & n10081;
  assign n10083 = ~n10078 & ~n10082;
  assign n10084 = ~n7474 & ~n10083;
  assign n10085 = ~n8886 & ~n10084;
  assign n10086 = n6263 & ~n8889;
  assign n10087 = ~n10078 & n10086;
  assign n10088 = ~n10085 & ~n10087;
  assign n10089 = n8887 & ~n10088;
  assign n10090 = ~n10073 & ~n10089;
  assign n10091 = n8882 & ~n10090;
  assign n10092 = ~pi0090 & n6138;
  assign n10093 = ~pi0093 & ~n10092;
  assign n10094 = ~n6157 & ~n10093;
  assign n10095 = ~pi0035 & ~n10094;
  assign n10096 = pi0035 & ~n2915;
  assign n10097 = n8938 & ~n10096;
  assign n10098 = ~n10095 & n10097;
  assign n10099 = ~pi0032 & n10098;
  assign n10100 = pi0032 & ~pi0093;
  assign n10101 = n8895 & n10100;
  assign n10102 = n7432 & n10101;
  assign n10103 = ~n10099 & ~n10102;
  assign n10104 = ~pi0095 & ~n6169;
  assign n10105 = ~n10103 & n10104;
  assign n10106 = n6169 & ~n10095;
  assign n10107 = ~pi0137 & ~n6169;
  assign n10108 = n2924 & n7479;
  assign n10109 = ~n7425 & ~n10107;
  assign n10110 = n10108 & n10109;
  assign n10111 = ~pi0122 & ~po0740;
  assign n10112 = n7425 & ~n10107;
  assign n10113 = n10111 & n10112;
  assign n10114 = ~n10110 & ~n10113;
  assign n10115 = ~n10106 & n10114;
  assign n10116 = n2704 & n8932;
  assign n10117 = n10095 & ~n10116;
  assign n10118 = n2518 & n10097;
  assign n10119 = ~n10117 & n10118;
  assign n10120 = ~n10115 & n10119;
  assign n10121 = ~n2743 & ~n10098;
  assign n10122 = pi1082 & n2518;
  assign n10123 = ~n10121 & n10122;
  assign n10124 = ~pi0038 & ~n10120;
  assign n10125 = ~n10123 & n10124;
  assign n10126 = ~n10105 & n10125;
  assign n10127 = pi0038 & ~n8962;
  assign n10128 = ~pi0039 & ~pi0100;
  assign n10129 = ~n10127 & n10128;
  assign n10130 = ~n10126 & n10129;
  assign n10131 = ~n10091 & ~n10130;
  assign n10132 = n2533 & ~n10131;
  assign n10133 = pi0137 & ~po0840;
  assign n10134 = ~n6282 & n10133;
  assign n10135 = ~n8964 & ~n10134;
  assign n10136 = n8967 & ~n10135;
  assign n10137 = n8962 & n10136;
  assign n10138 = ~n10132 & ~n10137;
  assign n10139 = ~pi0092 & ~n10138;
  assign n10140 = ~pi0054 & ~n10139;
  assign n10141 = n2529 & n8879;
  assign n10142 = ~n10072 & n10141;
  assign n10143 = ~n10140 & n10142;
  assign n10144 = ~pi0059 & ~n10143;
  assign n10145 = ~pi0057 & ~n10070;
  assign po0193 = ~n10144 & n10145;
  assign n10147 = n2717 & n2771;
  assign n10148 = ~pi0065 & n2462;
  assign n10149 = n2487 & n10148;
  assign n10150 = n9081 & n10149;
  assign n10151 = ~pi0069 & n10150;
  assign n10152 = ~pi0067 & ~pi0071;
  assign n10153 = ~pi0083 & n2802;
  assign n10154 = pi0036 & ~pi0103;
  assign n10155 = n10152 & n10154;
  assign n10156 = n10151 & n10155;
  assign n10157 = n10153 & n10156;
  assign n10158 = n10147 & n10157;
  assign n10159 = ~pi0058 & n7522;
  assign n10160 = ~n10158 & ~n10159;
  assign n10161 = n2704 & n6479;
  assign n10162 = n6170 & n10161;
  assign n10163 = n2532 & ~po1038;
  assign n10164 = n3373 & n10163;
  assign n10165 = ~pi0092 & n10164;
  assign n10166 = n10162 & n10165;
  assign n10167 = po0740 & n10166;
  assign po0194 = ~n10160 & n10167;
  assign n10169 = ~pi0081 & ~n2789;
  assign n10170 = ~pi0045 & ~pi0073;
  assign n10171 = n8920 & n10170;
  assign n10172 = ~pi0071 & n2487;
  assign n10173 = ~pi0104 & n2472;
  assign n10174 = n10172 & n10173;
  assign n10175 = ~pi0048 & ~pi0065;
  assign n10176 = ~pi0082 & ~pi0084;
  assign n10177 = pi0089 & n10176;
  assign n10178 = n10175 & n10177;
  assign n10179 = n10171 & n10178;
  assign n10180 = n9080 & n10179;
  assign n10181 = n10174 & n10180;
  assign n10182 = pi0332 & n10181;
  assign n10183 = ~pi0064 & ~n10182;
  assign n10184 = n6479 & n9468;
  assign n10185 = n2501 & n10184;
  assign n10186 = n2508 & n10185;
  assign n10187 = ~pi0039 & ~pi0841;
  assign n10188 = n2465 & n10187;
  assign n10189 = ~n10183 & n10188;
  assign n10190 = n10186 & n10189;
  assign n10191 = n10169 & n10190;
  assign n10192 = ~pi0038 & ~n10191;
  assign n10193 = ~pi0039 & n2519;
  assign n10194 = pi0024 & n10193;
  assign n10195 = n2709 & n10194;
  assign n10196 = pi0038 & ~n10195;
  assign n10197 = n2571 & ~po1038;
  assign n10198 = ~n10192 & n10197;
  assign po0196 = ~n10196 & n10198;
  assign n10200 = ~pi0038 & n10197;
  assign n10201 = pi0786 & ~pi1082;
  assign n10202 = ~pi0984 & ~n2932;
  assign n10203 = pi0835 & ~n10202;
  assign n10204 = n6183 & ~n10203;
  assign n10205 = n6217 & ~n10204;
  assign n10206 = pi1093 & n10205;
  assign n10207 = n6184 & n6380;
  assign n10208 = ~n10206 & n10207;
  assign n10209 = ~pi0223 & n10208;
  assign n10210 = n6198 & n10205;
  assign n10211 = n10207 & ~n10210;
  assign n10212 = n6205 & n10211;
  assign n10213 = ~n6227 & n10205;
  assign n10214 = n10207 & ~n10213;
  assign n10215 = ~n6205 & n10214;
  assign n10216 = ~pi0299 & ~n10212;
  assign n10217 = ~n10215 & n10216;
  assign n10218 = ~n10209 & n10217;
  assign n10219 = ~pi0215 & n10208;
  assign n10220 = n6242 & n10211;
  assign n10221 = ~n6242 & n10214;
  assign n10222 = pi0299 & ~n10220;
  assign n10223 = ~n10221 & n10222;
  assign n10224 = ~n10219 & n10223;
  assign n10225 = ~n10201 & ~n10218;
  assign n10226 = ~n10224 & n10225;
  assign n10227 = n5853 & ~n6244;
  assign n10228 = n3470 & ~n6207;
  assign n10229 = ~n10227 & ~n10228;
  assign n10230 = po0740 & n10201;
  assign n10231 = ~n10229 & n10230;
  assign n10232 = n6382 & n10231;
  assign n10233 = ~n10226 & ~n10232;
  assign n10234 = pi0039 & ~n10233;
  assign n10235 = ~pi0039 & ~pi0095;
  assign n10236 = n6169 & n6486;
  assign n10237 = ~pi0986 & ~po0740;
  assign n10238 = pi0252 & ~n10237;
  assign n10239 = pi0314 & ~n10238;
  assign n10240 = pi0108 & n2714;
  assign n10241 = n2773 & n10240;
  assign n10242 = ~pi0841 & n2494;
  assign n10243 = n2720 & n10242;
  assign n10244 = n2714 & ~n2774;
  assign n10245 = n8921 & n9076;
  assign n10246 = ~pi0065 & ~pi0069;
  assign n10247 = n10245 & n10246;
  assign n10248 = pi0048 & ~pi0049;
  assign n10249 = ~pi0068 & ~pi0082;
  assign n10250 = n10248 & n10249;
  assign n10251 = n10170 & n10250;
  assign n10252 = n8910 & n8914;
  assign n10253 = n9078 & n10252;
  assign n10254 = n10247 & n10251;
  assign n10255 = n10253 & n10254;
  assign n10256 = n10174 & n10255;
  assign n10257 = ~pi0097 & n10243;
  assign n10258 = n10256 & n10257;
  assign n10259 = n10244 & n10258;
  assign n10260 = ~pi0047 & ~n10241;
  assign n10261 = ~n10259 & n10260;
  assign n10262 = n6151 & n10239;
  assign n10263 = ~n10261 & n10262;
  assign n10264 = ~pi0047 & ~pi0841;
  assign n10265 = n10256 & n10264;
  assign n10266 = ~n2760 & ~n10265;
  assign n10267 = n2500 & n2700;
  assign n10268 = ~n10239 & n10267;
  assign n10269 = ~n10266 & n10268;
  assign n10270 = ~n10263 & ~n10269;
  assign n10271 = n2704 & ~n10270;
  assign n10272 = ~pi0035 & ~n10271;
  assign n10273 = pi0035 & ~n6483;
  assign n10274 = n2508 & ~n10273;
  assign n10275 = n2510 & n10274;
  assign n10276 = ~n10272 & n10275;
  assign n10277 = ~n10236 & ~n10276;
  assign n10278 = n10235 & ~n10277;
  assign n10279 = ~n10234 & ~n10278;
  assign po0197 = n10200 & ~n10279;
  assign n10281 = ~pi0093 & pi0102;
  assign n10282 = n2461 & n10281;
  assign n10283 = n2464 & n10282;
  assign n10284 = n6170 & n10283;
  assign n10285 = n2501 & n10284;
  assign n10286 = n2490 & n10285;
  assign n10287 = n6479 & n10286;
  assign n10288 = pi1082 & ~n10287;
  assign n10289 = n2518 & ~n3411;
  assign n10290 = ~pi0040 & ~n10286;
  assign n10291 = n10289 & ~n10290;
  assign n10292 = ~pi1082 & ~n10291;
  assign n10293 = n10165 & ~n10288;
  assign po0198 = ~n10292 & n10293;
  assign n10295 = ~pi0189 & n6197;
  assign n10296 = pi0144 & n10295;
  assign n10297 = ~pi0174 & n10296;
  assign n10298 = ~pi0299 & ~n10297;
  assign n10299 = ~pi0166 & n6197;
  assign n10300 = pi0161 & n10299;
  assign n10301 = ~pi0152 & n10300;
  assign n10302 = ~n7470 & ~n10301;
  assign n10303 = pi0232 & ~n10298;
  assign n10304 = ~n10302 & n10303;
  assign n10305 = ~pi0072 & ~n10304;
  assign n10306 = pi0039 & ~n10305;
  assign n10307 = ~pi0041 & ~pi0072;
  assign n10308 = ~pi0039 & ~n10307;
  assign n10309 = ~n10306 & ~n10308;
  assign n10310 = ~n2620 & n10309;
  assign n10311 = ~n7506 & ~n10307;
  assign n10312 = ~n2924 & n10307;
  assign n10313 = n7506 & ~n10312;
  assign n10314 = ~pi0041 & pi0072;
  assign n10315 = n2924 & ~n10314;
  assign n10316 = ~pi0044 & n2521;
  assign n10317 = ~pi0101 & n10316;
  assign n10318 = n7479 & n10317;
  assign n10319 = n7477 & n10318;
  assign n10320 = pi0041 & ~n10319;
  assign n10321 = ~pi0099 & n6272;
  assign n10322 = ~pi0072 & pi0101;
  assign n10323 = ~pi0041 & ~n10322;
  assign n10324 = pi0252 & n6479;
  assign n10325 = ~pi0024 & n2709;
  assign n10326 = n7479 & n10324;
  assign n10327 = n10325 & n10326;
  assign n10328 = ~pi0044 & n10327;
  assign n10329 = n10323 & n10328;
  assign n10330 = ~n10321 & n10329;
  assign n10331 = n10315 & ~n10330;
  assign n10332 = ~n10320 & n10331;
  assign n10333 = n10313 & ~n10332;
  assign n10334 = ~n10311 & ~n10333;
  assign n10335 = ~pi0039 & ~n10334;
  assign n10336 = n2620 & ~n10306;
  assign n10337 = ~n10335 & n10336;
  assign n10338 = pi0075 & ~n10310;
  assign n10339 = ~n10337 & n10338;
  assign n10340 = ~n2608 & n10308;
  assign n10341 = ~pi0228 & n10307;
  assign n10342 = n2709 & n6479;
  assign n10343 = ~pi0044 & n10342;
  assign n10344 = n10323 & n10343;
  assign n10345 = ~n10314 & ~n10344;
  assign n10346 = pi0041 & ~n10317;
  assign n10347 = pi0228 & n10345;
  assign n10348 = ~n10346 & n10347;
  assign n10349 = n2625 & ~n10341;
  assign n10350 = ~n10348 & n10349;
  assign n10351 = pi0087 & ~n10340;
  assign n10352 = ~n10306 & n10351;
  assign n10353 = ~n10350 & n10352;
  assign n10354 = pi0038 & ~n10309;
  assign n10355 = pi0041 & ~n10318;
  assign n10356 = n2924 & ~n10321;
  assign n10357 = ~n10315 & ~n10356;
  assign n10358 = ~pi0072 & ~n7479;
  assign n10359 = ~n10345 & ~n10358;
  assign n10360 = ~n10321 & n10359;
  assign n10361 = ~n10355 & ~n10357;
  assign n10362 = ~n10360 & n10361;
  assign n10363 = n10313 & ~n10362;
  assign n10364 = ~n10311 & ~n10363;
  assign n10365 = ~pi0039 & ~n10364;
  assign n10366 = ~n10306 & ~n10365;
  assign n10367 = n6285 & ~n10366;
  assign n10368 = pi0287 & n2521;
  assign n10369 = n10304 & n10368;
  assign n10370 = ~n10305 & ~n10369;
  assign n10371 = pi0039 & ~n10370;
  assign n10372 = pi0901 & ~pi0959;
  assign n10373 = ~pi0480 & pi0949;
  assign n10374 = n2717 & n2780;
  assign n10375 = n2708 & n10374;
  assign n10376 = ~n10373 & n10375;
  assign n10377 = n2708 & n10373;
  assign n10378 = n2700 & ~n2759;
  assign n10379 = ~pi0109 & n6451;
  assign n10380 = n2780 & n10379;
  assign n10381 = ~pi0110 & ~n10380;
  assign n10382 = ~pi0047 & n10377;
  assign n10383 = n10378 & n10382;
  assign n10384 = ~n10381 & n10383;
  assign n10385 = n10372 & ~n10376;
  assign n10386 = ~n10384 & n10385;
  assign n10387 = n2701 & n2758;
  assign n10388 = pi0110 & n10387;
  assign n10389 = n10377 & n10388;
  assign n10390 = ~n10372 & ~n10389;
  assign n10391 = ~pi0250 & pi0252;
  assign n10392 = n6479 & n10391;
  assign n10393 = ~n10390 & n10392;
  assign n10394 = ~n10386 & n10393;
  assign n10395 = ~pi0072 & n10394;
  assign n10396 = n10162 & n10388;
  assign n10397 = n10373 & ~n10391;
  assign n10398 = n10396 & n10397;
  assign n10399 = ~n10395 & ~n10398;
  assign n10400 = ~pi0044 & ~n10399;
  assign n10401 = ~pi0101 & n10400;
  assign n10402 = pi0041 & ~n10401;
  assign n10403 = pi0044 & pi0072;
  assign n10404 = n6479 & ~n10391;
  assign n10405 = n10389 & n10404;
  assign n10406 = ~pi0072 & ~n10405;
  assign n10407 = ~n10394 & n10406;
  assign n10408 = ~pi0044 & ~n10407;
  assign n10409 = ~n10403 & ~n10408;
  assign n10410 = ~pi0101 & n10409;
  assign n10411 = n10323 & ~n10410;
  assign n10412 = ~n10402 & ~n10411;
  assign n10413 = ~pi0228 & ~n10412;
  assign n10414 = ~pi0072 & ~n7451;
  assign n10415 = ~n7457 & n10414;
  assign n10416 = n6479 & ~n7455;
  assign n10417 = ~n7454 & n10416;
  assign n10418 = ~pi0072 & n7457;
  assign n10419 = ~n10417 & n10418;
  assign n10420 = ~pi1093 & ~n10415;
  assign n10421 = ~n10419 & n10420;
  assign n10422 = n10414 & ~n10421;
  assign n10423 = ~pi0044 & ~n10422;
  assign n10424 = ~n10403 & ~n10423;
  assign n10425 = ~pi0101 & n10424;
  assign n10426 = n10323 & ~n10425;
  assign n10427 = n7451 & ~n7457;
  assign n10428 = ~pi1093 & ~n7459;
  assign n10429 = ~n10427 & n10428;
  assign n10430 = ~pi0044 & ~n10429;
  assign n10431 = pi1093 & ~n7451;
  assign n10432 = n10430 & ~n10431;
  assign n10433 = ~pi0101 & n10432;
  assign n10434 = pi0041 & ~n10433;
  assign n10435 = ~n2924 & ~n10434;
  assign n10436 = ~n10426 & n10435;
  assign n10437 = n2935 & ~n7443;
  assign n10438 = n2937 & n10437;
  assign n10439 = ~n7522 & ~n10438;
  assign n10440 = n2461 & ~n10439;
  assign n10441 = n7434 & ~n10440;
  assign n10442 = n7431 & ~n10441;
  assign n10443 = ~pi0051 & ~n10442;
  assign n10444 = ~n2747 & ~n10443;
  assign n10445 = ~pi0096 & ~n10444;
  assign n10446 = n10416 & n10418;
  assign n10447 = ~n10445 & n10446;
  assign n10448 = ~n10427 & ~n10447;
  assign n10449 = pi1093 & n10448;
  assign n10450 = n10430 & ~n10449;
  assign n10451 = ~pi0101 & n10450;
  assign n10452 = pi0041 & ~n10451;
  assign n10453 = ~pi0072 & n10448;
  assign n10454 = pi1093 & ~n10453;
  assign n10455 = ~n10421 & ~n10454;
  assign n10456 = ~pi0044 & ~n10455;
  assign n10457 = ~n10403 & ~n10456;
  assign n10458 = ~pi0101 & n10457;
  assign n10459 = n10323 & ~n10458;
  assign n10460 = n2924 & ~n10459;
  assign n10461 = ~n10452 & n10460;
  assign n10462 = pi0228 & ~n10436;
  assign n10463 = ~n10461 & n10462;
  assign n10464 = ~pi0039 & ~n10413;
  assign n10465 = ~n10463 & n10464;
  assign n10466 = n2608 & ~n10371;
  assign n10467 = ~n10465 & n10466;
  assign n10468 = ~pi0087 & ~n10354;
  assign n10469 = ~n10367 & n10468;
  assign n10470 = ~n10467 & n10469;
  assign n10471 = ~pi0075 & ~n10353;
  assign n10472 = ~n10470 & n10471;
  assign n10473 = ~n10339 & ~n10472;
  assign n10474 = n7429 & ~n10473;
  assign n10475 = ~n7429 & ~n10309;
  assign n10476 = ~po1038 & ~n10475;
  assign n10477 = ~n10474 & n10476;
  assign n10478 = pi0039 & pi0232;
  assign n10479 = n10301 & n10478;
  assign n10480 = ~pi0072 & ~n10308;
  assign n10481 = po1038 & n10480;
  assign n10482 = ~n10479 & n10481;
  assign po0199 = ~n10477 & ~n10482;
  assign n10484 = pi0211 & pi0214;
  assign n10485 = pi0212 & n10484;
  assign n10486 = ~pi0219 & ~n10485;
  assign n10487 = pi0207 & pi0208;
  assign n10488 = pi0042 & ~pi0072;
  assign n10489 = ~n2620 & n10488;
  assign n10490 = ~n7506 & ~n10488;
  assign n10491 = ~pi0115 & n2924;
  assign n10492 = n10488 & ~n10491;
  assign n10493 = n7506 & ~n10492;
  assign n10494 = pi0114 & ~n10488;
  assign n10495 = n10491 & ~n10494;
  assign n10496 = n6266 & n10328;
  assign n10497 = ~pi0113 & n10496;
  assign n10498 = ~pi0116 & n10497;
  assign n10499 = n10488 & ~n10498;
  assign n10500 = n6265 & n10317;
  assign n10501 = n6269 & n10500;
  assign n10502 = n7479 & n10501;
  assign n10503 = ~pi0114 & ~n6268;
  assign n10504 = n10502 & n10503;
  assign n10505 = n7477 & n10504;
  assign n10506 = ~pi0042 & n10505;
  assign n10507 = ~pi0114 & ~n10499;
  assign n10508 = ~n10506 & n10507;
  assign n10509 = n10495 & ~n10508;
  assign n10510 = n10493 & ~n10509;
  assign n10511 = n2620 & ~n10490;
  assign n10512 = ~n10510 & n10511;
  assign n10513 = ~pi0039 & ~n10489;
  assign n10514 = ~n10512 & n10513;
  assign n10515 = ~pi0072 & pi0199;
  assign n10516 = ~pi0232 & ~n10515;
  assign n10517 = ~pi0299 & ~n10516;
  assign n10518 = ~pi0072 & ~n10295;
  assign n10519 = pi0199 & n10518;
  assign n10520 = pi0232 & ~n10519;
  assign n10521 = n10517 & ~n10520;
  assign n10522 = ~pi0166 & n7473;
  assign n10523 = ~pi0072 & ~n10522;
  assign n10524 = pi0299 & n10523;
  assign n10525 = pi0039 & ~n10524;
  assign n10526 = ~n10521 & n10525;
  assign n10527 = ~n10514 & ~n10526;
  assign n10528 = pi0075 & ~n10527;
  assign n10529 = ~pi0039 & ~n10488;
  assign n10530 = ~n2608 & n10529;
  assign n10531 = n6266 & n10343;
  assign n10532 = pi0228 & n10531;
  assign n10533 = n6271 & n10532;
  assign n10534 = n10488 & ~n10533;
  assign n10535 = pi0228 & n10501;
  assign n10536 = ~pi0115 & n10535;
  assign n10537 = ~pi0114 & n10536;
  assign n10538 = ~pi0042 & n10537;
  assign n10539 = n2625 & ~n10534;
  assign n10540 = ~n10538 & n10539;
  assign n10541 = pi0087 & ~n10530;
  assign n10542 = ~n10540 & n10541;
  assign n10543 = ~n10526 & n10542;
  assign n10544 = pi0115 & ~n10488;
  assign n10545 = pi0042 & ~pi0114;
  assign n10546 = pi0072 & pi0116;
  assign n10547 = pi0072 & pi0113;
  assign n10548 = pi0072 & ~n6265;
  assign n10549 = ~pi0099 & n10411;
  assign n10550 = ~n10548 & ~n10549;
  assign n10551 = ~pi0113 & ~n10550;
  assign n10552 = ~n10547 & ~n10551;
  assign n10553 = ~pi0116 & ~n10552;
  assign n10554 = ~n10546 & ~n10553;
  assign n10555 = n10545 & ~n10554;
  assign n10556 = n6265 & n10401;
  assign n10557 = ~pi0113 & n10556;
  assign n10558 = ~pi0116 & n10557;
  assign n10559 = ~pi0042 & ~n10558;
  assign n10560 = ~n10494 & ~n10559;
  assign n10561 = ~n10555 & n10560;
  assign n10562 = ~pi0115 & ~n10561;
  assign n10563 = ~pi0228 & ~n10544;
  assign n10564 = ~n10562 & n10563;
  assign n10565 = ~pi0099 & n10459;
  assign n10566 = ~n10548 & ~n10565;
  assign n10567 = ~pi0113 & ~n10566;
  assign n10568 = ~n10547 & ~n10567;
  assign n10569 = ~pi0116 & ~n10568;
  assign n10570 = ~n10546 & ~n10569;
  assign n10571 = n10545 & ~n10570;
  assign n10572 = n6265 & n10451;
  assign n10573 = n6269 & n10572;
  assign n10574 = ~pi0042 & ~n10573;
  assign n10575 = ~n10494 & ~n10574;
  assign n10576 = ~n10571 & n10575;
  assign n10577 = n10491 & ~n10576;
  assign n10578 = ~pi0115 & ~n2924;
  assign n10579 = n6265 & n10433;
  assign n10580 = n6269 & n10579;
  assign n10581 = ~pi0042 & n10580;
  assign n10582 = ~pi0099 & n10426;
  assign n10583 = ~n10548 & ~n10582;
  assign n10584 = ~pi0113 & ~n10583;
  assign n10585 = ~n10547 & ~n10584;
  assign n10586 = ~pi0116 & ~n10585;
  assign n10587 = ~n10546 & ~n10586;
  assign n10588 = pi0042 & n10587;
  assign n10589 = ~pi0114 & ~n10581;
  assign n10590 = ~n10588 & n10589;
  assign n10591 = ~n10494 & ~n10590;
  assign n10592 = n10578 & ~n10591;
  assign n10593 = pi0228 & ~n10544;
  assign n10594 = ~n10592 & n10593;
  assign n10595 = ~n10577 & n10594;
  assign n10596 = ~pi0039 & ~n10564;
  assign n10597 = ~n10595 & n10596;
  assign n10598 = pi0232 & pi0299;
  assign n10599 = n10299 & n10368;
  assign n10600 = ~n10523 & n10598;
  assign n10601 = ~n10599 & n10600;
  assign n10602 = pi0232 & ~pi0299;
  assign n10603 = n6197 & n10368;
  assign n10604 = ~pi0189 & n10603;
  assign n10605 = ~n10518 & ~n10604;
  assign n10606 = pi0199 & ~n10605;
  assign n10607 = n10602 & ~n10606;
  assign n10608 = pi0072 & ~pi0232;
  assign n10609 = pi0299 & ~n10608;
  assign n10610 = n10516 & ~n10609;
  assign n10611 = ~n10601 & ~n10610;
  assign n10612 = ~n10607 & n10611;
  assign n10613 = pi0039 & ~n10612;
  assign n10614 = ~n10597 & ~n10613;
  assign n10615 = n2608 & ~n10614;
  assign n10616 = n6269 & n10531;
  assign n10617 = ~pi0072 & ~n10616;
  assign n10618 = ~n10358 & ~n10617;
  assign n10619 = pi0042 & ~n10618;
  assign n10620 = ~pi0042 & n10504;
  assign n10621 = ~pi0114 & ~n10619;
  assign n10622 = ~n10620 & n10621;
  assign n10623 = n10495 & ~n10622;
  assign n10624 = n10493 & ~n10623;
  assign n10625 = ~n10490 & ~n10624;
  assign n10626 = ~pi0039 & ~n10625;
  assign n10627 = ~n10526 & ~n10626;
  assign n10628 = n6285 & ~n10627;
  assign n10629 = ~n10526 & ~n10529;
  assign n10630 = pi0038 & ~n10629;
  assign n10631 = ~pi0087 & ~n10630;
  assign n10632 = ~n10628 & n10631;
  assign n10633 = ~n10615 & n10632;
  assign n10634 = ~pi0075 & ~n10543;
  assign n10635 = ~n10633 & n10634;
  assign n10636 = n7429 & ~n10528;
  assign n10637 = ~n10635 & n10636;
  assign n10638 = ~n10487 & ~n10637;
  assign n10639 = ~pi0072 & pi0200;
  assign n10640 = ~pi0232 & ~n10639;
  assign n10641 = ~pi0299 & ~n10640;
  assign n10642 = pi0200 & n10518;
  assign n10643 = pi0232 & ~n10642;
  assign n10644 = n10641 & ~n10643;
  assign n10645 = pi0039 & ~n10644;
  assign n10646 = ~n10521 & n10645;
  assign n10647 = ~n10529 & ~n10646;
  assign n10648 = ~n7429 & n10647;
  assign n10649 = n10487 & ~n10648;
  assign n10650 = n10526 & n10645;
  assign n10651 = ~n10514 & ~n10650;
  assign n10652 = pi0075 & ~n10651;
  assign n10653 = ~n10626 & ~n10650;
  assign n10654 = n6285 & ~n10653;
  assign n10655 = pi0038 & ~n10647;
  assign n10656 = ~pi0087 & ~n10655;
  assign n10657 = ~n10631 & ~n10656;
  assign n10658 = pi0232 & ~n10606;
  assign n10659 = pi0200 & ~n10605;
  assign n10660 = n10658 & ~n10659;
  assign n10661 = ~pi0299 & n10660;
  assign n10662 = n10610 & ~n10639;
  assign n10663 = ~n10601 & ~n10662;
  assign n10664 = ~n10661 & n10663;
  assign n10665 = pi0039 & ~n10664;
  assign n10666 = ~n10597 & ~n10665;
  assign n10667 = n2608 & ~n10666;
  assign n10668 = ~n10654 & ~n10657;
  assign n10669 = ~n10667 & n10668;
  assign n10670 = n10541 & ~n10650;
  assign n10671 = ~n10540 & n10670;
  assign n10672 = ~pi0075 & ~n10671;
  assign n10673 = ~n10669 & n10672;
  assign n10674 = n7429 & ~n10652;
  assign n10675 = ~n10673 & n10674;
  assign n10676 = n10649 & ~n10675;
  assign n10677 = ~n10638 & ~n10676;
  assign n10678 = ~n7429 & n10629;
  assign n10679 = ~n10486 & ~n10678;
  assign n10680 = ~n10677 & n10679;
  assign n10681 = pi0039 & ~n10521;
  assign n10682 = ~n10514 & ~n10681;
  assign n10683 = pi0075 & ~n10682;
  assign n10684 = n10542 & ~n10681;
  assign n10685 = ~n10626 & ~n10681;
  assign n10686 = n6285 & ~n10685;
  assign n10687 = ~n10529 & ~n10681;
  assign n10688 = pi0038 & ~n10687;
  assign n10689 = n10517 & ~n10658;
  assign n10690 = pi0039 & ~n10689;
  assign n10691 = ~n10597 & ~n10690;
  assign n10692 = n2608 & ~n10691;
  assign n10693 = ~pi0087 & ~n10688;
  assign n10694 = ~n10686 & n10693;
  assign n10695 = ~n10692 & n10694;
  assign n10696 = ~pi0075 & ~n10684;
  assign n10697 = ~n10695 & n10696;
  assign n10698 = n7429 & ~n10683;
  assign n10699 = ~n10697 & n10698;
  assign n10700 = ~n7429 & n10687;
  assign n10701 = ~n10487 & ~n10700;
  assign n10702 = ~n10699 & n10701;
  assign n10703 = ~n10514 & ~n10646;
  assign n10704 = pi0075 & ~n10703;
  assign n10705 = n10542 & ~n10646;
  assign n10706 = ~n10517 & ~n10641;
  assign n10707 = ~n10660 & ~n10706;
  assign n10708 = pi0039 & ~n10707;
  assign n10709 = ~n10597 & ~n10708;
  assign n10710 = n2608 & ~n10709;
  assign n10711 = ~n10626 & ~n10646;
  assign n10712 = n6285 & ~n10711;
  assign n10713 = n10656 & ~n10712;
  assign n10714 = ~n10710 & n10713;
  assign n10715 = ~pi0075 & ~n10705;
  assign n10716 = ~n10714 & n10715;
  assign n10717 = n7429 & ~n10704;
  assign n10718 = ~n10716 & n10717;
  assign n10719 = n10649 & ~n10718;
  assign n10720 = ~n10702 & ~n10719;
  assign n10721 = n10486 & ~n10720;
  assign n10722 = ~po1038 & ~n10680;
  assign n10723 = ~n10721 & n10722;
  assign n10724 = ~n10486 & n10523;
  assign n10725 = pi0039 & ~n10724;
  assign n10726 = po1038 & ~n10529;
  assign n10727 = ~n10725 & n10726;
  assign po0200 = n10723 | n10727;
  assign n10729 = pi0043 & ~pi0072;
  assign n10730 = ~n7506 & ~n10729;
  assign n10731 = ~pi0042 & n6270;
  assign n10732 = n2924 & n10731;
  assign n10733 = n10729 & ~n10732;
  assign n10734 = n7506 & ~n10733;
  assign n10735 = ~pi0072 & ~n10498;
  assign n10736 = pi0043 & n10735;
  assign n10737 = ~pi0043 & pi0052;
  assign n10738 = n7477 & n10502;
  assign n10739 = n10737 & n10738;
  assign n10740 = ~n10736 & ~n10739;
  assign n10741 = n10732 & ~n10740;
  assign n10742 = n10734 & ~n10741;
  assign n10743 = ~n10730 & ~n10742;
  assign n10744 = ~pi0039 & ~n10743;
  assign n10745 = n2620 & ~n10744;
  assign n10746 = ~pi0039 & ~n10729;
  assign n10747 = ~n2620 & ~n10746;
  assign n10748 = ~n10745 & ~n10747;
  assign n10749 = ~n10645 & ~n10748;
  assign n10750 = pi0075 & ~n10749;
  assign n10751 = ~n2608 & n10746;
  assign n10752 = ~pi0043 & ~n10501;
  assign n10753 = pi0043 & ~n10617;
  assign n10754 = pi0228 & n10731;
  assign n10755 = ~n10753 & n10754;
  assign n10756 = ~n10752 & n10755;
  assign n10757 = n10729 & ~n10754;
  assign n10758 = n2625 & ~n10757;
  assign n10759 = ~n10756 & n10758;
  assign n10760 = pi0087 & ~n10751;
  assign n10761 = ~n10759 & n10760;
  assign n10762 = ~n10645 & n10761;
  assign n10763 = n10502 & n10737;
  assign n10764 = pi0043 & ~n10618;
  assign n10765 = ~n10763 & ~n10764;
  assign n10766 = n10732 & ~n10765;
  assign n10767 = n10734 & ~n10766;
  assign n10768 = ~n10730 & ~n10767;
  assign n10769 = ~pi0039 & ~n10768;
  assign n10770 = ~n10645 & ~n10769;
  assign n10771 = n6285 & ~n10770;
  assign n10772 = ~n10645 & ~n10746;
  assign n10773 = pi0038 & ~n10772;
  assign n10774 = pi0232 & ~n10659;
  assign n10775 = n10641 & ~n10774;
  assign n10776 = pi0039 & ~n10775;
  assign n10777 = ~pi0228 & ~n10558;
  assign n10778 = ~n2924 & ~n10579;
  assign n10779 = n2924 & ~n10572;
  assign n10780 = ~n10778 & ~n10779;
  assign n10781 = n6269 & n10780;
  assign n10782 = pi0228 & ~n10781;
  assign n10783 = ~n10777 & ~n10782;
  assign n10784 = ~pi0043 & ~n10783;
  assign n10785 = ~n10729 & ~n10731;
  assign n10786 = ~n2924 & ~n10587;
  assign n10787 = n2924 & ~n10570;
  assign n10788 = ~n10786 & ~n10787;
  assign n10789 = pi0228 & ~n10788;
  assign n10790 = ~pi0228 & ~n10554;
  assign n10791 = ~n10789 & ~n10790;
  assign n10792 = pi0043 & n10731;
  assign n10793 = ~n10791 & n10792;
  assign n10794 = ~n10784 & ~n10785;
  assign n10795 = ~n10793 & n10794;
  assign n10796 = ~pi0039 & ~n10795;
  assign n10797 = ~n10776 & ~n10796;
  assign n10798 = n2608 & ~n10797;
  assign n10799 = ~pi0087 & ~n10773;
  assign n10800 = ~n10771 & n10799;
  assign n10801 = ~n10798 & n10800;
  assign n10802 = ~pi0075 & ~n10762;
  assign n10803 = ~n10801 & n10802;
  assign n10804 = n7429 & ~n10750;
  assign n10805 = ~n10803 & n10804;
  assign n10806 = ~n7429 & n10772;
  assign n10807 = ~n10487 & ~n10806;
  assign n10808 = ~n10805 & n10807;
  assign n10809 = ~pi0199 & ~pi0200;
  assign n10810 = ~pi0299 & ~n10809;
  assign n10811 = ~pi0072 & ~n10810;
  assign n10812 = ~pi0232 & ~n10811;
  assign n10813 = ~pi0299 & ~n10812;
  assign n10814 = n10518 & n10809;
  assign n10815 = pi0232 & ~n10814;
  assign n10816 = n10813 & ~n10815;
  assign n10817 = pi0039 & ~n10816;
  assign n10818 = ~n10746 & ~n10817;
  assign n10819 = ~n7429 & n10818;
  assign n10820 = ~n10748 & ~n10817;
  assign n10821 = pi0075 & ~n10820;
  assign n10822 = ~n10769 & ~n10817;
  assign n10823 = n6285 & ~n10822;
  assign n10824 = pi0038 & ~n10818;
  assign n10825 = ~n10605 & n10809;
  assign n10826 = pi0232 & ~n10825;
  assign n10827 = n10813 & ~n10826;
  assign n10828 = pi0039 & ~n10827;
  assign n10829 = ~n10796 & ~n10828;
  assign n10830 = n2608 & ~n10829;
  assign n10831 = ~pi0087 & ~n10824;
  assign n10832 = ~n10823 & n10831;
  assign n10833 = ~n10830 & n10832;
  assign n10834 = ~n2531 & ~n10818;
  assign n10835 = n10761 & ~n10834;
  assign n10836 = ~pi0075 & ~n10835;
  assign n10837 = ~n10833 & n10836;
  assign n10838 = n7429 & ~n10821;
  assign n10839 = ~n10837 & n10838;
  assign n10840 = n10487 & ~n10819;
  assign n10841 = ~n10839 & n10840;
  assign n10842 = ~n10808 & ~n10841;
  assign n10843 = pi0212 & pi0214;
  assign n10844 = ~pi0211 & ~pi0219;
  assign n10845 = n10843 & ~n10844;
  assign n10846 = ~pi0211 & ~n10843;
  assign n10847 = ~n10845 & ~n10846;
  assign n10848 = ~n10842 & ~n10847;
  assign n10849 = n10525 & ~n10644;
  assign n10850 = ~n10748 & ~n10849;
  assign n10851 = pi0075 & ~n10850;
  assign n10852 = n10761 & ~n10849;
  assign n10853 = ~n10769 & ~n10849;
  assign n10854 = n6285 & ~n10853;
  assign n10855 = ~n10746 & ~n10849;
  assign n10856 = pi0038 & ~n10855;
  assign n10857 = n10602 & ~n10659;
  assign n10858 = ~n10609 & n10640;
  assign n10859 = ~n10601 & ~n10858;
  assign n10860 = ~n10857 & n10859;
  assign n10861 = pi0039 & ~n10860;
  assign n10862 = ~n10796 & ~n10861;
  assign n10863 = n2608 & ~n10862;
  assign n10864 = ~pi0087 & ~n10856;
  assign n10865 = ~n10854 & n10864;
  assign n10866 = ~n10863 & n10865;
  assign n10867 = ~pi0075 & ~n10852;
  assign n10868 = ~n10866 & n10867;
  assign n10869 = n7429 & ~n10851;
  assign n10870 = ~n10868 & n10869;
  assign n10871 = ~n7429 & n10855;
  assign n10872 = ~n10487 & ~n10871;
  assign n10873 = ~n10870 & n10872;
  assign n10874 = ~n10524 & n10817;
  assign n10875 = ~n10746 & ~n10874;
  assign n10876 = ~n7429 & n10875;
  assign n10877 = ~n10748 & ~n10874;
  assign n10878 = pi0075 & ~n10877;
  assign n10879 = n10761 & ~n10874;
  assign n10880 = ~n10769 & ~n10874;
  assign n10881 = n6285 & ~n10880;
  assign n10882 = pi0038 & ~n10875;
  assign n10883 = n10602 & ~n10825;
  assign n10884 = ~n10601 & ~n10812;
  assign n10885 = ~n10883 & n10884;
  assign n10886 = pi0039 & ~n10885;
  assign n10887 = ~n10796 & ~n10886;
  assign n10888 = n2608 & ~n10887;
  assign n10889 = ~pi0087 & ~n10882;
  assign n10890 = ~n10881 & n10889;
  assign n10891 = ~n10888 & n10890;
  assign n10892 = ~pi0075 & ~n10879;
  assign n10893 = ~n10891 & n10892;
  assign n10894 = n7429 & ~n10878;
  assign n10895 = ~n10893 & n10894;
  assign n10896 = n10487 & ~n10876;
  assign n10897 = ~n10895 & n10896;
  assign n10898 = ~n10873 & ~n10897;
  assign n10899 = n10847 & ~n10898;
  assign n10900 = ~po1038 & ~n10848;
  assign n10901 = ~n10899 & n10900;
  assign n10902 = n10523 & n10847;
  assign n10903 = pi0039 & ~n10902;
  assign n10904 = po1038 & ~n10746;
  assign n10905 = ~n10903 & n10904;
  assign po0201 = n10901 | n10905;
  assign n10907 = ~pi0072 & n7474;
  assign n10908 = pi0039 & ~n10907;
  assign n10909 = pi0044 & ~pi0072;
  assign n10910 = ~pi0039 & ~n10909;
  assign n10911 = ~n10908 & ~n10910;
  assign n10912 = ~n2620 & n10911;
  assign n10913 = ~n7506 & ~n10909;
  assign n10914 = ~pi0039 & ~n10913;
  assign n10915 = ~n2924 & n10909;
  assign n10916 = n7506 & ~n10915;
  assign n10917 = n7594 & ~n10403;
  assign n10918 = n7479 & n10316;
  assign n10919 = n7477 & n10918;
  assign n10920 = pi0044 & ~n10327;
  assign n10921 = ~n10919 & ~n10920;
  assign n10922 = n10917 & ~n10921;
  assign n10923 = n10916 & ~n10922;
  assign n10924 = n10914 & ~n10923;
  assign n10925 = pi0039 & n7474;
  assign n10926 = ~pi0072 & n10925;
  assign n10927 = ~n10924 & ~n10926;
  assign n10928 = n2620 & ~n10927;
  assign n10929 = pi0075 & ~n10912;
  assign n10930 = ~n10928 & n10929;
  assign n10931 = pi0228 & n2608;
  assign n10932 = n10316 & n10931;
  assign n10933 = n10342 & n10931;
  assign n10934 = n10909 & ~n10933;
  assign n10935 = ~pi0039 & ~n10934;
  assign n10936 = ~n10932 & n10935;
  assign n10937 = pi0087 & ~n10908;
  assign n10938 = ~n10936 & n10937;
  assign n10939 = pi0038 & ~n10911;
  assign n10940 = n7479 & n10342;
  assign n10941 = pi0044 & ~n10940;
  assign n10942 = ~n10918 & ~n10941;
  assign n10943 = n10917 & ~n10942;
  assign n10944 = n10916 & ~n10943;
  assign n10945 = n10914 & ~n10944;
  assign n10946 = n6285 & ~n10926;
  assign n10947 = ~n10945 & n10946;
  assign n10948 = pi0287 & n10342;
  assign n10949 = ~pi0072 & ~n10948;
  assign n10950 = n10925 & n10949;
  assign n10951 = pi0044 & n10407;
  assign n10952 = ~pi0228 & ~n10951;
  assign n10953 = ~n10400 & n10952;
  assign n10954 = pi0044 & n10455;
  assign n10955 = n2924 & ~n10450;
  assign n10956 = ~n10954 & n10955;
  assign n10957 = pi0044 & n10422;
  assign n10958 = ~n2924 & ~n10432;
  assign n10959 = ~n10957 & n10958;
  assign n10960 = ~n10956 & ~n10959;
  assign n10961 = pi0228 & ~n10960;
  assign n10962 = ~pi0039 & ~n10953;
  assign n10963 = ~n10961 & n10962;
  assign n10964 = n2608 & ~n10950;
  assign n10965 = ~n10963 & n10964;
  assign n10966 = ~pi0087 & ~n10939;
  assign n10967 = ~n10947 & n10966;
  assign n10968 = ~n10965 & n10967;
  assign n10969 = ~pi0075 & ~n10938;
  assign n10970 = ~n10968 & n10969;
  assign n10971 = ~n10930 & ~n10970;
  assign n10972 = n7429 & ~n10971;
  assign n10973 = ~n7429 & ~n10911;
  assign n10974 = ~po1038 & ~n10973;
  assign n10975 = ~n10972 & n10974;
  assign n10976 = n2639 & n7473;
  assign n10977 = ~pi0072 & n10976;
  assign n10978 = pi0039 & ~n10977;
  assign n10979 = po1038 & ~n10910;
  assign n10980 = ~n10978 & n10979;
  assign po0202 = n10975 | n10980;
  assign n10982 = ~pi0038 & pi0039;
  assign n10983 = n10197 & n10982;
  assign n10984 = pi0979 & n10983;
  assign po0203 = n6380 & n10984;
  assign n10986 = ~pi0102 & ~pi0104;
  assign n10987 = ~pi0111 & n10986;
  assign n10988 = ~pi0049 & ~pi0076;
  assign n10989 = n8909 & n10988;
  assign n10990 = pi0061 & ~pi0082;
  assign n10991 = ~pi0083 & ~pi0089;
  assign n10992 = n10990 & n10991;
  assign n10993 = n7438 & n8915;
  assign n10994 = n10992 & n10993;
  assign n10995 = n10172 & n10987;
  assign n10996 = n10989 & n10995;
  assign n10997 = n8912 & n10994;
  assign n10998 = n10247 & n10997;
  assign n10999 = n10996 & n10998;
  assign n11000 = n8935 & n10999;
  assign n11001 = ~pi0841 & n11000;
  assign n11002 = n2702 & n2888;
  assign n11003 = pi0024 & n11002;
  assign n11004 = ~n11001 & ~n11003;
  assign po0204 = n10166 & ~n11004;
  assign n11006 = ~pi0082 & n2474;
  assign n11007 = ~pi0084 & pi0104;
  assign n11008 = n2805 & n11007;
  assign n11009 = n10171 & n11008;
  assign n11010 = n11006 & n11009;
  assign n11011 = ~pi0036 & ~n11010;
  assign n11012 = n8916 & n9081;
  assign n11013 = ~pi0067 & ~pi0103;
  assign n11014 = n2487 & n11013;
  assign n11015 = ~pi0098 & n11014;
  assign n11016 = n11012 & n11015;
  assign n11017 = ~n11011 & n11016;
  assign n11018 = ~n2803 & n11017;
  assign n11019 = ~pi0088 & ~n11018;
  assign n11020 = ~n2871 & n7438;
  assign n11021 = n2754 & ~n11019;
  assign n11022 = n11020 & n11021;
  assign n11023 = n2700 & n11022;
  assign n11024 = ~n10159 & ~n11023;
  assign n11025 = n10162 & ~n11024;
  assign n11026 = n7490 & ~n11025;
  assign n11027 = ~pi0036 & n11017;
  assign n11028 = ~pi0088 & ~n11027;
  assign n11029 = n11020 & ~n11028;
  assign n11030 = n10186 & n11029;
  assign n11031 = ~pi0824 & n2932;
  assign n11032 = n11030 & n11031;
  assign n11033 = ~n2932 & n11025;
  assign n11034 = pi0829 & ~n11032;
  assign n11035 = ~n11033 & n11034;
  assign n11036 = ~n2923 & n11035;
  assign n11037 = ~n11026 & ~n11036;
  assign n11038 = pi1091 & ~n11037;
  assign n11039 = ~n7417 & n11025;
  assign n11040 = ~pi0829 & ~n11039;
  assign n11041 = ~n11035 & ~n11040;
  assign n11042 = ~pi1093 & ~n11041;
  assign n11043 = n7417 & n10162;
  assign n11044 = ~n10160 & n11043;
  assign n11045 = ~n6394 & ~n7626;
  assign n11046 = ~n11044 & ~n11045;
  assign n11047 = ~n11039 & n11046;
  assign n11048 = n10165 & ~n11047;
  assign n11049 = ~n11042 & n11048;
  assign po0205 = ~n11038 & n11049;
  assign n11051 = ~pi0072 & pi0841;
  assign n11052 = n2705 & n11051;
  assign n11053 = ~pi0051 & n11052;
  assign n11054 = n10256 & n11053;
  assign n11055 = n10165 & n11054;
  assign po0206 = n10185 & n11055;
  assign n11057 = n2464 & n2487;
  assign n11058 = ~pi0103 & n2804;
  assign n11059 = n10245 & n11058;
  assign n11060 = n8909 & n8916;
  assign n11061 = n11059 & n11060;
  assign n11062 = ~pi0045 & pi0049;
  assign n11063 = n10987 & n11062;
  assign n11064 = n11057 & n11063;
  assign n11065 = n11061 & n11064;
  assign n11066 = n11006 & n11065;
  assign n11067 = n2706 & n8935;
  assign n11068 = n11066 & n11067;
  assign n11069 = n10161 & n11052;
  assign n11070 = n11068 & n11069;
  assign n11071 = ~pi0074 & ~n11070;
  assign n11072 = pi0074 & ~n8962;
  assign n11073 = n7363 & ~po1038;
  assign n11074 = ~n11071 & n11073;
  assign po0207 = ~n11072 & n11074;
  assign n11076 = pi0024 & n8897;
  assign n11077 = ~n10374 & ~n11076;
  assign n11078 = ~pi0252 & ~n8888;
  assign n11079 = pi0252 & ~po0840;
  assign n11080 = ~n11078 & ~n11079;
  assign n11081 = pi0024 & ~pi0094;
  assign n11082 = ~n8899 & n11081;
  assign n11083 = n10162 & n11080;
  assign n11084 = ~n11082 & n11083;
  assign n11085 = ~n11077 & n11084;
  assign n11086 = n2962 & n7450;
  assign n11087 = pi0024 & ~pi0090;
  assign n11088 = n11086 & n11087;
  assign n11089 = ~n11080 & n11088;
  assign n11090 = n8901 & n11089;
  assign n11091 = ~n11085 & ~n11090;
  assign n11092 = ~pi0100 & ~n11091;
  assign n11093 = pi0100 & ~n6263;
  assign n11094 = n6353 & n11093;
  assign n11095 = ~n11092 & ~n11094;
  assign n11096 = n2530 & n2533;
  assign n11097 = ~n11095 & n11096;
  assign n11098 = n6282 & n8967;
  assign n11099 = n8963 & n11098;
  assign n11100 = ~n11097 & ~n11099;
  assign po0208 = n8881 & ~n11100;
  assign n11102 = n9082 & n11057;
  assign n11103 = n2467 & n11102;
  assign n11104 = ~pi0069 & n11103;
  assign n11105 = n2804 & n11104;
  assign n11106 = n2700 & n10166;
  assign n11107 = n2754 & n11106;
  assign n11108 = n2807 & n11105;
  assign po0209 = n11107 & n11108;
  assign n11110 = ~pi0219 & n10846;
  assign n11111 = pi0052 & ~pi0072;
  assign n11112 = ~pi0039 & ~n11111;
  assign n11113 = ~n10525 & ~n11112;
  assign n11114 = ~n7429 & ~n11113;
  assign n11115 = ~n10601 & n10609;
  assign n11116 = pi0039 & ~n11115;
  assign n11117 = n6267 & n6270;
  assign n11118 = ~n11111 & ~n11117;
  assign n11119 = ~pi0052 & n10558;
  assign n11120 = pi0052 & n10554;
  assign n11121 = n11117 & ~n11119;
  assign n11122 = ~n11120 & n11121;
  assign n11123 = ~pi0228 & ~n11118;
  assign n11124 = ~n11122 & n11123;
  assign n11125 = ~pi0114 & n6267;
  assign n11126 = ~pi0052 & n10573;
  assign n11127 = pi0052 & n10570;
  assign n11128 = n10491 & ~n11126;
  assign n11129 = ~n11127 & n11128;
  assign n11130 = ~pi0052 & n10580;
  assign n11131 = pi0052 & n10587;
  assign n11132 = n10578 & ~n11130;
  assign n11133 = ~n11131 & n11132;
  assign n11134 = ~n11129 & ~n11133;
  assign n11135 = n11125 & ~n11134;
  assign n11136 = pi0228 & ~n11118;
  assign n11137 = ~n11135 & n11136;
  assign n11138 = ~pi0039 & ~n11124;
  assign n11139 = ~n11137 & n11138;
  assign n11140 = ~n11116 & ~n11139;
  assign n11141 = n2608 & ~n11140;
  assign n11142 = pi0038 & ~n11113;
  assign n11143 = n7506 & n10491;
  assign n11144 = n11125 & n11143;
  assign n11145 = n7479 & n11144;
  assign n11146 = n10616 & n11145;
  assign n11147 = n11111 & ~n11146;
  assign n11148 = ~pi0039 & ~n11147;
  assign n11149 = ~n10525 & ~n11148;
  assign n11150 = n6285 & ~n11149;
  assign n11151 = ~n11142 & ~n11150;
  assign n11152 = ~n11141 & n11151;
  assign n11153 = ~pi0087 & ~n11152;
  assign n11154 = ~n2608 & n11113;
  assign n11155 = pi0087 & ~n11154;
  assign n11156 = pi0228 & n11117;
  assign n11157 = ~pi0052 & n10501;
  assign n11158 = pi0052 & n10617;
  assign n11159 = ~n11157 & ~n11158;
  assign n11160 = n11156 & ~n11159;
  assign n11161 = n11111 & ~n11156;
  assign n11162 = ~n11160 & ~n11161;
  assign n11163 = ~pi0039 & n11162;
  assign n11164 = n2608 & ~n10525;
  assign n11165 = ~n11163 & n11164;
  assign n11166 = n11155 & ~n11165;
  assign n11167 = n10487 & ~n11166;
  assign n11168 = ~n11153 & n11167;
  assign n11169 = ~n10817 & ~n11112;
  assign n11170 = ~n2608 & n11169;
  assign n11171 = n2608 & ~n10874;
  assign n11172 = ~n11163 & n11171;
  assign n11173 = n11155 & ~n11170;
  assign n11174 = ~n11172 & n11173;
  assign n11175 = ~n10886 & ~n11139;
  assign n11176 = n2608 & ~n11175;
  assign n11177 = ~n10874 & ~n11148;
  assign n11178 = n6285 & ~n11177;
  assign n11179 = pi0038 & ~n11169;
  assign n11180 = ~n11113 & n11179;
  assign n11181 = ~n11178 & ~n11180;
  assign n11182 = ~n11176 & n11181;
  assign n11183 = ~pi0087 & ~n11182;
  assign n11184 = ~n10487 & ~n11174;
  assign n11185 = ~n11183 & n11184;
  assign n11186 = ~n11168 & ~n11185;
  assign n11187 = ~pi0075 & ~n11186;
  assign n11188 = n10498 & n11144;
  assign n11189 = n2620 & n11188;
  assign n11190 = ~pi0039 & n11111;
  assign n11191 = ~n11189 & n11190;
  assign n11192 = ~pi0039 & ~n11191;
  assign n11193 = ~n10487 & n10874;
  assign n11194 = n10487 & n10525;
  assign n11195 = pi0075 & ~n11194;
  assign n11196 = ~n11193 & n11195;
  assign n11197 = ~n11192 & n11196;
  assign n11198 = n7429 & ~n11197;
  assign n11199 = ~n11187 & n11198;
  assign n11200 = n11110 & ~n11114;
  assign n11201 = ~n11199 & n11200;
  assign n11202 = ~n7429 & ~n10487;
  assign n11203 = n11169 & n11202;
  assign n11204 = ~n7429 & ~n11190;
  assign n11205 = pi0075 & n11191;
  assign n11206 = pi0100 & ~n11190;
  assign n11207 = pi0038 & ~n11190;
  assign n11208 = ~pi0038 & n11162;
  assign n11209 = ~n11207 & ~n11208;
  assign n11210 = ~pi0100 & ~n11209;
  assign n11211 = ~pi0100 & n10982;
  assign n11212 = pi0087 & ~n11211;
  assign n11213 = ~n11206 & n11212;
  assign n11214 = ~n11210 & n11213;
  assign n11215 = pi0100 & ~n11147;
  assign n11216 = ~pi0100 & n11139;
  assign n11217 = ~pi0039 & ~n11215;
  assign n11218 = ~n11216 & n11217;
  assign n11219 = ~pi0038 & ~n11218;
  assign n11220 = ~pi0087 & ~n11207;
  assign n11221 = ~n11219 & n11220;
  assign n11222 = ~n11214 & ~n11221;
  assign n11223 = ~pi0075 & ~n11222;
  assign n11224 = n7429 & ~n11205;
  assign n11225 = ~n11223 & n11224;
  assign n11226 = n10487 & ~n11204;
  assign n11227 = ~n11225 & n11226;
  assign n11228 = n2608 & ~n10817;
  assign n11229 = ~n11163 & n11228;
  assign n11230 = ~n11170 & ~n11229;
  assign n11231 = pi0087 & ~n11230;
  assign n11232 = ~n10828 & ~n11139;
  assign n11233 = n2608 & ~n11232;
  assign n11234 = ~n10817 & ~n11148;
  assign n11235 = n6285 & ~n11234;
  assign n11236 = ~pi0087 & ~n11179;
  assign n11237 = ~n11235 & n11236;
  assign n11238 = ~n11233 & n11237;
  assign n11239 = ~pi0075 & ~n11231;
  assign n11240 = ~n11238 & n11239;
  assign n11241 = ~n2620 & n11169;
  assign n11242 = n11111 & ~n11188;
  assign n11243 = ~pi0039 & ~n11242;
  assign n11244 = n2620 & ~n10817;
  assign n11245 = ~n11243 & n11244;
  assign n11246 = pi0075 & ~n11241;
  assign n11247 = ~n11245 & n11246;
  assign n11248 = n7429 & ~n10487;
  assign n11249 = ~n11247 & n11248;
  assign n11250 = ~n11240 & n11249;
  assign n11251 = ~n11227 & ~n11250;
  assign n11252 = ~n11110 & ~n11251;
  assign n11253 = ~po1038 & ~n11203;
  assign n11254 = ~n11201 & n11253;
  assign n11255 = ~n11252 & n11254;
  assign n11256 = pi0039 & n11110;
  assign n11257 = n10523 & n11256;
  assign n11258 = po1038 & ~n11190;
  assign n11259 = ~n11257 & n11258;
  assign po0210 = ~n11255 & ~n11259;
  assign n11261 = ~pi0287 & ~pi0979;
  assign n11262 = n6181 & n11261;
  assign n11263 = pi0039 & ~n11262;
  assign n11264 = pi0024 & n10162;
  assign n11265 = pi0053 & n2720;
  assign n11266 = n2717 & n11265;
  assign n11267 = n2721 & n11266;
  assign n11268 = n11264 & n11267;
  assign n11269 = ~pi0039 & ~n11268;
  assign n11270 = n10200 & ~n11263;
  assign n11271 = ~n11269 & n11270;
  assign po0211 = ~n3402 & n11271;
  assign n11273 = n8897 & n9254;
  assign n11274 = ~pi0060 & ~pi0085;
  assign n11275 = pi0106 & n11274;
  assign n11276 = n2479 & n8913;
  assign n11277 = n11275 & n11276;
  assign n11278 = n10989 & n11277;
  assign n11279 = n8919 & n11059;
  assign n11280 = n11278 & n11279;
  assign n11281 = n11057 & n11280;
  assign n11282 = n11273 & n11281;
  assign n11283 = ~pi0841 & n2704;
  assign n11284 = n8960 & n11283;
  assign n11285 = n2611 & n2706;
  assign n11286 = n11284 & n11285;
  assign n11287 = n11282 & n11286;
  assign n11288 = ~pi0054 & ~n11287;
  assign n11289 = n2621 & n10195;
  assign n11290 = pi0054 & ~n11289;
  assign n11291 = n8880 & ~n11288;
  assign po0212 = ~n11290 & n11291;
  assign n11293 = ~pi0054 & n11289;
  assign n11294 = ~pi0074 & n11293;
  assign n11295 = pi0055 & ~n11294;
  assign n11296 = pi0045 & n2479;
  assign n11297 = n2487 & n11296;
  assign n11298 = n11061 & n11297;
  assign n11299 = n2476 & n11298;
  assign n11300 = n6479 & n9500;
  assign n11301 = n2465 & n2572;
  assign n11302 = n11300 & n11301;
  assign n11303 = n11299 & n11302;
  assign n11304 = ~pi0055 & ~n11303;
  assign n11305 = n8878 & ~n11304;
  assign po0213 = ~n11295 & n11305;
  assign n11307 = n2518 & n2537;
  assign n11308 = n6172 & n11307;
  assign n11309 = pi0056 & ~n11308;
  assign n11310 = pi0056 & ~pi0062;
  assign n11311 = pi0055 & n10068;
  assign n11312 = ~n11310 & ~n11311;
  assign n11313 = n3328 & ~n11309;
  assign po0214 = ~n11312 & n11313;
  assign n11315 = n6304 & n11294;
  assign n11316 = pi0057 & ~n11315;
  assign n11317 = n6485 & n11307;
  assign n11318 = ~pi0056 & pi0062;
  assign n11319 = ~pi0924 & n11318;
  assign n11320 = ~n11310 & ~n11319;
  assign n11321 = n11317 & ~n11320;
  assign n11322 = ~pi0057 & ~n11321;
  assign n11323 = ~pi0059 & ~n11316;
  assign po0215 = ~n11322 & n11323;
  assign n11325 = ~pi0093 & n11086;
  assign n11326 = n10165 & n11325;
  assign po0216 = n7433 & n11326;
  assign n11328 = pi0059 & ~n11315;
  assign n11329 = pi0924 & n11318;
  assign n11330 = n11317 & n11329;
  assign n11331 = ~pi0059 & ~n11330;
  assign n11332 = ~pi0057 & ~n11328;
  assign po0217 = ~n11331 & n11332;
  assign n11334 = pi0039 & ~pi0979;
  assign n11335 = ~n6181 & n11334;
  assign n11336 = n6182 & n11335;
  assign n11337 = n6380 & n11336;
  assign n11338 = ~pi0039 & n11264;
  assign n11339 = n11273 & n11338;
  assign n11340 = n2718 & n11339;
  assign n11341 = ~n11337 & ~n11340;
  assign po0218 = n10200 & ~n11341;
  assign n11343 = pi0841 & n11000;
  assign n11344 = ~pi0024 & n11273;
  assign n11345 = n2718 & n11344;
  assign n11346 = ~n11343 & ~n11345;
  assign po0219 = n10166 & ~n11346;
  assign n11348 = pi0057 & ~n10069;
  assign n11349 = n11308 & n11318;
  assign n11350 = ~pi0057 & ~n11349;
  assign n11351 = ~pi0059 & ~n11348;
  assign po0220 = ~n11350 & n11351;
  assign n11353 = n2861 & n8935;
  assign n11354 = n9100 & n11353;
  assign n11355 = pi0999 & n11354;
  assign n11356 = ~pi0024 & n11002;
  assign n11357 = ~n11355 & ~n11356;
  assign po0221 = n10166 & ~n11357;
  assign n11359 = ~pi0063 & pi0107;
  assign n11360 = n9100 & n11359;
  assign n11361 = ~pi0841 & ~n11360;
  assign n11362 = n2486 & n11359;
  assign n11363 = ~pi0064 & ~n11362;
  assign n11364 = n2465 & ~n11363;
  assign n11365 = n10169 & n11364;
  assign n11366 = pi0841 & ~n11365;
  assign n11367 = n11107 & ~n11361;
  assign po0222 = ~n11366 & n11367;
  assign n11369 = pi0039 & n10201;
  assign n11370 = n10200 & n11369;
  assign n11371 = ~n10217 & n11370;
  assign po0223 = ~n10223 & n11371;
  assign n11373 = pi0199 & ~pi0299;
  assign n11374 = n2570 & n2608;
  assign n11375 = pi0314 & n2464;
  assign n11376 = n11300 & n11375;
  assign n11377 = pi0081 & ~pi0102;
  assign n11378 = n11376 & n11377;
  assign n11379 = n2489 & n11378;
  assign n11380 = n2609 & n11373;
  assign n11381 = n11374 & n11380;
  assign n11382 = n11379 & n11381;
  assign n11383 = ~pi0219 & ~n11382;
  assign n11384 = ~pi0199 & ~pi0299;
  assign n11385 = n2572 & n11379;
  assign n11386 = ~n11384 & n11385;
  assign n11387 = pi0219 & ~n11386;
  assign n11388 = ~po1038 & ~n11383;
  assign po0224 = ~n11387 & n11388;
  assign n11390 = pi0083 & ~pi0103;
  assign n11391 = n11102 & n11390;
  assign n11392 = n10165 & n11391;
  assign n11393 = n11376 & n11392;
  assign po0225 = n2484 & n11393;
  assign n11395 = ~n6244 & n6396;
  assign n11396 = n3310 & n5853;
  assign n11397 = n11395 & n11396;
  assign n11398 = ~n6207 & n6396;
  assign n11399 = n3351 & n3470;
  assign n11400 = n11398 & n11399;
  assign n11401 = ~n11397 & ~n11400;
  assign po0226 = n10983 & ~n11401;
  assign n11403 = pi0069 & n11058;
  assign n11404 = n10153 & n11403;
  assign n11405 = ~pi0071 & ~n11404;
  assign n11406 = ~pi0081 & ~pi0314;
  assign n11407 = n2465 & n11406;
  assign n11408 = n6438 & n11407;
  assign n11409 = ~n11405 & n11408;
  assign n11410 = pi0071 & pi0314;
  assign n11411 = n7438 & n11410;
  assign n11412 = n10150 & n11411;
  assign n11413 = n2485 & n11412;
  assign n11414 = ~n11409 & ~n11413;
  assign po0227 = n11107 & ~n11414;
  assign n11416 = n2505 & n2749;
  assign n11417 = ~pi0096 & n11416;
  assign n11418 = n10194 & n11417;
  assign n11419 = pi0198 & pi0589;
  assign n11420 = n3471 & ~n6207;
  assign n11421 = n11419 & n11420;
  assign n11422 = pi0210 & pi0589;
  assign n11423 = ~pi0221 & n5853;
  assign n11424 = ~pi0216 & n11423;
  assign n11425 = ~n6244 & n11424;
  assign n11426 = n11422 & n11425;
  assign n11427 = ~n11421 & ~n11426;
  assign n11428 = ~pi0593 & n6381;
  assign n11429 = ~n6389 & n11428;
  assign n11430 = ~n11427 & n11429;
  assign n11431 = ~pi0287 & ~n11430;
  assign n11432 = pi0039 & ~n11431;
  assign n11433 = n2521 & n11432;
  assign n11434 = ~n11418 & ~n11433;
  assign po0228 = n10200 & ~n11434;
  assign n11436 = n2469 & n2481;
  assign n11437 = n6424 & n11436;
  assign n11438 = n11014 & n11437;
  assign n11439 = ~pi0064 & n8916;
  assign n11440 = n11438 & n11439;
  assign n11441 = ~pi0081 & ~n11440;
  assign n11442 = ~pi0050 & n8935;
  assign n11443 = n6444 & n11442;
  assign n11444 = ~pi0199 & pi0200;
  assign n11445 = ~pi0299 & n11444;
  assign n11446 = pi0211 & ~pi0219;
  assign n11447 = pi0299 & n11446;
  assign n11448 = ~n11445 & ~n11447;
  assign n11449 = pi0314 & ~n11448;
  assign n11450 = n10162 & n11449;
  assign n11451 = ~n11441 & n11450;
  assign n11452 = n11443 & n11451;
  assign n11453 = n11012 & n11448;
  assign n11454 = n11376 & n11453;
  assign n11455 = n11438 & n11454;
  assign n11456 = ~n11452 & ~n11455;
  assign po0229 = n10165 & ~n11456;
  assign n11458 = pi0024 & n2709;
  assign n11459 = pi0072 & n11458;
  assign n11460 = pi0088 & n10147;
  assign n11461 = n6388 & n9141;
  assign n11462 = n11460 & n11461;
  assign n11463 = n2870 & n11462;
  assign n11464 = ~n11459 & ~n11463;
  assign n11465 = n6479 & ~n11464;
  assign n11466 = ~pi0039 & ~n11465;
  assign n11467 = n7604 & n11395;
  assign n11468 = n7608 & n11398;
  assign n11469 = pi0039 & ~n11467;
  assign n11470 = ~n11468 & n11469;
  assign n11471 = n10200 & ~n11470;
  assign po0230 = ~n11466 & n11471;
  assign n11473 = ~pi0314 & pi1050;
  assign n11474 = n9090 & n10162;
  assign n11475 = n11473 & n11474;
  assign n11476 = ~pi0039 & ~n11475;
  assign n11477 = n9051 & n11398;
  assign n11478 = ~pi0299 & ~n11477;
  assign n11479 = n9036 & n11395;
  assign n11480 = pi0299 & ~n11479;
  assign n11481 = ~n11478 & ~n11480;
  assign n11482 = pi0039 & ~n11481;
  assign n11483 = n10200 & ~n11476;
  assign po0231 = ~n11482 & n11483;
  assign n11485 = pi0074 & n11293;
  assign n11486 = n2964 & n7526;
  assign n11487 = ~pi0096 & ~n11486;
  assign n11488 = ~pi0096 & ~pi1093;
  assign n11489 = n7417 & n11488;
  assign n11490 = ~pi0096 & ~n6169;
  assign n11491 = pi0479 & ~n11490;
  assign n11492 = n3373 & n7429;
  assign n11493 = ~n11489 & n11492;
  assign n11494 = ~po0840 & ~n11491;
  assign n11495 = n11493 & n11494;
  assign n11496 = ~n11487 & n11495;
  assign n11497 = n7456 & n11496;
  assign n11498 = ~n11485 & ~n11497;
  assign po0232 = ~po1038 & ~n11498;
  assign n11500 = n2620 & n10195;
  assign n11501 = pi0075 & ~n11500;
  assign n11502 = pi0096 & ~pi1093;
  assign n11503 = n2931 & ~n11487;
  assign n11504 = ~n11502 & ~n11503;
  assign n11505 = n2610 & ~n11504;
  assign n11506 = n7534 & n11505;
  assign n11507 = ~pi0075 & ~n11506;
  assign n11508 = n8881 & ~n11501;
  assign po0233 = ~n11507 & n11508;
  assign n11510 = n8930 & n10186;
  assign n11511 = ~n10111 & n11510;
  assign n11512 = po1057 & ~n11511;
  assign n11513 = n2519 & n10375;
  assign n11514 = pi0252 & n2933;
  assign n11515 = n11513 & ~n11514;
  assign n11516 = ~pi0137 & n11515;
  assign n11517 = ~pi0137 & n2924;
  assign n11518 = ~pi0094 & ~n8931;
  assign n11519 = ~n8897 & ~n10374;
  assign n11520 = n10162 & ~n11518;
  assign n11521 = ~n11519 & n11520;
  assign n11522 = ~n2933 & ~n11521;
  assign n11523 = ~pi0252 & n11521;
  assign n11524 = pi0252 & n11510;
  assign n11525 = n2933 & ~n11524;
  assign n11526 = ~n11523 & n11525;
  assign n11527 = ~n11522 & ~n11526;
  assign n11528 = pi0122 & ~n11527;
  assign n11529 = n7417 & n11522;
  assign n11530 = ~n6277 & ~n11513;
  assign n11531 = ~n11526 & ~n11530;
  assign n11532 = ~n11529 & n11531;
  assign n11533 = ~pi0122 & ~n11532;
  assign n11534 = ~n11528 & ~n11533;
  assign n11535 = ~pi1093 & ~n11534;
  assign n11536 = ~pi0122 & ~n11515;
  assign n11537 = ~n11528 & ~n11536;
  assign n11538 = pi1093 & ~n11537;
  assign n11539 = ~n11535 & ~n11538;
  assign n11540 = n2924 & ~n11539;
  assign n11541 = ~n11517 & ~n11540;
  assign n11542 = ~n11516 & ~n11541;
  assign n11543 = ~pi0122 & n11513;
  assign n11544 = pi1093 & ~n11521;
  assign n11545 = ~n7418 & ~n11544;
  assign n11546 = ~n11543 & ~n11545;
  assign n11547 = ~n11535 & ~n11546;
  assign n11548 = ~n2924 & ~n11547;
  assign n11549 = ~pi0137 & ~n2924;
  assign n11550 = ~n11548 & ~n11549;
  assign n11551 = pi0252 & pi1092;
  assign n11552 = ~pi1093 & n11551;
  assign n11553 = n2925 & n11552;
  assign n11554 = ~pi0137 & ~n11553;
  assign n11555 = n11513 & n11554;
  assign n11556 = ~n11550 & ~n11555;
  assign n11557 = ~n11542 & ~n11556;
  assign n11558 = ~po1057 & ~n11557;
  assign n11559 = ~pi0137 & po1057;
  assign n11560 = ~n11512 & ~n11559;
  assign n11561 = ~n11558 & n11560;
  assign n11562 = ~pi0210 & ~n11561;
  assign n11563 = ~n11540 & ~n11548;
  assign n11564 = ~po1057 & ~n11563;
  assign n11565 = ~n11512 & ~n11564;
  assign n11566 = pi0210 & ~n11565;
  assign n11567 = ~n11562 & ~n11566;
  assign n11568 = n2638 & n10299;
  assign n11569 = ~n11567 & ~n11568;
  assign n11570 = ~pi0210 & ~n11557;
  assign n11571 = pi0210 & ~n11563;
  assign n11572 = ~n11570 & ~n11571;
  assign n11573 = n11568 & ~n11572;
  assign n11574 = pi0299 & ~n11573;
  assign n11575 = ~n11569 & n11574;
  assign n11576 = ~pi0198 & ~n11561;
  assign n11577 = pi0198 & ~n11565;
  assign n11578 = ~n11576 & ~n11577;
  assign n11579 = n2669 & n6197;
  assign n11580 = ~n11578 & ~n11579;
  assign n11581 = pi0198 & ~n11563;
  assign n11582 = ~pi0198 & ~n11557;
  assign n11583 = ~n11581 & ~n11582;
  assign n11584 = n11579 & ~n11583;
  assign n11585 = ~pi0299 & ~n11584;
  assign n11586 = ~n11580 & n11585;
  assign n11587 = ~n11575 & ~n11586;
  assign n11588 = pi0232 & ~n11587;
  assign n11589 = pi0299 & ~n11567;
  assign n11590 = ~pi0299 & ~n11578;
  assign n11591 = ~pi0232 & ~n11589;
  assign n11592 = ~n11590 & n11591;
  assign n11593 = ~n11588 & ~n11592;
  assign n11594 = n7425 & ~n11593;
  assign n11595 = ~n2924 & n11544;
  assign n11596 = n2933 & ~n11513;
  assign n11597 = ~n11514 & ~n11522;
  assign n11598 = ~n11596 & n11597;
  assign n11599 = n7418 & ~n11598;
  assign n11600 = ~n11528 & ~n11599;
  assign n11601 = n2924 & ~n11600;
  assign n11602 = ~pi1093 & ~n11527;
  assign n11603 = ~n11595 & ~n11602;
  assign n11604 = ~n11601 & n11603;
  assign n11605 = ~po1057 & n11604;
  assign n11606 = po1057 & n11510;
  assign n11607 = ~n10108 & n11606;
  assign n11608 = ~n11605 & ~n11607;
  assign n11609 = pi0210 & ~n11608;
  assign n11610 = n8904 & n11559;
  assign n11611 = pi0137 & n11602;
  assign n11612 = ~pi0137 & ~n11598;
  assign n11613 = ~pi1093 & n11612;
  assign n11614 = ~n11544 & ~n11611;
  assign n11615 = ~n11613 & n11614;
  assign n11616 = ~po1057 & n11615;
  assign n11617 = ~n11606 & ~n11616;
  assign n11618 = ~n2924 & ~n11610;
  assign n11619 = ~n11617 & n11618;
  assign n11620 = pi0137 & ~n7418;
  assign n11621 = n2933 & ~n11620;
  assign n11622 = n11510 & ~n11621;
  assign n11623 = po1057 & ~n11622;
  assign n11624 = pi0137 & ~n11600;
  assign n11625 = ~n11611 & ~n11612;
  assign n11626 = ~n11624 & n11625;
  assign n11627 = ~po1057 & ~n11626;
  assign n11628 = n2924 & ~n11623;
  assign n11629 = ~n11627 & n11628;
  assign n11630 = ~n11619 & ~n11629;
  assign n11631 = ~pi0210 & ~n11630;
  assign n11632 = ~n11609 & ~n11631;
  assign n11633 = ~n11568 & ~n11632;
  assign n11634 = ~n2924 & n11615;
  assign n11635 = n2924 & n11626;
  assign n11636 = ~n11634 & ~n11635;
  assign n11637 = ~pi0210 & n11636;
  assign n11638 = pi0210 & ~n11604;
  assign n11639 = n11568 & ~n11638;
  assign n11640 = ~n11637 & n11639;
  assign n11641 = pi0299 & ~n11640;
  assign n11642 = ~n11633 & n11641;
  assign n11643 = pi0198 & ~n11608;
  assign n11644 = ~pi0198 & ~n11630;
  assign n11645 = ~n11643 & ~n11644;
  assign n11646 = ~n11579 & ~n11645;
  assign n11647 = ~pi0198 & ~n11636;
  assign n11648 = pi0198 & n11604;
  assign n11649 = ~n11647 & ~n11648;
  assign n11650 = n11579 & ~n11649;
  assign n11651 = ~pi0299 & ~n11650;
  assign n11652 = ~n11646 & n11651;
  assign n11653 = ~n11642 & ~n11652;
  assign n11654 = pi0232 & ~n11653;
  assign n11655 = ~pi0299 & ~n11645;
  assign n11656 = pi0299 & ~n11632;
  assign n11657 = ~pi0232 & ~n11655;
  assign n11658 = ~n11656 & n11657;
  assign n11659 = ~n7425 & ~n11658;
  assign n11660 = ~n11654 & n11659;
  assign n11661 = ~n11594 & ~n11660;
  assign po0234 = n10165 & ~n11661;
  assign n11663 = pi0086 & n8897;
  assign n11664 = n2778 & n11663;
  assign n11665 = pi0314 & ~n11664;
  assign n11666 = n2769 & n2784;
  assign n11667 = ~pi0086 & ~n11666;
  assign n11668 = n6452 & ~n11667;
  assign n11669 = n2702 & n11668;
  assign n11670 = ~pi0314 & ~n11669;
  assign n11671 = n10166 & ~n11665;
  assign po0235 = ~n11670 & n11671;
  assign n11673 = pi0119 & pi0232;
  assign po0236 = ~pi0468 & n11673;
  assign n11675 = pi0163 & ~n9700;
  assign n11676 = ~pi0163 & ~n9696;
  assign n11677 = ~n9698 & n11676;
  assign n11678 = ~n11675 & ~n11677;
  assign n11679 = pi0232 & n11678;
  assign n11680 = ~n8989 & n11679;
  assign n11681 = pi0074 & ~n11680;
  assign n11682 = pi0075 & ~n11679;
  assign n11683 = pi0100 & ~n11679;
  assign n11684 = ~n11682 & ~n11683;
  assign n11685 = pi0147 & n7473;
  assign n11686 = n8989 & n11685;
  assign n11687 = n11684 & ~n11686;
  assign n11688 = ~n3328 & ~n11681;
  assign n11689 = n11687 & n11688;
  assign n11690 = pi0054 & ~n11687;
  assign n11691 = ~pi0038 & ~pi0040;
  assign n11692 = pi0038 & ~n11685;
  assign n11693 = ~pi0100 & ~n11692;
  assign n11694 = ~n11691 & n11693;
  assign n11695 = ~n11683 & ~n11694;
  assign n11696 = ~pi0075 & ~n11695;
  assign n11697 = ~n11682 & ~n11696;
  assign n11698 = ~pi0054 & ~n11697;
  assign n11699 = ~n11690 & ~n11698;
  assign n11700 = ~pi0074 & ~n11699;
  assign n11701 = ~n11681 & ~n11700;
  assign n11702 = ~n2529 & ~n11701;
  assign n11703 = n3328 & ~n11702;
  assign n11704 = ~n9722 & n9724;
  assign n11705 = ~pi0184 & n11704;
  assign n11706 = pi0184 & n6197;
  assign n11707 = ~n11704 & n11706;
  assign n11708 = ~pi0299 & ~n11705;
  assign n11709 = ~n11707 & n11708;
  assign n11710 = pi0299 & ~n11678;
  assign n11711 = pi0232 & ~n11709;
  assign n11712 = ~n11710 & n11711;
  assign n11713 = ~n8989 & n11712;
  assign n11714 = pi0074 & ~n11713;
  assign n11715 = ~pi0055 & ~n11714;
  assign n11716 = ~pi0187 & ~pi0299;
  assign n11717 = ~pi0147 & pi0299;
  assign n11718 = ~n11716 & ~n11717;
  assign n11719 = n7473 & n11718;
  assign n11720 = n8989 & ~n11719;
  assign n11721 = pi0054 & ~n11720;
  assign n11722 = ~n11713 & n11721;
  assign n11723 = pi0075 & ~n11712;
  assign n11724 = pi0100 & ~n11712;
  assign n11725 = pi0038 & ~n11719;
  assign n11726 = ~pi0100 & ~n11725;
  assign n11727 = ~pi0179 & ~pi0299;
  assign n11728 = ~pi0156 & pi0299;
  assign n11729 = ~n11727 & ~n11728;
  assign n11730 = n7473 & n11729;
  assign n11731 = n2518 & n2609;
  assign n11732 = n11730 & n11731;
  assign n11733 = n2509 & n11732;
  assign n11734 = n11691 & ~n11733;
  assign n11735 = n11726 & ~n11734;
  assign n11736 = ~n11724 & ~n11735;
  assign n11737 = n9205 & ~n11736;
  assign n11738 = ~pi0187 & ~n9187;
  assign n11739 = pi0187 & ~n9189;
  assign n11740 = pi0147 & ~n11739;
  assign n11741 = ~n11738 & n11740;
  assign n11742 = ~pi0147 & pi0187;
  assign n11743 = n9194 & n11742;
  assign n11744 = ~n11741 & ~n11743;
  assign n11745 = pi0038 & ~n11744;
  assign n11746 = n2509 & n9093;
  assign n11747 = ~n6242 & n9036;
  assign n11748 = pi0156 & n6188;
  assign n11749 = ~pi0166 & n9293;
  assign n11750 = ~n11748 & ~n11749;
  assign n11751 = n11747 & ~n11750;
  assign n11752 = n11746 & n11751;
  assign n11753 = ~pi0040 & pi0299;
  assign n11754 = ~n11752 & n11753;
  assign n11755 = ~pi0189 & n9293;
  assign n11756 = pi0179 & n6188;
  assign n11757 = ~n11755 & ~n11756;
  assign n11758 = ~n6205 & n9051;
  assign n11759 = ~n11757 & n11758;
  assign n11760 = n11746 & n11759;
  assign n11761 = ~pi0040 & ~pi0299;
  assign n11762 = ~n11760 & n11761;
  assign n11763 = pi0039 & ~n11754;
  assign n11764 = ~n11762 & n11763;
  assign n11765 = ~pi0175 & ~pi0299;
  assign n11766 = pi0184 & n9147;
  assign n11767 = ~pi0184 & ~n9143;
  assign n11768 = ~pi0189 & ~n11767;
  assign n11769 = ~n11766 & n11768;
  assign n11770 = ~pi0032 & pi0095;
  assign n11771 = ~pi0479 & n11770;
  assign n11772 = n2509 & n11771;
  assign n11773 = pi0182 & n11772;
  assign n11774 = pi0184 & pi0189;
  assign n11775 = ~n9150 & n11774;
  assign n11776 = ~n11773 & ~n11775;
  assign n11777 = ~n11769 & n11776;
  assign n11778 = n6197 & ~n11777;
  assign n11779 = ~pi0040 & ~n11778;
  assign n11780 = n11765 & ~n11779;
  assign n11781 = n6197 & n11772;
  assign n11782 = pi0153 & n9093;
  assign n11783 = n9133 & n11782;
  assign n11784 = n9143 & n10299;
  assign n11785 = ~pi0040 & ~pi0163;
  assign n11786 = ~n11784 & n11785;
  assign n11787 = ~n11783 & n11786;
  assign n11788 = ~n11781 & n11787;
  assign n11789 = pi0040 & ~n6197;
  assign n11790 = pi0166 & n6197;
  assign n11791 = ~pi0040 & ~n11772;
  assign n11792 = n9166 & n11791;
  assign n11793 = n11790 & ~n11792;
  assign n11794 = n9162 & n11791;
  assign n11795 = n10299 & ~n11794;
  assign n11796 = ~pi0153 & ~n11793;
  assign n11797 = ~n11795 & n11796;
  assign n11798 = ~pi0210 & ~n9120;
  assign n11799 = ~n9118 & n11791;
  assign n11800 = ~n11798 & n11799;
  assign n11801 = n10299 & ~n11800;
  assign n11802 = ~n9129 & n11792;
  assign n11803 = n11790 & ~n11802;
  assign n11804 = pi0153 & ~n11803;
  assign n11805 = ~n11801 & n11804;
  assign n11806 = ~n11797 & ~n11805;
  assign n11807 = pi0163 & ~n11789;
  assign n11808 = ~n11806 & n11807;
  assign n11809 = pi0160 & ~n11808;
  assign n11810 = pi0153 & n9118;
  assign n11811 = n9162 & ~n11810;
  assign n11812 = n10299 & ~n11811;
  assign n11813 = pi0153 & n9129;
  assign n11814 = n9166 & ~n11813;
  assign n11815 = n11790 & ~n11814;
  assign n11816 = ~pi0040 & pi0163;
  assign n11817 = ~n11815 & n11816;
  assign n11818 = ~n11812 & n11817;
  assign n11819 = ~pi0160 & ~n11787;
  assign n11820 = ~n11818 & n11819;
  assign n11821 = ~n11809 & ~n11820;
  assign n11822 = pi0299 & ~n11788;
  assign n11823 = ~n11821 & n11822;
  assign n11824 = ~n9121 & n11799;
  assign n11825 = n10295 & ~n11824;
  assign n11826 = pi0189 & n6197;
  assign n11827 = n9130 & n11791;
  assign n11828 = n11826 & ~n11827;
  assign n11829 = pi0182 & pi0184;
  assign n11830 = ~n11789 & n11829;
  assign n11831 = ~n11828 & n11830;
  assign n11832 = ~n11825 & n11831;
  assign n11833 = pi0175 & ~pi0299;
  assign n11834 = pi0189 & ~n9133;
  assign n11835 = ~pi0189 & ~n9092;
  assign n11836 = n2518 & ~n11834;
  assign n11837 = ~n11835 & n11836;
  assign n11838 = ~n11773 & ~n11837;
  assign n11839 = n6197 & ~n11838;
  assign n11840 = ~pi0184 & ~n11839;
  assign n11841 = pi0189 & n9131;
  assign n11842 = ~n9122 & n10295;
  assign n11843 = ~pi0182 & pi0184;
  assign n11844 = ~n11841 & n11843;
  assign n11845 = ~n11842 & n11844;
  assign n11846 = ~n11840 & ~n11845;
  assign n11847 = ~pi0040 & ~n11846;
  assign n11848 = ~n11832 & n11833;
  assign n11849 = ~n11847 & n11848;
  assign n11850 = ~n11780 & ~n11849;
  assign n11851 = ~n11823 & n11850;
  assign n11852 = ~pi0039 & ~n11851;
  assign n11853 = pi0232 & ~n11764;
  assign n11854 = ~n11852 & n11853;
  assign n11855 = ~pi0040 & ~pi0232;
  assign n11856 = ~pi0038 & ~n11855;
  assign n11857 = ~n11854 & n11856;
  assign n11858 = ~n11745 & ~n11857;
  assign n11859 = n2568 & ~n11858;
  assign n11860 = pi0087 & ~n11691;
  assign n11861 = n11726 & n11860;
  assign n11862 = ~n11724 & ~n11861;
  assign n11863 = ~n11859 & n11862;
  assign n11864 = n2569 & ~n11863;
  assign n11865 = ~n11723 & ~n11737;
  assign n11866 = ~n11864 & n11865;
  assign n11867 = ~pi0054 & ~n11866;
  assign n11868 = ~n11722 & ~n11867;
  assign n11869 = ~pi0074 & ~n11868;
  assign n11870 = n11715 & ~n11869;
  assign n11871 = pi0055 & ~n11681;
  assign n11872 = pi0163 & pi0232;
  assign n11873 = ~pi0092 & n2609;
  assign n11874 = n11872 & n11873;
  assign n11875 = n11746 & n11874;
  assign n11876 = n11691 & ~n11875;
  assign n11877 = ~pi0075 & n11693;
  assign n11878 = ~n11876 & n11877;
  assign n11879 = n11684 & ~n11878;
  assign n11880 = ~pi0054 & ~n11879;
  assign n11881 = ~n11690 & ~n11880;
  assign n11882 = ~pi0074 & ~n11881;
  assign n11883 = n11871 & ~n11882;
  assign n11884 = n2529 & ~n11883;
  assign n11885 = ~n11870 & n11884;
  assign n11886 = n11703 & ~n11885;
  assign n11887 = ~n11689 & ~n11886;
  assign n11888 = pi0079 & n11887;
  assign n11889 = n2487 & ~n9260;
  assign n11890 = ~pi0040 & ~n11889;
  assign n11891 = ~n6197 & n9260;
  assign n11892 = n9248 & ~n11891;
  assign n11893 = n11872 & n11892;
  assign n11894 = n11890 & ~n11893;
  assign n11895 = ~pi0039 & ~n11894;
  assign n11896 = pi0039 & ~n9466;
  assign n11897 = n9208 & ~n11896;
  assign n11898 = ~n11895 & n11897;
  assign n11899 = pi0087 & ~n2487;
  assign n11900 = n11691 & n11899;
  assign n11901 = n11693 & ~n11900;
  assign n11902 = ~n11898 & n11901;
  assign n11903 = ~n11683 & ~n11902;
  assign n11904 = n2569 & ~n11903;
  assign n11905 = ~n9284 & n11695;
  assign n11906 = n9205 & ~n11905;
  assign n11907 = ~n11682 & ~n11906;
  assign n11908 = ~n11904 & n11907;
  assign n11909 = ~pi0054 & ~n11908;
  assign n11910 = ~n11690 & ~n11909;
  assign n11911 = ~pi0074 & ~n11910;
  assign n11912 = n11871 & ~n11911;
  assign n11913 = n11726 & ~n11900;
  assign n11914 = n2487 & n11730;
  assign n11915 = n11890 & ~n11914;
  assign n11916 = ~pi0039 & ~n11915;
  assign n11917 = n11897 & ~n11916;
  assign n11918 = n11913 & ~n11917;
  assign n11919 = ~n11724 & ~n11918;
  assign n11920 = n9205 & ~n11919;
  assign n11921 = pi0087 & n11913;
  assign n11922 = ~pi0040 & ~n9297;
  assign n11923 = n6242 & ~n11922;
  assign n11924 = n6227 & n9466;
  assign n11925 = n2487 & ~n9295;
  assign n11926 = ~pi0040 & ~n11925;
  assign n11927 = ~n6227 & n11926;
  assign n11928 = ~n11924 & ~n11927;
  assign n11929 = ~n6242 & n11928;
  assign n11930 = ~n11923 & ~n11929;
  assign n11931 = n9291 & n11930;
  assign n11932 = n6205 & ~n11922;
  assign n11933 = ~n6205 & n11928;
  assign n11934 = ~n11932 & ~n11933;
  assign n11935 = n9051 & ~n11934;
  assign n11936 = ~n9051 & ~n9466;
  assign n11937 = ~pi0299 & ~n11936;
  assign n11938 = ~n11935 & n11937;
  assign n11939 = ~pi0232 & ~n11931;
  assign n11940 = ~n11938 & n11939;
  assign n11941 = ~pi0189 & ~n11922;
  assign n11942 = n2487 & ~n9311;
  assign n11943 = n9140 & ~n11942;
  assign n11944 = n6198 & n11926;
  assign n11945 = ~n11924 & ~n11944;
  assign n11946 = ~n11943 & n11945;
  assign n11947 = pi0189 & ~n6205;
  assign n11948 = n11946 & n11947;
  assign n11949 = ~n11941 & ~n11948;
  assign n11950 = pi0179 & ~n11949;
  assign n11951 = pi0189 & ~n11928;
  assign n11952 = n9140 & n9324;
  assign n11953 = ~n2487 & n9140;
  assign n11954 = ~n11952 & ~n11953;
  assign n11955 = n11945 & n11954;
  assign n11956 = ~pi0189 & ~n11955;
  assign n11957 = ~pi0179 & ~n6205;
  assign n11958 = ~n11951 & n11957;
  assign n11959 = ~n11956 & n11958;
  assign n11960 = ~n11932 & ~n11959;
  assign n11961 = ~n11950 & n11960;
  assign n11962 = n9051 & ~n11961;
  assign n11963 = ~n11936 & ~n11962;
  assign n11964 = ~pi0299 & ~n11963;
  assign n11965 = ~n9036 & n9466;
  assign n11966 = pi0299 & ~n11965;
  assign n11967 = ~pi0166 & ~n6242;
  assign n11968 = ~n11930 & ~n11967;
  assign n11969 = n11955 & n11967;
  assign n11970 = n9036 & ~n11969;
  assign n11971 = ~n11968 & n11970;
  assign n11972 = n11966 & ~n11971;
  assign n11973 = ~n11964 & ~n11972;
  assign n11974 = ~pi0156 & pi0232;
  assign n11975 = ~n11973 & n11974;
  assign n11976 = pi0166 & ~n6242;
  assign n11977 = n11946 & n11976;
  assign n11978 = ~n11922 & ~n11976;
  assign n11979 = n9036 & ~n11978;
  assign n11980 = ~n11977 & n11979;
  assign n11981 = n11966 & ~n11980;
  assign n11982 = ~n11964 & ~n11981;
  assign n11983 = pi0156 & pi0232;
  assign n11984 = ~n11982 & n11983;
  assign n11985 = pi0039 & ~n11940;
  assign n11986 = ~n11975 & n11985;
  assign n11987 = ~n11984 & n11986;
  assign n11988 = ~n2442 & ~n9485;
  assign n11989 = n9348 & ~n9349;
  assign n11990 = ~n11988 & ~n11989;
  assign n11991 = ~pi0040 & ~n9456;
  assign n11992 = ~pi0095 & ~n11991;
  assign n11993 = ~n11990 & ~n11992;
  assign n11994 = ~pi0299 & n11993;
  assign n11995 = ~pi0040 & ~n9581;
  assign n11996 = ~pi0095 & ~n11995;
  assign n11997 = ~n11990 & ~n11996;
  assign n11998 = pi0299 & n11997;
  assign n11999 = ~pi0232 & ~n11994;
  assign n12000 = ~n11998 & n11999;
  assign n12001 = ~n6197 & n11993;
  assign n12002 = ~pi0040 & ~n9427;
  assign n12003 = ~pi0095 & ~n12002;
  assign n12004 = ~pi0040 & ~n9442;
  assign n12005 = pi0189 & n12004;
  assign n12006 = n12003 & ~n12005;
  assign n12007 = ~pi0182 & n11990;
  assign n12008 = pi0182 & n9485;
  assign n12009 = n6197 & ~n12008;
  assign n12010 = ~n12007 & n12009;
  assign n12011 = ~n12006 & n12010;
  assign n12012 = pi0184 & ~n12011;
  assign n12013 = ~pi0040 & n9403;
  assign n12014 = ~pi0032 & ~n12013;
  assign n12015 = ~n9487 & ~n12014;
  assign n12016 = ~pi0095 & ~n12015;
  assign n12017 = ~n9485 & ~n12016;
  assign n12018 = ~pi0198 & ~n12017;
  assign n12019 = ~n9467 & ~n12014;
  assign n12020 = ~pi0095 & ~n12019;
  assign n12021 = ~n9485 & ~n12020;
  assign n12022 = pi0198 & ~n12021;
  assign n12023 = n10295 & ~n12018;
  assign n12024 = ~n12022 & n12023;
  assign n12025 = n11826 & n11991;
  assign n12026 = pi0182 & ~pi0184;
  assign n12027 = ~n12024 & n12026;
  assign n12028 = ~n12025 & n12027;
  assign n12029 = ~n12012 & ~n12028;
  assign n12030 = n11765 & ~n12029;
  assign n12031 = pi0095 & ~pi0182;
  assign n12032 = ~pi0040 & ~n9503;
  assign n12033 = ~pi0095 & pi0189;
  assign n12034 = n2487 & ~n12033;
  assign n12035 = n12032 & ~n12034;
  assign n12036 = ~n12031 & ~n12035;
  assign n12037 = n11706 & ~n12036;
  assign n12038 = ~n12007 & n12037;
  assign n12039 = n9560 & n10295;
  assign n12040 = ~pi0198 & ~n9490;
  assign n12041 = ~pi0095 & ~n9479;
  assign n12042 = ~n9485 & ~n12041;
  assign n12043 = pi0198 & ~n12042;
  assign n12044 = n11826 & ~n12040;
  assign n12045 = ~n12043 & n12044;
  assign n12046 = pi0182 & ~n12039;
  assign n12047 = ~n12045 & n12046;
  assign n12048 = ~n9489 & ~n11990;
  assign n12049 = ~pi0198 & ~n12048;
  assign n12050 = ~n11990 & ~n12041;
  assign n12051 = pi0198 & ~n12050;
  assign n12052 = n11826 & ~n12049;
  assign n12053 = ~n12051 & n12052;
  assign n12054 = ~pi0182 & ~n12053;
  assign n12055 = ~n12047 & ~n12054;
  assign n12056 = ~n9560 & ~n12031;
  assign n12057 = n10295 & ~n11990;
  assign n12058 = ~n12056 & n12057;
  assign n12059 = ~n12055 & ~n12058;
  assign n12060 = ~pi0184 & ~n12059;
  assign n12061 = n11833 & ~n12038;
  assign n12062 = ~n12060 & n12061;
  assign n12063 = ~n12030 & ~n12062;
  assign n12064 = ~n12001 & ~n12063;
  assign n12065 = ~n6197 & n11997;
  assign n12066 = ~pi0095 & ~n12032;
  assign n12067 = pi0166 & ~n12066;
  assign n12068 = ~n11474 & ~n12066;
  assign n12069 = pi0153 & ~n12067;
  assign n12070 = ~n12068 & n12069;
  assign n12071 = pi0166 & n12004;
  assign n12072 = n12003 & ~n12071;
  assign n12073 = ~pi0153 & n12072;
  assign n12074 = ~pi0160 & n6197;
  assign n12075 = ~n12070 & n12074;
  assign n12076 = ~n11990 & n12075;
  assign n12077 = ~n12073 & n12076;
  assign n12078 = n6197 & ~n9485;
  assign n12079 = n12067 & n12078;
  assign n12080 = n9466 & n10299;
  assign n12081 = pi0153 & ~n12080;
  assign n12082 = ~n12079 & n12081;
  assign n12083 = ~n12072 & n12078;
  assign n12084 = ~pi0153 & ~n12083;
  assign n12085 = pi0160 & ~n12082;
  assign n12086 = ~n12084 & n12085;
  assign n12087 = pi0163 & ~n12077;
  assign n12088 = ~n12086 & n12087;
  assign n12089 = pi0210 & ~n12050;
  assign n12090 = ~pi0210 & ~n12048;
  assign n12091 = n11790 & ~n12089;
  assign n12092 = ~n12090 & n12091;
  assign n12093 = ~n9557 & ~n11990;
  assign n12094 = ~pi0210 & ~n12093;
  assign n12095 = ~n9553 & ~n11990;
  assign n12096 = pi0210 & ~n12095;
  assign n12097 = n10299 & ~n12094;
  assign n12098 = ~n12096 & n12097;
  assign n12099 = pi0153 & ~n12092;
  assign n12100 = ~n12098 & n12099;
  assign n12101 = pi0166 & n11997;
  assign n12102 = ~n11990 & ~n12020;
  assign n12103 = pi0210 & ~n12102;
  assign n12104 = ~n11990 & ~n12016;
  assign n12105 = ~pi0210 & ~n12104;
  assign n12106 = n10299 & ~n12103;
  assign n12107 = ~n12105 & n12106;
  assign n12108 = ~pi0153 & ~n12107;
  assign n12109 = ~n12101 & n12108;
  assign n12110 = ~pi0160 & ~n12100;
  assign n12111 = ~n12109 & n12110;
  assign n12112 = pi0210 & ~n9554;
  assign n12113 = ~pi0210 & ~n9558;
  assign n12114 = n10299 & ~n12112;
  assign n12115 = ~n12113 & n12114;
  assign n12116 = ~pi0210 & ~n9490;
  assign n12117 = pi0210 & ~n12042;
  assign n12118 = n11790 & ~n12116;
  assign n12119 = ~n12117 & n12118;
  assign n12120 = pi0153 & ~n12115;
  assign n12121 = ~n12119 & n12120;
  assign n12122 = n11790 & n11995;
  assign n12123 = ~pi0210 & ~n12017;
  assign n12124 = pi0210 & ~n12021;
  assign n12125 = n10299 & ~n12123;
  assign n12126 = ~n12124 & n12125;
  assign n12127 = ~pi0153 & ~n12126;
  assign n12128 = ~n12122 & n12127;
  assign n12129 = pi0160 & ~n12121;
  assign n12130 = ~n12128 & n12129;
  assign n12131 = ~pi0163 & ~n12130;
  assign n12132 = ~n12111 & n12131;
  assign n12133 = ~n12088 & ~n12132;
  assign n12134 = pi0299 & ~n12065;
  assign n12135 = ~n12133 & n12134;
  assign n12136 = ~n10295 & n11993;
  assign n12137 = pi0198 & ~n12102;
  assign n12138 = ~pi0198 & ~n12104;
  assign n12139 = n10295 & ~n12137;
  assign n12140 = ~n12138 & n12139;
  assign n12141 = ~pi0182 & ~pi0184;
  assign n12142 = n11765 & n12141;
  assign n12143 = ~n12140 & n12142;
  assign n12144 = ~n12136 & n12143;
  assign n12145 = ~n12064 & ~n12144;
  assign n12146 = ~n12135 & n12145;
  assign n12147 = pi0232 & ~n12146;
  assign n12148 = ~pi0039 & ~n12000;
  assign n12149 = ~n12147 & n12148;
  assign n12150 = ~pi0038 & ~n11987;
  assign n12151 = ~n12149 & n12150;
  assign n12152 = ~n11745 & ~n12151;
  assign n12153 = n2568 & ~n12152;
  assign n12154 = ~n11724 & ~n11921;
  assign n12155 = ~n12153 & n12154;
  assign n12156 = n2569 & ~n12155;
  assign n12157 = ~n11723 & ~n11920;
  assign n12158 = ~n12156 & n12157;
  assign n12159 = ~pi0054 & ~n12158;
  assign n12160 = ~n11722 & ~n12159;
  assign n12161 = ~pi0074 & ~n12160;
  assign n12162 = n11715 & ~n12161;
  assign n12163 = n2529 & ~n11912;
  assign n12164 = ~n12162 & n12163;
  assign n12165 = ~n9252 & n11703;
  assign n12166 = ~n12164 & n12165;
  assign n12167 = ~n11689 & ~n12166;
  assign n12168 = ~pi0079 & n12167;
  assign n12169 = ~pi0034 & n10058;
  assign n12170 = ~n11888 & ~n12169;
  assign n12171 = ~n12168 & n12170;
  assign n12172 = ~pi0079 & ~n8977;
  assign n12173 = n11887 & n12172;
  assign n12174 = n12167 & ~n12172;
  assign n12175 = n12169 & ~n12173;
  assign n12176 = ~n12174 & n12175;
  assign po0237 = n12171 | n12176;
  assign n12178 = pi0098 & pi1092;
  assign n12179 = pi1093 & n12178;
  assign n12180 = ~pi0567 & n2926;
  assign n12181 = ~n12179 & ~n12180;
  assign n12182 = ~pi0080 & ~n12181;
  assign n12183 = pi0217 & ~n12182;
  assign n12184 = n7425 & n12181;
  assign n12185 = ~n8041 & n12181;
  assign n12186 = pi0588 & ~n12185;
  assign n12187 = pi0592 & ~n8093;
  assign n12188 = n7422 & ~n8119;
  assign n12189 = ~n12187 & n12188;
  assign n12190 = n12181 & ~n12189;
  assign n12191 = ~pi1199 & ~n12190;
  assign n12192 = pi0428 & ~n12190;
  assign n12193 = ~n7644 & n12181;
  assign n12194 = ~pi0428 & ~n12193;
  assign n12195 = ~n12192 & ~n12194;
  assign n12196 = ~pi0427 & ~n12195;
  assign n12197 = ~pi0428 & ~n12190;
  assign n12198 = pi0428 & ~n12193;
  assign n12199 = ~n12197 & ~n12198;
  assign n12200 = pi0427 & ~n12199;
  assign n12201 = ~n12196 & ~n12200;
  assign n12202 = ~pi0430 & ~n12201;
  assign n12203 = ~pi0427 & ~n12199;
  assign n12204 = pi0427 & ~n12195;
  assign n12205 = ~n12203 & ~n12204;
  assign n12206 = pi0430 & ~n12205;
  assign n12207 = ~n12202 & ~n12206;
  assign n12208 = ~pi0426 & ~n12207;
  assign n12209 = ~pi0430 & ~n12205;
  assign n12210 = pi0430 & ~n12201;
  assign n12211 = ~n12209 & ~n12210;
  assign n12212 = pi0426 & ~n12211;
  assign n12213 = ~n12208 & ~n12212;
  assign n12214 = ~pi0445 & ~n12213;
  assign n12215 = ~pi0426 & ~n12211;
  assign n12216 = pi0426 & ~n12207;
  assign n12217 = ~n12215 & ~n12216;
  assign n12218 = pi0445 & ~n12217;
  assign n12219 = ~n12214 & ~n12218;
  assign n12220 = pi0448 & ~n12219;
  assign n12221 = ~pi0445 & ~n12217;
  assign n12222 = pi0445 & ~n12213;
  assign n12223 = ~n12221 & ~n12222;
  assign n12224 = ~pi0448 & ~n12223;
  assign n12225 = n8128 & ~n12220;
  assign n12226 = ~n12224 & n12225;
  assign n12227 = ~pi0448 & ~n12219;
  assign n12228 = pi0448 & ~n12223;
  assign n12229 = ~n8128 & ~n12227;
  assign n12230 = ~n12228 & n12229;
  assign n12231 = pi1199 & ~n12226;
  assign n12232 = ~n12230 & n12231;
  assign n12233 = n8041 & ~n12191;
  assign n12234 = ~n12232 & n12233;
  assign n12235 = n12186 & ~n12234;
  assign n12236 = pi0591 & ~n12181;
  assign n12237 = pi0590 & ~n12236;
  assign n12238 = ~n7645 & n12181;
  assign n12239 = n7854 & n12238;
  assign n12240 = ~n7757 & n12239;
  assign n12241 = ~n12193 & ~n12240;
  assign n12242 = pi0461 & ~n12241;
  assign n12243 = ~n7862 & n12239;
  assign n12244 = ~n12193 & ~n12243;
  assign n12245 = ~pi0461 & ~n12244;
  assign n12246 = ~n12242 & ~n12245;
  assign n12247 = pi0357 & ~n12246;
  assign n12248 = pi0461 & ~n12244;
  assign n12249 = ~pi0461 & ~n12241;
  assign n12250 = ~n12248 & ~n12249;
  assign n12251 = ~pi0357 & ~n12250;
  assign n12252 = ~n12247 & ~n12251;
  assign n12253 = pi0356 & ~n12252;
  assign n12254 = pi0357 & ~n12250;
  assign n12255 = ~pi0357 & ~n12246;
  assign n12256 = ~n12254 & ~n12255;
  assign n12257 = ~pi0356 & ~n12256;
  assign n12258 = ~n12253 & ~n12257;
  assign n12259 = pi0354 & n12258;
  assign n12260 = pi0356 & ~n12256;
  assign n12261 = ~pi0356 & ~n12252;
  assign n12262 = ~n12260 & ~n12261;
  assign n12263 = ~pi0354 & n12262;
  assign n12264 = ~n7887 & ~n12259;
  assign n12265 = ~n12263 & n12264;
  assign n12266 = pi0354 & n12262;
  assign n12267 = ~pi0354 & n12258;
  assign n12268 = n7887 & ~n12266;
  assign n12269 = ~n12267 & n12268;
  assign n12270 = ~pi0591 & ~n12265;
  assign n12271 = ~n12269 & n12270;
  assign n12272 = n12237 & ~n12271;
  assign n12273 = ~pi1197 & ~n8395;
  assign n12274 = ~n12193 & ~n12273;
  assign n12275 = pi0592 & ~n12181;
  assign n12276 = ~pi1196 & ~n12181;
  assign n12277 = ~n12275 & ~n12276;
  assign n12278 = pi0397 & ~pi0404;
  assign n12279 = ~pi0397 & pi0404;
  assign n12280 = ~n12278 & ~n12279;
  assign n12281 = pi0411 & ~n12280;
  assign n12282 = ~pi0411 & n12280;
  assign n12283 = ~n12281 & ~n12282;
  assign n12284 = ~n7932 & n12283;
  assign n12285 = n7932 & ~n12283;
  assign n12286 = ~n12284 & ~n12285;
  assign n12287 = n7417 & ~n12286;
  assign n12288 = ~n12178 & ~n12287;
  assign n12289 = ~pi0412 & ~n12288;
  assign n12290 = n7417 & n12286;
  assign n12291 = ~n12178 & ~n12290;
  assign n12292 = pi0412 & ~n12291;
  assign n12293 = n7944 & ~n12289;
  assign n12294 = ~n12292 & n12293;
  assign n12295 = pi0412 & ~n12288;
  assign n12296 = ~pi0412 & ~n12291;
  assign n12297 = ~n7944 & ~n12295;
  assign n12298 = ~n12296 & n12297;
  assign n12299 = ~pi0122 & ~n12294;
  assign n12300 = ~n12298 & n12299;
  assign n12301 = ~n12178 & ~n12300;
  assign n12302 = n7626 & ~n12301;
  assign n12303 = pi1091 & n12179;
  assign n12304 = ~n12302 & ~n12303;
  assign n12305 = pi0567 & ~n12304;
  assign n12306 = ~n12180 & ~n12305;
  assign n12307 = n7958 & ~n12306;
  assign n12308 = n12277 & ~n12307;
  assign n12309 = ~pi1199 & ~n12308;
  assign n12310 = ~pi0122 & n7417;
  assign n12311 = ~n12178 & ~n12310;
  assign n12312 = ~n7626 & ~n12303;
  assign n12313 = n7417 & n7926;
  assign n12314 = ~pi0122 & ~n12178;
  assign n12315 = ~n12313 & n12314;
  assign n12316 = ~n12312 & ~n12315;
  assign n12317 = ~n12311 & n12316;
  assign n12318 = pi0567 & n12317;
  assign n12319 = ~n12180 & ~n12318;
  assign n12320 = ~n12305 & n12319;
  assign n12321 = n7958 & ~n12320;
  assign n12322 = n8668 & ~n12319;
  assign n12323 = ~n12275 & ~n12322;
  assign n12324 = ~n12321 & n12323;
  assign n12325 = pi1199 & ~n12324;
  assign n12326 = ~n12309 & ~n12325;
  assign n12327 = n12273 & ~n12326;
  assign n12328 = ~n12274 & ~n12327;
  assign n12329 = pi0333 & ~n12328;
  assign n12330 = n8395 & ~n12193;
  assign n12331 = ~n8395 & ~n12326;
  assign n12332 = ~n12330 & ~n12331;
  assign n12333 = ~pi0333 & ~n12332;
  assign n12334 = ~n12329 & ~n12333;
  assign n12335 = pi0391 & ~n12334;
  assign n12336 = ~pi0333 & ~n12328;
  assign n12337 = pi0333 & ~n12332;
  assign n12338 = ~n12336 & ~n12337;
  assign n12339 = ~pi0391 & ~n12338;
  assign n12340 = pi0392 & n8801;
  assign n12341 = ~pi0392 & ~n8801;
  assign n12342 = ~n12340 & ~n12341;
  assign n12343 = ~n12335 & ~n12342;
  assign n12344 = ~n12339 & n12343;
  assign n12345 = pi0391 & ~n12338;
  assign n12346 = ~pi0391 & ~n12334;
  assign n12347 = n12342 & ~n12345;
  assign n12348 = ~n12346 & n12347;
  assign n12349 = pi0591 & ~n12344;
  assign n12350 = ~n12348 & n12349;
  assign n12351 = ~n7644 & ~n7755;
  assign n12352 = n7422 & ~n7726;
  assign n12353 = ~pi1198 & ~n12352;
  assign n12354 = ~n7970 & ~n12353;
  assign n12355 = ~n12351 & n12354;
  assign n12356 = n12181 & ~n12355;
  assign n12357 = ~pi0591 & ~n12356;
  assign n12358 = ~pi0590 & ~n12357;
  assign n12359 = ~n12350 & n12358;
  assign n12360 = ~pi0588 & ~n12272;
  assign n12361 = ~n12359 & n12360;
  assign n12362 = ~n7425 & ~n12235;
  assign n12363 = ~n12361 & n12362;
  assign n12364 = ~pi0080 & po1038;
  assign n12365 = ~n12184 & n12364;
  assign n12366 = ~n12363 & n12365;
  assign n12367 = pi0567 & n7429;
  assign n12368 = ~n7420 & ~n12179;
  assign n12369 = ~pi0122 & n12368;
  assign n12370 = n7626 & ~n12369;
  assign n12371 = n2625 & ~n12303;
  assign n12372 = ~n12370 & n12371;
  assign n12373 = pi0824 & pi0950;
  assign n12374 = ~pi0110 & n2701;
  assign n12375 = ~pi0088 & n2495;
  assign n12376 = n10379 & n12375;
  assign n12377 = n12374 & n12376;
  assign n12378 = n7440 & n12377;
  assign n12379 = n7446 & n12378;
  assign n12380 = pi0051 & n12379;
  assign n12381 = pi0090 & pi0093;
  assign n12382 = ~pi0841 & ~n2704;
  assign n12383 = ~n12381 & n12382;
  assign n12384 = n2962 & n12383;
  assign n12385 = n12378 & n12384;
  assign n12386 = ~n12380 & ~n12385;
  assign n12387 = n7450 & n12373;
  assign n12388 = ~n12386 & n12387;
  assign n12389 = ~pi0098 & ~n12388;
  assign n12390 = pi1092 & ~n12389;
  assign n12391 = ~pi0087 & n12371;
  assign n12392 = ~n12390 & n12391;
  assign n12393 = n2520 & n12373;
  assign n12394 = n12379 & n12393;
  assign n12395 = ~pi0098 & ~n12394;
  assign n12396 = pi1092 & ~n12395;
  assign n12397 = pi0087 & n12371;
  assign n12398 = ~n12396 & n12397;
  assign n12399 = ~n12392 & ~n12398;
  assign n12400 = pi0122 & ~n12399;
  assign n12401 = ~n12372 & ~n12400;
  assign n12402 = ~pi0075 & ~n12401;
  assign n12403 = ~n7465 & n12368;
  assign n12404 = n12367 & ~n12403;
  assign n12405 = ~n12402 & n12404;
  assign n12406 = ~n7429 & ~n12368;
  assign n12407 = ~n12180 & ~n12406;
  assign n12408 = ~n12405 & n12407;
  assign n12409 = ~pi0592 & ~n12408;
  assign n12410 = ~n12275 & ~n12409;
  assign n12411 = ~n8093 & n12410;
  assign n12412 = n8093 & ~n12276;
  assign n12413 = ~pi0443 & ~n12181;
  assign n12414 = pi0443 & ~n12410;
  assign n12415 = ~n12413 & ~n12414;
  assign n12416 = n8249 & n12415;
  assign n12417 = pi0443 & ~n12181;
  assign n12418 = ~pi0443 & ~n12410;
  assign n12419 = ~n12417 & ~n12418;
  assign n12420 = ~n8249 & n12419;
  assign n12421 = ~n12416 & ~n12420;
  assign n12422 = pi0435 & ~n12421;
  assign n12423 = ~pi0444 & n12419;
  assign n12424 = pi0444 & n12415;
  assign n12425 = ~pi0436 & ~n12423;
  assign n12426 = ~n12424 & n12425;
  assign n12427 = ~pi0444 & n12415;
  assign n12428 = pi0444 & n12419;
  assign n12429 = pi0436 & ~n12427;
  assign n12430 = ~n12428 & n12429;
  assign n12431 = ~n12426 & ~n12430;
  assign n12432 = ~pi0435 & n12431;
  assign n12433 = ~n12422 & ~n12432;
  assign n12434 = ~pi0429 & n12433;
  assign n12435 = ~pi0435 & ~n12421;
  assign n12436 = pi0435 & n12431;
  assign n12437 = ~n12435 & ~n12436;
  assign n12438 = pi0429 & n12437;
  assign n12439 = n8105 & ~n12434;
  assign n12440 = ~n12438 & n12439;
  assign n12441 = ~pi0429 & n12437;
  assign n12442 = pi0429 & n12433;
  assign n12443 = ~n8105 & ~n12441;
  assign n12444 = ~n12442 & n12443;
  assign n12445 = pi1196 & ~n12440;
  assign n12446 = ~n12444 & n12445;
  assign n12447 = n12412 & ~n12446;
  assign n12448 = ~n12411 & ~n12447;
  assign n12449 = ~pi1199 & n12448;
  assign n12450 = pi0428 & ~n12448;
  assign n12451 = ~pi0428 & n12410;
  assign n12452 = ~n12450 & ~n12451;
  assign n12453 = ~pi0427 & ~n12452;
  assign n12454 = ~pi0428 & ~n12448;
  assign n12455 = pi0428 & n12410;
  assign n12456 = ~n12454 & ~n12455;
  assign n12457 = pi0427 & ~n12456;
  assign n12458 = ~n12453 & ~n12457;
  assign n12459 = pi0430 & ~n12458;
  assign n12460 = ~pi0427 & ~n12456;
  assign n12461 = pi0427 & ~n12452;
  assign n12462 = ~n12460 & ~n12461;
  assign n12463 = ~pi0430 & ~n12462;
  assign n12464 = ~n12459 & ~n12463;
  assign n12465 = pi0426 & ~n12464;
  assign n12466 = pi0430 & ~n12462;
  assign n12467 = ~pi0430 & ~n12458;
  assign n12468 = ~n12466 & ~n12467;
  assign n12469 = ~pi0426 & ~n12468;
  assign n12470 = ~n12465 & ~n12469;
  assign n12471 = pi0445 & ~n12470;
  assign n12472 = pi0426 & ~n12468;
  assign n12473 = ~pi0426 & ~n12464;
  assign n12474 = ~n12472 & ~n12473;
  assign n12475 = ~pi0445 & ~n12474;
  assign n12476 = ~n12471 & ~n12475;
  assign n12477 = pi0448 & n12476;
  assign n12478 = pi0445 & ~n12474;
  assign n12479 = ~pi0445 & ~n12470;
  assign n12480 = ~n12478 & ~n12479;
  assign n12481 = ~pi0448 & n12480;
  assign n12482 = ~n8128 & ~n12477;
  assign n12483 = ~n12481 & n12482;
  assign n12484 = ~pi0448 & n12476;
  assign n12485 = pi0448 & n12480;
  assign n12486 = n8128 & ~n12484;
  assign n12487 = ~n12485 & n12486;
  assign n12488 = pi1199 & ~n12483;
  assign n12489 = ~n12487 & n12488;
  assign n12490 = n8041 & ~n12449;
  assign n12491 = ~n12489 & n12490;
  assign n12492 = n12186 & ~n12491;
  assign n12493 = n7850 & n12181;
  assign n12494 = ~n7850 & n12410;
  assign n12495 = ~n12493 & ~n12494;
  assign n12496 = pi1198 & ~n12495;
  assign n12497 = ~pi1198 & ~n12276;
  assign n12498 = n7791 & n12181;
  assign n12499 = ~n7791 & n12410;
  assign n12500 = ~n12498 & ~n12499;
  assign n12501 = ~pi0355 & ~n12500;
  assign n12502 = pi0455 & ~n12181;
  assign n12503 = ~pi0455 & ~n12410;
  assign n12504 = ~n12502 & ~n12503;
  assign n12505 = ~pi0452 & ~n12504;
  assign n12506 = ~pi0455 & ~n12181;
  assign n12507 = pi0455 & ~n12410;
  assign n12508 = ~n12506 & ~n12507;
  assign n12509 = pi0452 & ~n12508;
  assign n12510 = ~n12505 & ~n12509;
  assign n12511 = pi0355 & n12510;
  assign n12512 = ~n12501 & ~n12511;
  assign n12513 = ~pi0458 & n12512;
  assign n12514 = pi0355 & ~n12500;
  assign n12515 = ~pi0355 & n12510;
  assign n12516 = ~n12514 & ~n12515;
  assign n12517 = pi0458 & n12516;
  assign n12518 = n7812 & ~n12513;
  assign n12519 = ~n12517 & n12518;
  assign n12520 = ~pi0458 & n12516;
  assign n12521 = pi0458 & n12512;
  assign n12522 = ~n7812 & ~n12520;
  assign n12523 = ~n12521 & n12522;
  assign n12524 = pi1196 & ~n12519;
  assign n12525 = ~n12523 & n12524;
  assign n12526 = n12497 & ~n12525;
  assign n12527 = ~n12496 & ~n12526;
  assign n12528 = ~n7782 & ~n12527;
  assign n12529 = n7782 & n12410;
  assign n12530 = ~n12528 & ~n12529;
  assign n12531 = ~n7757 & n12530;
  assign n12532 = pi1199 & ~n12410;
  assign n12533 = pi0351 & n12532;
  assign n12534 = ~n12531 & ~n12533;
  assign n12535 = ~pi0461 & ~n12534;
  assign n12536 = ~n7862 & n12530;
  assign n12537 = ~pi0351 & n12532;
  assign n12538 = ~n12536 & ~n12537;
  assign n12539 = pi0461 & ~n12538;
  assign n12540 = ~n12535 & ~n12539;
  assign n12541 = ~pi0357 & ~n12540;
  assign n12542 = ~pi0461 & ~n12538;
  assign n12543 = pi0461 & ~n12534;
  assign n12544 = ~n12542 & ~n12543;
  assign n12545 = pi0357 & ~n12544;
  assign n12546 = ~n12541 & ~n12545;
  assign n12547 = ~pi0356 & ~n12546;
  assign n12548 = ~pi0357 & ~n12544;
  assign n12549 = pi0357 & ~n12540;
  assign n12550 = ~n12548 & ~n12549;
  assign n12551 = pi0356 & ~n12550;
  assign n12552 = ~n12547 & ~n12551;
  assign n12553 = ~pi0354 & ~n12552;
  assign n12554 = ~pi0356 & ~n12550;
  assign n12555 = pi0356 & ~n12546;
  assign n12556 = ~n12554 & ~n12555;
  assign n12557 = pi0354 & ~n12556;
  assign n12558 = ~n7887 & ~n12553;
  assign n12559 = ~n12557 & n12558;
  assign n12560 = ~pi0354 & ~n12556;
  assign n12561 = pi0354 & ~n12552;
  assign n12562 = n7887 & ~n12560;
  assign n12563 = ~n12561 & n12562;
  assign n12564 = ~pi0591 & ~n12559;
  assign n12565 = ~n12563 & n12564;
  assign n12566 = n12237 & ~n12565;
  assign n12567 = ~n12273 & n12410;
  assign n12568 = n7429 & ~n12180;
  assign n12569 = ~n12306 & ~n12568;
  assign n12570 = pi0075 & n12304;
  assign n12571 = ~pi0411 & n12178;
  assign n12572 = n7950 & ~n12571;
  assign n12573 = pi0411 & n12396;
  assign n12574 = n12572 & ~n12573;
  assign n12575 = ~pi0411 & n12396;
  assign n12576 = ~n7950 & ~n12178;
  assign n12577 = ~n7952 & ~n12576;
  assign n12578 = ~n12575 & ~n12577;
  assign n12579 = ~n12574 & ~n12578;
  assign n12580 = pi0122 & n12579;
  assign n12581 = ~n12300 & ~n12580;
  assign n12582 = n7626 & ~n12581;
  assign n12583 = n12397 & ~n12582;
  assign n12584 = pi0411 & n12390;
  assign n12585 = n12572 & ~n12584;
  assign n12586 = ~pi0411 & n12390;
  assign n12587 = ~n12577 & ~n12586;
  assign n12588 = ~n12585 & ~n12587;
  assign n12589 = pi0122 & n12588;
  assign n12590 = ~n12300 & ~n12589;
  assign n12591 = n7626 & ~n12590;
  assign n12592 = n12391 & ~n12591;
  assign n12593 = ~n2625 & n12304;
  assign n12594 = ~n12583 & ~n12593;
  assign n12595 = ~n12592 & n12594;
  assign n12596 = ~pi0075 & ~n12595;
  assign n12597 = n12367 & ~n12570;
  assign n12598 = ~n12596 & n12597;
  assign n12599 = ~n12569 & ~n12598;
  assign n12600 = n7958 & ~n12599;
  assign n12601 = ~n12276 & ~n12600;
  assign n12602 = ~pi1199 & ~n12601;
  assign n12603 = ~n12320 & ~n12568;
  assign n12604 = ~n7465 & ~n12317;
  assign n12605 = ~n12302 & n12604;
  assign n12606 = n2625 & ~n12316;
  assign n12607 = ~n12302 & n12606;
  assign n12608 = ~pi0122 & n12313;
  assign n12609 = n7926 & n12390;
  assign n12610 = ~n7926 & n12178;
  assign n12611 = ~n12609 & ~n12610;
  assign n12612 = n12391 & n12611;
  assign n12613 = ~n7950 & ~n12586;
  assign n12614 = ~n12585 & ~n12613;
  assign n12615 = n12612 & ~n12614;
  assign n12616 = n7926 & n12396;
  assign n12617 = n12397 & ~n12616;
  assign n12618 = ~n12579 & n12617;
  assign n12619 = ~n12615 & ~n12618;
  assign n12620 = ~n12300 & ~n12608;
  assign n12621 = ~n12619 & n12620;
  assign n12622 = ~n12607 & ~n12621;
  assign n12623 = ~pi0075 & ~n12622;
  assign n12624 = n12367 & ~n12605;
  assign n12625 = ~n12623 & n12624;
  assign n12626 = ~n12603 & ~n12625;
  assign n12627 = n7958 & ~n12626;
  assign n12628 = ~n12319 & ~n12568;
  assign n12629 = ~n12610 & ~n12616;
  assign n12630 = n12397 & n12629;
  assign n12631 = ~n12612 & ~n12630;
  assign n12632 = pi0122 & ~n12631;
  assign n12633 = ~n12606 & ~n12632;
  assign n12634 = ~pi0075 & ~n12633;
  assign n12635 = n12367 & ~n12604;
  assign n12636 = ~n12634 & n12635;
  assign n12637 = ~n12628 & ~n12636;
  assign n12638 = n8668 & ~n12637;
  assign n12639 = ~n12627 & ~n12638;
  assign n12640 = pi1199 & ~n12639;
  assign n12641 = ~n12275 & ~n12640;
  assign n12642 = ~n12602 & n12641;
  assign n12643 = n12273 & n12642;
  assign n12644 = ~n12567 & ~n12643;
  assign n12645 = pi0333 & ~n12644;
  assign n12646 = n8395 & ~n12410;
  assign n12647 = ~n8395 & ~n12642;
  assign n12648 = ~n12646 & ~n12647;
  assign n12649 = ~pi0333 & n12648;
  assign n12650 = ~n12645 & ~n12649;
  assign n12651 = pi0391 & ~n12650;
  assign n12652 = pi0333 & ~n12648;
  assign n12653 = ~pi0333 & n12644;
  assign n12654 = ~n12652 & ~n12653;
  assign n12655 = ~pi0391 & n12654;
  assign n12656 = ~n12651 & ~n12655;
  assign n12657 = pi0392 & ~n12656;
  assign n12658 = ~pi0391 & n12650;
  assign n12659 = pi0391 & ~n12654;
  assign n12660 = ~n12658 & ~n12659;
  assign n12661 = ~pi0392 & n12660;
  assign n12662 = ~n12657 & ~n12661;
  assign n12663 = pi0393 & ~n12662;
  assign n12664 = ~pi0392 & ~n12656;
  assign n12665 = pi0392 & n12660;
  assign n12666 = ~n12664 & ~n12665;
  assign n12667 = ~pi0393 & ~n12666;
  assign n12668 = ~n12663 & ~n12667;
  assign n12669 = ~n8028 & ~n12668;
  assign n12670 = pi0393 & ~n12666;
  assign n12671 = ~pi0393 & ~n12662;
  assign n12672 = ~n12670 & ~n12671;
  assign n12673 = n8028 & ~n12672;
  assign n12674 = pi0591 & ~n12669;
  assign n12675 = ~n12673 & n12674;
  assign n12676 = ~pi0592 & ~n12181;
  assign n12677 = pi0592 & ~n12408;
  assign n12678 = ~n12676 & ~n12677;
  assign n12679 = ~n7722 & n12678;
  assign n12680 = n7722 & n12181;
  assign n12681 = ~n12679 & ~n12680;
  assign n12682 = pi1199 & n12681;
  assign n12683 = n7670 & n12678;
  assign n12684 = ~pi1197 & ~n12181;
  assign n12685 = ~n7670 & ~n12684;
  assign n12686 = pi0367 & ~n12181;
  assign n12687 = ~pi0367 & ~n12678;
  assign n12688 = ~n12686 & ~n12687;
  assign n12689 = n7673 & ~n12688;
  assign n12690 = ~pi0367 & ~n12181;
  assign n12691 = pi0367 & ~n12678;
  assign n12692 = ~n12690 & ~n12691;
  assign n12693 = ~n7673 & ~n12692;
  assign n12694 = ~n12689 & ~n12693;
  assign n12695 = n7676 & ~n12694;
  assign n12696 = ~n7673 & n12688;
  assign n12697 = n7673 & n12692;
  assign n12698 = ~n12696 & ~n12697;
  assign n12699 = ~n7676 & n12698;
  assign n12700 = ~n7685 & ~n12695;
  assign n12701 = ~n12699 & n12700;
  assign n12702 = ~n7676 & ~n12694;
  assign n12703 = n7676 & n12698;
  assign n12704 = n7685 & ~n12702;
  assign n12705 = ~n12703 & n12704;
  assign n12706 = pi1197 & ~n12701;
  assign n12707 = ~n12705 & n12706;
  assign n12708 = n12685 & ~n12707;
  assign n12709 = ~pi1199 & ~n12683;
  assign n12710 = ~n12708 & n12709;
  assign n12711 = ~n12682 & ~n12710;
  assign n12712 = ~pi0374 & ~n12711;
  assign n12713 = n8499 & n12681;
  assign n12714 = ~pi1198 & n12710;
  assign n12715 = pi1198 & ~n12678;
  assign n12716 = ~n12713 & ~n12715;
  assign n12717 = ~n12714 & n12716;
  assign n12718 = pi0374 & ~n12717;
  assign n12719 = ~n12712 & ~n12718;
  assign n12720 = pi0369 & ~n12719;
  assign n12721 = ~pi0374 & ~n12717;
  assign n12722 = pi0374 & ~n12711;
  assign n12723 = ~n12721 & ~n12722;
  assign n12724 = ~pi0369 & ~n12723;
  assign n12725 = pi0371 & n8853;
  assign n12726 = ~pi0371 & ~n8853;
  assign n12727 = ~n12725 & ~n12726;
  assign n12728 = pi0370 & ~n12727;
  assign n12729 = ~pi0370 & n12727;
  assign n12730 = ~n12728 & ~n12729;
  assign n12731 = ~n12720 & n12730;
  assign n12732 = ~n12724 & n12731;
  assign n12733 = ~pi0369 & ~n12719;
  assign n12734 = pi0369 & ~n12723;
  assign n12735 = ~n12730 & ~n12733;
  assign n12736 = ~n12734 & n12735;
  assign n12737 = ~pi0591 & ~n12732;
  assign n12738 = ~n12736 & n12737;
  assign n12739 = ~pi0590 & ~n12675;
  assign n12740 = ~n12738 & n12739;
  assign n12741 = ~pi0588 & ~n12740;
  assign n12742 = ~n12566 & n12741;
  assign n12743 = ~n7425 & ~n12742;
  assign n12744 = ~n12492 & n12743;
  assign n12745 = ~n7429 & n12181;
  assign n12746 = pi0075 & n12179;
  assign n12747 = ~n12303 & ~n12396;
  assign n12748 = n8162 & ~n12312;
  assign n12749 = ~n12747 & n12748;
  assign n12750 = ~n12303 & ~n12390;
  assign n12751 = n2610 & ~n12312;
  assign n12752 = ~n12750 & n12751;
  assign n12753 = ~n2625 & n12179;
  assign n12754 = ~n12749 & ~n12753;
  assign n12755 = ~n12752 & n12754;
  assign n12756 = ~pi0075 & ~n12755;
  assign n12757 = ~n12746 & ~n12756;
  assign n12758 = pi0567 & ~n12757;
  assign n12759 = n12568 & ~n12758;
  assign n12760 = ~n12745 & ~n12759;
  assign n12761 = ~pi0592 & n12760;
  assign n12762 = ~n12275 & ~n12761;
  assign n12763 = ~n8093 & n12762;
  assign n12764 = pi0443 & ~n12762;
  assign n12765 = ~n12413 & ~n12764;
  assign n12766 = n8249 & n12765;
  assign n12767 = ~pi0443 & ~n12762;
  assign n12768 = ~n12417 & ~n12767;
  assign n12769 = ~n8249 & n12768;
  assign n12770 = ~n12766 & ~n12769;
  assign n12771 = pi0435 & ~n12770;
  assign n12772 = ~pi0444 & n12768;
  assign n12773 = pi0444 & n12765;
  assign n12774 = ~pi0436 & ~n12772;
  assign n12775 = ~n12773 & n12774;
  assign n12776 = ~pi0444 & n12765;
  assign n12777 = pi0444 & n12768;
  assign n12778 = pi0436 & ~n12776;
  assign n12779 = ~n12777 & n12778;
  assign n12780 = ~n12775 & ~n12779;
  assign n12781 = ~pi0435 & n12780;
  assign n12782 = ~n12771 & ~n12781;
  assign n12783 = ~pi0429 & n12782;
  assign n12784 = ~pi0435 & ~n12770;
  assign n12785 = pi0435 & n12780;
  assign n12786 = ~n12784 & ~n12785;
  assign n12787 = pi0429 & n12786;
  assign n12788 = n8105 & ~n12783;
  assign n12789 = ~n12787 & n12788;
  assign n12790 = ~pi0429 & n12786;
  assign n12791 = pi0429 & n12782;
  assign n12792 = ~n8105 & ~n12790;
  assign n12793 = ~n12791 & n12792;
  assign n12794 = pi1196 & ~n12789;
  assign n12795 = ~n12793 & n12794;
  assign n12796 = n12412 & ~n12795;
  assign n12797 = ~n12763 & ~n12796;
  assign n12798 = ~pi1199 & n12797;
  assign n12799 = ~pi0428 & ~n12797;
  assign n12800 = pi0428 & n12762;
  assign n12801 = ~n12799 & ~n12800;
  assign n12802 = ~pi0427 & ~n12801;
  assign n12803 = pi0428 & ~n12797;
  assign n12804 = ~pi0428 & n12762;
  assign n12805 = ~n12803 & ~n12804;
  assign n12806 = pi0427 & ~n12805;
  assign n12807 = ~n12802 & ~n12806;
  assign n12808 = pi0430 & ~n12807;
  assign n12809 = ~pi0427 & ~n12805;
  assign n12810 = pi0427 & ~n12801;
  assign n12811 = ~n12809 & ~n12810;
  assign n12812 = ~pi0430 & ~n12811;
  assign n12813 = ~n12808 & ~n12812;
  assign n12814 = pi0426 & ~n12813;
  assign n12815 = pi0430 & ~n12811;
  assign n12816 = ~pi0430 & ~n12807;
  assign n12817 = ~n12815 & ~n12816;
  assign n12818 = ~pi0426 & ~n12817;
  assign n12819 = ~n12814 & ~n12818;
  assign n12820 = pi0445 & ~n12819;
  assign n12821 = pi0426 & ~n12817;
  assign n12822 = ~pi0426 & ~n12813;
  assign n12823 = ~n12821 & ~n12822;
  assign n12824 = ~pi0445 & ~n12823;
  assign n12825 = ~n12820 & ~n12824;
  assign n12826 = pi0448 & n12825;
  assign n12827 = pi0445 & ~n12823;
  assign n12828 = ~pi0445 & ~n12819;
  assign n12829 = ~n12827 & ~n12828;
  assign n12830 = ~pi0448 & n12829;
  assign n12831 = n8128 & ~n12826;
  assign n12832 = ~n12830 & n12831;
  assign n12833 = pi0448 & n12829;
  assign n12834 = ~pi0448 & n12825;
  assign n12835 = ~n8128 & ~n12833;
  assign n12836 = ~n12834 & n12835;
  assign n12837 = pi1199 & ~n12832;
  assign n12838 = ~n12836 & n12837;
  assign n12839 = n8041 & ~n12798;
  assign n12840 = ~n12838 & n12839;
  assign n12841 = n12186 & ~n12840;
  assign n12842 = ~n12273 & ~n12762;
  assign n12843 = n8410 & n12568;
  assign n12844 = ~n12181 & ~n12843;
  assign n12845 = n7958 & ~n12745;
  assign n12846 = ~n12303 & ~n12579;
  assign n12847 = n12748 & ~n12846;
  assign n12848 = ~n12303 & ~n12588;
  assign n12849 = n12751 & ~n12848;
  assign n12850 = ~n12753 & ~n12847;
  assign n12851 = ~n12849 & n12850;
  assign n12852 = n7926 & n12749;
  assign n12853 = ~n12611 & n12752;
  assign n12854 = ~n12852 & ~n12853;
  assign n12855 = n12851 & n12854;
  assign n12856 = n12845 & ~n12855;
  assign n12857 = ~n12629 & n12749;
  assign n12858 = ~n12753 & ~n12857;
  assign n12859 = ~n12853 & n12858;
  assign n12860 = n8668 & ~n12745;
  assign n12861 = ~n12859 & n12860;
  assign n12862 = ~n12856 & ~n12861;
  assign n12863 = ~pi0075 & pi0567;
  assign n12864 = ~n12862 & n12863;
  assign n12865 = pi1199 & ~n12844;
  assign n12866 = ~n12864 & n12865;
  assign n12867 = ~pi0075 & ~n12851;
  assign n12868 = ~n12746 & ~n12867;
  assign n12869 = pi0567 & ~n12868;
  assign n12870 = n12568 & ~n12869;
  assign n12871 = n12845 & ~n12870;
  assign n12872 = ~pi1199 & n12277;
  assign n12873 = ~n12871 & n12872;
  assign n12874 = ~n8395 & ~n12866;
  assign n12875 = ~n12873 & n12874;
  assign n12876 = ~pi1197 & n12875;
  assign n12877 = ~n12842 & ~n12876;
  assign n12878 = ~pi0333 & ~n12877;
  assign n12879 = n8395 & ~n12762;
  assign n12880 = ~n12875 & ~n12879;
  assign n12881 = pi0333 & ~n12880;
  assign n12882 = ~n12878 & ~n12881;
  assign n12883 = ~pi0391 & ~n12882;
  assign n12884 = pi0333 & ~n12877;
  assign n12885 = ~pi0333 & ~n12880;
  assign n12886 = ~n12884 & ~n12885;
  assign n12887 = pi0391 & ~n12886;
  assign n12888 = ~n12883 & ~n12887;
  assign n12889 = ~pi0392 & ~n12888;
  assign n12890 = ~pi0391 & ~n12886;
  assign n12891 = pi0391 & ~n12882;
  assign n12892 = ~n12890 & ~n12891;
  assign n12893 = pi0392 & ~n12892;
  assign n12894 = ~n12889 & ~n12893;
  assign n12895 = ~pi0393 & ~n12894;
  assign n12896 = ~pi0392 & ~n12892;
  assign n12897 = pi0392 & ~n12888;
  assign n12898 = ~n12896 & ~n12897;
  assign n12899 = pi0393 & ~n12898;
  assign n12900 = ~n8028 & ~n12895;
  assign n12901 = ~n12899 & n12900;
  assign n12902 = ~pi0393 & ~n12898;
  assign n12903 = pi0393 & ~n12894;
  assign n12904 = n8028 & ~n12902;
  assign n12905 = ~n12903 & n12904;
  assign n12906 = pi0591 & ~n12901;
  assign n12907 = ~n12905 & n12906;
  assign n12908 = pi0592 & n12760;
  assign n12909 = ~n12676 & ~n12908;
  assign n12910 = ~n7722 & n12909;
  assign n12911 = pi1199 & ~n12680;
  assign n12912 = ~n12910 & n12911;
  assign n12913 = n7673 & n7688;
  assign n12914 = ~n7673 & ~n7688;
  assign n12915 = ~n12913 & ~n12914;
  assign n12916 = pi0367 & ~n12915;
  assign n12917 = ~pi0367 & n12915;
  assign n12918 = ~n12916 & ~n12917;
  assign n12919 = n12181 & ~n12918;
  assign n12920 = n12909 & n12918;
  assign n12921 = pi1197 & ~n12919;
  assign n12922 = ~n12920 & n12921;
  assign n12923 = n12685 & ~n12922;
  assign n12924 = n7670 & n12909;
  assign n12925 = ~pi1199 & ~n12924;
  assign n12926 = ~n12923 & n12925;
  assign n12927 = ~n12912 & ~n12926;
  assign n12928 = ~pi0374 & ~n12927;
  assign n12929 = ~pi1198 & ~n12927;
  assign n12930 = pi1198 & ~n12909;
  assign n12931 = ~n12929 & ~n12930;
  assign n12932 = pi0374 & ~n12931;
  assign n12933 = ~n12928 & ~n12932;
  assign n12934 = ~pi0369 & ~n12933;
  assign n12935 = ~pi0374 & ~n12931;
  assign n12936 = pi0374 & ~n12927;
  assign n12937 = ~n12935 & ~n12936;
  assign n12938 = pi0369 & ~n12937;
  assign n12939 = ~n12730 & ~n12934;
  assign n12940 = ~n12938 & n12939;
  assign n12941 = pi0369 & ~n12933;
  assign n12942 = ~pi0369 & ~n12937;
  assign n12943 = n12730 & ~n12941;
  assign n12944 = ~n12942 & n12943;
  assign n12945 = ~pi0591 & ~n12940;
  assign n12946 = ~n12944 & n12945;
  assign n12947 = ~pi0590 & ~n12946;
  assign n12948 = ~n12907 & n12947;
  assign n12949 = ~n7850 & n12762;
  assign n12950 = ~n12493 & ~n12949;
  assign n12951 = pi1198 & ~n12950;
  assign n12952 = ~n7791 & n12762;
  assign n12953 = ~n12498 & ~n12952;
  assign n12954 = pi0355 & ~n12953;
  assign n12955 = ~pi0455 & ~n12762;
  assign n12956 = ~n12502 & ~n12955;
  assign n12957 = ~pi0452 & ~n12956;
  assign n12958 = pi0455 & ~n12762;
  assign n12959 = ~n12506 & ~n12958;
  assign n12960 = pi0452 & ~n12959;
  assign n12961 = ~n12957 & ~n12960;
  assign n12962 = ~pi0355 & n12961;
  assign n12963 = ~n12954 & ~n12962;
  assign n12964 = ~pi0458 & n12963;
  assign n12965 = ~pi0355 & ~n12953;
  assign n12966 = pi0355 & n12961;
  assign n12967 = ~n12965 & ~n12966;
  assign n12968 = pi0458 & n12967;
  assign n12969 = ~n7812 & ~n12964;
  assign n12970 = ~n12968 & n12969;
  assign n12971 = ~pi0458 & n12967;
  assign n12972 = pi0458 & n12963;
  assign n12973 = n7812 & ~n12971;
  assign n12974 = ~n12972 & n12973;
  assign n12975 = pi1196 & ~n12970;
  assign n12976 = ~n12974 & n12975;
  assign n12977 = n12497 & ~n12976;
  assign n12978 = ~n12951 & ~n12977;
  assign n12979 = ~n7782 & ~n12978;
  assign n12980 = n7782 & n12762;
  assign n12981 = ~n12979 & ~n12980;
  assign n12982 = ~n7757 & n12981;
  assign n12983 = pi1199 & ~n12762;
  assign n12984 = pi0351 & n12983;
  assign n12985 = ~n12982 & ~n12984;
  assign n12986 = ~pi0461 & ~n12985;
  assign n12987 = ~n7862 & n12981;
  assign n12988 = ~pi0351 & n12983;
  assign n12989 = ~n12987 & ~n12988;
  assign n12990 = pi0461 & ~n12989;
  assign n12991 = ~n12986 & ~n12990;
  assign n12992 = ~pi0357 & ~n12991;
  assign n12993 = ~pi0461 & ~n12989;
  assign n12994 = pi0461 & ~n12985;
  assign n12995 = ~n12993 & ~n12994;
  assign n12996 = pi0357 & ~n12995;
  assign n12997 = ~n12992 & ~n12996;
  assign n12998 = ~pi0356 & ~n12997;
  assign n12999 = ~pi0357 & ~n12995;
  assign n13000 = pi0357 & ~n12991;
  assign n13001 = ~n12999 & ~n13000;
  assign n13002 = pi0356 & ~n13001;
  assign n13003 = ~n12998 & ~n13002;
  assign n13004 = ~pi0354 & ~n13003;
  assign n13005 = ~pi0356 & ~n13001;
  assign n13006 = pi0356 & ~n12997;
  assign n13007 = ~n13005 & ~n13006;
  assign n13008 = pi0354 & ~n13007;
  assign n13009 = ~n7887 & ~n13004;
  assign n13010 = ~n13008 & n13009;
  assign n13011 = ~pi0354 & ~n13007;
  assign n13012 = pi0354 & ~n13003;
  assign n13013 = n7887 & ~n13011;
  assign n13014 = ~n13012 & n13013;
  assign n13015 = ~pi0591 & ~n13010;
  assign n13016 = ~n13014 & n13015;
  assign n13017 = n12237 & ~n13016;
  assign n13018 = ~pi0588 & ~n12948;
  assign n13019 = ~n13017 & n13018;
  assign n13020 = n7425 & ~n13019;
  assign n13021 = ~n12841 & n13020;
  assign n13022 = ~pi0080 & ~po1038;
  assign n13023 = ~n12744 & n13022;
  assign n13024 = ~n13021 & n13023;
  assign n13025 = ~pi0217 & ~n12366;
  assign n13026 = ~n13024 & n13025;
  assign n13027 = n7643 & ~n12183;
  assign po0238 = ~n13026 & n13027;
  assign n13029 = ~po1038 & n11302;
  assign n13030 = pi0081 & ~pi0314;
  assign n13031 = n2489 & n13030;
  assign n13032 = pi0068 & ~pi0081;
  assign n13033 = n2480 & n13032;
  assign n13034 = n11014 & n13033;
  assign n13035 = n11439 & n13034;
  assign n13036 = n2800 & n13035;
  assign n13037 = ~n13031 & ~n13036;
  assign po0239 = n13029 & ~n13037;
  assign n13039 = pi0069 & pi0314;
  assign n13040 = n2792 & n13039;
  assign n13041 = pi0066 & ~pi0073;
  assign n13042 = n2468 & n13041;
  assign n13043 = n2482 & n13042;
  assign n13044 = ~n13040 & ~n13043;
  assign n13045 = n11103 & n11107;
  assign po0240 = ~n13044 & n13045;
  assign n13047 = n2480 & n2799;
  assign n13048 = pi0084 & n9077;
  assign n13049 = n13047 & n13048;
  assign n13050 = n2467 & n13049;
  assign n13051 = n2499 & n11102;
  assign n13052 = n2702 & n13051;
  assign n13053 = n13050 & n13052;
  assign n13054 = pi0314 & ~n13053;
  assign n13055 = ~pi0083 & ~n13049;
  assign n13056 = n13052 & ~n13055;
  assign n13057 = n2795 & n13056;
  assign n13058 = ~pi0314 & ~n13057;
  assign n13059 = n10166 & ~n13054;
  assign po0241 = ~n13058 & n13059;
  assign n13061 = pi0211 & pi0299;
  assign n13062 = pi0219 & pi0299;
  assign n13063 = ~n13061 & ~n13062;
  assign n13064 = ~n10810 & n13063;
  assign n13065 = ~po1038 & n13064;
  assign po0242 = n11385 & n13065;
  assign n13067 = n6423 & n11104;
  assign n13068 = ~pi0314 & n11105;
  assign n13069 = n11437 & n13068;
  assign n13070 = ~n13067 & ~n13069;
  assign po0243 = n11107 & ~n13070;
  assign n13072 = n7603 & n11396;
  assign n13073 = n7606 & n11399;
  assign n13074 = ~n13072 & ~n13073;
  assign po0244 = n10983 & ~n13074;
  assign n13076 = n2845 & n13051;
  assign n13077 = pi0314 & n10166;
  assign n13078 = n2702 & n13077;
  assign po0245 = n13076 & n13078;
  assign n13080 = n2708 & n7417;
  assign n13081 = ~pi1093 & n2519;
  assign n13082 = n2572 & n13081;
  assign n13083 = n13080 & n13082;
  assign n13084 = n11460 & n13083;
  assign n13085 = n2870 & n13084;
  assign n13086 = ~n7425 & ~n13085;
  assign n13087 = n7417 & n11030;
  assign n13088 = ~pi1093 & ~n13087;
  assign n13089 = n7439 & n12376;
  assign n13090 = n11027 & n13089;
  assign n13091 = n11043 & n12374;
  assign n13092 = n13090 & n13091;
  assign n13093 = pi1093 & ~n13092;
  assign n13094 = n2572 & ~n10074;
  assign n13095 = ~n13093 & n13094;
  assign n13096 = ~n13088 & n13095;
  assign n13097 = n7425 & ~n13096;
  assign n13098 = ~po1038 & ~n13086;
  assign po0246 = ~n13097 & n13098;
  assign n13100 = n2465 & n8921;
  assign n13101 = n8935 & n13100;
  assign n13102 = n10181 & n13101;
  assign n13103 = pi0841 & n7445;
  assign n13104 = n13102 & n13103;
  assign n13105 = ~pi0070 & ~n13104;
  assign n13106 = pi0070 & ~n8959;
  assign n13107 = n2520 & n10165;
  assign n13108 = ~n13105 & n13107;
  assign po0247 = ~n13106 & n13108;
  assign n13110 = ~pi1050 & n9090;
  assign n13111 = ~pi0090 & ~n13110;
  assign n13112 = n11326 & ~n13111;
  assign n13113 = ~n2896 & n13112;
  assign po0248 = ~n7433 & n13113;
  assign n13115 = ~pi0058 & n2756;
  assign n13116 = ~n10158 & ~n13115;
  assign n13117 = n2928 & n10162;
  assign n13118 = ~n13116 & n13117;
  assign n13119 = pi0024 & n2938;
  assign n13120 = ~n2928 & n13119;
  assign n13121 = n11086 & n13120;
  assign n13122 = n2756 & n13121;
  assign n13123 = ~pi0039 & ~n13122;
  assign n13124 = ~n13118 & n13123;
  assign n13125 = n10197 & ~n13124;
  assign po0249 = n7612 & n13125;
  assign n13127 = pi0092 & n2521;
  assign n13128 = n3373 & n11473;
  assign n13129 = n13127 & n13128;
  assign n13130 = n5853 & n6235;
  assign n13131 = n7603 & n13130;
  assign n13132 = n3470 & n6189;
  assign n13133 = n7606 & n13132;
  assign n13134 = ~n13131 & ~n13133;
  assign n13135 = n2534 & n11211;
  assign n13136 = ~n13134 & n13135;
  assign n13137 = ~n13129 & ~n13136;
  assign po0250 = n10163 & ~n13137;
  assign n13139 = pi0093 & n11086;
  assign n13140 = n2914 & n13139;
  assign n13141 = ~pi0092 & ~n13140;
  assign n13142 = ~pi1050 & n2521;
  assign n13143 = pi0092 & ~n13142;
  assign n13144 = n10164 & ~n13141;
  assign po0251 = ~n13143 & n13144;
  assign n13146 = n11068 & n11284;
  assign n13147 = ~n8888 & ~n13146;
  assign n13148 = n2924 & n13146;
  assign n13149 = pi1093 & ~n13148;
  assign n13150 = n2933 & ~n13149;
  assign n13151 = n10243 & n11066;
  assign n13152 = ~n2780 & ~n13151;
  assign n13153 = n2717 & n10162;
  assign n13154 = pi0252 & n13153;
  assign n13155 = ~n13152 & n13154;
  assign n13156 = ~n13150 & ~n13155;
  assign n13157 = ~po0840 & ~n13156;
  assign n13158 = ~n13146 & ~n13157;
  assign n13159 = pi0252 & n13156;
  assign n13160 = ~n13158 & ~n13159;
  assign n13161 = n8888 & ~n13160;
  assign n13162 = n10165 & ~n13147;
  assign po0252 = ~n13161 & n13162;
  assign n13164 = n2517 & n11770;
  assign n13165 = n11458 & n13164;
  assign n13166 = ~pi0332 & n10162;
  assign n13167 = n11283 & n13166;
  assign n13168 = n13102 & n13167;
  assign n13169 = ~pi0039 & ~n13168;
  assign n13170 = ~n13165 & n13169;
  assign n13171 = ~n11422 & n11425;
  assign n13172 = ~n6392 & n13171;
  assign n13173 = ~n6207 & ~n6392;
  assign n13174 = n3471 & ~n11419;
  assign n13175 = n13173 & n13174;
  assign n13176 = pi0039 & ~n13172;
  assign n13177 = ~n13175 & n13176;
  assign n13178 = n10200 & ~n13170;
  assign po0253 = ~n13177 & n13178;
  assign n13180 = n10325 & n13164;
  assign n13181 = pi0479 & ~po0840;
  assign n13182 = n3183 & n13181;
  assign n13183 = pi0096 & n2510;
  assign n13184 = n2961 & n13183;
  assign n13185 = ~n13181 & n13184;
  assign n13186 = n2916 & n13185;
  assign n13187 = ~n13182 & ~n13186;
  assign n13188 = ~pi0095 & ~n13187;
  assign n13189 = ~n13180 & ~n13188;
  assign po0254 = n10165 & ~n13189;
  assign n13191 = pi0039 & pi0593;
  assign n13192 = ~n11427 & n13191;
  assign n13193 = ~n6392 & n13192;
  assign n13194 = n6169 & n13181;
  assign n13195 = ~po0740 & ~n13194;
  assign n13196 = ~pi0096 & n10193;
  assign n13197 = ~n13195 & n13196;
  assign n13198 = n11486 & n13197;
  assign n13199 = ~n13193 & ~n13198;
  assign po0255 = n10200 & ~n13199;
  assign n13201 = ~pi0092 & n11474;
  assign n13202 = ~n13127 & ~n13201;
  assign n13203 = pi0314 & pi1050;
  assign n13204 = n10164 & n13203;
  assign po0256 = ~n13202 & n13204;
  assign n13206 = ~pi0072 & pi0152;
  assign n13207 = n10300 & n13206;
  assign n13208 = pi0299 & n13207;
  assign n13209 = ~pi0072 & pi0174;
  assign n13210 = ~pi0299 & n13209;
  assign n13211 = n10296 & n13210;
  assign n13212 = ~n13208 & ~n13211;
  assign n13213 = pi0232 & ~n13212;
  assign n13214 = pi0039 & ~n13213;
  assign n13215 = ~pi0072 & pi0099;
  assign n13216 = ~pi0039 & ~n13215;
  assign n13217 = ~n13214 & ~n13216;
  assign n13218 = ~n2620 & n13217;
  assign n13219 = ~n7506 & ~n13215;
  assign n13220 = ~n2924 & n13215;
  assign n13221 = n7506 & ~n13220;
  assign n13222 = ~n10329 & n13215;
  assign n13223 = n6266 & n10919;
  assign n13224 = ~n13222 & ~n13223;
  assign n13225 = n10356 & ~n13224;
  assign n13226 = n13221 & ~n13225;
  assign n13227 = ~n13219 & ~n13226;
  assign n13228 = ~pi0039 & ~n13227;
  assign n13229 = n2620 & ~n13214;
  assign n13230 = ~n13228 & n13229;
  assign n13231 = pi0075 & ~n13218;
  assign n13232 = ~n13230 & n13231;
  assign n13233 = pi0228 & n10500;
  assign n13234 = pi0228 & n10344;
  assign n13235 = n13215 & ~n13234;
  assign n13236 = n2531 & ~n13235;
  assign n13237 = ~n13233 & n13236;
  assign n13238 = ~n2531 & ~n13217;
  assign n13239 = pi0087 & ~n13238;
  assign n13240 = ~n13237 & n13239;
  assign n13241 = pi0038 & ~n13217;
  assign n13242 = n10478 & ~n13212;
  assign n13243 = ~n10948 & n13242;
  assign n13244 = pi0041 & pi0072;
  assign n13245 = pi0099 & ~n13244;
  assign n13246 = ~n10411 & n13245;
  assign n13247 = ~pi0228 & ~n10556;
  assign n13248 = ~n13246 & n13247;
  assign n13249 = ~n10459 & n13245;
  assign n13250 = n10779 & ~n13249;
  assign n13251 = ~n10426 & n13245;
  assign n13252 = n10778 & ~n13251;
  assign n13253 = ~n13250 & ~n13252;
  assign n13254 = pi0228 & ~n13253;
  assign n13255 = ~pi0039 & ~n13248;
  assign n13256 = ~n13254 & n13255;
  assign n13257 = n2608 & ~n13243;
  assign n13258 = ~n13256 & n13257;
  assign n13259 = ~n10359 & n13215;
  assign n13260 = n6265 & n10318;
  assign n13261 = ~n13259 & ~n13260;
  assign n13262 = n10356 & ~n13261;
  assign n13263 = n13221 & ~n13262;
  assign n13264 = ~n13219 & ~n13263;
  assign n13265 = ~pi0039 & ~n13264;
  assign n13266 = ~n13214 & ~n13265;
  assign n13267 = n6285 & ~n13266;
  assign n13268 = ~pi0087 & ~n13241;
  assign n13269 = ~n13267 & n13268;
  assign n13270 = ~n13258 & n13269;
  assign n13271 = ~pi0075 & ~n13240;
  assign n13272 = ~n13270 & n13271;
  assign n13273 = ~n13232 & ~n13272;
  assign n13274 = n7429 & ~n13273;
  assign n13275 = ~n7429 & ~n13217;
  assign n13276 = ~po1038 & ~n13275;
  assign n13277 = ~n13274 & n13276;
  assign n13278 = pi0232 & n13207;
  assign n13279 = pi0039 & ~n13278;
  assign n13280 = po1038 & ~n13216;
  assign n13281 = ~n13279 & n13280;
  assign po0257 = n13277 | n13281;
  assign n13283 = ~n6263 & ~n6281;
  assign n13284 = ~n7473 & n10078;
  assign n13285 = pi0129 & ~n13284;
  assign n13286 = n7472 & ~n13285;
  assign n13287 = pi0129 & ~n10078;
  assign n13288 = ~n10081 & ~n13287;
  assign n13289 = ~n13283 & ~n13288;
  assign n13290 = ~n13286 & n13289;
  assign n13291 = ~pi0075 & n2609;
  assign n13292 = n6285 & n13291;
  assign n13293 = ~n13290 & n13292;
  assign n13294 = ~pi0024 & n8967;
  assign n13295 = po0840 & n13294;
  assign n13296 = ~n8964 & n13295;
  assign n13297 = ~n13293 & ~n13296;
  assign n13298 = n8881 & ~n13297;
  assign po0258 = n2521 & n13298;
  assign n13300 = ~pi0039 & ~n10322;
  assign n13301 = pi0152 & n3389;
  assign n13302 = n6197 & n13301;
  assign n13303 = ~pi0072 & n13302;
  assign n13304 = pi0299 & ~n13303;
  assign n13305 = ~pi0144 & pi0174;
  assign n13306 = n10295 & n13305;
  assign n13307 = ~pi0072 & n13306;
  assign n13308 = ~pi0299 & ~n13307;
  assign n13309 = pi0232 & ~n13304;
  assign n13310 = ~n13308 & n13309;
  assign n13311 = pi0039 & ~n13310;
  assign n13312 = ~n13300 & ~n13311;
  assign n13313 = ~n2620 & n13312;
  assign n13314 = ~n7506 & ~n10322;
  assign n13315 = ~n2924 & n10322;
  assign n13316 = n7506 & ~n13315;
  assign n13317 = n2924 & ~n6273;
  assign n13318 = n10322 & ~n10328;
  assign n13319 = ~n10319 & ~n13318;
  assign n13320 = n13317 & ~n13319;
  assign n13321 = n13316 & ~n13320;
  assign n13322 = ~n13314 & ~n13321;
  assign n13323 = ~pi0039 & ~n13322;
  assign n13324 = n2620 & ~n13311;
  assign n13325 = ~n13323 & n13324;
  assign n13326 = pi0075 & ~n13313;
  assign n13327 = ~n13325 & n13326;
  assign n13328 = n10343 & n10931;
  assign n13329 = n10322 & ~n13328;
  assign n13330 = ~pi0101 & n10932;
  assign n13331 = ~pi0039 & ~n13329;
  assign n13332 = ~n13330 & n13331;
  assign n13333 = pi0087 & ~n13311;
  assign n13334 = ~n13332 & n13333;
  assign n13335 = pi0038 & ~n13312;
  assign n13336 = n10949 & n13302;
  assign n13337 = pi0299 & ~n13336;
  assign n13338 = n10949 & n13306;
  assign n13339 = ~pi0299 & ~n13338;
  assign n13340 = n10478 & ~n13337;
  assign n13341 = ~n13339 & n13340;
  assign n13342 = pi0101 & n10409;
  assign n13343 = ~pi0228 & ~n10401;
  assign n13344 = ~n13342 & n13343;
  assign n13345 = pi0101 & n10457;
  assign n13346 = n2924 & ~n10451;
  assign n13347 = ~n13345 & n13346;
  assign n13348 = pi0101 & n10424;
  assign n13349 = ~n2924 & ~n10433;
  assign n13350 = ~n13348 & n13349;
  assign n13351 = ~n13347 & ~n13350;
  assign n13352 = pi0228 & ~n13351;
  assign n13353 = ~pi0039 & ~n13344;
  assign n13354 = ~n13352 & n13353;
  assign n13355 = n2608 & ~n13341;
  assign n13356 = ~n13354 & n13355;
  assign n13357 = ~pi0044 & n10940;
  assign n13358 = n10322 & ~n13357;
  assign n13359 = ~n10318 & ~n13358;
  assign n13360 = n13317 & ~n13359;
  assign n13361 = n13316 & ~n13360;
  assign n13362 = ~n13314 & ~n13361;
  assign n13363 = ~pi0039 & ~n13362;
  assign n13364 = ~n13311 & ~n13363;
  assign n13365 = n6285 & ~n13364;
  assign n13366 = ~pi0087 & ~n13335;
  assign n13367 = ~n13365 & n13366;
  assign n13368 = ~n13356 & n13367;
  assign n13369 = ~pi0075 & ~n13334;
  assign n13370 = ~n13368 & n13369;
  assign n13371 = ~n13327 & ~n13370;
  assign n13372 = n7429 & ~n13371;
  assign n13373 = ~n7429 & ~n13312;
  assign n13374 = ~po1038 & ~n13373;
  assign n13375 = ~n13372 & n13374;
  assign n13376 = pi0232 & n13303;
  assign n13377 = pi0039 & ~n13376;
  assign n13378 = po1038 & ~n13300;
  assign n13379 = ~n13377 & n13378;
  assign po0259 = n13375 | n13379;
  assign n13381 = n2851 & n8922;
  assign po0260 = n13029 & n13381;
  assign n13383 = pi0109 & n2765;
  assign n13384 = n2699 & n13383;
  assign n13385 = pi0314 & ~n13384;
  assign n13386 = ~pi0109 & ~n13076;
  assign n13387 = n6422 & ~n13386;
  assign n13388 = ~pi0314 & ~n13387;
  assign n13389 = n11106 & ~n13385;
  assign po0261 = ~n13388 & n13389;
  assign n13391 = n7425 & ~n8888;
  assign n13392 = n10075 & ~n13391;
  assign n13393 = n10396 & ~n13392;
  assign n13394 = po1057 & ~n13092;
  assign n13395 = ~pi0110 & ~n13090;
  assign n13396 = ~pi0047 & n11043;
  assign n13397 = ~n13395 & n13396;
  assign n13398 = n10378 & n13397;
  assign n13399 = ~po1057 & ~n13398;
  assign n13400 = ~n7474 & ~n10074;
  assign n13401 = ~n13394 & n13400;
  assign n13402 = ~n13399 & n13401;
  assign n13403 = n7474 & ~n10074;
  assign n13404 = n13398 & n13403;
  assign n13405 = ~n13402 & ~n13404;
  assign n13406 = ~n7425 & ~n13405;
  assign n13407 = ~n13393 & ~n13406;
  assign po0262 = n10165 & ~n13407;
  assign n13409 = pi0024 & n11282;
  assign n13410 = ~pi0053 & ~n11281;
  assign n13411 = n2723 & ~n13410;
  assign n13412 = ~pi0024 & n2717;
  assign n13413 = n13411 & n13412;
  assign n13414 = ~n13409 & ~n13413;
  assign n13415 = pi0841 & ~n13414;
  assign n13416 = n8946 & n11267;
  assign n13417 = ~n13415 & ~n13416;
  assign po0264 = n10166 & ~n13417;
  assign n13419 = ~pi0999 & n10166;
  assign po0265 = n11354 & n13419;
  assign n13421 = ~pi0097 & n7442;
  assign n13422 = ~pi0108 & ~n13421;
  assign n13423 = n2701 & ~n13422;
  assign n13424 = n10244 & n13423;
  assign n13425 = ~pi0314 & ~n13424;
  assign n13426 = pi0314 & ~n7444;
  assign n13427 = n7446 & ~n10238;
  assign n13428 = ~n13426 & n13427;
  assign n13429 = ~n13425 & n13428;
  assign n13430 = n7446 & n10238;
  assign n13431 = n13424 & n13430;
  assign n13432 = ~pi0051 & ~n13431;
  assign n13433 = ~n13429 & n13432;
  assign n13434 = n2625 & n7518;
  assign n13435 = ~n13433 & n13434;
  assign n13436 = ~pi0087 & ~n13435;
  assign n13437 = n6133 & n8881;
  assign po0266 = ~n13436 & n13437;
  assign n13439 = n2784 & n11442;
  assign po0267 = n13077 & n13439;
  assign n13441 = ~pi0082 & ~pi0109;
  assign n13442 = pi0111 & n13441;
  assign n13443 = n12374 & n13442;
  assign n13444 = n2499 & n13443;
  assign n13445 = n11105 & n13444;
  assign n13446 = n2801 & n13445;
  assign n13447 = pi0314 & n13446;
  assign n13448 = n8888 & n10075;
  assign n13449 = n10388 & n13448;
  assign n13450 = ~n13447 & ~n13449;
  assign po0268 = n10166 & ~n13450;
  assign n13452 = pi0072 & n10325;
  assign n13453 = ~pi0314 & n13446;
  assign n13454 = n9141 & n13453;
  assign n13455 = ~n13452 & ~n13454;
  assign n13456 = n6479 & n10165;
  assign po0269 = ~n13455 & n13456;
  assign po0270 = ~pi0124 | pi0468;
  assign n13459 = ~pi0072 & pi0113;
  assign n13460 = ~pi0039 & n13459;
  assign n13461 = pi0038 & ~n13460;
  assign n13462 = n2924 & n7506;
  assign n13463 = n7479 & n10531;
  assign n13464 = ~n6272 & ~n13463;
  assign n13465 = n13462 & ~n13464;
  assign n13466 = n13459 & ~n13465;
  assign n13467 = ~n6272 & n13462;
  assign n13468 = ~pi0113 & n13467;
  assign n13469 = n13260 & n13468;
  assign n13470 = ~n13466 & ~n13469;
  assign n13471 = ~pi0039 & ~n13470;
  assign n13472 = n6285 & ~n13471;
  assign n13473 = pi0113 & n10550;
  assign n13474 = ~pi0228 & ~n10557;
  assign n13475 = ~n13473 & n13474;
  assign n13476 = ~pi0113 & n10780;
  assign n13477 = ~n2924 & ~n10426;
  assign n13478 = ~pi0099 & ~n13477;
  assign n13479 = ~n10460 & n13478;
  assign n13480 = pi0113 & ~n10548;
  assign n13481 = ~n13479 & n13480;
  assign n13482 = pi0228 & ~n13476;
  assign n13483 = ~n13481 & n13482;
  assign n13484 = ~pi0039 & ~n13475;
  assign n13485 = ~n13483 & n13484;
  assign n13486 = n2608 & ~n13485;
  assign n13487 = ~n13461 & ~n13472;
  assign n13488 = ~n13486 & n13487;
  assign n13489 = ~pi0087 & ~n13488;
  assign n13490 = ~n2608 & n13460;
  assign n13491 = ~n10532 & n13459;
  assign n13492 = ~pi0113 & n13233;
  assign n13493 = ~n13491 & ~n13492;
  assign n13494 = n2531 & ~n13493;
  assign n13495 = pi0087 & ~n13490;
  assign n13496 = ~n13494 & n13495;
  assign n13497 = ~n13489 & ~n13496;
  assign n13498 = ~pi0075 & ~n13497;
  assign n13499 = n7477 & n13469;
  assign n13500 = ~n6272 & ~n10496;
  assign n13501 = n13462 & ~n13500;
  assign n13502 = n13459 & ~n13501;
  assign n13503 = ~n13499 & ~n13502;
  assign n13504 = n2610 & ~n13503;
  assign n13505 = ~n2620 & n13460;
  assign n13506 = pi0075 & ~n13505;
  assign n13507 = ~n13504 & n13506;
  assign n13508 = ~n13498 & ~n13507;
  assign n13509 = n8881 & ~n13508;
  assign n13510 = ~n8881 & ~n13460;
  assign po0271 = ~n13509 & ~n13510;
  assign n13512 = ~pi0072 & pi0114;
  assign n13513 = ~pi0039 & n13512;
  assign n13514 = ~n2620 & n13513;
  assign n13515 = ~n11143 & ~n13512;
  assign n13516 = pi0114 & n10735;
  assign n13517 = n11143 & ~n13516;
  assign n13518 = ~n10505 & n13517;
  assign n13519 = n2610 & ~n13515;
  assign n13520 = ~n13518 & n13519;
  assign n13521 = pi0075 & ~n13514;
  assign n13522 = ~n13520 & n13521;
  assign n13523 = ~n2608 & ~n13513;
  assign n13524 = pi0228 & n10616;
  assign n13525 = ~pi0115 & n13524;
  assign n13526 = n13512 & ~n13525;
  assign n13527 = n2608 & ~n13526;
  assign n13528 = ~n10537 & n13527;
  assign n13529 = n11212 & ~n13523;
  assign n13530 = ~n13528 & n13529;
  assign n13531 = pi0038 & ~n13513;
  assign n13532 = pi0114 & ~n10618;
  assign n13533 = n11143 & ~n13532;
  assign n13534 = ~n10504 & n13533;
  assign n13535 = ~pi0039 & ~n13515;
  assign n13536 = ~n13534 & n13535;
  assign n13537 = n6285 & ~n13536;
  assign n13538 = ~pi0114 & ~n10783;
  assign n13539 = pi0114 & ~n10791;
  assign n13540 = ~n13538 & ~n13539;
  assign n13541 = ~pi0115 & ~n13540;
  assign n13542 = pi0115 & ~n13512;
  assign n13543 = ~pi0039 & ~n13542;
  assign n13544 = ~n13541 & n13543;
  assign n13545 = n2608 & ~n13544;
  assign n13546 = ~pi0087 & ~n13531;
  assign n13547 = ~n13537 & n13546;
  assign n13548 = ~n13545 & n13547;
  assign n13549 = ~pi0075 & ~n13530;
  assign n13550 = ~n13548 & n13549;
  assign n13551 = ~n13522 & ~n13550;
  assign n13552 = n8881 & ~n13551;
  assign n13553 = ~n8881 & ~n13513;
  assign po0272 = ~n13552 & ~n13553;
  assign n13555 = ~pi0072 & pi0115;
  assign n13556 = ~pi0039 & n13555;
  assign n13557 = ~n2620 & n13556;
  assign n13558 = ~n13462 & ~n13555;
  assign n13559 = pi0115 & n10735;
  assign n13560 = ~pi0052 & n11125;
  assign n13561 = ~pi0115 & ~n13560;
  assign n13562 = n10502 & n13561;
  assign n13563 = n7477 & n13562;
  assign n13564 = n13462 & ~n13559;
  assign n13565 = ~n13563 & n13564;
  assign n13566 = n2610 & ~n13558;
  assign n13567 = ~n13565 & n13566;
  assign n13568 = pi0075 & ~n13557;
  assign n13569 = ~n13567 & n13568;
  assign n13570 = ~n2608 & ~n13556;
  assign n13571 = ~n13524 & n13555;
  assign n13572 = n2608 & ~n13571;
  assign n13573 = ~n10536 & n13572;
  assign n13574 = n11212 & ~n13570;
  assign n13575 = ~n13573 & n13574;
  assign n13576 = pi0038 & ~n13556;
  assign n13577 = pi0115 & ~n10618;
  assign n13578 = n13462 & ~n13577;
  assign n13579 = ~n13562 & n13578;
  assign n13580 = ~pi0039 & ~n13558;
  assign n13581 = ~n13579 & n13580;
  assign n13582 = n6285 & ~n13581;
  assign n13583 = ~pi0115 & ~n10783;
  assign n13584 = pi0115 & ~n10791;
  assign n13585 = ~pi0039 & ~n13583;
  assign n13586 = ~n13584 & n13585;
  assign n13587 = n2608 & ~n13586;
  assign n13588 = ~pi0087 & ~n13576;
  assign n13589 = ~n13582 & n13588;
  assign n13590 = ~n13587 & n13589;
  assign n13591 = ~pi0075 & ~n13575;
  assign n13592 = ~n13590 & n13591;
  assign n13593 = ~n13569 & ~n13592;
  assign n13594 = n8881 & ~n13593;
  assign n13595 = ~n8881 & ~n13556;
  assign po0273 = ~n13594 & ~n13595;
  assign n13597 = ~pi0072 & pi0116;
  assign n13598 = ~pi0039 & n13597;
  assign n13599 = pi0038 & ~n13598;
  assign n13600 = ~pi0113 & n10532;
  assign n13601 = n13597 & ~n13600;
  assign n13602 = ~pi0038 & ~n13601;
  assign n13603 = ~n10535 & n13602;
  assign n13604 = ~n13599 & ~n13603;
  assign n13605 = ~pi0100 & ~n13604;
  assign n13606 = pi0100 & ~n13598;
  assign n13607 = n11212 & ~n13606;
  assign n13608 = ~n13605 & n13607;
  assign n13609 = ~n2924 & n10580;
  assign n13610 = pi0116 & n10585;
  assign n13611 = ~n2924 & ~n13610;
  assign n13612 = n2924 & ~n10568;
  assign n13613 = pi0116 & ~n13612;
  assign n13614 = ~n10573 & ~n13613;
  assign n13615 = ~n13611 & ~n13614;
  assign n13616 = pi0228 & ~n13609;
  assign n13617 = ~n13615 & n13616;
  assign n13618 = pi0116 & n10552;
  assign n13619 = n10777 & ~n13618;
  assign n13620 = ~pi0039 & ~n13619;
  assign n13621 = ~n13617 & n13620;
  assign n13622 = n2608 & ~n13621;
  assign n13623 = ~n13462 & n13597;
  assign n13624 = ~pi0113 & n13463;
  assign n13625 = n13597 & ~n13624;
  assign n13626 = ~n10502 & ~n13625;
  assign n13627 = n13467 & ~n13626;
  assign n13628 = ~n13623 & ~n13627;
  assign n13629 = ~pi0039 & ~n13628;
  assign n13630 = n6285 & ~n13629;
  assign n13631 = ~pi0087 & ~n13599;
  assign n13632 = ~n13630 & n13631;
  assign n13633 = ~n13622 & n13632;
  assign n13634 = ~pi0075 & ~n13608;
  assign n13635 = ~n13633 & n13634;
  assign n13636 = ~n10497 & n13597;
  assign n13637 = ~n10738 & ~n13636;
  assign n13638 = n13467 & ~n13637;
  assign n13639 = ~n13623 & ~n13638;
  assign n13640 = n2610 & ~n13639;
  assign n13641 = ~n2620 & n13598;
  assign n13642 = pi0075 & ~n13641;
  assign n13643 = ~n13640 & n13642;
  assign n13644 = ~n13635 & ~n13643;
  assign n13645 = n8881 & ~n13644;
  assign n13646 = ~n8881 & ~n13598;
  assign po0274 = ~n13645 & ~n13646;
  assign n13648 = n3686 & n7379;
  assign n13649 = ~n3685 & ~n13648;
  assign n13650 = ~pi0038 & ~n13649;
  assign n13651 = ~pi0087 & ~n13650;
  assign n13652 = n6133 & ~n13651;
  assign n13653 = ~pi0092 & ~n13652;
  assign n13654 = ~pi0054 & ~n7305;
  assign n13655 = ~pi0074 & n13654;
  assign n13656 = ~n13653 & n13655;
  assign n13657 = ~pi0055 & ~n13656;
  assign n13658 = ~n7347 & ~n13657;
  assign n13659 = ~pi0056 & ~n13658;
  assign n13660 = ~n6127 & ~n13659;
  assign n13661 = ~pi0062 & ~n13660;
  assign n13662 = ~pi0057 & n6300;
  assign po0275 = ~n13661 & n13662;
  assign n13664 = ~pi0079 & n12169;
  assign n13665 = pi0163 & n6197;
  assign n13666 = ~n11678 & ~n13665;
  assign n13667 = ~pi0150 & ~n13666;
  assign n13668 = pi0150 & n9699;
  assign n13669 = n11676 & n13668;
  assign n13670 = ~n13667 & ~n13669;
  assign n13671 = pi0232 & ~n13670;
  assign n13672 = ~n8989 & n13671;
  assign n13673 = pi0074 & ~n13672;
  assign n13674 = pi0165 & n7473;
  assign n13675 = ~pi0038 & ~pi0054;
  assign n13676 = ~n13674 & ~n13675;
  assign n13677 = n8989 & n13676;
  assign n13678 = ~pi0074 & ~n13672;
  assign n13679 = ~n13677 & n13678;
  assign n13680 = ~n13673 & ~n13679;
  assign n13681 = ~n2529 & ~n13680;
  assign n13682 = n3328 & ~n13681;
  assign n13683 = ~n9883 & ~n13682;
  assign n13684 = pi0055 & ~n13673;
  assign n13685 = pi0150 & n7473;
  assign n13686 = ~pi0092 & n9282;
  assign n13687 = n13685 & n13686;
  assign n13688 = n9248 & n13675;
  assign n13689 = ~n13687 & n13688;
  assign n13690 = ~n13676 & ~n13689;
  assign n13691 = n8989 & ~n13690;
  assign n13692 = n13678 & ~n13691;
  assign n13693 = n13684 & ~n13692;
  assign n13694 = ~pi0184 & ~n11704;
  assign n13695 = pi0185 & ~n13694;
  assign n13696 = ~pi0185 & n13694;
  assign n13697 = n6197 & ~n13695;
  assign n13698 = ~n13696 & n13697;
  assign n13699 = ~pi0299 & ~n13698;
  assign n13700 = pi0299 & n13670;
  assign n13701 = pi0232 & ~n13699;
  assign n13702 = ~n13700 & n13701;
  assign n13703 = ~n8989 & n13702;
  assign n13704 = pi0074 & ~n13703;
  assign n13705 = ~pi0055 & ~n13704;
  assign n13706 = ~pi0143 & ~pi0299;
  assign n13707 = ~pi0165 & pi0299;
  assign n13708 = ~n13706 & ~n13707;
  assign n13709 = n7473 & n13708;
  assign n13710 = n8989 & ~n13709;
  assign n13711 = pi0054 & ~n13710;
  assign n13712 = ~n13703 & n13711;
  assign n13713 = pi0075 & ~n13702;
  assign n13714 = pi0100 & ~n13702;
  assign n13715 = pi0038 & ~n13709;
  assign n13716 = ~pi0100 & ~n13715;
  assign n13717 = ~pi0157 & pi0299;
  assign n13718 = ~pi0178 & ~pi0299;
  assign n13719 = ~n13717 & ~n13718;
  assign n13720 = n7473 & n13719;
  assign n13721 = n9282 & n13720;
  assign n13722 = n9249 & ~n13721;
  assign n13723 = n13716 & ~n13722;
  assign n13724 = ~n13714 & ~n13723;
  assign n13725 = n9205 & ~n13724;
  assign n13726 = ~pi0143 & ~n9187;
  assign n13727 = pi0143 & ~n9189;
  assign n13728 = pi0165 & ~n13727;
  assign n13729 = ~n13726 & n13728;
  assign n13730 = pi0143 & ~pi0165;
  assign n13731 = n9194 & n13730;
  assign n13732 = pi0038 & ~n13731;
  assign n13733 = ~n13729 & n13732;
  assign n13734 = n2568 & ~n13733;
  assign n13735 = ~pi0232 & n9532;
  assign n13736 = ~n6197 & ~n9532;
  assign n13737 = n6197 & ~n9574;
  assign n13738 = ~n13736 & ~n13737;
  assign n13739 = pi0151 & pi0168;
  assign n13740 = ~n13738 & n13739;
  assign n13741 = ~n6197 & n9532;
  assign n13742 = pi0151 & ~pi0168;
  assign n13743 = ~n9606 & n13742;
  assign n13744 = ~pi0168 & n9615;
  assign n13745 = pi0168 & n9612;
  assign n13746 = ~pi0151 & ~n13744;
  assign n13747 = ~n13745 & n13746;
  assign n13748 = ~n13743 & ~n13747;
  assign n13749 = ~n13741 & ~n13748;
  assign n13750 = pi0150 & ~n13740;
  assign n13751 = ~n13749 & n13750;
  assign n13752 = pi0168 & n6197;
  assign n13753 = n9532 & ~n13752;
  assign n13754 = pi0168 & n9506;
  assign n13755 = ~pi0151 & ~n13753;
  assign n13756 = ~n13754 & n13755;
  assign n13757 = ~n9645 & ~n13736;
  assign n13758 = ~pi0168 & n13757;
  assign n13759 = ~n9445 & ~n13736;
  assign n13760 = pi0168 & n13759;
  assign n13761 = pi0151 & ~n13758;
  assign n13762 = ~n13760 & n13761;
  assign n13763 = ~pi0150 & ~n13756;
  assign n13764 = ~n13762 & n13763;
  assign n13765 = pi0299 & ~n13764;
  assign n13766 = ~n13751 & n13765;
  assign n13767 = ~n9506 & ~n13741;
  assign n13768 = ~pi0173 & ~n13767;
  assign n13769 = pi0173 & n13759;
  assign n13770 = ~pi0185 & ~n13768;
  assign n13771 = ~n13769 & n13770;
  assign n13772 = n6197 & ~n9391;
  assign n13773 = pi0173 & ~n13736;
  assign n13774 = ~n13772 & n13773;
  assign n13775 = ~n9496 & ~n13741;
  assign n13776 = ~pi0173 & ~n13775;
  assign n13777 = pi0185 & ~n13774;
  assign n13778 = ~n13776 & n13777;
  assign n13779 = pi0190 & ~n13771;
  assign n13780 = ~n13778 & n13779;
  assign n13781 = ~pi0173 & ~n9527;
  assign n13782 = pi0173 & ~n9949;
  assign n13783 = n6197 & ~n13781;
  assign n13784 = ~n13782 & n13783;
  assign n13785 = pi0185 & ~n13741;
  assign n13786 = ~n13784 & n13785;
  assign n13787 = pi0173 & n13757;
  assign n13788 = ~pi0173 & n9532;
  assign n13789 = ~pi0185 & ~n13788;
  assign n13790 = ~n13787 & n13789;
  assign n13791 = ~pi0190 & ~n13790;
  assign n13792 = ~n13786 & n13791;
  assign n13793 = ~pi0299 & ~n13792;
  assign n13794 = ~n13780 & n13793;
  assign n13795 = pi0232 & ~n13794;
  assign n13796 = ~n13766 & n13795;
  assign n13797 = ~pi0039 & ~n13735;
  assign n13798 = ~n13796 & n13797;
  assign n13799 = pi0168 & n9311;
  assign n13800 = pi0157 & n9324;
  assign n13801 = ~n13799 & ~n13800;
  assign n13802 = n6197 & n11747;
  assign n13803 = ~n13801 & n13802;
  assign n13804 = pi0299 & ~n13803;
  assign n13805 = ~n13718 & ~n13804;
  assign n13806 = n9248 & ~n13805;
  assign n13807 = pi0178 & ~n9338;
  assign n13808 = ~pi0190 & ~n13807;
  assign n13809 = ~pi0299 & ~n13808;
  assign n13810 = ~n13806 & ~n13809;
  assign n13811 = n6205 & ~n9248;
  assign n13812 = n9051 & ~n13811;
  assign n13813 = ~pi0178 & n13812;
  assign n13814 = ~n9314 & n13813;
  assign n13815 = ~pi0299 & ~n9303;
  assign n13816 = pi0178 & n13812;
  assign n13817 = ~n9305 & n13816;
  assign n13818 = pi0190 & n13815;
  assign n13819 = ~n13814 & n13818;
  assign n13820 = ~n13817 & n13819;
  assign n13821 = pi0232 & ~n13820;
  assign n13822 = ~n13810 & n13821;
  assign n13823 = ~pi0232 & n9248;
  assign n13824 = pi0039 & ~n13823;
  assign n13825 = ~n13822 & n13824;
  assign n13826 = ~pi0038 & ~n13825;
  assign n13827 = ~n13798 & n13826;
  assign n13828 = n13734 & ~n13827;
  assign n13829 = n8161 & ~n13715;
  assign n13830 = ~n9249 & n13829;
  assign n13831 = ~n13714 & ~n13830;
  assign n13832 = ~n13828 & n13831;
  assign n13833 = n2569 & ~n13832;
  assign n13834 = ~n13713 & ~n13725;
  assign n13835 = ~n13833 & n13834;
  assign n13836 = ~pi0054 & ~n13835;
  assign n13837 = ~n13712 & ~n13836;
  assign n13838 = ~pi0074 & ~n13837;
  assign n13839 = n13705 & ~n13838;
  assign n13840 = n2529 & ~n13693;
  assign n13841 = ~n13839 & n13840;
  assign n13842 = ~n13683 & ~n13841;
  assign n13843 = n8989 & n13674;
  assign n13844 = ~n8989 & ~n13671;
  assign n13845 = ~n3328 & ~n13843;
  assign n13846 = ~n13844 & n13845;
  assign n13847 = ~n13673 & n13846;
  assign n13848 = ~n13842 & ~n13847;
  assign n13849 = pi0118 & n13848;
  assign n13850 = n8965 & ~n13720;
  assign n13851 = n2521 & n13850;
  assign n13852 = n13716 & ~n13851;
  assign n13853 = ~n13714 & ~n13852;
  assign n13854 = n9205 & ~n13853;
  assign n13855 = n7309 & n9061;
  assign n13856 = ~n6244 & n13130;
  assign n13857 = ~n6392 & n13856;
  assign n13858 = ~pi0232 & ~n13857;
  assign n13859 = ~n13855 & n13858;
  assign n13860 = n6198 & ~n6392;
  assign n13861 = pi0157 & ~n9039;
  assign n13862 = ~pi0157 & n9044;
  assign n13863 = pi0168 & ~n13862;
  assign n13864 = ~pi0157 & ~pi0168;
  assign n13865 = ~n9037 & n13864;
  assign n13866 = ~n13861 & ~n13865;
  assign n13867 = ~n13863 & n13866;
  assign n13868 = ~n13860 & ~n13867;
  assign n13869 = n13130 & ~n13868;
  assign n13870 = ~pi0178 & ~n6205;
  assign n13871 = n9043 & n13870;
  assign n13872 = ~n13860 & ~n13871;
  assign n13873 = pi0190 & ~n13872;
  assign n13874 = pi0178 & ~n9052;
  assign n13875 = ~n13860 & n13874;
  assign n13876 = ~pi0178 & ~n13173;
  assign n13877 = ~pi0190 & ~n13875;
  assign n13878 = ~n13876 & n13877;
  assign n13879 = ~n13873 & ~n13878;
  assign n13880 = n13132 & ~n13879;
  assign n13881 = pi0232 & ~n13880;
  assign n13882 = ~n13869 & n13881;
  assign n13883 = pi0039 & ~n13859;
  assign n13884 = ~n13882 & n13883;
  assign n13885 = ~n6169 & ~n9120;
  assign n13886 = ~pi0232 & ~n9118;
  assign n13887 = ~n13885 & n13886;
  assign n13888 = ~n9118 & ~n11798;
  assign n13889 = ~n6197 & ~n13888;
  assign n13890 = n9142 & n13742;
  assign n13891 = pi0168 & ~n9133;
  assign n13892 = ~pi0168 & ~n9092;
  assign n13893 = ~pi0151 & ~n13891;
  assign n13894 = ~n13892 & n13893;
  assign n13895 = ~n13890 & ~n13894;
  assign n13896 = n9094 & ~n13895;
  assign n13897 = pi0150 & ~n13896;
  assign n13898 = ~pi0151 & n9129;
  assign n13899 = n9166 & ~n13898;
  assign n13900 = n13752 & ~n13899;
  assign n13901 = ~pi0151 & n9118;
  assign n13902 = n9162 & ~n13901;
  assign n13903 = ~pi0168 & ~n13902;
  assign n13904 = ~pi0150 & ~n13900;
  assign n13905 = ~n13903 & n13904;
  assign n13906 = ~n13897 & ~n13905;
  assign n13907 = pi0299 & ~n13889;
  assign n13908 = ~n13906 & n13907;
  assign n13909 = ~n6197 & ~n9122;
  assign n13910 = n6479 & n9142;
  assign n13911 = pi0173 & n13910;
  assign n13912 = ~pi0173 & n6479;
  assign n13913 = n9092 & n13912;
  assign n13914 = ~n13911 & ~n13913;
  assign n13915 = ~pi0190 & n6197;
  assign n13916 = ~n13914 & n13915;
  assign n13917 = ~pi0173 & pi0190;
  assign n13918 = n9134 & n13917;
  assign n13919 = pi0185 & ~n13918;
  assign n13920 = ~n13916 & n13919;
  assign n13921 = pi0173 & n9150;
  assign n13922 = pi0190 & n9131;
  assign n13923 = ~n13921 & n13922;
  assign n13924 = ~pi0173 & n9118;
  assign n13925 = n9147 & ~n13924;
  assign n13926 = ~pi0190 & ~n13925;
  assign n13927 = ~pi0185 & ~n13923;
  assign n13928 = ~n13926 & n13927;
  assign n13929 = ~n13920 & ~n13928;
  assign n13930 = ~pi0299 & ~n13909;
  assign n13931 = ~n13929 & n13930;
  assign n13932 = ~n13908 & ~n13931;
  assign n13933 = pi0232 & ~n13932;
  assign n13934 = ~pi0039 & ~n13887;
  assign n13935 = ~n13933 & n13934;
  assign n13936 = ~n13884 & ~n13935;
  assign n13937 = ~pi0038 & ~n13936;
  assign n13938 = n13734 & ~n13937;
  assign n13939 = ~n13714 & ~n13829;
  assign n13940 = ~n13938 & n13939;
  assign n13941 = n2569 & ~n13940;
  assign n13942 = ~n13713 & ~n13854;
  assign n13943 = ~n13941 & n13942;
  assign n13944 = ~pi0054 & ~n13943;
  assign n13945 = ~n13712 & ~n13944;
  assign n13946 = ~pi0074 & ~n13945;
  assign n13947 = n13705 & ~n13946;
  assign n13948 = pi0054 & n13674;
  assign n13949 = ~pi0092 & n8989;
  assign n13950 = n8965 & n13949;
  assign n13951 = ~n13685 & n13950;
  assign n13952 = ~n13948 & n13951;
  assign n13953 = n2521 & n13952;
  assign n13954 = n13679 & ~n13953;
  assign n13955 = n13684 & ~n13954;
  assign n13956 = n2529 & ~n13955;
  assign n13957 = ~n13947 & n13956;
  assign n13958 = n13682 & ~n13957;
  assign n13959 = ~n13847 & ~n13958;
  assign n13960 = ~pi0118 & n13959;
  assign n13961 = ~n13664 & ~n13960;
  assign n13962 = ~n13849 & n13961;
  assign n13963 = ~pi0118 & ~n8976;
  assign n13964 = n13959 & ~n13963;
  assign n13965 = n13848 & n13963;
  assign n13966 = n13664 & ~n13964;
  assign n13967 = ~n13965 & n13966;
  assign po0276 = n13962 | n13967;
  assign n13969 = pi0128 & pi0228;
  assign n13970 = ~n10163 & n13969;
  assign n13971 = n7384 & n8965;
  assign n13972 = ~n13969 & ~n13971;
  assign n13973 = pi0075 & ~n13972;
  assign n13974 = pi0087 & ~n13969;
  assign n13975 = n2530 & n3335;
  assign n13976 = ~n13969 & ~n13975;
  assign n13977 = pi0100 & ~n13976;
  assign n13978 = ~n2603 & n3470;
  assign n13979 = n7606 & n13978;
  assign n13980 = ~n3448 & n5853;
  assign n13981 = n7603 & n13980;
  assign n13982 = ~n13979 & ~n13981;
  assign n13983 = pi0039 & ~n13982;
  assign n13984 = pi0299 & n6418;
  assign n13985 = ~n6528 & ~n13984;
  assign n13986 = n7473 & ~n13985;
  assign n13987 = pi0109 & ~n13986;
  assign n13988 = ~n2928 & n11668;
  assign n13989 = n2770 & n10157;
  assign n13990 = n11667 & ~n13989;
  assign n13991 = n2783 & ~n13990;
  assign n13992 = ~pi0097 & ~n13991;
  assign n13993 = ~pi0046 & n2928;
  assign n13994 = n2936 & n13993;
  assign n13995 = ~n13992 & n13994;
  assign n13996 = ~n13987 & ~n13988;
  assign n13997 = ~n13995 & n13996;
  assign n13998 = ~n6422 & ~n13986;
  assign n13999 = ~n6491 & n13986;
  assign n14000 = ~n13998 & ~n13999;
  assign n14001 = ~n13997 & n14000;
  assign n14002 = ~pi0091 & ~n14001;
  assign n14003 = n2938 & ~n6419;
  assign n14004 = ~n14002 & n14003;
  assign n14005 = ~n2752 & ~n14004;
  assign n14006 = ~pi0039 & n11086;
  assign n14007 = ~n14005 & n14006;
  assign n14008 = ~n13983 & ~n14007;
  assign n14009 = ~pi0038 & ~n14008;
  assign n14010 = ~pi0228 & n14009;
  assign n14011 = ~n13969 & ~n14010;
  assign n14012 = ~pi0100 & ~n14011;
  assign n14013 = ~pi0087 & ~n13977;
  assign n14014 = ~n14012 & n14013;
  assign n14015 = ~pi0075 & ~n13974;
  assign n14016 = ~n14014 & n14015;
  assign n14017 = ~pi0092 & ~n13973;
  assign n14018 = ~n14016 & n14017;
  assign n14019 = pi0092 & ~n13969;
  assign n14020 = ~n7369 & n14019;
  assign n14021 = n10163 & ~n14020;
  assign n14022 = ~n14018 & n14021;
  assign po0277 = n13970 | n14022;
  assign n14024 = ~pi0031 & ~pi0080;
  assign n14025 = pi0818 & n14024;
  assign n14026 = n7420 & ~n7429;
  assign n14027 = ~n7425 & ~n14026;
  assign n14028 = ~pi0120 & ~n7429;
  assign n14029 = ~pi1093 & n14028;
  assign n14030 = n14027 & ~n14029;
  assign n14031 = pi0120 & ~n7420;
  assign n14032 = ~pi0120 & pi1093;
  assign n14033 = ~pi1091 & n12310;
  assign n14034 = n14032 & ~n14033;
  assign n14035 = ~n14031 & ~n14034;
  assign n14036 = n2521 & n7595;
  assign n14037 = ~n7619 & n14031;
  assign n14038 = n14036 & ~n14037;
  assign n14039 = n7619 & ~n14032;
  assign n14040 = ~n14038 & ~n14039;
  assign n14041 = n2530 & n7506;
  assign n14042 = ~n14040 & n14041;
  assign n14043 = pi0100 & ~n14035;
  assign n14044 = ~n14042 & n14043;
  assign n14045 = pi0038 & n7420;
  assign n14046 = ~pi1093 & n7460;
  assign n14047 = pi0120 & n14046;
  assign n14048 = ~pi0039 & ~n14047;
  assign n14049 = pi0122 & ~n7452;
  assign n14050 = n7534 & ~n10445;
  assign n14051 = n7417 & n7451;
  assign n14052 = ~pi0829 & n14051;
  assign n14053 = ~pi0122 & ~n14052;
  assign n14054 = ~n14050 & n14053;
  assign n14055 = ~n2923 & ~n14049;
  assign n14056 = ~n14054 & n14055;
  assign n14057 = n2930 & ~n14056;
  assign n14058 = n7626 & ~n14051;
  assign n14059 = ~n12310 & n14058;
  assign n14060 = ~n14057 & ~n14059;
  assign n14061 = n14048 & n14060;
  assign n14062 = ~n7570 & n14035;
  assign n14063 = ~n6198 & n14035;
  assign n14064 = ~n7602 & n14031;
  assign n14065 = pi1091 & pi1092;
  assign n14066 = n7554 & n14065;
  assign n14067 = n14034 & ~n14066;
  assign n14068 = ~n14064 & ~n14067;
  assign n14069 = n6198 & n14068;
  assign n14070 = ~n14063 & ~n14069;
  assign n14071 = n6242 & n14070;
  assign n14072 = n6227 & ~n14035;
  assign n14073 = ~n6227 & ~n14068;
  assign n14074 = ~n14072 & ~n14073;
  assign n14075 = ~n6242 & ~n14074;
  assign n14076 = n7570 & ~n14071;
  assign n14077 = ~n14075 & n14076;
  assign n14078 = pi0299 & ~n14062;
  assign n14079 = ~n14077 & n14078;
  assign n14080 = n6205 & n14070;
  assign n14081 = ~n6205 & ~n14074;
  assign n14082 = n7551 & ~n14080;
  assign n14083 = ~n14081 & n14082;
  assign n14084 = ~n7551 & n14035;
  assign n14085 = ~pi0299 & ~n14084;
  assign n14086 = ~n14083 & n14085;
  assign n14087 = pi0039 & ~n14079;
  assign n14088 = ~n14086 & n14087;
  assign n14089 = ~n14061 & ~n14088;
  assign n14090 = ~pi0038 & ~n14089;
  assign n14091 = ~pi0120 & ~pi1093;
  assign n14092 = pi0038 & n14091;
  assign n14093 = ~pi0100 & ~n14092;
  assign n14094 = ~n14045 & n14093;
  assign n14095 = ~n14090 & n14094;
  assign n14096 = ~n14044 & ~n14095;
  assign n14097 = ~pi0087 & ~n14096;
  assign n14098 = n7631 & ~n14091;
  assign n14099 = ~n2625 & n7420;
  assign n14100 = n7626 & ~n12310;
  assign n14101 = ~n7496 & n14100;
  assign n14102 = n7629 & ~n14101;
  assign n14103 = pi0087 & ~n14099;
  assign n14104 = ~n14102 & n14103;
  assign n14105 = n14098 & n14104;
  assign n14106 = ~n14097 & ~n14105;
  assign n14107 = ~pi0075 & ~n14106;
  assign n14108 = n7474 & n14035;
  assign n14109 = ~n7596 & n14034;
  assign n14110 = ~pi1091 & ~n7419;
  assign n14111 = ~n7482 & ~n14110;
  assign n14112 = pi0120 & ~n14111;
  assign n14113 = ~n7474 & ~n14112;
  assign n14114 = ~n14109 & n14113;
  assign n14115 = ~n14108 & ~n14114;
  assign n14116 = n2610 & ~n14115;
  assign n14117 = ~n2610 & n14035;
  assign n14118 = pi0075 & ~n14117;
  assign n14119 = ~n14116 & n14118;
  assign n14120 = n7429 & ~n14119;
  assign n14121 = ~n14107 & n14120;
  assign n14122 = n14030 & ~n14121;
  assign n14123 = n7599 & ~n14091;
  assign n14124 = ~n14057 & ~n14058;
  assign n14125 = n14048 & n14124;
  assign n14126 = pi1093 & ~n6198;
  assign n14127 = n6242 & n14126;
  assign n14128 = n6227 & ~n6242;
  assign n14129 = n7570 & ~n14128;
  assign n14130 = ~n14127 & n14129;
  assign n14131 = n7602 & n14130;
  assign n14132 = pi0299 & ~n14091;
  assign n14133 = ~n14131 & n14132;
  assign n14134 = n6205 & n14126;
  assign n14135 = ~n6205 & n6227;
  assign n14136 = n7551 & ~n14135;
  assign n14137 = ~n14134 & n14136;
  assign n14138 = n7602 & n14137;
  assign n14139 = ~pi0299 & ~n14091;
  assign n14140 = ~n14138 & n14139;
  assign n14141 = pi0039 & ~n14133;
  assign n14142 = ~n14140 & n14141;
  assign n14143 = ~n14125 & ~n14142;
  assign n14144 = ~pi0038 & ~n14143;
  assign n14145 = n14093 & ~n14144;
  assign n14146 = pi0120 & n7619;
  assign n14147 = ~pi0120 & n14036;
  assign n14148 = ~n14146 & ~n14147;
  assign n14149 = n14041 & ~n14148;
  assign n14150 = pi0100 & ~n14091;
  assign n14151 = ~n14149 & n14150;
  assign n14152 = ~n14145 & ~n14151;
  assign n14153 = ~pi0087 & ~n14152;
  assign n14154 = ~n14098 & ~n14153;
  assign n14155 = ~pi0075 & ~n14154;
  assign n14156 = n7429 & ~n14123;
  assign n14157 = ~n14155 & n14156;
  assign n14158 = n7425 & ~n14029;
  assign n14159 = ~n14157 & n14158;
  assign n14160 = ~n14122 & ~n14159;
  assign n14161 = n14025 & ~n14160;
  assign n14162 = ~po1038 & ~n14161;
  assign n14163 = ~n7425 & n14035;
  assign n14164 = pi0120 & ~n14163;
  assign n14165 = n14025 & ~n14091;
  assign n14166 = ~n14163 & n14165;
  assign n14167 = po1038 & ~n14166;
  assign n14168 = ~n14164 & n14167;
  assign n14169 = ~n7643 & ~n14168;
  assign n14170 = pi0951 & pi0982;
  assign n14171 = pi1092 & n14170;
  assign n14172 = pi1093 & n14171;
  assign n14173 = ~pi0120 & ~n14172;
  assign n14174 = ~n14163 & ~n14173;
  assign n14175 = n14167 & ~n14174;
  assign n14176 = n7643 & ~n14175;
  assign n14177 = ~n14169 & ~n14176;
  assign n14178 = ~n14162 & ~n14177;
  assign n14179 = n14028 & ~n14172;
  assign n14180 = ~n2610 & ~n14173;
  assign n14181 = pi0120 & n7597;
  assign n14182 = ~pi1091 & n14172;
  assign n14183 = ~pi0120 & ~n14182;
  assign n14184 = n2930 & n14171;
  assign n14185 = ~pi0093 & ~pi0122;
  assign n14186 = n2506 & n14185;
  assign n14187 = n2925 & n8894;
  assign n14188 = n14186 & n14187;
  assign n14189 = n2962 & n14188;
  assign n14190 = n10324 & n14189;
  assign n14191 = n7478 & n14190;
  assign n14192 = n2703 & n14191;
  assign n14193 = n14184 & ~n14192;
  assign n14194 = n14183 & ~n14193;
  assign n14195 = ~n14181 & ~n14194;
  assign n14196 = ~n7474 & ~n14195;
  assign n14197 = n7474 & n14173;
  assign n14198 = n2610 & ~n14197;
  assign n14199 = ~n14196 & n14198;
  assign n14200 = pi0075 & ~n14180;
  assign n14201 = ~n14199 & n14200;
  assign n14202 = ~n2625 & n14173;
  assign n14203 = pi0087 & ~n14202;
  assign n14204 = pi0950 & n2521;
  assign n14205 = ~n2923 & ~n6213;
  assign n14206 = n14204 & n14205;
  assign n14207 = n14184 & ~n14206;
  assign n14208 = pi0824 & n14204;
  assign n14209 = n14182 & ~n14208;
  assign n14210 = ~n14207 & ~n14209;
  assign n14211 = ~pi0120 & ~n14210;
  assign n14212 = ~n7627 & ~n7628;
  assign n14213 = pi0120 & ~n14212;
  assign n14214 = n2625 & ~n14213;
  assign n14215 = ~n14211 & n14214;
  assign n14216 = n14203 & ~n14215;
  assign n14217 = n7430 & n7478;
  assign n14218 = n14204 & n14217;
  assign n14219 = n14184 & ~n14218;
  assign n14220 = n14183 & ~n14219;
  assign n14221 = ~n14146 & ~n14220;
  assign n14222 = ~pi0039 & n7506;
  assign n14223 = ~n14221 & n14222;
  assign n14224 = pi0100 & ~n14223;
  assign n14225 = ~pi0038 & ~n14224;
  assign n14226 = ~n14041 & n14173;
  assign n14227 = ~n14225 & ~n14226;
  assign n14228 = ~n7551 & n14173;
  assign n14229 = ~pi0299 & ~n14228;
  assign n14230 = ~n8621 & ~n14173;
  assign n14231 = ~n6205 & n14230;
  assign n14232 = ~n8624 & ~n14173;
  assign n14233 = n6205 & n14232;
  assign n14234 = n7551 & ~n14231;
  assign n14235 = ~n14233 & n14234;
  assign n14236 = n14229 & ~n14235;
  assign n14237 = ~n7570 & n14173;
  assign n14238 = pi0299 & ~n14237;
  assign n14239 = ~n6242 & n14230;
  assign n14240 = n6242 & n14232;
  assign n14241 = n7570 & ~n14239;
  assign n14242 = ~n14240 & n14241;
  assign n14243 = n14238 & ~n14242;
  assign n14244 = ~n14236 & ~n14243;
  assign n14245 = pi0039 & ~n14244;
  assign n14246 = n2771 & n7437;
  assign n14247 = n2767 & n14246;
  assign n14248 = n9110 & n14247;
  assign n14249 = n7431 & n14248;
  assign n14250 = n7436 & ~n14249;
  assign n14251 = pi0950 & n7518;
  assign n14252 = ~n14250 & n14251;
  assign n14253 = pi0824 & n14252;
  assign n14254 = n14171 & ~n14253;
  assign n14255 = ~pi0829 & n14254;
  assign n14256 = ~pi0097 & ~n14247;
  assign n14257 = n2935 & ~n14256;
  assign n14258 = n2937 & n14257;
  assign n14259 = ~n7522 & ~n14258;
  assign n14260 = n2461 & ~n14259;
  assign n14261 = n7434 & ~n14260;
  assign n14262 = n7431 & ~n14261;
  assign n14263 = ~pi0051 & ~n14262;
  assign n14264 = ~n2747 & ~n14263;
  assign n14265 = ~pi0096 & ~n14264;
  assign n14266 = ~pi0072 & pi0950;
  assign n14267 = n10416 & n14266;
  assign n14268 = ~n14265 & n14267;
  assign n14269 = n7430 & n14171;
  assign n14270 = ~n14268 & n14269;
  assign n14271 = pi0829 & pi1092;
  assign n14272 = pi0122 & n14170;
  assign n14273 = n14271 & n14272;
  assign n14274 = ~n14252 & n14273;
  assign n14275 = ~n14255 & ~n14274;
  assign n14276 = ~n14270 & n14275;
  assign n14277 = n7517 & ~n14276;
  assign n14278 = n2923 & n14172;
  assign n14279 = ~n14277 & ~n14278;
  assign n14280 = pi1091 & ~n14279;
  assign n14281 = n14182 & ~n14253;
  assign n14282 = ~pi0120 & ~n14281;
  assign n14283 = ~n14280 & n14282;
  assign n14284 = ~n14046 & n14124;
  assign n14285 = pi0120 & n14284;
  assign n14286 = ~pi0039 & ~n14283;
  assign n14287 = ~n14285 & n14286;
  assign n14288 = ~n14245 & ~n14287;
  assign n14289 = n2608 & ~n14288;
  assign n14290 = ~n14227 & ~n14289;
  assign n14291 = ~pi0087 & ~n14290;
  assign n14292 = ~pi0075 & ~n14216;
  assign n14293 = ~n14291 & n14292;
  assign n14294 = ~n14201 & ~n14293;
  assign n14295 = n7429 & ~n14294;
  assign n14296 = n7425 & ~n14295;
  assign n14297 = ~n14035 & ~n14173;
  assign n14298 = ~n2530 & ~n14297;
  assign n14299 = ~n7506 & n14297;
  assign n14300 = ~n12310 & n14182;
  assign n14301 = ~n14219 & ~n14300;
  assign n14302 = ~pi0120 & ~n14301;
  assign n14303 = ~n14037 & ~n14302;
  assign n14304 = n7506 & ~n14303;
  assign n14305 = n2530 & ~n14299;
  assign n14306 = ~n14304 & n14305;
  assign n14307 = pi0100 & ~n14298;
  assign n14308 = ~n14306 & n14307;
  assign n14309 = pi0038 & ~n14297;
  assign n14310 = ~n14046 & n14060;
  assign n14311 = pi0120 & n14310;
  assign n14312 = n14100 & n14254;
  assign n14313 = ~pi0120 & ~n14312;
  assign n14314 = ~n14280 & n14313;
  assign n14315 = ~n14311 & ~n14314;
  assign n14316 = ~pi0039 & ~n14315;
  assign n14317 = ~n7554 & n14184;
  assign n14318 = ~n14300 & ~n14317;
  assign n14319 = ~pi0120 & ~n14318;
  assign n14320 = ~n14064 & ~n14319;
  assign n14321 = n6198 & ~n14320;
  assign n14322 = ~n6198 & n14297;
  assign n14323 = ~n14321 & ~n14322;
  assign n14324 = n6205 & ~n14323;
  assign n14325 = ~n6227 & ~n14320;
  assign n14326 = n6227 & n14297;
  assign n14327 = ~n14325 & ~n14326;
  assign n14328 = ~n6205 & ~n14327;
  assign n14329 = n7551 & ~n14324;
  assign n14330 = ~n14328 & n14329;
  assign n14331 = ~n14084 & n14229;
  assign n14332 = ~n14330 & n14331;
  assign n14333 = n6242 & ~n14323;
  assign n14334 = ~n6242 & ~n14327;
  assign n14335 = n7570 & ~n14333;
  assign n14336 = ~n14334 & n14335;
  assign n14337 = n7420 & ~n7570;
  assign n14338 = n14238 & ~n14337;
  assign n14339 = ~n14336 & n14338;
  assign n14340 = pi0039 & ~n14332;
  assign n14341 = ~n14339 & n14340;
  assign n14342 = ~n14316 & ~n14341;
  assign n14343 = ~pi0038 & ~n14342;
  assign n14344 = ~pi0100 & ~n14309;
  assign n14345 = ~n14343 & n14344;
  assign n14346 = ~n14308 & ~n14345;
  assign n14347 = ~pi0087 & ~n14346;
  assign n14348 = ~n14102 & ~n14214;
  assign n14349 = ~n14207 & ~n14300;
  assign n14350 = n14211 & ~n14349;
  assign n14351 = ~n14348 & ~n14350;
  assign n14352 = ~n14099 & n14203;
  assign n14353 = ~n14351 & n14352;
  assign n14354 = ~n14347 & ~n14353;
  assign n14355 = ~pi0075 & ~n14354;
  assign n14356 = n7474 & ~n14297;
  assign n14357 = ~n14193 & ~n14300;
  assign n14358 = ~pi0120 & ~n14357;
  assign n14359 = n14113 & ~n14358;
  assign n14360 = ~n14356 & ~n14359;
  assign n14361 = n2610 & ~n14360;
  assign n14362 = ~n2610 & ~n14297;
  assign n14363 = pi0075 & ~n14362;
  assign n14364 = ~n14361 & n14363;
  assign n14365 = n7429 & ~n14364;
  assign n14366 = ~n14355 & n14365;
  assign n14367 = n14030 & ~n14366;
  assign n14368 = ~n14296 & ~n14367;
  assign n14369 = n14176 & ~n14179;
  assign n14370 = ~n14368 & n14369;
  assign n14371 = ~n7420 & n7623;
  assign n14372 = ~pi0039 & ~n14310;
  assign n14373 = n7420 & ~n7551;
  assign n14374 = ~n7556 & ~n14110;
  assign n14375 = n6198 & ~n14374;
  assign n14376 = ~n6198 & ~n7420;
  assign n14377 = ~n14375 & ~n14376;
  assign n14378 = n6205 & ~n14377;
  assign n14379 = ~n6227 & ~n14374;
  assign n14380 = n6227 & ~n7420;
  assign n14381 = ~n14379 & ~n14380;
  assign n14382 = ~n6205 & ~n14381;
  assign n14383 = n7551 & ~n14378;
  assign n14384 = ~n14382 & n14383;
  assign n14385 = ~pi0299 & ~n14373;
  assign n14386 = ~n14384 & n14385;
  assign n14387 = n6242 & ~n14377;
  assign n14388 = ~n6242 & ~n14381;
  assign n14389 = n7570 & ~n14387;
  assign n14390 = ~n14388 & n14389;
  assign n14391 = pi0299 & ~n14337;
  assign n14392 = ~n14390 & n14391;
  assign n14393 = ~n14386 & ~n14392;
  assign n14394 = pi0039 & ~n14393;
  assign n14395 = ~pi0038 & ~n14394;
  assign n14396 = ~n14372 & n14395;
  assign n14397 = ~pi0100 & ~n14045;
  assign n14398 = ~n14396 & n14397;
  assign n14399 = ~n14371 & ~n14398;
  assign n14400 = ~pi0087 & ~n14399;
  assign n14401 = ~n14104 & ~n14400;
  assign n14402 = ~pi0075 & ~n14401;
  assign n14403 = n7420 & ~n7475;
  assign n14404 = n7475 & n14111;
  assign n14405 = pi0075 & ~n14403;
  assign n14406 = ~n14404 & n14405;
  assign n14407 = ~n14402 & ~n14406;
  assign n14408 = n14027 & ~n14407;
  assign n14409 = ~n7429 & ~n14163;
  assign n14410 = ~pi0039 & ~n14284;
  assign n14411 = n7612 & ~n14410;
  assign n14412 = ~pi0100 & ~n14411;
  assign n14413 = ~n7623 & ~n14412;
  assign n14414 = ~pi0087 & ~n14413;
  assign n14415 = ~n7631 & ~n14414;
  assign n14416 = ~pi0075 & ~n14415;
  assign n14417 = ~n7599 & ~n14416;
  assign n14418 = n7425 & ~n14028;
  assign n14419 = ~n14417 & n14418;
  assign n14420 = ~n14408 & ~n14409;
  assign n14421 = ~n14419 & n14420;
  assign n14422 = pi0120 & n14169;
  assign n14423 = ~n14421 & n14422;
  assign n14424 = ~n14370 & ~n14423;
  assign n14425 = ~n14025 & ~n14424;
  assign po0278 = n14178 | n14425;
  assign n14427 = ~pi0134 & ~pi0135;
  assign n14428 = ~pi0136 & n14427;
  assign n14429 = ~pi0130 & n14428;
  assign n14430 = ~pi0132 & n14429;
  assign n14431 = ~pi0126 & n14430;
  assign n14432 = ~pi0121 & n14431;
  assign n14433 = ~pi0125 & ~pi0133;
  assign n14434 = pi0121 & ~n14433;
  assign n14435 = ~pi0121 & n14433;
  assign n14436 = ~n14434 & ~n14435;
  assign n14437 = ~n14432 & ~n14436;
  assign n14438 = n2478 & n10152;
  assign n14439 = ~pi0051 & n14438;
  assign n14440 = ~pi0087 & n14439;
  assign n14441 = ~n14437 & n14440;
  assign n14442 = pi0051 & pi0146;
  assign n14443 = pi0051 & n6197;
  assign n14444 = ~pi0146 & n14443;
  assign n14445 = pi0161 & ~n14444;
  assign n14446 = n6197 & ~n14439;
  assign n14447 = ~n14442 & ~n14445;
  assign n14448 = n14446 & n14447;
  assign n14449 = ~pi0087 & ~n14448;
  assign n14450 = pi0087 & ~n13665;
  assign n14451 = pi0232 & ~n14450;
  assign n14452 = ~n14449 & n14451;
  assign n14453 = po1038 & ~n14441;
  assign n14454 = ~n14452 & n14453;
  assign n14455 = ~pi0087 & ~n2570;
  assign n14456 = ~n14439 & n14455;
  assign n14457 = ~pi0142 & n14443;
  assign n14458 = pi0144 & ~n14457;
  assign n14459 = pi0051 & pi0142;
  assign n14460 = n14446 & ~n14459;
  assign n14461 = ~n14458 & n14460;
  assign n14462 = ~pi0299 & ~n14461;
  assign n14463 = pi0299 & ~n14448;
  assign n14464 = pi0232 & ~n14462;
  assign n14465 = ~n14463 & n14464;
  assign n14466 = n14456 & ~n14465;
  assign n14467 = pi0100 & n14439;
  assign n14468 = n2535 & ~n14467;
  assign n14469 = pi0100 & n14465;
  assign n14470 = pi0038 & ~n14465;
  assign n14471 = ~pi0100 & ~n14470;
  assign n14472 = pi0038 & ~n14439;
  assign n14473 = ~pi0100 & ~n14472;
  assign n14474 = ~n14471 & ~n14473;
  assign n14475 = ~pi0161 & ~n14444;
  assign n14476 = n2705 & n7445;
  assign n14477 = ~pi0024 & pi0314;
  assign n14478 = n14476 & n14477;
  assign n14479 = n2467 & n10151;
  assign n14480 = n13047 & n14479;
  assign n14481 = ~pi0050 & pi0077;
  assign n14482 = n2495 & n14481;
  assign n14483 = n14480 & n14482;
  assign n14484 = n8897 & n14478;
  assign n14485 = n14483 & n14484;
  assign n14486 = n2519 & n14485;
  assign n14487 = n2770 & n14480;
  assign n14488 = ~pi0058 & n14476;
  assign n14489 = n9253 & n14488;
  assign n14490 = n14487 & n14489;
  assign n14491 = pi0072 & n6479;
  assign n14492 = n14490 & n14491;
  assign n14493 = n14438 & ~n14476;
  assign n14494 = ~pi0051 & ~n14493;
  assign n14495 = ~pi0024 & n11663;
  assign n14496 = n14487 & n14495;
  assign n14497 = pi0086 & n14487;
  assign n14498 = ~n14483 & ~n14497;
  assign n14499 = n11076 & ~n14498;
  assign n14500 = n14438 & ~n14496;
  assign n14501 = ~n14499 & n14500;
  assign n14502 = n14494 & ~n14501;
  assign n14503 = n2519 & n14502;
  assign n14504 = n14439 & ~n14503;
  assign n14505 = ~n14492 & n14504;
  assign n14506 = ~n14486 & n14505;
  assign n14507 = ~n6197 & ~n14506;
  assign n14508 = pi0072 & n10342;
  assign n14509 = ~n14443 & ~n14508;
  assign n14510 = n6197 & ~n14509;
  assign n14511 = ~n14507 & ~n14510;
  assign n14512 = n14475 & ~n14511;
  assign n14513 = n14439 & ~n14486;
  assign n14514 = ~n14503 & n14513;
  assign n14515 = ~n6197 & ~n14514;
  assign n14516 = ~n14446 & ~n14515;
  assign n14517 = ~n14492 & n14516;
  assign n14518 = pi0146 & n14517;
  assign n14519 = ~pi0051 & n6197;
  assign n14520 = n14438 & ~n14492;
  assign n14521 = n14519 & ~n14520;
  assign n14522 = ~pi0146 & ~n14521;
  assign n14523 = ~n14507 & n14522;
  assign n14524 = pi0161 & ~n14518;
  assign n14525 = ~n14523 & n14524;
  assign n14526 = ~n14512 & ~n14525;
  assign n14527 = n9572 & ~n14526;
  assign n14528 = ~n6197 & n14506;
  assign n14529 = ~pi0051 & n14478;
  assign n14530 = n13439 & n14529;
  assign n14531 = ~pi0072 & ~n14530;
  assign n14532 = n6480 & ~n14531;
  assign n14533 = n6197 & ~n14532;
  assign n14534 = ~n14528 & ~n14533;
  assign n14535 = ~pi0146 & ~n14534;
  assign n14536 = n2519 & n6197;
  assign n14537 = n14530 & n14536;
  assign n14538 = n14511 & ~n14537;
  assign n14539 = pi0146 & n14538;
  assign n14540 = ~pi0161 & ~n14535;
  assign n14541 = ~n14539 & n14540;
  assign n14542 = n14519 & n14520;
  assign n14543 = ~n14486 & n14542;
  assign n14544 = ~n14443 & ~n14543;
  assign n14545 = pi0146 & ~n14439;
  assign n14546 = ~n14544 & ~n14545;
  assign n14547 = pi0161 & ~n14546;
  assign n14548 = ~n14528 & n14547;
  assign n14549 = ~n14541 & ~n14548;
  assign n14550 = n9603 & ~n14549;
  assign n14551 = ~n14527 & ~n14550;
  assign n14552 = pi0156 & ~n14551;
  assign n14553 = pi0144 & ~n14517;
  assign n14554 = ~pi0144 & ~n14511;
  assign n14555 = ~n14553 & ~n14554;
  assign n14556 = ~n14457 & ~n14555;
  assign n14557 = pi0180 & ~n14556;
  assign n14558 = ~pi0142 & ~n14534;
  assign n14559 = pi0142 & n14538;
  assign n14560 = ~pi0144 & ~n14558;
  assign n14561 = ~n14559 & n14560;
  assign n14562 = ~n14486 & n14517;
  assign n14563 = n14458 & ~n14562;
  assign n14564 = ~pi0180 & ~n14563;
  assign n14565 = ~n14561 & n14564;
  assign n14566 = pi0179 & ~n14557;
  assign n14567 = ~n14565 & n14566;
  assign n14568 = n14458 & ~n14506;
  assign n14569 = ~pi0024 & ~n11664;
  assign n14570 = pi0024 & ~n11669;
  assign n14571 = ~n14569 & ~n14570;
  assign n14572 = ~pi0314 & ~n14571;
  assign n14573 = pi0314 & ~n11669;
  assign n14574 = ~n14572 & ~n14573;
  assign n14575 = n7445 & n8960;
  assign n14576 = n14574 & n14575;
  assign n14577 = ~pi0051 & ~n14576;
  assign n14578 = ~n14508 & n14577;
  assign n14579 = n6197 & ~n14578;
  assign n14580 = ~n14507 & ~n14579;
  assign n14581 = pi0142 & n14580;
  assign n14582 = n2708 & n14574;
  assign n14583 = ~pi0072 & ~n14582;
  assign n14584 = n6480 & ~n14583;
  assign n14585 = n6197 & ~n14584;
  assign n14586 = ~n14528 & ~n14585;
  assign n14587 = ~pi0142 & ~n14586;
  assign n14588 = ~pi0144 & ~n14581;
  assign n14589 = ~n14587 & n14588;
  assign n14590 = ~pi0180 & ~n14568;
  assign n14591 = ~n14589 & n14590;
  assign n14592 = ~n14505 & n14519;
  assign n14593 = ~n14507 & ~n14592;
  assign n14594 = n6197 & ~n14504;
  assign n14595 = ~pi0142 & ~n14594;
  assign n14596 = ~pi0051 & ~n14438;
  assign n14597 = n6197 & n14596;
  assign n14598 = ~n14536 & ~n14597;
  assign n14599 = n2519 & ~n14502;
  assign n14600 = ~n14598 & ~n14599;
  assign n14601 = pi0142 & ~n14600;
  assign n14602 = ~n14595 & ~n14601;
  assign n14603 = ~n14516 & ~n14602;
  assign n14604 = n14593 & ~n14603;
  assign n14605 = pi0144 & ~n14604;
  assign n14606 = n2708 & n14571;
  assign n14607 = ~pi0072 & ~n14606;
  assign n14608 = n6480 & ~n14607;
  assign n14609 = n6197 & ~n14608;
  assign n14610 = ~n14528 & ~n14609;
  assign n14611 = ~pi0142 & ~n14610;
  assign n14612 = n14536 & n14606;
  assign n14613 = ~n14510 & ~n14612;
  assign n14614 = ~n14507 & n14613;
  assign n14615 = pi0142 & n14614;
  assign n14616 = ~pi0144 & ~n14615;
  assign n14617 = ~n14611 & n14616;
  assign n14618 = pi0180 & ~n14605;
  assign n14619 = ~n14617 & n14618;
  assign n14620 = ~pi0179 & ~n14619;
  assign n14621 = ~n14591 & n14620;
  assign n14622 = ~n14567 & ~n14621;
  assign n14623 = ~pi0299 & ~n14622;
  assign n14624 = pi0146 & n14614;
  assign n14625 = ~pi0146 & ~n14610;
  assign n14626 = n9572 & ~n14624;
  assign n14627 = ~n14625 & n14626;
  assign n14628 = ~pi0146 & ~n14586;
  assign n14629 = pi0146 & n14580;
  assign n14630 = n9603 & ~n14628;
  assign n14631 = ~n14629 & n14630;
  assign n14632 = ~pi0161 & ~n14627;
  assign n14633 = ~n14631 & n14632;
  assign n14634 = ~pi0146 & ~n14594;
  assign n14635 = pi0146 & ~n14600;
  assign n14636 = ~n14634 & ~n14635;
  assign n14637 = ~n14516 & ~n14636;
  assign n14638 = n14593 & ~n14637;
  assign n14639 = n9572 & ~n14638;
  assign n14640 = n9603 & ~n14444;
  assign n14641 = ~n14506 & n14640;
  assign n14642 = pi0161 & ~n14641;
  assign n14643 = ~n14639 & n14642;
  assign n14644 = ~pi0156 & ~n14643;
  assign n14645 = ~n14633 & n14644;
  assign n14646 = ~n14552 & ~n14645;
  assign n14647 = ~n14623 & n14646;
  assign n14648 = n9159 & ~n14647;
  assign n14649 = n2519 & n14490;
  assign n14650 = ~n6640 & ~n7607;
  assign n14651 = n14649 & ~n14650;
  assign n14652 = ~pi0232 & n14439;
  assign n14653 = ~n14651 & n14652;
  assign n14654 = n14439 & ~n14649;
  assign n14655 = ~pi0051 & ~n14654;
  assign n14656 = ~pi0287 & ~n14655;
  assign n14657 = ~pi0287 & n6197;
  assign n14658 = ~n14597 & ~n14657;
  assign n14659 = ~n14656 & ~n14658;
  assign n14660 = ~n14460 & ~n14659;
  assign n14661 = n9051 & ~n14660;
  assign n14662 = n14438 & n14661;
  assign n14663 = ~n14439 & ~n14457;
  assign n14664 = ~n6405 & ~n14663;
  assign n14665 = pi0144 & ~n14664;
  assign n14666 = pi0051 & ~n6197;
  assign n14667 = ~n14655 & ~n14666;
  assign n14668 = n6405 & ~n14459;
  assign n14669 = n14667 & n14668;
  assign n14670 = n14665 & ~n14669;
  assign n14671 = ~n14662 & n14670;
  assign n14672 = ~n6197 & ~n14654;
  assign n14673 = ~n6222 & ~n14672;
  assign n14674 = ~pi0142 & ~n14673;
  assign n14675 = n2515 & n7450;
  assign n14676 = ~pi0051 & ~n14675;
  assign n14677 = n6197 & ~n14676;
  assign n14678 = ~n14672 & ~n14677;
  assign n14679 = pi0142 & ~n14678;
  assign n14680 = n6405 & ~n14674;
  assign n14681 = ~n14679 & n14680;
  assign n14682 = ~n9051 & ~n14681;
  assign n14683 = ~pi0051 & n14657;
  assign n14684 = ~n14678 & ~n14683;
  assign n14685 = pi0224 & ~n14457;
  assign n14686 = n14684 & n14685;
  assign n14687 = ~n14682 & ~n14686;
  assign n14688 = ~n6405 & n14597;
  assign n14689 = ~n14664 & ~n14688;
  assign n14690 = ~n14665 & n14689;
  assign n14691 = ~n14687 & n14690;
  assign n14692 = pi0181 & ~n14671;
  assign n14693 = ~n14691 & n14692;
  assign n14694 = ~n14681 & n14690;
  assign n14695 = ~pi0181 & ~n14670;
  assign n14696 = ~n14694 & n14695;
  assign n14697 = ~pi0299 & ~n14696;
  assign n14698 = ~n14693 & n14697;
  assign n14699 = ~n14444 & ~n14654;
  assign n14700 = pi0161 & ~n14699;
  assign n14701 = ~pi0146 & ~n14673;
  assign n14702 = pi0146 & ~n14678;
  assign n14703 = ~pi0161 & ~n14701;
  assign n14704 = ~n14702 & n14703;
  assign n14705 = ~n14700 & ~n14704;
  assign n14706 = n6379 & ~n14705;
  assign n14707 = ~n14439 & ~n14448;
  assign n14708 = ~n6379 & ~n14707;
  assign n14709 = n9793 & ~n14708;
  assign n14710 = ~n14706 & n14709;
  assign n14711 = ~n9036 & ~n14706;
  assign n14712 = n14475 & n14684;
  assign n14713 = n14649 & ~n14657;
  assign n14714 = n14439 & ~n14713;
  assign n14715 = n14445 & ~n14714;
  assign n14716 = ~n14712 & ~n14715;
  assign n14717 = pi0216 & ~n14716;
  assign n14718 = ~n14711 & ~n14717;
  assign n14719 = n9794 & ~n14708;
  assign n14720 = ~n14718 & n14719;
  assign n14721 = pi0232 & ~n14710;
  assign n14722 = ~n14698 & n14721;
  assign n14723 = ~n14720 & n14722;
  assign n14724 = pi0039 & ~n14653;
  assign n14725 = ~n14723 & n14724;
  assign n14726 = ~pi0039 & ~pi0232;
  assign n14727 = ~n14506 & n14726;
  assign n14728 = ~n14725 & ~n14727;
  assign n14729 = ~n14648 & n14728;
  assign n14730 = ~pi0038 & ~n14729;
  assign n14731 = ~n14474 & ~n14730;
  assign n14732 = n14468 & ~n14469;
  assign n14733 = ~n14731 & n14732;
  assign n14734 = ~pi0184 & ~pi0299;
  assign n14735 = ~pi0163 & pi0299;
  assign n14736 = ~n14734 & ~n14735;
  assign n14737 = n7473 & n14736;
  assign n14738 = pi0087 & ~n14737;
  assign n14739 = ~n14437 & ~n14738;
  assign n14740 = ~n14466 & n14739;
  assign n14741 = ~n14733 & n14740;
  assign n14742 = n14455 & ~n14465;
  assign n14743 = ~pi0158 & n14463;
  assign n14744 = n14445 & ~n14537;
  assign n14745 = n6197 & ~n14513;
  assign n14746 = ~pi0146 & n14745;
  assign n14747 = n14438 & ~n14485;
  assign n14748 = ~pi0051 & ~n14747;
  assign n14749 = n2519 & ~n14748;
  assign n14750 = ~n14598 & ~n14749;
  assign n14751 = pi0146 & n14750;
  assign n14752 = ~pi0161 & ~n14746;
  assign n14753 = ~n14751 & n14752;
  assign n14754 = ~n14744 & ~n14753;
  assign n14755 = n9572 & ~n14754;
  assign n14756 = pi0232 & ~n14743;
  assign n14757 = ~n14755 & n14756;
  assign n14758 = ~pi0156 & n2530;
  assign n14759 = ~n14757 & n14758;
  assign n14760 = ~pi0159 & n14463;
  assign n14761 = ~pi0181 & n14461;
  assign n14762 = ~pi0144 & ~n14460;
  assign n14763 = ~n14661 & n14762;
  assign n14764 = n9051 & n14657;
  assign n14765 = pi0142 & ~n2521;
  assign n14766 = ~pi0142 & ~n14675;
  assign n14767 = n14764 & ~n14765;
  assign n14768 = ~n14766 & n14767;
  assign n14769 = n14458 & ~n14768;
  assign n14770 = pi0181 & ~n14763;
  assign n14771 = ~n14769 & n14770;
  assign n14772 = ~pi0299 & ~n14761;
  assign n14773 = ~n14771 & n14772;
  assign n14774 = ~n9036 & n14448;
  assign n14775 = n14475 & ~n14659;
  assign n14776 = n6197 & n6380;
  assign n14777 = n14445 & ~n14776;
  assign n14778 = n9036 & ~n14775;
  assign n14779 = ~n14777 & n14778;
  assign n14780 = n9794 & ~n14774;
  assign n14781 = ~n14779 & n14780;
  assign n14782 = n10478 & ~n14760;
  assign n14783 = ~n14781 & n14782;
  assign n14784 = ~n14773 & n14783;
  assign n14785 = n6197 & ~n14577;
  assign n14786 = ~n14442 & n14785;
  assign n14787 = pi0161 & ~n14786;
  assign n14788 = n6197 & ~n14514;
  assign n14789 = ~pi0146 & n14788;
  assign n14790 = n14476 & n14747;
  assign n14791 = n14501 & n14790;
  assign n14792 = n14494 & ~n14791;
  assign n14793 = n2519 & ~n14792;
  assign n14794 = ~n14598 & ~n14793;
  assign n14795 = pi0146 & n14794;
  assign n14796 = ~pi0161 & ~n14789;
  assign n14797 = ~n14795 & n14796;
  assign n14798 = ~n14787 & ~n14797;
  assign n14799 = n9572 & ~n14798;
  assign n14800 = n14445 & ~n14612;
  assign n14801 = ~pi0161 & ~n14636;
  assign n14802 = ~n14800 & ~n14801;
  assign n14803 = n9603 & ~n14802;
  assign n14804 = pi0232 & ~n14803;
  assign n14805 = ~n14799 & n14804;
  assign n14806 = pi0156 & ~n14805;
  assign n14807 = ~pi0142 & n14788;
  assign n14808 = pi0142 & n14794;
  assign n14809 = ~pi0144 & ~n14807;
  assign n14810 = ~n14808 & n14809;
  assign n14811 = ~n14459 & n14785;
  assign n14812 = pi0144 & ~n14811;
  assign n14813 = pi0180 & ~n14810;
  assign n14814 = ~n14812 & n14813;
  assign n14815 = n14458 & ~n14612;
  assign n14816 = ~pi0144 & ~n14602;
  assign n14817 = ~pi0180 & ~n14816;
  assign n14818 = ~n14815 & n14817;
  assign n14819 = pi0179 & ~n14818;
  assign n14820 = ~n14814 & n14819;
  assign n14821 = ~pi0180 & n14461;
  assign n14822 = ~pi0142 & n14745;
  assign n14823 = pi0142 & n14750;
  assign n14824 = ~pi0144 & ~n14822;
  assign n14825 = ~n14823 & n14824;
  assign n14826 = n14458 & ~n14537;
  assign n14827 = pi0180 & ~n14825;
  assign n14828 = ~n14826 & n14827;
  assign n14829 = ~pi0179 & ~n14821;
  assign n14830 = ~n14828 & n14829;
  assign n14831 = ~n14820 & ~n14830;
  assign n14832 = ~pi0299 & ~n14831;
  assign n14833 = ~pi0039 & ~n14806;
  assign n14834 = ~n14832 & n14833;
  assign n14835 = ~pi0038 & ~n14784;
  assign n14836 = ~n14834 & n14835;
  assign n14837 = n14471 & ~n14759;
  assign n14838 = ~n14836 & n14837;
  assign n14839 = n2535 & ~n14469;
  assign n14840 = ~n14838 & n14839;
  assign n14841 = n14437 & ~n14738;
  assign n14842 = ~n14742 & n14841;
  assign n14843 = ~n14840 & n14842;
  assign n14844 = ~po1038 & ~n14843;
  assign n14845 = ~n14741 & n14844;
  assign po0279 = n14454 | n14845;
  assign n14847 = n7420 & n7427;
  assign n14848 = n7429 & n14407;
  assign n14849 = n14027 & ~n14848;
  assign n14850 = n7429 & n14417;
  assign n14851 = n7425 & ~n14850;
  assign n14852 = ~po1038 & ~n14849;
  assign n14853 = ~n14851 & n14852;
  assign po0280 = n14847 | n14853;
  assign n14855 = pi0110 & n10075;
  assign n14856 = ~n10976 & n14855;
  assign n14857 = po1057 & n14856;
  assign n14858 = ~pi0039 & ~n14857;
  assign n14859 = ~pi0110 & n9293;
  assign n14860 = ~n6244 & n6379;
  assign n14861 = n14859 & n14860;
  assign n14862 = pi0039 & ~n14861;
  assign n14863 = po1038 & ~n14858;
  assign n14864 = ~n14862 & n14863;
  assign n14865 = pi0110 & n13448;
  assign n14866 = ~pi0039 & ~n14865;
  assign n14867 = ~n6207 & n7607;
  assign n14868 = n14859 & n14867;
  assign n14869 = pi0299 & n14861;
  assign n14870 = pi0039 & ~n14868;
  assign n14871 = ~n14869 & n14870;
  assign n14872 = ~n14866 & ~n14871;
  assign n14873 = ~pi0038 & n2571;
  assign n14874 = ~n14872 & ~n14873;
  assign n14875 = pi0090 & ~n10387;
  assign n14876 = ~pi0111 & ~n6429;
  assign n14877 = ~pi0036 & n2809;
  assign n14878 = ~n14876 & n14877;
  assign n14879 = n2468 & ~n14878;
  assign n14880 = ~n2793 & ~n2798;
  assign n14881 = ~n14879 & n14880;
  assign n14882 = ~pi0083 & ~n14881;
  assign n14883 = n2795 & ~n14882;
  assign n14884 = ~pi0071 & ~n14883;
  assign n14885 = n6438 & ~n14884;
  assign n14886 = ~pi0081 & ~n14885;
  assign n14887 = n11443 & ~n14886;
  assign n14888 = ~pi0090 & ~n14887;
  assign n14889 = n2707 & ~n14888;
  assign n14890 = n9073 & ~n14875;
  assign n14891 = n14889 & n14890;
  assign n14892 = pi0072 & n2708;
  assign n14893 = n10387 & n14892;
  assign n14894 = ~n14891 & ~n14893;
  assign n14895 = n6479 & ~n14894;
  assign n14896 = ~pi0110 & ~n14895;
  assign n14897 = n13448 & ~n14896;
  assign n14898 = n2897 & n14889;
  assign n14899 = ~pi0072 & ~n14898;
  assign n14900 = n6480 & ~n13448;
  assign n14901 = ~n14899 & n14900;
  assign n14902 = ~pi0039 & ~n14901;
  assign n14903 = ~n14897 & n14902;
  assign n14904 = ~n14871 & ~n14903;
  assign n14905 = n14873 & ~n14904;
  assign n14906 = ~po1038 & ~n14874;
  assign n14907 = ~n14905 & n14906;
  assign po0281 = ~n14864 & ~n14907;
  assign n14909 = ~pi0125 & n14432;
  assign n14910 = pi0125 & pi0133;
  assign n14911 = ~n14433 & ~n14910;
  assign n14912 = ~n14909 & ~n14911;
  assign n14913 = n14439 & ~n14912;
  assign n14914 = pi0172 & n14443;
  assign n14915 = ~pi0152 & n14597;
  assign n14916 = ~n14914 & ~n14915;
  assign n14917 = pi0232 & ~n14916;
  assign n14918 = ~n14913 & ~n14917;
  assign n14919 = ~pi0087 & ~n14918;
  assign n14920 = pi0087 & n7473;
  assign n14921 = pi0162 & n14920;
  assign n14922 = po1038 & ~n14921;
  assign n14923 = ~n14919 & n14922;
  assign n14924 = pi0193 & n14443;
  assign n14925 = ~pi0174 & n14597;
  assign n14926 = ~pi0299 & ~n14924;
  assign n14927 = ~n14925 & n14926;
  assign n14928 = pi0299 & n14916;
  assign n14929 = pi0232 & ~n14927;
  assign n14930 = ~n14928 & n14929;
  assign n14931 = n14455 & ~n14930;
  assign n14932 = pi0140 & ~pi0299;
  assign n14933 = pi0162 & pi0299;
  assign n14934 = ~n14932 & ~n14933;
  assign n14935 = n7473 & ~n14934;
  assign n14936 = pi0087 & ~n14935;
  assign n14937 = pi0100 & n14930;
  assign n14938 = ~pi0232 & ~n14508;
  assign n14939 = ~pi0039 & ~n14938;
  assign n14940 = ~pi0299 & ~n7551;
  assign n14941 = pi0299 & ~n7570;
  assign n14942 = ~n14940 & ~n14941;
  assign n14943 = n2521 & n14942;
  assign n14944 = ~pi0232 & ~n14943;
  assign n14945 = pi0039 & ~n14944;
  assign n14946 = ~n7570 & n14916;
  assign n14947 = n2521 & ~n6197;
  assign n14948 = n6197 & ~n14654;
  assign n14949 = ~n14947 & ~n14948;
  assign n14950 = ~pi0152 & ~n14949;
  assign n14951 = ~n14677 & ~n14947;
  assign n14952 = pi0152 & ~n14951;
  assign n14953 = ~n14950 & ~n14952;
  assign n14954 = pi0051 & ~pi0172;
  assign n14955 = ~n14953 & ~n14954;
  assign n14956 = ~pi0216 & ~n14955;
  assign n14957 = n6379 & n14956;
  assign n14958 = ~n14946 & ~n14957;
  assign n14959 = n9603 & ~n14958;
  assign n14960 = ~n6379 & ~n14916;
  assign n14961 = n14649 & n14657;
  assign n14962 = ~n14446 & ~n14961;
  assign n14963 = ~pi0152 & n14962;
  assign n14964 = n14657 & n14675;
  assign n14965 = ~n14443 & ~n14964;
  assign n14966 = pi0152 & n14965;
  assign n14967 = pi0172 & ~n14963;
  assign n14968 = ~n14966 & n14967;
  assign n14969 = ~pi0152 & ~n14659;
  assign n14970 = pi0152 & ~n14776;
  assign n14971 = ~pi0172 & ~n14969;
  assign n14972 = ~n14970 & n14971;
  assign n14973 = pi0216 & ~n14968;
  assign n14974 = ~n14972 & n14973;
  assign n14975 = n6379 & ~n14974;
  assign n14976 = ~n14956 & n14975;
  assign n14977 = n9572 & ~n14960;
  assign n14978 = ~n14976 & n14977;
  assign n14979 = ~n7551 & ~n14446;
  assign n14980 = n6197 & n14655;
  assign n14981 = ~n14947 & ~n14980;
  assign n14982 = ~n14979 & ~n14981;
  assign n14983 = ~pi0174 & n14982;
  assign n14984 = n2521 & n7551;
  assign n14985 = pi0174 & n14984;
  assign n14986 = ~n14924 & ~n14985;
  assign n14987 = ~n14983 & n14986;
  assign n14988 = ~pi0180 & ~n14987;
  assign n14989 = n7551 & n14949;
  assign n14990 = pi0224 & ~n14961;
  assign n14991 = n6405 & ~n14990;
  assign n14992 = ~n14446 & ~n14991;
  assign n14993 = ~n14989 & ~n14992;
  assign n14994 = ~pi0174 & n14993;
  assign n14995 = pi0224 & n14965;
  assign n14996 = n6405 & ~n14995;
  assign n14997 = n7551 & n14951;
  assign n14998 = n14996 & ~n14997;
  assign n14999 = ~n14443 & ~n14998;
  assign n15000 = pi0174 & ~n14999;
  assign n15001 = pi0193 & ~n14994;
  assign n15002 = ~n15000 & n15001;
  assign n15003 = ~n7551 & ~n14764;
  assign n15004 = n2521 & ~n15003;
  assign n15005 = pi0174 & n15004;
  assign n15006 = pi0224 & ~n14659;
  assign n15007 = ~pi0224 & n14981;
  assign n15008 = n6405 & ~n15006;
  assign n15009 = ~n15007 & n15008;
  assign n15010 = ~n14688 & ~n15009;
  assign n15011 = ~pi0174 & ~n15010;
  assign n15012 = ~pi0193 & ~n15005;
  assign n15013 = ~n15011 & n15012;
  assign n15014 = pi0180 & ~n15013;
  assign n15015 = ~n15002 & n15014;
  assign n15016 = ~pi0299 & ~n14988;
  assign n15017 = ~n15015 & n15016;
  assign n15018 = ~n14959 & ~n14978;
  assign n15019 = ~n15017 & n15018;
  assign n15020 = pi0232 & ~n15019;
  assign n15021 = n14945 & ~n15020;
  assign n15022 = ~pi0038 & ~n14939;
  assign n15023 = ~n15021 & n15022;
  assign n15024 = pi0038 & ~n14930;
  assign n15025 = ~pi0100 & ~n15024;
  assign n15026 = ~pi0152 & n14521;
  assign n15027 = ~pi0152 & n6197;
  assign n15028 = n14508 & ~n15027;
  assign n15029 = ~pi0197 & ~n15026;
  assign n15030 = ~n15028 & n15029;
  assign n15031 = ~n6197 & n14508;
  assign n15032 = ~n14519 & ~n15031;
  assign n15033 = ~n14543 & ~n15032;
  assign n15034 = ~pi0152 & pi0197;
  assign n15035 = ~n15033 & n15034;
  assign n15036 = ~n15030 & ~n15035;
  assign n15037 = ~n14914 & ~n15036;
  assign n15038 = ~n6197 & ~n14508;
  assign n15039 = ~n14533 & ~n15038;
  assign n15040 = ~pi0172 & n15039;
  assign n15041 = ~n14443 & ~n14537;
  assign n15042 = ~n14508 & n15041;
  assign n15043 = pi0172 & ~n15042;
  assign n15044 = pi0152 & pi0197;
  assign n15045 = ~n15043 & n15044;
  assign n15046 = ~n15040 & n15045;
  assign n15047 = ~n15037 & ~n15046;
  assign n15048 = n9766 & ~n15047;
  assign n15049 = n14505 & n14542;
  assign n15050 = ~n15038 & ~n15049;
  assign n15051 = ~pi0152 & n15050;
  assign n15052 = n14509 & ~n14612;
  assign n15053 = pi0152 & ~n15052;
  assign n15054 = pi0172 & ~n15051;
  assign n15055 = ~n15053 & n15054;
  assign n15056 = ~n14609 & ~n15038;
  assign n15057 = pi0152 & n15056;
  assign n15058 = ~n14592 & ~n15031;
  assign n15059 = ~pi0152 & ~n15058;
  assign n15060 = ~pi0172 & ~n15059;
  assign n15061 = ~n15057 & n15060;
  assign n15062 = ~pi0197 & ~n15055;
  assign n15063 = ~n15061 & n15062;
  assign n15064 = ~n14585 & ~n15038;
  assign n15065 = ~pi0172 & n15064;
  assign n15066 = ~n14578 & ~n15038;
  assign n15067 = pi0172 & n15066;
  assign n15068 = pi0152 & ~n15067;
  assign n15069 = ~n15065 & n15068;
  assign n15070 = n6197 & n14506;
  assign n15071 = ~n15032 & ~n15070;
  assign n15072 = ~pi0152 & ~n14914;
  assign n15073 = ~n15071 & n15072;
  assign n15074 = pi0197 & ~n15073;
  assign n15075 = ~n15069 & n15074;
  assign n15076 = n9760 & ~n15063;
  assign n15077 = ~n15075 & n15076;
  assign n15078 = ~n15048 & ~n15077;
  assign n15079 = pi0299 & ~n15078;
  assign n15080 = ~pi0145 & n14508;
  assign n15081 = pi0145 & n15039;
  assign n15082 = pi0174 & ~n15080;
  assign n15083 = ~n15081 & n15082;
  assign n15084 = ~n14521 & ~n15031;
  assign n15085 = ~pi0145 & ~n15084;
  assign n15086 = pi0145 & n15033;
  assign n15087 = ~pi0174 & ~n15085;
  assign n15088 = ~n15086 & n15087;
  assign n15089 = ~n15083 & ~n15088;
  assign n15090 = ~pi0193 & ~n15089;
  assign n15091 = ~pi0145 & n14537;
  assign n15092 = ~n15041 & ~n15091;
  assign n15093 = ~n14508 & ~n15092;
  assign n15094 = pi0174 & ~n15093;
  assign n15095 = ~n14443 & ~n14486;
  assign n15096 = pi0145 & ~n15095;
  assign n15097 = n14542 & ~n15096;
  assign n15098 = ~pi0174 & ~n15097;
  assign n15099 = ~n15038 & n15098;
  assign n15100 = pi0193 & ~n15099;
  assign n15101 = ~n15094 & n15100;
  assign n15102 = ~n15090 & ~n15101;
  assign n15103 = n9772 & ~n15102;
  assign n15104 = pi0193 & n15050;
  assign n15105 = ~pi0193 & ~n15058;
  assign n15106 = ~pi0145 & ~n15104;
  assign n15107 = ~n15105 & n15106;
  assign n15108 = pi0145 & ~n14924;
  assign n15109 = ~n15071 & n15108;
  assign n15110 = ~pi0174 & ~n15109;
  assign n15111 = ~n15107 & n15110;
  assign n15112 = pi0145 & n15066;
  assign n15113 = ~pi0145 & ~n15052;
  assign n15114 = pi0193 & ~n15113;
  assign n15115 = ~n15112 & n15114;
  assign n15116 = ~pi0145 & n15056;
  assign n15117 = pi0145 & n15064;
  assign n15118 = ~pi0193 & ~n15116;
  assign n15119 = ~n15117 & n15118;
  assign n15120 = pi0174 & ~n15115;
  assign n15121 = ~n15119 & n15120;
  assign n15122 = n9776 & ~n15111;
  assign n15123 = ~n15121 & n15122;
  assign n15124 = ~n15103 & ~n15123;
  assign n15125 = ~pi0038 & ~n15124;
  assign n15126 = ~n15079 & ~n15125;
  assign n15127 = n9159 & ~n15126;
  assign n15128 = ~n15023 & n15025;
  assign n15129 = ~n15127 & n15128;
  assign n15130 = n2535 & ~n14937;
  assign n15131 = ~n15129 & n15130;
  assign n15132 = n14912 & ~n14936;
  assign n15133 = ~n14931 & n15132;
  assign n15134 = ~n15131 & n15133;
  assign n15135 = n14456 & ~n14930;
  assign n15136 = ~n14473 & ~n15025;
  assign n15137 = ~n14515 & ~n14612;
  assign n15138 = pi0145 & n15137;
  assign n15139 = n14536 & n14582;
  assign n15140 = ~n14515 & ~n15139;
  assign n15141 = ~pi0145 & n15140;
  assign n15142 = ~pi0174 & ~n15138;
  assign n15143 = ~n15141 & n15142;
  assign n15144 = ~n14515 & ~n14794;
  assign n15145 = ~pi0145 & ~n14513;
  assign n15146 = ~n6197 & ~n14513;
  assign n15147 = ~n14446 & ~n15146;
  assign n15148 = ~n14503 & n15147;
  assign n15149 = ~n15145 & n15148;
  assign n15150 = n2519 & n15149;
  assign n15151 = pi0174 & ~n15144;
  assign n15152 = ~n15150 & n15151;
  assign n15153 = pi0193 & ~n15152;
  assign n15154 = ~n15143 & n15153;
  assign n15155 = pi0174 & ~n15149;
  assign n15156 = ~pi0051 & n15138;
  assign n15157 = ~pi0145 & ~n14515;
  assign n15158 = ~n14785 & n15157;
  assign n15159 = ~pi0174 & ~n15156;
  assign n15160 = ~n15158 & n15159;
  assign n15161 = ~pi0193 & ~n15155;
  assign n15162 = ~n15160 & n15161;
  assign n15163 = n9772 & ~n15154;
  assign n15164 = ~n15162 & n15163;
  assign n15165 = pi0145 & ~n14597;
  assign n15166 = ~pi0174 & ~n15091;
  assign n15167 = ~pi0145 & pi0174;
  assign n15168 = ~n14750 & n15167;
  assign n15169 = ~n15165 & ~n15168;
  assign n15170 = ~n15166 & n15169;
  assign n15171 = pi0193 & ~n14515;
  assign n15172 = ~n15170 & n15171;
  assign n15173 = ~n14443 & ~n14515;
  assign n15174 = pi0145 & n14438;
  assign n15175 = ~n15166 & ~n15174;
  assign n15176 = n15173 & ~n15175;
  assign n15177 = ~n14515 & ~n14745;
  assign n15178 = pi0174 & n15177;
  assign n15179 = ~n15176 & ~n15178;
  assign n15180 = ~pi0193 & ~n15179;
  assign n15181 = n9776 & ~n15172;
  assign n15182 = ~n15180 & n15181;
  assign n15183 = ~n15164 & ~n15182;
  assign n15184 = ~pi0038 & ~n15183;
  assign n15185 = ~pi0172 & n14443;
  assign n15186 = ~pi0172 & n15148;
  assign n15187 = ~n14515 & ~n14600;
  assign n15188 = pi0172 & n15187;
  assign n15189 = pi0152 & ~n15186;
  assign n15190 = ~n15188 & n15189;
  assign n15191 = ~pi0152 & ~n15137;
  assign n15192 = pi0197 & ~n15185;
  assign n15193 = ~n15190 & n15192;
  assign n15194 = ~n15191 & n15193;
  assign n15195 = ~pi0152 & ~n15140;
  assign n15196 = pi0152 & ~n15144;
  assign n15197 = pi0172 & ~n15196;
  assign n15198 = ~n15195 & n15197;
  assign n15199 = ~pi0152 & n14785;
  assign n15200 = ~n14514 & ~n15027;
  assign n15201 = ~pi0172 & ~n15200;
  assign n15202 = ~n15199 & n15201;
  assign n15203 = ~n15198 & ~n15202;
  assign n15204 = ~pi0197 & ~n15203;
  assign n15205 = pi0299 & n9766;
  assign n15206 = ~n15194 & n15205;
  assign n15207 = ~n15204 & n15206;
  assign n15208 = pi0152 & n14597;
  assign n15209 = ~n14515 & ~n15208;
  assign n15210 = pi0172 & ~n15209;
  assign n15211 = ~pi0172 & ~n14915;
  assign n15212 = ~n14516 & n15211;
  assign n15213 = pi0197 & ~n15210;
  assign n15214 = ~n15212 & n15213;
  assign n15215 = pi0152 & n15177;
  assign n15216 = ~n14515 & ~n14537;
  assign n15217 = ~pi0152 & n15216;
  assign n15218 = ~n14443 & n15217;
  assign n15219 = ~pi0172 & ~n15215;
  assign n15220 = ~n15218 & n15219;
  assign n15221 = ~n14515 & ~n14750;
  assign n15222 = pi0152 & n15221;
  assign n15223 = pi0172 & ~n15222;
  assign n15224 = ~n15217 & n15223;
  assign n15225 = ~pi0197 & ~n15224;
  assign n15226 = ~n15220 & n15225;
  assign n15227 = pi0299 & n9760;
  assign n15228 = ~n15214 & n15227;
  assign n15229 = ~n15226 & n15228;
  assign n15230 = ~n15207 & ~n15229;
  assign n15231 = ~n15184 & n15230;
  assign n15232 = n9159 & ~n15231;
  assign n15233 = ~n14439 & n14916;
  assign n15234 = ~n9036 & ~n15233;
  assign n15235 = ~n14654 & ~n15027;
  assign n15236 = ~pi0152 & n14677;
  assign n15237 = ~n15235 & ~n15236;
  assign n15238 = ~pi0172 & ~n15237;
  assign n15239 = ~pi0152 & n14673;
  assign n15240 = pi0152 & n14667;
  assign n15241 = pi0172 & ~n15240;
  assign n15242 = ~n15239 & n15241;
  assign n15243 = n9036 & ~n15238;
  assign n15244 = ~n15242 & n15243;
  assign n15245 = n9603 & ~n15244;
  assign n15246 = pi0152 & ~n14914;
  assign n15247 = ~n14714 & n15246;
  assign n15248 = n14684 & n15072;
  assign n15249 = n9036 & ~n15247;
  assign n15250 = ~n15248 & n15249;
  assign n15251 = n9572 & ~n15250;
  assign n15252 = ~n15245 & ~n15251;
  assign n15253 = ~n15234 & ~n15252;
  assign n15254 = pi0180 & n14714;
  assign n15255 = n9051 & n14649;
  assign n15256 = n14439 & ~n15255;
  assign n15257 = pi0174 & ~n15256;
  assign n15258 = ~n15254 & n15257;
  assign n15259 = n9051 & n14678;
  assign n15260 = ~n6197 & ~n14438;
  assign n15261 = ~n9051 & ~n15260;
  assign n15262 = ~pi0051 & n15261;
  assign n15263 = ~n15259 & ~n15262;
  assign n15264 = pi0180 & n14683;
  assign n15265 = ~pi0174 & ~n15264;
  assign n15266 = n15263 & n15265;
  assign n15267 = ~pi0193 & ~n15258;
  assign n15268 = ~n15266 & n15267;
  assign n15269 = ~n14666 & n15261;
  assign n15270 = n9051 & n14673;
  assign n15271 = ~n15269 & ~n15270;
  assign n15272 = ~pi0174 & ~n15271;
  assign n15273 = ~n14443 & ~n15256;
  assign n15274 = pi0174 & ~n15273;
  assign n15275 = ~pi0180 & ~n15274;
  assign n15276 = ~n15272 & n15275;
  assign n15277 = n9051 & ~n14672;
  assign n15278 = ~n10603 & n15277;
  assign n15279 = ~n15269 & ~n15278;
  assign n15280 = ~pi0174 & ~n15279;
  assign n15281 = ~pi0051 & ~n14714;
  assign n15282 = n6197 & ~n15281;
  assign n15283 = ~n15256 & ~n15282;
  assign n15284 = pi0174 & ~n15283;
  assign n15285 = pi0180 & ~n15284;
  assign n15286 = ~n15280 & n15285;
  assign n15287 = pi0193 & ~n15286;
  assign n15288 = ~n15276 & n15287;
  assign n15289 = ~pi0299 & ~n15268;
  assign n15290 = ~n15288 & n15289;
  assign n15291 = ~n15253 & ~n15290;
  assign n15292 = pi0232 & ~n15291;
  assign n15293 = ~pi0299 & ~n15256;
  assign n15294 = n9036 & n14649;
  assign n15295 = n14439 & ~n15294;
  assign n15296 = pi0299 & ~n15295;
  assign n15297 = ~n15293 & ~n15296;
  assign n15298 = ~pi0232 & ~n15297;
  assign n15299 = pi0039 & ~n15298;
  assign n15300 = ~n15292 & n15299;
  assign n15301 = ~pi0232 & ~n14514;
  assign n15302 = ~pi0039 & ~n15301;
  assign n15303 = ~pi0038 & ~n15302;
  assign n15304 = ~n15300 & n15303;
  assign n15305 = ~n15136 & ~n15304;
  assign n15306 = ~n15232 & n15305;
  assign n15307 = n14468 & ~n14937;
  assign n15308 = ~n15306 & n15307;
  assign n15309 = ~n14912 & ~n14936;
  assign n15310 = ~n15135 & n15309;
  assign n15311 = ~n15308 & n15310;
  assign n15312 = ~po1038 & ~n15311;
  assign n15313 = ~n15134 & n15312;
  assign po0282 = n14923 | n15313;
  assign n15315 = pi0175 & n14443;
  assign n15316 = ~pi0189 & n14597;
  assign n15317 = ~pi0299 & ~n15315;
  assign n15318 = ~n15316 & n15317;
  assign n15319 = ~pi0051 & ~n14597;
  assign n15320 = ~n10299 & ~n14438;
  assign n15321 = ~pi0051 & ~n15320;
  assign n15322 = pi0153 & n14443;
  assign n15323 = ~n15321 & ~n15322;
  assign n15324 = ~n15319 & ~n15323;
  assign n15325 = pi0299 & ~n15324;
  assign n15326 = pi0232 & ~n15318;
  assign n15327 = ~n15325 & n15326;
  assign n15328 = ~n2608 & n15327;
  assign n15329 = ~pi0126 & n14435;
  assign n15330 = pi0126 & ~n14435;
  assign n15331 = ~n15329 & ~n15330;
  assign n15332 = ~n14431 & ~n15331;
  assign n15333 = ~n2608 & n14439;
  assign n15334 = ~n15332 & n15333;
  assign n15335 = pi0182 & n14714;
  assign n15336 = pi0189 & ~n15256;
  assign n15337 = ~n15335 & n15336;
  assign n15338 = pi0182 & n14683;
  assign n15339 = ~pi0189 & ~n15338;
  assign n15340 = n15263 & n15339;
  assign n15341 = ~n15337 & ~n15340;
  assign n15342 = n11765 & ~n15341;
  assign n15343 = ~pi0189 & ~n15271;
  assign n15344 = pi0189 & ~n15273;
  assign n15345 = ~pi0182 & ~n15344;
  assign n15346 = ~n15343 & n15345;
  assign n15347 = ~pi0189 & ~n15279;
  assign n15348 = pi0189 & ~n15283;
  assign n15349 = pi0182 & ~n15348;
  assign n15350 = ~n15347 & n15349;
  assign n15351 = ~n15346 & ~n15350;
  assign n15352 = n11833 & ~n15351;
  assign n15353 = ~n9036 & ~n15323;
  assign n15354 = ~pi0166 & n14684;
  assign n15355 = pi0166 & ~n14714;
  assign n15356 = ~n15354 & ~n15355;
  assign n15357 = pi0160 & ~n15322;
  assign n15358 = ~n15356 & n15357;
  assign n15359 = ~n10299 & ~n14654;
  assign n15360 = ~pi0166 & n14677;
  assign n15361 = ~n15359 & ~n15360;
  assign n15362 = ~pi0153 & ~n15361;
  assign n15363 = ~pi0166 & n14673;
  assign n15364 = pi0166 & n14667;
  assign n15365 = pi0153 & ~n15364;
  assign n15366 = ~n15363 & n15365;
  assign n15367 = ~n15362 & ~n15366;
  assign n15368 = ~pi0160 & ~n15367;
  assign n15369 = n9036 & ~n15358;
  assign n15370 = ~n15368 & n15369;
  assign n15371 = pi0299 & ~n15353;
  assign n15372 = ~n15370 & n15371;
  assign n15373 = ~n15342 & ~n15352;
  assign n15374 = ~n15372 & n15373;
  assign n15375 = pi0232 & ~n15374;
  assign n15376 = n15299 & ~n15375;
  assign n15377 = ~pi0189 & n15173;
  assign n15378 = pi0178 & ~n15377;
  assign n15379 = pi0189 & n14516;
  assign n15380 = n15378 & ~n15379;
  assign n15381 = pi0189 & n15148;
  assign n15382 = ~n14612 & n15377;
  assign n15383 = ~pi0178 & ~n15381;
  assign n15384 = ~n15382 & n15383;
  assign n15385 = pi0181 & ~n15380;
  assign n15386 = ~n15384 & n15385;
  assign n15387 = pi0189 & n15177;
  assign n15388 = ~pi0189 & n15216;
  assign n15389 = pi0178 & ~n15388;
  assign n15390 = ~n15378 & ~n15389;
  assign n15391 = ~n15387 & ~n15390;
  assign n15392 = ~n10295 & ~n14514;
  assign n15393 = ~pi0189 & n14785;
  assign n15394 = ~n15392 & ~n15393;
  assign n15395 = ~pi0178 & ~n15394;
  assign n15396 = ~pi0181 & ~n15391;
  assign n15397 = ~n15395 & n15396;
  assign n15398 = n11765 & ~n15386;
  assign n15399 = ~n15397 & n15398;
  assign n15400 = ~pi0189 & ~n14612;
  assign n15401 = pi0189 & ~n14600;
  assign n15402 = ~pi0178 & ~n15401;
  assign n15403 = ~n15400 & n15402;
  assign n15404 = pi0178 & n11826;
  assign n15405 = n14596 & n15404;
  assign n15406 = pi0181 & ~n15405;
  assign n15407 = ~n14515 & n15406;
  assign n15408 = ~n15403 & n15407;
  assign n15409 = pi0189 & n15221;
  assign n15410 = n15389 & ~n15409;
  assign n15411 = ~pi0189 & n15140;
  assign n15412 = pi0189 & n15144;
  assign n15413 = ~pi0178 & ~n15412;
  assign n15414 = ~n15411 & n15413;
  assign n15415 = ~pi0181 & ~n15410;
  assign n15416 = ~n15414 & n15415;
  assign n15417 = n11833 & ~n15408;
  assign n15418 = ~n15416 & n15417;
  assign n15419 = pi0166 & n14597;
  assign n15420 = ~n14515 & ~n15419;
  assign n15421 = pi0153 & ~n15420;
  assign n15422 = ~pi0153 & ~n15324;
  assign n15423 = ~n14516 & n15422;
  assign n15424 = pi0157 & ~n15421;
  assign n15425 = ~n15423 & n15424;
  assign n15426 = pi0153 & pi0166;
  assign n15427 = ~n15187 & n15426;
  assign n15428 = ~pi0166 & ~n15137;
  assign n15429 = pi0166 & ~n15148;
  assign n15430 = pi0051 & n10299;
  assign n15431 = ~n15429 & ~n15430;
  assign n15432 = ~pi0153 & ~n15431;
  assign n15433 = ~pi0157 & ~n15427;
  assign n15434 = ~n15432 & n15433;
  assign n15435 = ~n15428 & n15434;
  assign n15436 = n9794 & ~n15425;
  assign n15437 = ~n15435 & n15436;
  assign n15438 = ~pi0166 & ~n15216;
  assign n15439 = pi0166 & ~n15177;
  assign n15440 = ~n15430 & ~n15439;
  assign n15441 = ~pi0153 & ~n15440;
  assign n15442 = ~n15221 & n15426;
  assign n15443 = pi0157 & ~n15442;
  assign n15444 = ~n15438 & n15443;
  assign n15445 = ~n15441 & n15444;
  assign n15446 = ~pi0166 & ~n15140;
  assign n15447 = pi0166 & ~n15144;
  assign n15448 = pi0153 & ~n15447;
  assign n15449 = ~n15446 & n15448;
  assign n15450 = ~pi0166 & n14785;
  assign n15451 = ~n10299 & ~n14514;
  assign n15452 = ~pi0153 & ~n15451;
  assign n15453 = ~n15450 & n15452;
  assign n15454 = ~n15449 & ~n15453;
  assign n15455 = ~pi0157 & ~n15454;
  assign n15456 = n9793 & ~n15445;
  assign n15457 = ~n15455 & n15456;
  assign n15458 = ~n15418 & ~n15437;
  assign n15459 = ~n15399 & n15458;
  assign n15460 = ~n15457 & n15459;
  assign n15461 = pi0232 & ~n15460;
  assign n15462 = n15302 & ~n15461;
  assign n15463 = ~n15332 & ~n15376;
  assign n15464 = ~n15462 & n15463;
  assign n15465 = ~pi0189 & n14982;
  assign n15466 = pi0189 & n14984;
  assign n15467 = ~pi0182 & ~n15466;
  assign n15468 = ~n15465 & n15467;
  assign n15469 = ~n14443 & n15468;
  assign n15470 = ~pi0189 & n14993;
  assign n15471 = pi0189 & ~n14999;
  assign n15472 = pi0182 & ~n15470;
  assign n15473 = ~n15471 & n15472;
  assign n15474 = ~n15469 & ~n15473;
  assign n15475 = n11833 & ~n15474;
  assign n15476 = ~pi0189 & ~n15010;
  assign n15477 = pi0189 & n15004;
  assign n15478 = pi0182 & ~n15477;
  assign n15479 = ~n15476 & n15478;
  assign n15480 = ~n15468 & ~n15479;
  assign n15481 = n11765 & ~n15480;
  assign n15482 = ~pi0160 & pi0216;
  assign n15483 = n6379 & ~n15482;
  assign n15484 = n15324 & ~n15483;
  assign n15485 = ~pi0166 & n14659;
  assign n15486 = pi0166 & n14776;
  assign n15487 = ~pi0153 & ~n15485;
  assign n15488 = ~n15486 & n15487;
  assign n15489 = pi0166 & ~n14965;
  assign n15490 = ~pi0166 & ~n14962;
  assign n15491 = pi0153 & ~n15490;
  assign n15492 = ~n15489 & n15491;
  assign n15493 = pi0160 & ~n15488;
  assign n15494 = ~n15492 & n15493;
  assign n15495 = pi0216 & ~n15494;
  assign n15496 = ~pi0166 & ~n14949;
  assign n15497 = pi0166 & ~n14951;
  assign n15498 = ~n15496 & ~n15497;
  assign n15499 = pi0051 & ~pi0153;
  assign n15500 = ~n15498 & ~n15499;
  assign n15501 = ~pi0216 & ~n15500;
  assign n15502 = n6379 & ~n15495;
  assign n15503 = ~n15501 & n15502;
  assign n15504 = pi0299 & ~n15484;
  assign n15505 = ~n15503 & n15504;
  assign n15506 = ~n15475 & ~n15481;
  assign n15507 = ~n15505 & n15506;
  assign n15508 = pi0232 & ~n15507;
  assign n15509 = n14945 & ~n15508;
  assign n15510 = ~pi0153 & n15064;
  assign n15511 = pi0153 & n15066;
  assign n15512 = pi0157 & ~n15511;
  assign n15513 = ~n15510 & n15512;
  assign n15514 = ~pi0153 & n15039;
  assign n15515 = pi0153 & ~n15042;
  assign n15516 = ~pi0157 & ~n15515;
  assign n15517 = ~n15514 & n15516;
  assign n15518 = ~n15513 & ~n15517;
  assign n15519 = pi0166 & ~n15518;
  assign n15520 = pi0157 & n15071;
  assign n15521 = ~pi0157 & n15033;
  assign n15522 = ~pi0166 & ~n15322;
  assign n15523 = ~n15520 & n15522;
  assign n15524 = ~n15521 & n15523;
  assign n15525 = ~n15519 & ~n15524;
  assign n15526 = n9794 & ~n15525;
  assign n15527 = ~pi0166 & n15050;
  assign n15528 = pi0166 & ~n15052;
  assign n15529 = pi0153 & ~n15527;
  assign n15530 = ~n15528 & n15529;
  assign n15531 = pi0166 & n15056;
  assign n15532 = ~pi0166 & ~n15058;
  assign n15533 = ~pi0153 & ~n15532;
  assign n15534 = ~n15531 & n15533;
  assign n15535 = ~n15530 & ~n15534;
  assign n15536 = pi0157 & ~n15535;
  assign n15537 = pi0166 & n14508;
  assign n15538 = ~pi0166 & ~n15084;
  assign n15539 = ~pi0157 & ~n15322;
  assign n15540 = ~n15537 & n15539;
  assign n15541 = ~n15538 & n15540;
  assign n15542 = ~n15536 & ~n15541;
  assign n15543 = n9793 & ~n15542;
  assign n15544 = ~pi0189 & ~n15084;
  assign n15545 = pi0189 & n14508;
  assign n15546 = ~pi0178 & ~n15545;
  assign n15547 = ~n14443 & n15546;
  assign n15548 = ~n15544 & n15547;
  assign n15549 = ~pi0181 & ~n15548;
  assign n15550 = pi0189 & ~n15052;
  assign n15551 = ~pi0189 & n15050;
  assign n15552 = pi0178 & ~n15551;
  assign n15553 = ~n15550 & n15552;
  assign n15554 = n15549 & ~n15553;
  assign n15555 = pi0189 & n15042;
  assign n15556 = ~pi0189 & ~n15033;
  assign n15557 = ~n14443 & n15556;
  assign n15558 = ~n15555 & ~n15557;
  assign n15559 = ~pi0178 & ~n15558;
  assign n15560 = ~pi0189 & n15071;
  assign n15561 = n15066 & ~n15377;
  assign n15562 = pi0178 & ~n15560;
  assign n15563 = ~n15561 & n15562;
  assign n15564 = pi0181 & ~n15559;
  assign n15565 = ~n15563 & n15564;
  assign n15566 = n11833 & ~n15554;
  assign n15567 = ~n15565 & n15566;
  assign n15568 = n15084 & n15546;
  assign n15569 = ~pi0189 & ~n15058;
  assign n15570 = pi0189 & n15056;
  assign n15571 = pi0178 & ~n15569;
  assign n15572 = ~n15570 & n15571;
  assign n15573 = n15549 & ~n15568;
  assign n15574 = ~n15572 & n15573;
  assign n15575 = pi0189 & n15064;
  assign n15576 = ~n15560 & ~n15575;
  assign n15577 = pi0178 & ~n15576;
  assign n15578 = pi0189 & ~n15039;
  assign n15579 = ~pi0178 & ~n15556;
  assign n15580 = ~n15578 & n15579;
  assign n15581 = ~n15577 & ~n15580;
  assign n15582 = pi0181 & ~n15581;
  assign n15583 = n11765 & ~n15574;
  assign n15584 = ~n15582 & n15583;
  assign n15585 = ~n15543 & ~n15567;
  assign n15586 = ~n15526 & n15585;
  assign n15587 = ~n15584 & n15586;
  assign n15588 = pi0232 & ~n15587;
  assign n15589 = n14939 & ~n15588;
  assign n15590 = n15332 & ~n15509;
  assign n15591 = ~n15589 & n15590;
  assign n15592 = n2608 & ~n15464;
  assign n15593 = ~n15591 & n15592;
  assign n15594 = n2535 & ~n15334;
  assign n15595 = ~n15328 & n15594;
  assign n15596 = ~n15593 & n15595;
  assign n15597 = n14455 & ~n15327;
  assign n15598 = ~pi0150 & pi0299;
  assign n15599 = ~pi0185 & ~pi0299;
  assign n15600 = ~n15598 & ~n15599;
  assign n15601 = n7473 & n15600;
  assign n15602 = pi0087 & ~n15601;
  assign n15603 = ~n15597 & ~n15602;
  assign n15604 = n14440 & ~n15332;
  assign n15605 = ~n15603 & ~n15604;
  assign n15606 = ~po1038 & ~n15605;
  assign n15607 = ~n15596 & n15606;
  assign n15608 = pi0232 & ~n15319;
  assign n15609 = n15332 & ~n15608;
  assign n15610 = ~pi0232 & ~n14439;
  assign n15611 = ~n15323 & ~n15610;
  assign n15612 = ~n15609 & n15611;
  assign n15613 = ~pi0087 & ~n15612;
  assign n15614 = pi0087 & ~n13685;
  assign n15615 = po1038 & ~n15614;
  assign n15616 = ~n15613 & n15615;
  assign po0283 = ~n15607 & ~n15616;
  assign n15618 = n2537 & n8887;
  assign n15619 = n2529 & n15618;
  assign n15620 = ~n3328 & ~n15619;
  assign n15621 = ~n2529 & ~n15618;
  assign n15622 = pi0129 & n7301;
  assign n15623 = n6323 & n15622;
  assign n15624 = pi0074 & ~n15623;
  assign n15625 = pi0054 & n2611;
  assign n15626 = n8887 & n15625;
  assign n15627 = pi0092 & ~pi0129;
  assign n15628 = pi0075 & n15622;
  assign n15629 = ~n2625 & ~n8965;
  assign n15630 = n8887 & ~n15629;
  assign n15631 = ~n2568 & ~n15630;
  assign n15632 = pi0129 & n6135;
  assign n15633 = pi0038 & ~n15632;
  assign n15634 = pi0039 & n8887;
  assign n15635 = ~n2729 & ~n3106;
  assign n15636 = n2788 & ~n2859;
  assign n15637 = n2462 & ~n15636;
  assign n15638 = n2873 & ~n15637;
  assign n15639 = n2785 & ~n15638;
  assign n15640 = n2877 & ~n15639;
  assign n15641 = n2719 & ~n15640;
  assign n15642 = ~n2722 & ~n15641;
  assign n15643 = ~pi0086 & ~n15642;
  assign n15644 = n2783 & ~n15643;
  assign n15645 = ~pi0097 & ~n15644;
  assign n15646 = ~n2776 & ~n15645;
  assign n15647 = ~pi0108 & ~n15646;
  assign n15648 = n2775 & ~n15647;
  assign n15649 = n2889 & ~n15648;
  assign n15650 = ~n2766 & ~n15649;
  assign n15651 = n2765 & ~n15650;
  assign n15652 = n2764 & ~n15651;
  assign n15653 = po0740 & n15652;
  assign n15654 = pi0250 & ~n7474;
  assign n15655 = n10077 & n15654;
  assign n15656 = n2781 & ~n15644;
  assign n15657 = ~n2776 & ~n15656;
  assign n15658 = ~pi0108 & ~n15657;
  assign n15659 = n2775 & ~n15658;
  assign n15660 = n2889 & ~n15659;
  assign n15661 = ~n2766 & ~n15660;
  assign n15662 = n2765 & ~n15661;
  assign n15663 = n2764 & ~n15662;
  assign n15664 = ~po0740 & n15663;
  assign n15665 = ~n15653 & n15655;
  assign n15666 = ~n15664 & n15665;
  assign n15667 = ~pi0127 & n15652;
  assign n15668 = pi0127 & n15663;
  assign n15669 = ~n15655 & ~n15667;
  assign n15670 = ~n15668 & n15669;
  assign n15671 = ~n15666 & ~n15670;
  assign n15672 = n2757 & ~n15671;
  assign n15673 = n3108 & ~n15672;
  assign n15674 = n2504 & ~n15673;
  assign n15675 = n15635 & ~n15674;
  assign n15676 = ~pi0070 & ~n15675;
  assign n15677 = ~n3099 & ~n15676;
  assign n15678 = ~pi0051 & ~n15677;
  assign n15679 = n2748 & ~n15678;
  assign n15680 = n3168 & ~n15679;
  assign n15681 = ~n2745 & ~n15680;
  assign n15682 = n2510 & ~n15681;
  assign n15683 = n3413 & ~n15682;
  assign n15684 = ~pi0095 & ~n15683;
  assign n15685 = ~pi0039 & pi0129;
  assign n15686 = ~n2741 & n15685;
  assign n15687 = ~n15684 & n15686;
  assign n15688 = ~pi0038 & ~n15634;
  assign n15689 = ~n15687 & n15688;
  assign n15690 = ~n15633 & ~n15689;
  assign n15691 = n2568 & ~n15690;
  assign n15692 = ~pi0075 & ~n15631;
  assign n15693 = ~n15691 & n15692;
  assign n15694 = ~pi0092 & ~n15628;
  assign n15695 = ~n15693 & n15694;
  assign n15696 = n13654 & ~n15627;
  assign n15697 = ~n15695 & n15696;
  assign n15698 = ~pi0074 & ~n15626;
  assign n15699 = ~n15697 & n15698;
  assign n15700 = ~pi0055 & ~n15624;
  assign n15701 = ~n15699 & n15700;
  assign n15702 = pi0055 & n2570;
  assign n15703 = n15622 & n15702;
  assign n15704 = ~n15701 & ~n15703;
  assign n15705 = ~pi0056 & ~n15704;
  assign n15706 = ~n11310 & ~n11318;
  assign n15707 = ~n15705 & n15706;
  assign n15708 = ~n15621 & ~n15707;
  assign n15709 = n3328 & ~n15708;
  assign n15710 = ~n6120 & ~n15620;
  assign po0284 = ~n15709 & n15710;
  assign n15712 = ~n6130 & ~n7347;
  assign n15713 = n8888 & n10391;
  assign n15714 = po0740 & n15713;
  assign n15715 = ~pi0129 & ~n15713;
  assign n15716 = n8967 & ~n15714;
  assign n15717 = ~n15715 & n15716;
  assign n15718 = n2521 & n15717;
  assign n15719 = ~pi0038 & ~n3418;
  assign n15720 = n6137 & ~n15719;
  assign n15721 = ~n6280 & n6286;
  assign n15722 = ~pi0087 & ~n15721;
  assign n15723 = ~n15720 & n15722;
  assign n15724 = n6133 & ~n15723;
  assign n15725 = n6134 & ~n15718;
  assign n15726 = ~n15724 & n15725;
  assign n15727 = ~n7305 & ~n7341;
  assign n15728 = ~n15726 & n15727;
  assign n15729 = n8879 & ~n15728;
  assign n15730 = n15712 & ~n15729;
  assign n15731 = ~pi0056 & ~n15730;
  assign n15732 = ~n6127 & ~n15731;
  assign n15733 = ~pi0062 & ~n15732;
  assign n15734 = ~n6299 & ~n15733;
  assign n15735 = n3328 & ~n15734;
  assign po0286 = n6123 & ~n15735;
  assign n15737 = pi0087 & ~n9747;
  assign n15738 = n7473 & ~n9022;
  assign n15739 = n14596 & ~n15738;
  assign n15740 = ~n15319 & ~n15739;
  assign n15741 = n14455 & ~n15740;
  assign n15742 = ~n15737 & ~n15741;
  assign n15743 = ~n14440 & ~n15742;
  assign n15744 = ~pi0132 & n15329;
  assign n15745 = pi0130 & ~n15744;
  assign n15746 = ~pi0130 & n15744;
  assign n15747 = ~n15745 & ~n15746;
  assign n15748 = ~n14429 & ~n15747;
  assign n15749 = pi0100 & n15740;
  assign n15750 = n2535 & ~n15749;
  assign n15751 = ~n10982 & n15739;
  assign n15752 = ~pi0051 & ~n15297;
  assign n15753 = ~pi0232 & ~n15752;
  assign n15754 = n10982 & ~n15753;
  assign n15755 = ~pi0191 & ~pi0299;
  assign n15756 = ~pi0051 & ~n15256;
  assign n15757 = pi0140 & n15282;
  assign n15758 = n15756 & ~n15757;
  assign n15759 = n15755 & ~n15758;
  assign n15760 = ~pi0051 & n15263;
  assign n15761 = pi0140 & n14657;
  assign n15762 = n15760 & ~n15761;
  assign n15763 = n9020 & ~n15762;
  assign n15764 = pi0169 & n6197;
  assign n15765 = ~n9036 & n14596;
  assign n15766 = ~n15764 & n15765;
  assign n15767 = pi0162 & n9036;
  assign n15768 = ~pi0051 & ~n14678;
  assign n15769 = ~n14657 & n15768;
  assign n15770 = pi0169 & ~n15769;
  assign n15771 = ~pi0169 & ~n15281;
  assign n15772 = n15767 & ~n15771;
  assign n15773 = ~n15770 & n15772;
  assign n15774 = ~n2521 & n15764;
  assign n15775 = ~n14655 & ~n15764;
  assign n15776 = ~pi0162 & n9036;
  assign n15777 = ~n15775 & n15776;
  assign n15778 = ~n15774 & n15777;
  assign n15779 = pi0299 & ~n15766;
  assign n15780 = ~n15778 & n15779;
  assign n15781 = ~n15773 & n15780;
  assign n15782 = ~n15759 & ~n15763;
  assign n15783 = ~n15781 & n15782;
  assign n15784 = pi0232 & ~n15783;
  assign n15785 = n15754 & ~n15784;
  assign n15786 = ~pi0100 & ~n15751;
  assign n15787 = ~n15785 & n15786;
  assign n15788 = ~n14467 & n15750;
  assign n15789 = ~n15787 & n15788;
  assign n15790 = ~n15743 & ~n15748;
  assign n15791 = ~n15789 & n15790;
  assign n15792 = ~n14676 & ~n15764;
  assign n15793 = pi0169 & n14948;
  assign n15794 = ~n15792 & ~n15793;
  assign n15795 = ~pi0216 & ~n15794;
  assign n15796 = ~n14666 & n14962;
  assign n15797 = pi0169 & n15796;
  assign n15798 = ~pi0051 & ~n14964;
  assign n15799 = ~pi0169 & n15798;
  assign n15800 = pi0162 & pi0216;
  assign n15801 = ~n15797 & n15800;
  assign n15802 = ~n15799 & n15801;
  assign n15803 = ~n15795 & ~n15802;
  assign n15804 = n6379 & ~n15803;
  assign n15805 = pi0169 & n14597;
  assign n15806 = ~pi0051 & ~n15805;
  assign n15807 = ~n7570 & ~n15767;
  assign n15808 = ~n15806 & n15807;
  assign n15809 = ~n15804 & ~n15808;
  assign n15810 = pi0299 & ~n15809;
  assign n15811 = n7551 & n14675;
  assign n15812 = ~pi0051 & ~n15811;
  assign n15813 = ~pi0140 & n15812;
  assign n15814 = n14675 & n14996;
  assign n15815 = ~pi0051 & ~n15814;
  assign n15816 = pi0140 & n15815;
  assign n15817 = n15755 & ~n15813;
  assign n15818 = ~n15816 & n15817;
  assign n15819 = ~n6197 & ~n14676;
  assign n15820 = ~n14948 & ~n15819;
  assign n15821 = n7551 & ~n15820;
  assign n15822 = ~n7551 & ~n15319;
  assign n15823 = ~n15821 & ~n15822;
  assign n15824 = ~pi0140 & n15823;
  assign n15825 = pi0224 & ~n15796;
  assign n15826 = ~pi0224 & ~n15820;
  assign n15827 = ~n15825 & ~n15826;
  assign n15828 = n6405 & ~n15827;
  assign n15829 = ~n6405 & ~n15319;
  assign n15830 = ~n15828 & ~n15829;
  assign n15831 = pi0140 & n15830;
  assign n15832 = n9020 & ~n15824;
  assign n15833 = ~n15831 & n15832;
  assign n15834 = ~n15810 & ~n15818;
  assign n15835 = ~n15833 & n15834;
  assign n15836 = pi0232 & ~n15835;
  assign n15837 = n14675 & n14942;
  assign n15838 = ~pi0051 & ~n15837;
  assign n15839 = ~pi0232 & ~n15838;
  assign n15840 = pi0039 & ~n15839;
  assign n15841 = ~n15836 & n15840;
  assign n15842 = ~pi0232 & ~n14578;
  assign n15843 = ~pi0039 & ~n15842;
  assign n15844 = ~n6197 & n14578;
  assign n15845 = ~n15070 & ~n15844;
  assign n15846 = ~n9022 & ~n15845;
  assign n15847 = n9022 & n14578;
  assign n15848 = pi0232 & ~n15847;
  assign n15849 = ~n15846 & n15848;
  assign n15850 = n15843 & ~n15849;
  assign n15851 = ~n15841 & ~n15850;
  assign n15852 = ~pi0038 & ~n15851;
  assign n15853 = pi0038 & ~n15740;
  assign n15854 = ~pi0100 & ~n15853;
  assign n15855 = ~n15852 & n15854;
  assign n15856 = n15750 & ~n15855;
  assign n15857 = n15742 & n15748;
  assign n15858 = ~n15856 & n15857;
  assign n15859 = ~n15791 & ~n15858;
  assign n15860 = ~po1038 & ~n15859;
  assign n15861 = pi0087 & ~n9705;
  assign n15862 = pi0169 & n7473;
  assign n15863 = ~pi0087 & n14596;
  assign n15864 = ~n15862 & n15863;
  assign n15865 = ~pi0051 & ~pi0087;
  assign n15866 = ~n15805 & n15865;
  assign n15867 = n15748 & n15866;
  assign n15868 = po1038 & ~n15861;
  assign n15869 = ~n15864 & n15868;
  assign n15870 = ~n15867 & n15869;
  assign po0287 = ~n15860 & ~n15870;
  assign n15872 = ~pi0100 & ~n14009;
  assign n15873 = ~pi0087 & ~n7334;
  assign n15874 = ~n15872 & n15873;
  assign n15875 = ~pi0075 & ~n15874;
  assign n15876 = ~n7302 & ~n15875;
  assign n15877 = ~pi0092 & ~n15876;
  assign n15878 = n8880 & n13654;
  assign po0288 = ~n15877 & n15878;
  assign n15880 = pi0164 & n14920;
  assign n15881 = pi0051 & ~pi0151;
  assign n15882 = ~n13752 & ~n14443;
  assign n15883 = ~n15881 & ~n15882;
  assign n15884 = n14446 & n15883;
  assign n15885 = pi0232 & n15884;
  assign n15886 = pi0132 & ~n15329;
  assign n15887 = ~n15744 & ~n15886;
  assign n15888 = ~n14430 & ~n15887;
  assign n15889 = n14439 & ~n15888;
  assign n15890 = ~n15885 & ~n15889;
  assign n15891 = ~pi0087 & ~n15890;
  assign n15892 = po1038 & ~n15880;
  assign n15893 = ~n15891 & n15892;
  assign n15894 = pi0173 & n14443;
  assign n15895 = pi0190 & n14597;
  assign n15896 = ~pi0299 & ~n15894;
  assign n15897 = ~n15895 & n15896;
  assign n15898 = pi0299 & ~n15884;
  assign n15899 = pi0232 & ~n15897;
  assign n15900 = ~n15898 & n15899;
  assign n15901 = n14455 & ~n15900;
  assign n15902 = pi0087 & ~n9030;
  assign n15903 = ~n2608 & n15900;
  assign n15904 = ~n13752 & n14608;
  assign n15905 = pi0168 & n14592;
  assign n15906 = ~pi0151 & ~n15905;
  assign n15907 = ~n15904 & n15906;
  assign n15908 = ~n6197 & ~n14608;
  assign n15909 = pi0168 & ~n15049;
  assign n15910 = ~n15908 & n15909;
  assign n15911 = ~n6197 & n14608;
  assign n15912 = n14613 & ~n15911;
  assign n15913 = ~pi0168 & ~n15912;
  assign n15914 = pi0151 & ~n15910;
  assign n15915 = ~n15913 & n15914;
  assign n15916 = ~pi0160 & ~n15907;
  assign n15917 = ~n15915 & n15916;
  assign n15918 = pi0151 & n14578;
  assign n15919 = ~pi0151 & ~n14584;
  assign n15920 = ~pi0168 & ~n15918;
  assign n15921 = ~n15919 & n15920;
  assign n15922 = pi0168 & ~n15881;
  assign n15923 = ~n14506 & n15922;
  assign n15924 = n6197 & ~n15923;
  assign n15925 = ~n15921 & n15924;
  assign n15926 = pi0160 & ~n15908;
  assign n15927 = ~n15925 & n15926;
  assign n15928 = pi0299 & ~n15917;
  assign n15929 = ~n15927 & n15928;
  assign n15930 = pi0190 & ~pi0299;
  assign n15931 = pi0051 & ~pi0173;
  assign n15932 = pi0182 & n14486;
  assign n15933 = n14505 & ~n15932;
  assign n15934 = n6197 & ~n15931;
  assign n15935 = ~n15933 & n15934;
  assign n15936 = n15930 & ~n15935;
  assign n15937 = ~n15911 & n15936;
  assign n15938 = ~pi0190 & ~pi0299;
  assign n15939 = ~pi0182 & n14608;
  assign n15940 = pi0182 & ~n15908;
  assign n15941 = ~n14585 & n15940;
  assign n15942 = ~pi0173 & ~n15939;
  assign n15943 = ~n15941 & n15942;
  assign n15944 = ~pi0182 & ~n15912;
  assign n15945 = ~n14579 & ~n15911;
  assign n15946 = pi0182 & ~n15945;
  assign n15947 = pi0173 & ~n15944;
  assign n15948 = ~n15946 & n15947;
  assign n15949 = ~n15943 & ~n15948;
  assign n15950 = n15938 & ~n15949;
  assign n15951 = pi0232 & ~n15937;
  assign n15952 = ~n15929 & n15951;
  assign n15953 = ~n15950 & n15952;
  assign n15954 = ~pi0232 & n14608;
  assign n15955 = ~n15953 & ~n15954;
  assign n15956 = ~pi0039 & ~n15955;
  assign n15957 = ~pi0183 & n14979;
  assign n15958 = pi0183 & ~n15010;
  assign n15959 = ~pi0183 & ~n14981;
  assign n15960 = ~pi0173 & ~n15959;
  assign n15961 = ~n15958 & n15960;
  assign n15962 = ~pi0183 & ~n14989;
  assign n15963 = pi0173 & ~n14993;
  assign n15964 = ~n15962 & n15963;
  assign n15965 = ~n15957 & ~n15964;
  assign n15966 = ~n15961 & n15965;
  assign n15967 = n15930 & ~n15966;
  assign n15968 = ~pi0183 & ~n7551;
  assign n15969 = ~pi0173 & ~n15968;
  assign n15970 = n15004 & n15969;
  assign n15971 = pi0183 & n14999;
  assign n15972 = ~pi0183 & ~n14443;
  assign n15973 = ~n14984 & n15972;
  assign n15974 = pi0173 & ~n15973;
  assign n15975 = ~n15971 & n15974;
  assign n15976 = n15938 & ~n15970;
  assign n15977 = ~n15975 & n15976;
  assign n15978 = ~pi0149 & pi0216;
  assign n15979 = n6379 & ~n15978;
  assign n15980 = n15884 & ~n15979;
  assign n15981 = ~pi0168 & n14776;
  assign n15982 = pi0168 & n14659;
  assign n15983 = ~pi0151 & ~n15982;
  assign n15984 = ~n15981 & n15983;
  assign n15985 = ~pi0168 & ~n14965;
  assign n15986 = pi0168 & ~n14962;
  assign n15987 = pi0151 & ~n15986;
  assign n15988 = ~n15985 & n15987;
  assign n15989 = pi0149 & ~n15984;
  assign n15990 = ~n15988 & n15989;
  assign n15991 = pi0216 & ~n15990;
  assign n15992 = pi0168 & ~n14949;
  assign n15993 = ~pi0168 & ~n14951;
  assign n15994 = ~n15992 & ~n15993;
  assign n15995 = ~n15881 & ~n15994;
  assign n15996 = ~pi0216 & ~n15995;
  assign n15997 = n6379 & ~n15991;
  assign n15998 = ~n15996 & n15997;
  assign n15999 = pi0299 & ~n15980;
  assign n16000 = ~n15998 & n15999;
  assign n16001 = ~n15967 & ~n15977;
  assign n16002 = ~n16000 & n16001;
  assign n16003 = pi0232 & ~n16002;
  assign n16004 = n14945 & ~n16003;
  assign n16005 = ~n15956 & ~n16004;
  assign n16006 = n2608 & ~n16005;
  assign n16007 = n2535 & ~n15903;
  assign n16008 = ~n16006 & n16007;
  assign n16009 = n15888 & ~n15902;
  assign n16010 = ~n15901 & n16009;
  assign n16011 = ~n16008 & n16010;
  assign n16012 = n14456 & ~n15900;
  assign n16013 = ~n14439 & n15898;
  assign n16014 = ~n13130 & ~n16013;
  assign n16015 = ~pi0168 & ~n14667;
  assign n16016 = pi0168 & ~n14673;
  assign n16017 = pi0151 & ~n16015;
  assign n16018 = ~n16016 & n16017;
  assign n16019 = pi0168 & n14677;
  assign n16020 = ~n13752 & ~n14654;
  assign n16021 = ~pi0151 & ~n16020;
  assign n16022 = ~n16019 & n16021;
  assign n16023 = ~pi0149 & ~n16022;
  assign n16024 = ~n16018 & n16023;
  assign n16025 = ~n14714 & ~n15883;
  assign n16026 = ~pi0168 & ~n16025;
  assign n16027 = ~n14965 & ~n15881;
  assign n16028 = ~n14678 & ~n16027;
  assign n16029 = pi0168 & ~n16028;
  assign n16030 = pi0149 & ~n16026;
  assign n16031 = ~n16029 & n16030;
  assign n16032 = n9036 & ~n16024;
  assign n16033 = ~n16031 & n16032;
  assign n16034 = ~n16014 & ~n16033;
  assign n16035 = ~pi0183 & ~n15271;
  assign n16036 = pi0183 & ~n15279;
  assign n16037 = pi0173 & ~n16036;
  assign n16038 = ~n16035 & n16037;
  assign n16039 = pi0183 & n14683;
  assign n16040 = ~pi0173 & ~n16039;
  assign n16041 = n15263 & n16040;
  assign n16042 = ~n16038 & ~n16041;
  assign n16043 = n15930 & ~n16042;
  assign n16044 = pi0183 & n14714;
  assign n16045 = ~n15894 & n15938;
  assign n16046 = ~n15256 & n16045;
  assign n16047 = ~n16044 & n16046;
  assign n16048 = ~n16034 & ~n16047;
  assign n16049 = ~n16043 & n16048;
  assign n16050 = pi0232 & ~n16049;
  assign n16051 = ~n15298 & ~n16050;
  assign n16052 = pi0039 & ~n16051;
  assign n16053 = ~pi0232 & n14513;
  assign n16054 = pi0182 & n15147;
  assign n16055 = ~n14513 & n16045;
  assign n16056 = ~n16054 & n16055;
  assign n16057 = ~pi0182 & n14537;
  assign n16058 = ~n15146 & ~n15931;
  assign n16059 = ~n16057 & n16058;
  assign n16060 = n15930 & ~n16059;
  assign n16061 = ~pi0168 & n14597;
  assign n16062 = ~n15146 & ~n16061;
  assign n16063 = pi0151 & ~n16062;
  assign n16064 = ~pi0151 & ~n15884;
  assign n16065 = ~n15147 & n16064;
  assign n16066 = pi0160 & ~n16063;
  assign n16067 = ~n16065 & n16066;
  assign n16068 = ~pi0151 & ~n14513;
  assign n16069 = pi0151 & n14750;
  assign n16070 = ~pi0168 & ~n16068;
  assign n16071 = ~n16069 & n16070;
  assign n16072 = ~pi0151 & n14443;
  assign n16073 = pi0168 & ~n16072;
  assign n16074 = ~n14537 & n16073;
  assign n16075 = ~n16071 & ~n16074;
  assign n16076 = ~pi0160 & ~n15146;
  assign n16077 = ~n16075 & n16076;
  assign n16078 = pi0299 & ~n16067;
  assign n16079 = ~n16077 & n16078;
  assign n16080 = pi0232 & ~n16056;
  assign n16081 = ~n16060 & n16080;
  assign n16082 = ~n16079 & n16081;
  assign n16083 = ~pi0039 & ~n16053;
  assign n16084 = ~n16082 & n16083;
  assign n16085 = n2608 & ~n16084;
  assign n16086 = ~n16052 & n16085;
  assign n16087 = n2535 & ~n15333;
  assign n16088 = ~n15903 & n16087;
  assign n16089 = ~n16086 & n16088;
  assign n16090 = ~n15888 & ~n15902;
  assign n16091 = ~n16012 & n16090;
  assign n16092 = ~n16089 & n16091;
  assign n16093 = ~po1038 & ~n16092;
  assign n16094 = ~n16011 & n16093;
  assign po0289 = n15893 | n16094;
  assign n16096 = ~pi0133 & ~n14909;
  assign n16097 = pi0145 & n14714;
  assign n16098 = n15293 & ~n16097;
  assign n16099 = pi0197 & n14657;
  assign n16100 = n15294 & ~n16099;
  assign n16101 = n14439 & ~n16100;
  assign n16102 = pi0299 & ~n16101;
  assign n16103 = ~n16098 & ~n16102;
  assign n16104 = pi0232 & ~n16103;
  assign n16105 = n15299 & ~n16104;
  assign n16106 = ~n9212 & n14503;
  assign n16107 = ~pi0039 & n14439;
  assign n16108 = ~n16106 & n16107;
  assign n16109 = ~pi0038 & ~n16108;
  assign n16110 = ~n16105 & n16109;
  assign n16111 = n14473 & ~n16110;
  assign n16112 = n14468 & ~n16111;
  assign n16113 = ~n14456 & ~n16112;
  assign n16114 = ~n16096 & ~n16113;
  assign n16115 = ~pi0183 & ~pi0299;
  assign n16116 = ~pi0149 & pi0299;
  assign n16117 = ~n16115 & ~n16116;
  assign n16118 = n7473 & n16117;
  assign n16119 = pi0087 & ~n16118;
  assign n16120 = ~n9209 & n14532;
  assign n16121 = ~n6197 & ~n14532;
  assign n16122 = ~n14585 & ~n16121;
  assign n16123 = n9209 & n16122;
  assign n16124 = ~pi0039 & pi0176;
  assign n16125 = ~n16120 & n16124;
  assign n16126 = ~n16123 & n16125;
  assign n16127 = ~n5777 & ~n16099;
  assign n16128 = n6640 & ~n16127;
  assign n16129 = ~pi0145 & ~n7551;
  assign n16130 = ~pi0299 & ~n16129;
  assign n16131 = ~n15003 & n16130;
  assign n16132 = ~n16128 & ~n16131;
  assign n16133 = n2521 & ~n16132;
  assign n16134 = pi0232 & ~n16133;
  assign n16135 = ~n14944 & ~n16134;
  assign n16136 = pi0039 & ~n16135;
  assign n16137 = pi0154 & pi0232;
  assign n16138 = pi0299 & n16137;
  assign n16139 = n14532 & ~n16138;
  assign n16140 = n16122 & n16138;
  assign n16141 = ~pi0039 & ~pi0176;
  assign n16142 = ~n16139 & n16141;
  assign n16143 = ~n16140 & n16142;
  assign n16144 = n11374 & ~n16136;
  assign n16145 = ~n16126 & n16144;
  assign n16146 = ~n16143 & n16145;
  assign n16147 = ~pi0087 & n16096;
  assign n16148 = ~n16146 & n16147;
  assign n16149 = ~n16114 & ~n16119;
  assign n16150 = ~n16148 & n16149;
  assign n16151 = ~po1038 & ~n16150;
  assign n16152 = pi0149 & n14920;
  assign n16153 = n14440 & ~n16096;
  assign n16154 = po1038 & ~n16152;
  assign n16155 = ~n16153 & n16154;
  assign po0290 = n16151 | n16155;
  assign n16157 = po1038 & n15865;
  assign n16158 = ~pi0136 & n15746;
  assign n16159 = ~pi0135 & n16158;
  assign n16160 = pi0134 & ~n16159;
  assign n16161 = n14438 & ~n16160;
  assign n16162 = pi0171 & n6197;
  assign n16163 = ~n14438 & n16162;
  assign n16164 = pi0232 & n16163;
  assign n16165 = n16157 & ~n16164;
  assign n16166 = ~n16161 & n16165;
  assign n16167 = pi0192 & ~pi0299;
  assign n16168 = pi0171 & pi0299;
  assign n16169 = ~n16167 & ~n16168;
  assign n16170 = n7473 & ~n16169;
  assign n16171 = n14596 & ~n16170;
  assign n16172 = ~n15319 & ~n16171;
  assign n16173 = n14455 & ~n16172;
  assign n16174 = ~n2608 & n16172;
  assign n16175 = n2535 & ~n16174;
  assign n16176 = ~pi0051 & ~n16163;
  assign n16177 = ~pi0164 & pi0216;
  assign n16178 = n6379 & ~n16177;
  assign n16179 = ~n16176 & ~n16178;
  assign n16180 = ~n14676 & ~n16162;
  assign n16181 = pi0171 & n14948;
  assign n16182 = ~n16180 & ~n16181;
  assign n16183 = ~pi0216 & ~n16182;
  assign n16184 = pi0171 & n15796;
  assign n16185 = ~pi0171 & n15798;
  assign n16186 = pi0164 & pi0216;
  assign n16187 = ~n16184 & n16186;
  assign n16188 = ~n16185 & n16187;
  assign n16189 = ~n16183 & ~n16188;
  assign n16190 = n6379 & ~n16189;
  assign n16191 = ~n16179 & ~n16190;
  assign n16192 = pi0299 & ~n16191;
  assign n16193 = ~pi0192 & ~pi0299;
  assign n16194 = ~n15812 & n16193;
  assign n16195 = pi0039 & pi0186;
  assign n16196 = ~n15823 & n16167;
  assign n16197 = ~n16194 & ~n16195;
  assign n16198 = ~n16196 & n16197;
  assign n16199 = ~n15815 & n16193;
  assign n16200 = ~n15830 & n16167;
  assign n16201 = pi0186 & ~n16199;
  assign n16202 = ~n16200 & n16201;
  assign n16203 = ~n16198 & ~n16202;
  assign n16204 = ~n16192 & ~n16203;
  assign n16205 = pi0232 & ~n16204;
  assign n16206 = n15840 & ~n16205;
  assign n16207 = pi0232 & ~n16169;
  assign n16208 = ~n14578 & ~n16207;
  assign n16209 = n15845 & n16207;
  assign n16210 = ~pi0039 & ~n16208;
  assign n16211 = ~n16209 & n16210;
  assign n16212 = n2608 & ~n16206;
  assign n16213 = ~n16211 & n16212;
  assign n16214 = n16175 & ~n16213;
  assign n16215 = n16160 & ~n16173;
  assign n16216 = ~n16214 & n16215;
  assign n16217 = n14455 & n16171;
  assign n16218 = pi0039 & ~pi0186;
  assign n16219 = ~n15760 & n16167;
  assign n16220 = ~n15756 & n16193;
  assign n16221 = ~n16219 & ~n16220;
  assign n16222 = n15765 & ~n16162;
  assign n16223 = pi0299 & ~n16222;
  assign n16224 = ~n14655 & ~n16162;
  assign n16225 = n4192 & n6197;
  assign n16226 = n9036 & ~n16224;
  assign n16227 = ~n16225 & n16226;
  assign n16228 = n16223 & ~n16227;
  assign n16229 = n16221 & ~n16228;
  assign n16230 = pi0232 & ~n16229;
  assign n16231 = ~n15753 & ~n16230;
  assign n16232 = n16218 & ~n16231;
  assign n16233 = ~pi0039 & ~n16171;
  assign n16234 = ~n14657 & n15760;
  assign n16235 = n16167 & ~n16234;
  assign n16236 = ~n15282 & n15756;
  assign n16237 = n16193 & ~n16236;
  assign n16238 = ~n16235 & ~n16237;
  assign n16239 = ~n16228 & n16238;
  assign n16240 = pi0232 & ~n16239;
  assign n16241 = ~n15753 & ~n16240;
  assign n16242 = n16195 & ~n16241;
  assign n16243 = ~pi0164 & ~n16233;
  assign n16244 = ~n16232 & n16243;
  assign n16245 = ~n16242 & n16244;
  assign n16246 = ~pi0171 & ~n15281;
  assign n16247 = pi0171 & ~n15769;
  assign n16248 = n9036 & ~n16246;
  assign n16249 = ~n16247 & n16248;
  assign n16250 = n16223 & ~n16249;
  assign n16251 = n16221 & ~n16250;
  assign n16252 = pi0232 & ~n16251;
  assign n16253 = ~n15753 & ~n16252;
  assign n16254 = n16218 & ~n16253;
  assign n16255 = n16238 & ~n16250;
  assign n16256 = pi0232 & ~n16255;
  assign n16257 = ~n15753 & ~n16256;
  assign n16258 = n16195 & ~n16257;
  assign n16259 = pi0164 & ~n16233;
  assign n16260 = ~n16254 & n16259;
  assign n16261 = ~n16258 & n16260;
  assign n16262 = n2608 & ~n16245;
  assign n16263 = ~n16261 & n16262;
  assign n16264 = ~n15333 & n16175;
  assign n16265 = ~n16263 & n16264;
  assign n16266 = ~n16160 & ~n16217;
  assign n16267 = ~n16265 & n16266;
  assign n16268 = ~po1038 & ~n16216;
  assign n16269 = ~n16267 & n16268;
  assign po0291 = n16166 | n16269;
  assign n16271 = pi0135 & ~n16158;
  assign n16272 = pi0134 & n16159;
  assign n16273 = ~n16271 & ~n16272;
  assign n16274 = pi0170 & n6197;
  assign n16275 = n10598 & n16274;
  assign n16276 = n14596 & ~n16275;
  assign n16277 = pi0194 & n9193;
  assign n16278 = n16276 & ~n16277;
  assign n16279 = n14455 & n16278;
  assign n16280 = pi0185 & n15282;
  assign n16281 = n15756 & ~n16280;
  assign n16282 = ~n10982 & n16276;
  assign n16283 = ~pi0194 & ~n16282;
  assign n16284 = ~n16281 & n16283;
  assign n16285 = ~pi0185 & n15760;
  assign n16286 = pi0170 & n7473;
  assign n16287 = ~n9193 & ~n16286;
  assign n16288 = n14596 & n16287;
  assign n16289 = ~n10982 & n16288;
  assign n16290 = pi0194 & ~n16289;
  assign n16291 = ~n16234 & n16290;
  assign n16292 = ~n16285 & n16291;
  assign n16293 = ~n16284 & ~n16292;
  assign n16294 = ~pi0299 & ~n16293;
  assign n16295 = n15765 & ~n16274;
  assign n16296 = pi0150 & pi0299;
  assign n16297 = ~pi0170 & ~n15281;
  assign n16298 = pi0170 & ~n15769;
  assign n16299 = n9036 & ~n16297;
  assign n16300 = ~n16298 & n16299;
  assign n16301 = n16296 & ~n16300;
  assign n16302 = ~n14655 & ~n16274;
  assign n16303 = n4415 & n6197;
  assign n16304 = n9036 & ~n16302;
  assign n16305 = ~n16303 & n16304;
  assign n16306 = n15598 & ~n16305;
  assign n16307 = ~n16301 & ~n16306;
  assign n16308 = ~n16283 & ~n16290;
  assign n16309 = ~n16295 & ~n16308;
  assign n16310 = ~n16307 & n16309;
  assign n16311 = ~n16294 & ~n16310;
  assign n16312 = pi0232 & ~n16311;
  assign n16313 = ~n15754 & ~n16308;
  assign n16314 = ~n16312 & ~n16313;
  assign n16315 = ~pi0100 & ~n16314;
  assign n16316 = ~n15319 & ~n16278;
  assign n16317 = pi0100 & n16316;
  assign n16318 = n2535 & ~n16317;
  assign n16319 = ~n14467 & n16318;
  assign n16320 = ~n16315 & n16319;
  assign n16321 = n16273 & ~n16279;
  assign n16322 = ~n16320 & n16321;
  assign n16323 = ~n15319 & ~n16276;
  assign n16324 = pi0038 & ~n16323;
  assign n16325 = ~n14438 & n16274;
  assign n16326 = ~pi0051 & ~n16325;
  assign n16327 = ~n6379 & n16326;
  assign n16328 = pi0170 & n14948;
  assign n16329 = ~n14676 & ~n16274;
  assign n16330 = n7570 & ~n16328;
  assign n16331 = ~n16329 & n16330;
  assign n16332 = ~n9036 & ~n16331;
  assign n16333 = ~pi0170 & n15798;
  assign n16334 = pi0170 & n15796;
  assign n16335 = pi0216 & ~n16334;
  assign n16336 = ~n16333 & n16335;
  assign n16337 = ~n16332 & ~n16336;
  assign n16338 = n16296 & ~n16327;
  assign n16339 = ~n16337 & n16338;
  assign n16340 = ~n7570 & n16326;
  assign n16341 = n15598 & ~n16340;
  assign n16342 = ~n16331 & n16341;
  assign n16343 = ~n16339 & ~n16342;
  assign n16344 = ~pi0185 & n15812;
  assign n16345 = pi0185 & n15815;
  assign n16346 = ~pi0299 & ~n16344;
  assign n16347 = ~n16345 & n16346;
  assign n16348 = n16343 & ~n16347;
  assign n16349 = pi0232 & ~n16348;
  assign n16350 = n15840 & ~n16349;
  assign n16351 = ~pi0299 & ~n14578;
  assign n16352 = pi0170 & ~n15845;
  assign n16353 = ~pi0170 & n14578;
  assign n16354 = n10598 & ~n16353;
  assign n16355 = ~n16352 & n16354;
  assign n16356 = n15843 & ~n16355;
  assign n16357 = ~n16351 & n16356;
  assign n16358 = ~n16350 & ~n16357;
  assign n16359 = ~pi0038 & ~n16358;
  assign n16360 = ~pi0194 & ~n16324;
  assign n16361 = ~n16359 & n16360;
  assign n16362 = ~n15319 & ~n16288;
  assign n16363 = pi0038 & ~n16362;
  assign n16364 = ~pi0185 & n15823;
  assign n16365 = pi0185 & n15830;
  assign n16366 = ~pi0299 & ~n16364;
  assign n16367 = ~n16365 & n16366;
  assign n16368 = n16343 & ~n16367;
  assign n16369 = pi0232 & ~n16368;
  assign n16370 = n15840 & ~n16369;
  assign n16371 = n10602 & n15845;
  assign n16372 = n16356 & ~n16371;
  assign n16373 = ~n16370 & ~n16372;
  assign n16374 = ~pi0038 & ~n16373;
  assign n16375 = pi0194 & ~n16363;
  assign n16376 = ~n16374 & n16375;
  assign n16377 = ~n16361 & ~n16376;
  assign n16378 = ~pi0100 & ~n16377;
  assign n16379 = n16318 & ~n16378;
  assign n16380 = n14455 & ~n16316;
  assign n16381 = ~n16273 & ~n16380;
  assign n16382 = ~n16379 & n16381;
  assign n16383 = ~po1038 & ~n16322;
  assign n16384 = ~n16382 & n16383;
  assign n16385 = n14438 & n16273;
  assign n16386 = ~n14438 & n16286;
  assign n16387 = n16157 & ~n16386;
  assign n16388 = ~n16385 & n16387;
  assign po0292 = n16384 | n16388;
  assign n16390 = pi0136 & ~n15746;
  assign n16391 = ~n16158 & ~n16390;
  assign n16392 = ~n14428 & ~n16391;
  assign n16393 = ~n14596 & n16392;
  assign n16394 = pi0148 & n7473;
  assign n16395 = ~n14438 & ~n16394;
  assign n16396 = ~n16393 & ~n16395;
  assign n16397 = n16157 & ~n16396;
  assign n16398 = n9739 & ~n14438;
  assign n16399 = ~pi0051 & ~n16398;
  assign n16400 = n14455 & n16399;
  assign n16401 = ~n2608 & ~n16399;
  assign n16402 = ~n9738 & ~n15845;
  assign n16403 = n9738 & n14578;
  assign n16404 = pi0232 & ~n16403;
  assign n16405 = ~n16402 & n16404;
  assign n16406 = n15843 & ~n16405;
  assign n16407 = ~pi0184 & n15823;
  assign n16408 = pi0184 & n15830;
  assign n16409 = n9736 & ~n16407;
  assign n16410 = ~n16408 & n16409;
  assign n16411 = ~pi0141 & ~pi0299;
  assign n16412 = ~pi0184 & n15812;
  assign n16413 = pi0184 & n15815;
  assign n16414 = n16411 & ~n16412;
  assign n16415 = ~n16413 & n16414;
  assign n16416 = ~pi0287 & n13665;
  assign n16417 = pi0216 & ~n16416;
  assign n16418 = n6379 & ~n16417;
  assign n16419 = n14675 & n16418;
  assign n16420 = ~pi0051 & ~pi0148;
  assign n16421 = ~n16419 & n16420;
  assign n16422 = ~n6379 & n15319;
  assign n16423 = ~n7570 & ~n15319;
  assign n16424 = ~pi0163 & ~n16423;
  assign n16425 = pi0163 & n6379;
  assign n16426 = n15796 & n16425;
  assign n16427 = ~n16422 & ~n16424;
  assign n16428 = ~n16426 & n16427;
  assign n16429 = n7570 & ~n15820;
  assign n16430 = pi0148 & ~n16428;
  assign n16431 = ~n16429 & n16430;
  assign n16432 = pi0299 & ~n16421;
  assign n16433 = ~n16431 & n16432;
  assign n16434 = ~n16415 & ~n16433;
  assign n16435 = ~n16410 & n16434;
  assign n16436 = pi0232 & ~n16435;
  assign n16437 = n15840 & ~n16436;
  assign n16438 = n2608 & ~n16437;
  assign n16439 = ~n16406 & n16438;
  assign n16440 = n2535 & ~n16401;
  assign n16441 = ~n16439 & n16440;
  assign n16442 = n16392 & ~n16400;
  assign n16443 = ~n16441 & n16442;
  assign n16444 = ~n14438 & n16400;
  assign n16445 = ~n11211 & ~n14438;
  assign n16446 = n16399 & n16445;
  assign n16447 = pi0184 & n15282;
  assign n16448 = n15756 & ~n16447;
  assign n16449 = n16411 & ~n16448;
  assign n16450 = pi0184 & n14657;
  assign n16451 = n15760 & ~n16450;
  assign n16452 = n9736 & ~n16451;
  assign n16453 = ~n6197 & n15765;
  assign n16454 = n9036 & n15768;
  assign n16455 = pi0148 & ~n16453;
  assign n16456 = ~n16454 & n16455;
  assign n16457 = ~pi0051 & n15294;
  assign n16458 = ~pi0148 & ~n16457;
  assign n16459 = ~n16416 & ~n16458;
  assign n16460 = ~pi0148 & n14596;
  assign n16461 = ~n16459 & ~n16460;
  assign n16462 = ~n16456 & ~n16461;
  assign n16463 = pi0299 & ~n16462;
  assign n16464 = ~n16449 & ~n16452;
  assign n16465 = ~n16463 & n16464;
  assign n16466 = pi0232 & ~n16465;
  assign n16467 = ~pi0100 & n15754;
  assign n16468 = ~n16466 & n16467;
  assign n16469 = ~n16446 & ~n16468;
  assign n16470 = n2535 & ~n16469;
  assign n16471 = ~n16392 & ~n16444;
  assign n16472 = ~n16470 & n16471;
  assign n16473 = ~po1038 & ~n16472;
  assign n16474 = ~n16443 & n16473;
  assign po0293 = n16397 | n16474;
  assign n16476 = ~pi0039 & pi0137;
  assign n16477 = n10368 & n14873;
  assign n16478 = n6168 & n11568;
  assign n16479 = ~pi0299 & ~po1038;
  assign n16480 = ~pi0198 & n11579;
  assign n16481 = n16479 & n16480;
  assign n16482 = ~n16478 & ~n16481;
  assign n16483 = ~n16477 & ~n16482;
  assign n16484 = ~pi0210 & n11568;
  assign n16485 = po1038 & n16484;
  assign n16486 = ~n16483 & ~n16485;
  assign n16487 = n10478 & ~n16486;
  assign po0294 = n16476 | n16487;
  assign n16489 = ~n9739 & n13910;
  assign n16490 = ~pi0039 & ~n16489;
  assign n16491 = ~pi0232 & ~n11481;
  assign n16492 = n6198 & n6396;
  assign n16493 = n9051 & n16492;
  assign n16494 = n9736 & ~n16493;
  assign n16495 = ~n6198 & n9737;
  assign n16496 = ~n9736 & ~n11481;
  assign n16497 = ~n16494 & ~n16495;
  assign n16498 = ~n16496 & n16497;
  assign n16499 = pi0232 & ~n16498;
  assign n16500 = ~n16491 & ~n16499;
  assign n16501 = pi0039 & ~n16500;
  assign n16502 = n10200 & ~n16490;
  assign n16503 = ~n16501 & n16502;
  assign n16504 = ~pi0138 & n16503;
  assign n16505 = n9250 & ~n9282;
  assign n16506 = pi0092 & ~n16505;
  assign n16507 = n2532 & ~n16506;
  assign n16508 = ~pi0075 & ~n9288;
  assign n16509 = ~n9326 & ~n11892;
  assign n16510 = n9337 & ~n16509;
  assign n16511 = n13815 & ~n16510;
  assign n16512 = ~n6242 & ~n9326;
  assign n16513 = n9036 & ~n16509;
  assign n16514 = ~n16512 & n16513;
  assign n16515 = n9291 & ~n16514;
  assign n16516 = ~n16511 & ~n16515;
  assign n16517 = ~pi0232 & ~n16516;
  assign n16518 = ~pi0141 & n16511;
  assign n16519 = ~n9305 & n16510;
  assign n16520 = n13815 & ~n16519;
  assign n16521 = pi0141 & n16520;
  assign n16522 = ~n9300 & ~n16509;
  assign n16523 = ~n9290 & ~n16522;
  assign n16524 = pi0148 & ~n16523;
  assign n16525 = ~n9737 & ~n16515;
  assign n16526 = ~n16524 & ~n16525;
  assign n16527 = ~n16518 & ~n16521;
  assign n16528 = ~n16526 & n16527;
  assign n16529 = pi0232 & ~n16528;
  assign n16530 = ~n16517 & ~n16529;
  assign n16531 = pi0039 & ~n16530;
  assign n16532 = pi0299 & ~n9605;
  assign n16533 = ~pi0299 & ~n9949;
  assign n16534 = ~pi0232 & ~n16532;
  assign n16535 = ~n16533 & n16534;
  assign n16536 = ~pi0039 & ~n16535;
  assign n16537 = ~n6197 & ~n9949;
  assign n16538 = ~n13772 & ~n16537;
  assign n16539 = ~pi0299 & ~n16538;
  assign n16540 = pi0141 & n16539;
  assign n16541 = pi0148 & n6197;
  assign n16542 = ~n9605 & ~n16541;
  assign n16543 = pi0148 & n13737;
  assign n16544 = ~n16542 & ~n16543;
  assign n16545 = pi0299 & ~n16544;
  assign n16546 = ~pi0141 & n16533;
  assign n16547 = pi0232 & ~n16546;
  assign n16548 = ~n16540 & n16547;
  assign n16549 = ~n16545 & n16548;
  assign n16550 = n16536 & ~n16549;
  assign n16551 = n2608 & ~n16531;
  assign n16552 = ~n16550 & n16551;
  assign n16553 = ~pi0087 & ~n16552;
  assign n16554 = n16508 & ~n16553;
  assign n16555 = ~pi0092 & ~n16554;
  assign n16556 = n16507 & ~n16555;
  assign n16557 = ~pi0055 & ~n16556;
  assign n16558 = n9251 & ~n13686;
  assign n16559 = pi0055 & ~n16558;
  assign n16560 = ~n16557 & ~n16559;
  assign n16561 = n2529 & ~n16560;
  assign n16562 = n9883 & ~n16561;
  assign n16563 = pi0138 & n16562;
  assign n16564 = ~pi0118 & n13664;
  assign n16565 = ~pi0139 & n16564;
  assign n16566 = ~n16504 & ~n16565;
  assign n16567 = ~n16563 & n16566;
  assign n16568 = ~pi0138 & ~n8974;
  assign n16569 = n16503 & ~n16568;
  assign n16570 = n16562 & n16568;
  assign n16571 = n16565 & ~n16569;
  assign n16572 = ~n16570 & n16571;
  assign po0295 = ~n16567 & ~n16572;
  assign n16574 = n13910 & ~n15738;
  assign n16575 = ~pi0039 & ~n16574;
  assign n16576 = ~n11477 & n15755;
  assign n16577 = ~n6198 & n9021;
  assign n16578 = n9020 & ~n16493;
  assign n16579 = ~n11480 & ~n16577;
  assign n16580 = ~n16576 & ~n16578;
  assign n16581 = n16579 & n16580;
  assign n16582 = pi0232 & ~n16581;
  assign n16583 = ~n16491 & ~n16582;
  assign n16584 = pi0039 & ~n16583;
  assign n16585 = n10200 & ~n16575;
  assign n16586 = ~n16584 & n16585;
  assign n16587 = ~pi0139 & n16586;
  assign n16588 = ~pi0169 & n9326;
  assign n16589 = ~n16522 & ~n16588;
  assign n16590 = n9036 & ~n16589;
  assign n16591 = n9291 & ~n16590;
  assign n16592 = ~pi0191 & n16511;
  assign n16593 = pi0191 & n16520;
  assign n16594 = ~n16591 & ~n16592;
  assign n16595 = ~n16593 & n16594;
  assign n16596 = pi0232 & ~n16595;
  assign n16597 = ~n16517 & ~n16596;
  assign n16598 = pi0039 & ~n16597;
  assign n16599 = pi0191 & n16539;
  assign n16600 = ~n9605 & ~n15764;
  assign n16601 = pi0169 & n13737;
  assign n16602 = ~n16600 & ~n16601;
  assign n16603 = pi0299 & ~n16602;
  assign n16604 = ~pi0191 & n16533;
  assign n16605 = pi0232 & ~n16604;
  assign n16606 = ~n16599 & n16605;
  assign n16607 = ~n16603 & n16606;
  assign n16608 = n16536 & ~n16607;
  assign n16609 = n2608 & ~n16598;
  assign n16610 = ~n16608 & n16609;
  assign n16611 = ~pi0087 & ~n16610;
  assign n16612 = n16508 & ~n16611;
  assign n16613 = ~pi0092 & ~n16612;
  assign n16614 = n16507 & ~n16613;
  assign n16615 = ~pi0055 & ~n16614;
  assign n16616 = ~n16559 & ~n16615;
  assign n16617 = n2529 & ~n16616;
  assign n16618 = n9883 & ~n16617;
  assign n16619 = pi0139 & n16618;
  assign n16620 = ~n16564 & ~n16587;
  assign n16621 = ~n16619 & n16620;
  assign n16622 = ~pi0139 & ~n8975;
  assign n16623 = n16586 & ~n16622;
  assign n16624 = n16618 & n16622;
  assign n16625 = n16564 & ~n16623;
  assign n16626 = ~n16624 & n16625;
  assign po0296 = ~n16621 & ~n16626;
  assign n16628 = ~pi0641 & pi1158;
  assign n16629 = pi0641 & ~pi1158;
  assign n16630 = ~n16628 & ~n16629;
  assign n16631 = pi0788 & ~n16630;
  assign n16632 = ~pi0648 & pi1159;
  assign n16633 = pi0648 & ~pi1159;
  assign n16634 = ~n16632 & ~n16633;
  assign n16635 = pi0789 & ~n16634;
  assign n16636 = pi0627 & pi1154;
  assign n16637 = ~pi0627 & ~pi1154;
  assign n16638 = pi0781 & ~n16636;
  assign n16639 = ~n16637 & n16638;
  assign n16640 = pi0140 & ~n2571;
  assign n16641 = n2926 & n6284;
  assign n16642 = ~pi0140 & ~n16641;
  assign n16643 = pi0665 & pi1091;
  assign n16644 = pi0680 & ~n16643;
  assign n16645 = n2926 & n16644;
  assign n16646 = n6284 & n16645;
  assign n16647 = pi0038 & ~n16646;
  assign n16648 = ~n16642 & n16647;
  assign n16649 = ~n6184 & n6380;
  assign n16650 = ~pi0120 & ~n16649;
  assign n16651 = pi0120 & ~n2521;
  assign n16652 = ~n16650 & ~n16651;
  assign n16653 = n2926 & n16652;
  assign n16654 = n2603 & n16653;
  assign n16655 = n16644 & n16654;
  assign n16656 = ~pi0661 & ~pi0681;
  assign n16657 = ~pi0662 & n16656;
  assign n16658 = ~n16643 & n16653;
  assign n16659 = ~n6192 & n16658;
  assign n16660 = ~pi0824 & ~n16649;
  assign n16661 = n6380 & ~n10204;
  assign n16662 = pi1092 & n16661;
  assign n16663 = ~n11031 & ~n16662;
  assign n16664 = ~n16660 & ~n16663;
  assign n16665 = pi1093 & n16664;
  assign n16666 = ~pi0120 & ~n16665;
  assign n16667 = n2521 & n2926;
  assign n16668 = pi0120 & ~n16667;
  assign n16669 = ~pi1091 & ~n16668;
  assign n16670 = ~n16666 & n16669;
  assign n16671 = n2926 & n16649;
  assign n16672 = n2923 & n16671;
  assign n16673 = pi0829 & ~n16662;
  assign n16674 = ~pi0829 & ~n16664;
  assign n16675 = n7517 & ~n16673;
  assign n16676 = ~n16674 & n16675;
  assign n16677 = ~n16672 & ~n16676;
  assign n16678 = pi1091 & ~n16677;
  assign n16679 = ~pi0120 & ~n16678;
  assign n16680 = ~n16668 & ~n16679;
  assign n16681 = ~n16670 & ~n16680;
  assign n16682 = ~n6197 & n16681;
  assign n16683 = n6197 & ~n16653;
  assign n16684 = ~n16682 & ~n16683;
  assign n16685 = pi0665 & ~n16670;
  assign n16686 = ~n16681 & ~n16685;
  assign n16687 = ~n16658 & ~n16686;
  assign n16688 = n16684 & ~n16687;
  assign n16689 = n6192 & n16688;
  assign n16690 = ~n16659 & ~n16689;
  assign n16691 = ~n16657 & n16690;
  assign n16692 = n16657 & ~n16688;
  assign n16693 = pi0680 & ~n16692;
  assign n16694 = ~n16691 & n16693;
  assign n16695 = n6205 & ~n16694;
  assign n16696 = n6195 & n16686;
  assign n16697 = n6197 & ~n16681;
  assign n16698 = ~n6197 & n16653;
  assign n16699 = ~n16697 & ~n16698;
  assign n16700 = ~n6192 & n16699;
  assign n16701 = n6192 & n16681;
  assign n16702 = ~n16700 & ~n16701;
  assign n16703 = n16644 & n16702;
  assign n16704 = ~n16657 & n16703;
  assign n16705 = ~n16696 & ~n16704;
  assign n16706 = ~n6205 & n16705;
  assign n16707 = ~n2603 & ~n16695;
  assign n16708 = ~n16706 & n16707;
  assign n16709 = ~n16655 & ~n16708;
  assign n16710 = ~pi0223 & ~n16709;
  assign n16711 = n6187 & n14205;
  assign n16712 = n16667 & ~n16711;
  assign n16713 = pi0120 & ~n16712;
  assign n16714 = ~pi0120 & ~n16671;
  assign n16715 = pi1091 & ~n16713;
  assign n16716 = ~n16714 & n16715;
  assign n16717 = pi0120 & pi0824;
  assign n16718 = n6187 & n16717;
  assign n16719 = n16669 & ~n16718;
  assign n16720 = ~n16714 & n16719;
  assign n16721 = ~n16716 & ~n16720;
  assign n16722 = n6197 & ~n16721;
  assign n16723 = ~n16698 & ~n16722;
  assign n16724 = ~n6205 & n16723;
  assign n16725 = ~n6197 & n16721;
  assign n16726 = n16658 & ~n16725;
  assign n16727 = ~n16659 & ~n16726;
  assign n16728 = pi0680 & ~n16727;
  assign n16729 = ~n16724 & n16728;
  assign n16730 = n16657 & ~n16726;
  assign n16731 = pi0223 & ~n16730;
  assign n16732 = n16729 & n16731;
  assign n16733 = ~n16710 & ~n16732;
  assign n16734 = ~pi0299 & ~n16733;
  assign n16735 = ~n6242 & n16705;
  assign n16736 = n6242 & ~n16694;
  assign n16737 = ~n3448 & ~n16735;
  assign n16738 = ~n16736 & n16737;
  assign n16739 = n16644 & n16653;
  assign n16740 = n3448 & n16739;
  assign n16741 = ~n16738 & ~n16740;
  assign n16742 = ~pi0215 & ~n16741;
  assign n16743 = ~n6242 & n16723;
  assign n16744 = n16728 & ~n16743;
  assign n16745 = pi0215 & ~n16730;
  assign n16746 = n16744 & n16745;
  assign n16747 = ~n16742 & ~n16746;
  assign n16748 = pi0299 & ~n16747;
  assign n16749 = ~n16734 & ~n16748;
  assign n16750 = pi0140 & ~n16749;
  assign n16751 = pi0039 & pi0140;
  assign n16752 = ~n16644 & n16654;
  assign n16753 = ~pi0680 & ~n16702;
  assign n16754 = n16643 & n16680;
  assign n16755 = ~n6226 & n16754;
  assign n16756 = n16643 & n16698;
  assign n16757 = ~n6192 & n16756;
  assign n16758 = ~n16755 & ~n16757;
  assign n16759 = ~n16657 & ~n16758;
  assign n16760 = n16657 & n16754;
  assign n16761 = pi0680 & ~n16760;
  assign n16762 = ~n16759 & n16761;
  assign n16763 = ~n16753 & ~n16762;
  assign n16764 = ~n6205 & ~n16763;
  assign n16765 = pi0616 & ~n16653;
  assign n16766 = pi0614 & ~n16653;
  assign n16767 = ~pi0603 & ~n16653;
  assign n16768 = pi0603 & ~n16684;
  assign n16769 = ~n16767 & ~n16768;
  assign n16770 = ~pi0642 & ~n16769;
  assign n16771 = ~n6190 & ~n16653;
  assign n16772 = ~n16770 & ~n16771;
  assign n16773 = ~pi0614 & ~n16772;
  assign n16774 = ~n16766 & ~n16773;
  assign n16775 = ~pi0616 & ~n16774;
  assign n16776 = ~n16765 & ~n16775;
  assign n16777 = ~pi0680 & ~n16776;
  assign n16778 = n16643 & n16653;
  assign n16779 = n6197 & ~n16778;
  assign n16780 = ~n6197 & ~n16754;
  assign n16781 = ~n16779 & ~n16780;
  assign n16782 = n6192 & n16781;
  assign n16783 = ~n6192 & n16778;
  assign n16784 = pi0680 & ~n16783;
  assign n16785 = ~n16782 & n16784;
  assign n16786 = ~n16777 & ~n16785;
  assign n16787 = ~n16657 & n16786;
  assign n16788 = pi0680 & ~n16781;
  assign n16789 = n16657 & ~n16788;
  assign n16790 = ~n16777 & n16789;
  assign n16791 = ~n16787 & ~n16790;
  assign n16792 = n6205 & n16791;
  assign n16793 = ~n2603 & ~n16764;
  assign n16794 = ~n16792 & n16793;
  assign n16795 = ~pi0223 & ~n16752;
  assign n16796 = ~n16794 & n16795;
  assign n16797 = ~n16683 & ~n16725;
  assign n16798 = n6190 & ~n16797;
  assign n16799 = ~n16771 & ~n16798;
  assign n16800 = ~pi0614 & ~n16799;
  assign n16801 = ~n16766 & ~n16800;
  assign n16802 = ~pi0616 & ~n16801;
  assign n16803 = ~n16765 & ~n16802;
  assign n16804 = ~pi0680 & ~n16803;
  assign n16805 = pi0665 & n16716;
  assign n16806 = ~n6197 & ~n16805;
  assign n16807 = ~n16779 & ~n16806;
  assign n16808 = n6195 & ~n16807;
  assign n16809 = n16784 & ~n16807;
  assign n16810 = ~n16808 & ~n16809;
  assign n16811 = ~n16804 & n16810;
  assign n16812 = n6205 & n16811;
  assign n16813 = ~pi0616 & n16800;
  assign n16814 = ~n16723 & ~n16813;
  assign n16815 = ~pi0680 & ~n16814;
  assign n16816 = pi0680 & ~n16805;
  assign n16817 = ~n16757 & n16816;
  assign n16818 = ~n16815 & ~n16817;
  assign n16819 = n16810 & n16818;
  assign n16820 = ~n6205 & n16819;
  assign n16821 = pi0223 & ~n16812;
  assign n16822 = ~n16820 & n16821;
  assign n16823 = ~n16796 & ~n16822;
  assign n16824 = ~pi0299 & ~n16823;
  assign n16825 = n3448 & n16652;
  assign n16826 = n2926 & ~n16644;
  assign n16827 = n16825 & n16826;
  assign n16828 = ~n6242 & ~n16763;
  assign n16829 = n6242 & n16791;
  assign n16830 = ~n3448 & ~n16828;
  assign n16831 = ~n16829 & n16830;
  assign n16832 = ~pi0215 & ~n16827;
  assign n16833 = ~n16831 & n16832;
  assign n16834 = n6242 & n16811;
  assign n16835 = ~n6242 & n16819;
  assign n16836 = pi0215 & ~n16834;
  assign n16837 = ~n16835 & n16836;
  assign n16838 = ~n16833 & ~n16837;
  assign n16839 = pi0299 & ~n16838;
  assign n16840 = ~n16824 & ~n16839;
  assign n16841 = pi0039 & n16840;
  assign n16842 = ~n16751 & ~n16841;
  assign n16843 = ~n16750 & ~n16842;
  assign n16844 = ~pi0102 & ~n11299;
  assign n16845 = ~pi0098 & ~n2787;
  assign n16846 = ~n16844 & n16845;
  assign n16847 = n7438 & n12375;
  assign n16848 = n16846 & n16847;
  assign n16849 = n8897 & n9141;
  assign n16850 = n16848 & n16849;
  assign n16851 = ~pi0040 & ~n16850;
  assign n16852 = n10289 & ~n16851;
  assign n16853 = ~pi0252 & ~n16852;
  assign n16854 = n2763 & n2938;
  assign n16855 = n8896 & n16848;
  assign n16856 = ~pi0047 & ~n16855;
  assign n16857 = pi0314 & n10241;
  assign n16858 = n16856 & ~n16857;
  assign n16859 = n16854 & ~n16858;
  assign n16860 = ~pi0035 & ~n16859;
  assign n16861 = ~pi0040 & n10274;
  assign n16862 = ~n16860 & n16861;
  assign n16863 = pi0252 & ~n2743;
  assign n16864 = ~n16862 & n16863;
  assign n16865 = ~n16853 & ~n16864;
  assign n16866 = n2518 & n16865;
  assign n16867 = pi1092 & ~n12373;
  assign n16868 = n16866 & n16867;
  assign n16869 = ~pi0088 & ~n16846;
  assign n16870 = n11020 & ~n16869;
  assign n16871 = ~pi0252 & n9500;
  assign n16872 = n16870 & n16871;
  assign n16873 = n2500 & n16870;
  assign n16874 = ~pi0047 & ~n16857;
  assign n16875 = ~n16873 & n16874;
  assign n16876 = n16854 & ~n16875;
  assign n16877 = ~pi0035 & ~n16876;
  assign n16878 = pi0252 & n10274;
  assign n16879 = ~n16877 & n16878;
  assign n16880 = ~pi0040 & ~n16872;
  assign n16881 = ~n16879 & n16880;
  assign n16882 = n7417 & n10289;
  assign n16883 = ~n16881 & n16882;
  assign n16884 = ~n16868 & ~n16883;
  assign n16885 = pi1093 & ~n16884;
  assign n16886 = ~n2923 & ~n16885;
  assign n16887 = pi1092 & n2930;
  assign po1106 = n2923 & n16887;
  assign n16889 = n16866 & po1106;
  assign n16890 = ~n2924 & ~n16889;
  assign n16891 = ~n16886 & ~n16890;
  assign n16892 = ~pi1091 & n16885;
  assign n16893 = ~n16891 & ~n16892;
  assign n16894 = pi0665 & ~n16892;
  assign n16895 = ~n16893 & ~n16894;
  assign n16896 = ~pi0198 & ~n16895;
  assign n16897 = ~n3411 & ~n16881;
  assign n16898 = ~pi0032 & ~n16897;
  assign n16899 = pi0032 & ~n6485;
  assign n16900 = ~pi0095 & n2932;
  assign n16901 = ~n16899 & n16900;
  assign n16902 = ~n16898 & n16901;
  assign n16903 = pi0824 & n16902;
  assign n16904 = ~n16868 & ~n16903;
  assign n16905 = n7626 & ~n16904;
  assign n16906 = ~pi0032 & ~n16865;
  assign n16907 = n16901 & ~n16906;
  assign n16908 = ~pi0824 & pi0829;
  assign n16909 = n16907 & n16908;
  assign n16910 = n16904 & ~n16909;
  assign n16911 = pi1093 & ~n16910;
  assign n16912 = ~n2923 & ~n16911;
  assign n16913 = ~n16890 & ~n16912;
  assign n16914 = ~n16905 & ~n16913;
  assign n16915 = pi0665 & ~n16905;
  assign n16916 = ~n16914 & ~n16915;
  assign n16917 = pi0198 & ~n16916;
  assign n16918 = ~n16896 & ~n16917;
  assign n16919 = pi0680 & n16918;
  assign n16920 = ~pi0299 & ~n16919;
  assign n16921 = pi0210 & ~n16916;
  assign n16922 = ~pi0210 & ~n16895;
  assign n16923 = ~n16921 & ~n16922;
  assign n16924 = pi0680 & n16923;
  assign n16925 = pi0299 & ~n16924;
  assign n16926 = ~n16920 & ~n16925;
  assign n16927 = pi0140 & n16926;
  assign n16928 = ~pi0198 & n16893;
  assign n16929 = pi0198 & n16914;
  assign n16930 = ~n16928 & ~n16929;
  assign n16931 = pi0665 & n16913;
  assign n16932 = pi0198 & ~n16931;
  assign n16933 = pi0665 & n16891;
  assign n16934 = ~pi0198 & ~n16933;
  assign n16935 = ~n16932 & ~n16934;
  assign n16936 = pi0680 & ~n16935;
  assign n16937 = n16930 & ~n16936;
  assign n16938 = ~pi0299 & ~n16937;
  assign n16939 = ~pi0210 & n16893;
  assign n16940 = pi0210 & n16914;
  assign n16941 = ~n16939 & ~n16940;
  assign n16942 = ~pi0210 & ~n16933;
  assign n16943 = pi0210 & ~n16931;
  assign n16944 = ~n16942 & ~n16943;
  assign n16945 = pi0680 & ~n16944;
  assign n16946 = n16941 & ~n16945;
  assign n16947 = pi0299 & ~n16946;
  assign n16948 = ~n16938 & ~n16947;
  assign n16949 = ~pi0140 & ~n16948;
  assign n16950 = ~pi0039 & ~n16927;
  assign n16951 = ~n16949 & n16950;
  assign n16952 = ~n16843 & ~n16951;
  assign n16953 = ~pi0038 & ~n16952;
  assign n16954 = ~pi0738 & ~n16648;
  assign n16955 = ~n16953 & n16954;
  assign n16956 = pi0299 & ~n16941;
  assign n16957 = ~pi0299 & ~n16930;
  assign n16958 = ~n16956 & ~n16957;
  assign n16959 = ~pi0039 & ~n16958;
  assign n16960 = pi0681 & ~n16814;
  assign n16961 = pi0661 & n16814;
  assign n16962 = ~n6193 & ~n16803;
  assign n16963 = n6193 & n16721;
  assign n16964 = ~n6197 & ~n16963;
  assign n16965 = ~n16962 & n16964;
  assign n16966 = ~n16722 & ~n16965;
  assign n16967 = ~pi0661 & ~n16966;
  assign n16968 = ~pi0681 & ~n16961;
  assign n16969 = ~n16967 & n16968;
  assign n16970 = ~n16960 & ~n16969;
  assign n16971 = ~n6205 & ~n16970;
  assign n16972 = pi0681 & ~n16803;
  assign n16973 = pi0680 & ~n16797;
  assign n16974 = ~pi0680 & ~n16653;
  assign n16975 = pi0616 & n16657;
  assign n16976 = ~n16974 & n16975;
  assign n16977 = ~n16973 & n16976;
  assign n16978 = pi0616 & n16653;
  assign n16979 = ~n16657 & n16978;
  assign n16980 = ~n16977 & ~n16979;
  assign n16981 = ~pi0616 & ~n16657;
  assign n16982 = n16801 & n16981;
  assign n16983 = ~pi0680 & n16802;
  assign n16984 = ~pi0616 & n16657;
  assign n16985 = ~n16973 & n16984;
  assign n16986 = ~n16983 & n16985;
  assign n16987 = ~n16982 & ~n16986;
  assign n16988 = ~pi0681 & n16980;
  assign n16989 = n16987 & n16988;
  assign n16990 = ~n16972 & ~n16989;
  assign n16991 = n6205 & ~n16990;
  assign n16992 = ~n16971 & ~n16991;
  assign n16993 = pi0223 & ~n16992;
  assign n16994 = pi0681 & ~n16776;
  assign n16995 = pi0680 & ~n16684;
  assign n16996 = pi0614 & n16657;
  assign n16997 = ~n16974 & n16996;
  assign n16998 = ~n16995 & n16997;
  assign n16999 = pi0614 & n16653;
  assign n17000 = ~n16657 & n16999;
  assign n17001 = ~n16998 & ~n17000;
  assign n17002 = ~pi0614 & ~n6195;
  assign n17003 = ~pi0616 & ~n16772;
  assign n17004 = ~n16765 & n17002;
  assign n17005 = ~n17003 & n17004;
  assign n17006 = ~pi0614 & n6195;
  assign n17007 = n16684 & n17006;
  assign n17008 = ~n17005 & ~n17007;
  assign n17009 = ~pi0681 & n17001;
  assign n17010 = n17008 & n17009;
  assign n17011 = ~n16994 & ~n17010;
  assign n17012 = n6205 & ~n17011;
  assign n17013 = pi0681 & ~n16702;
  assign n17014 = n6194 & ~n16681;
  assign n17015 = ~n6194 & n16702;
  assign n17016 = ~pi0681 & ~n17014;
  assign n17017 = ~n17015 & n17016;
  assign n17018 = ~n17013 & ~n17017;
  assign n17019 = ~n6205 & ~n17018;
  assign n17020 = ~n17012 & ~n17019;
  assign n17021 = ~n2603 & n17020;
  assign n17022 = ~pi0223 & ~n16654;
  assign n17023 = ~n17021 & n17022;
  assign n17024 = ~n16993 & ~n17023;
  assign n17025 = ~pi0299 & ~n17024;
  assign n17026 = n3448 & n16653;
  assign n17027 = n6241 & ~n17011;
  assign n17028 = ~n6241 & ~n17018;
  assign n17029 = n6236 & ~n17028;
  assign n17030 = ~n17027 & n17029;
  assign n17031 = ~n3448 & n17030;
  assign n17032 = ~n6236 & n17018;
  assign n17033 = ~n3448 & n17032;
  assign n17034 = ~pi0215 & ~n17026;
  assign n17035 = ~n17033 & n17034;
  assign n17036 = ~n17031 & n17035;
  assign n17037 = ~n6236 & n16970;
  assign n17038 = ~n6241 & ~n16970;
  assign n17039 = n6241 & ~n16990;
  assign n17040 = n6236 & ~n17039;
  assign n17041 = ~n17038 & n17040;
  assign n17042 = ~n17037 & ~n17041;
  assign n17043 = pi0215 & n17042;
  assign n17044 = ~n17036 & ~n17043;
  assign n17045 = pi0299 & ~n17044;
  assign n17046 = ~n17025 & ~n17045;
  assign n17047 = pi0039 & ~n17046;
  assign n17048 = ~n16959 & ~n17047;
  assign n17049 = ~pi0038 & ~n17048;
  assign n17050 = n2926 & n6135;
  assign n17051 = pi0038 & ~n17050;
  assign n17052 = ~n17049 & ~n17051;
  assign n17053 = ~pi0140 & pi0738;
  assign n17054 = ~n17052 & n17053;
  assign n17055 = n2571 & ~n17054;
  assign n17056 = ~n16955 & n17055;
  assign n17057 = ~n16640 & ~n17056;
  assign n17058 = ~pi0778 & ~n17057;
  assign n17059 = n2571 & n17052;
  assign n17060 = ~pi0140 & ~n17059;
  assign n17061 = ~pi0625 & n17060;
  assign n17062 = pi0625 & n17057;
  assign n17063 = pi1153 & ~n17061;
  assign n17064 = ~n17062 & n17063;
  assign n17065 = ~pi0625 & n17057;
  assign n17066 = pi0625 & n17060;
  assign n17067 = ~pi1153 & ~n17066;
  assign n17068 = ~n17065 & n17067;
  assign n17069 = ~n17064 & ~n17068;
  assign n17070 = pi0778 & ~n17069;
  assign n17071 = ~n17058 & ~n17070;
  assign n17072 = pi0660 & pi1155;
  assign n17073 = ~pi0660 & ~pi1155;
  assign n17074 = pi0785 & ~n17072;
  assign n17075 = ~n17073 & n17074;
  assign n17076 = ~n17071 & ~n17075;
  assign n17077 = ~n17060 & n17075;
  assign n17078 = ~n17076 & ~n17077;
  assign n17079 = ~n16639 & n17078;
  assign n17080 = n16639 & n17060;
  assign n17081 = ~n17079 & ~n17080;
  assign n17082 = ~n16635 & n17081;
  assign n17083 = n16635 & ~n17060;
  assign n17084 = ~n17082 & ~n17083;
  assign n17085 = ~n16631 & n17084;
  assign n17086 = n16631 & n17060;
  assign n17087 = ~n17085 & ~n17086;
  assign n17088 = ~pi0792 & n17087;
  assign n17089 = ~pi0628 & n17060;
  assign n17090 = pi0628 & ~n17087;
  assign n17091 = pi1156 & ~n17089;
  assign n17092 = ~n17090 & n17091;
  assign n17093 = pi0628 & n17060;
  assign n17094 = ~pi0628 & ~n17087;
  assign n17095 = ~pi1156 & ~n17093;
  assign n17096 = ~n17094 & n17095;
  assign n17097 = ~n17092 & ~n17096;
  assign n17098 = pi0792 & ~n17097;
  assign n17099 = ~n17088 & ~n17098;
  assign n17100 = ~pi0787 & ~n17099;
  assign n17101 = ~pi0647 & n17060;
  assign n17102 = pi0647 & n17099;
  assign n17103 = pi1157 & ~n17101;
  assign n17104 = ~n17102 & n17103;
  assign n17105 = ~pi0647 & n17099;
  assign n17106 = pi0647 & n17060;
  assign n17107 = ~pi1157 & ~n17106;
  assign n17108 = ~n17105 & n17107;
  assign n17109 = ~n17104 & ~n17108;
  assign n17110 = pi0787 & ~n17109;
  assign n17111 = ~n17100 & ~n17110;
  assign n17112 = ~pi0644 & n17111;
  assign n17113 = ~pi0619 & n17060;
  assign n17114 = ~pi0608 & pi1153;
  assign n17115 = pi0608 & ~pi1153;
  assign n17116 = ~n17114 & ~n17115;
  assign n17117 = pi0778 & ~n17116;
  assign n17118 = pi0621 & n16891;
  assign n17119 = ~pi0210 & ~n17118;
  assign n17120 = pi0621 & n16913;
  assign n17121 = pi0210 & ~n17120;
  assign n17122 = ~n17119 & ~n17121;
  assign n17123 = pi0603 & ~n17122;
  assign n17124 = n16941 & ~n17123;
  assign n17125 = pi0299 & ~n17124;
  assign n17126 = ~pi0198 & ~n17118;
  assign n17127 = pi0198 & ~n17120;
  assign n17128 = ~n17126 & ~n17127;
  assign n17129 = pi0621 & ~n16892;
  assign n17130 = ~n16893 & ~n17129;
  assign n17131 = ~pi0198 & n17130;
  assign n17132 = pi0621 & ~n16905;
  assign n17133 = ~n16914 & ~n17132;
  assign n17134 = pi0198 & n17133;
  assign n17135 = ~n17131 & ~n17134;
  assign n17136 = ~pi0603 & ~n17135;
  assign n17137 = ~n17128 & ~n17136;
  assign n17138 = ~pi0299 & n17137;
  assign n17139 = ~n17125 & ~n17138;
  assign n17140 = ~pi0039 & ~n17139;
  assign n17141 = ~n6195 & ~n16702;
  assign n17142 = n6195 & n16681;
  assign n17143 = ~n17141 & ~n17142;
  assign n17144 = pi0621 & pi1091;
  assign n17145 = n16680 & n17144;
  assign n17146 = pi0621 & ~n16670;
  assign n17147 = ~n16681 & ~n17146;
  assign n17148 = ~pi0603 & n17147;
  assign n17149 = ~pi0603 & n16699;
  assign n17150 = n6197 & n17145;
  assign n17151 = n16698 & n17144;
  assign n17152 = pi0603 & ~n17151;
  assign n17153 = ~n17150 & n17152;
  assign n17154 = ~n17149 & ~n17153;
  assign n17155 = ~n17145 & ~n17148;
  assign n17156 = ~n17154 & n17155;
  assign n17157 = n17143 & ~n17156;
  assign n17158 = ~n6242 & ~n17157;
  assign n17159 = n16653 & n17144;
  assign n17160 = n6197 & ~n17159;
  assign n17161 = ~n6197 & ~n17145;
  assign n17162 = ~n17160 & ~n17161;
  assign n17163 = pi0603 & ~n17162;
  assign n17164 = n16684 & ~n17163;
  assign n17165 = n6195 & ~n17164;
  assign n17166 = ~pi0614 & ~pi0642;
  assign n17167 = ~pi0616 & n17166;
  assign n17168 = pi0603 & ~n17144;
  assign n17169 = n16653 & ~n17168;
  assign n17170 = ~n17167 & n17169;
  assign n17171 = ~n16767 & n17167;
  assign n17172 = ~n17163 & n17171;
  assign n17173 = ~n17170 & ~n17172;
  assign n17174 = ~n6195 & n17173;
  assign n17175 = ~n17165 & ~n17174;
  assign n17176 = n6242 & ~n17175;
  assign n17177 = ~n3448 & ~n17158;
  assign n17178 = ~n17176 & n17177;
  assign n17179 = n3448 & n17169;
  assign n17180 = ~n17178 & ~n17179;
  assign n17181 = ~pi0215 & ~n17180;
  assign n17182 = n2926 & ~n17168;
  assign n17183 = ~n16723 & n17182;
  assign n17184 = n6192 & ~n16716;
  assign n17185 = n17183 & ~n17184;
  assign n17186 = ~n6195 & ~n17185;
  assign n17187 = ~n16721 & n17182;
  assign n17188 = n6195 & ~n17187;
  assign n17189 = ~n17186 & ~n17188;
  assign n17190 = ~n6242 & ~n17189;
  assign n17191 = pi0621 & n16716;
  assign n17192 = ~n6197 & ~n17191;
  assign n17193 = ~n17160 & ~n17192;
  assign n17194 = pi0603 & ~n17193;
  assign n17195 = n17171 & ~n17194;
  assign n17196 = ~n17170 & ~n17195;
  assign n17197 = ~n6195 & ~n17196;
  assign n17198 = n6195 & n16797;
  assign n17199 = ~n17194 & n17198;
  assign n17200 = ~n17197 & ~n17199;
  assign n17201 = n6242 & n17200;
  assign n17202 = pi0215 & ~n17190;
  assign n17203 = ~n17201 & n17202;
  assign n17204 = ~n17181 & ~n17203;
  assign n17205 = pi0299 & ~n17204;
  assign n17206 = ~n6205 & ~n17157;
  assign n17207 = n6205 & ~n17175;
  assign n17208 = ~n2603 & ~n17206;
  assign n17209 = ~n17207 & n17208;
  assign n17210 = n2603 & n17169;
  assign n17211 = ~n17209 & ~n17210;
  assign n17212 = ~pi0223 & ~n17211;
  assign n17213 = ~n6205 & ~n17189;
  assign n17214 = n6205 & n17200;
  assign n17215 = pi0223 & ~n17213;
  assign n17216 = ~n17214 & n17215;
  assign n17217 = ~n17212 & ~n17216;
  assign n17218 = ~pi0299 & ~n17217;
  assign n17219 = ~n17205 & ~n17218;
  assign n17220 = pi0039 & n17219;
  assign n17221 = ~n17140 & ~n17220;
  assign n17222 = ~pi0761 & n17221;
  assign n17223 = pi0761 & n17048;
  assign n17224 = ~pi0140 & ~n17222;
  assign n17225 = ~n17223 & n17224;
  assign n17226 = pi0603 & ~n17135;
  assign n17227 = ~pi0299 & ~n17226;
  assign n17228 = ~pi0210 & ~n17130;
  assign n17229 = pi0210 & ~n17133;
  assign n17230 = ~n17228 & ~n17229;
  assign n17231 = pi0603 & n17230;
  assign n17232 = pi0299 & ~n17231;
  assign n17233 = ~n17227 & ~n17232;
  assign n17234 = ~pi0039 & ~n17233;
  assign n17235 = n16653 & n17168;
  assign n17236 = ~n16725 & n17235;
  assign n17237 = ~n16723 & n17235;
  assign n17238 = n16725 & n17167;
  assign n17239 = n17237 & ~n17238;
  assign n17240 = ~n6195 & n17239;
  assign n17241 = ~n17236 & ~n17240;
  assign n17242 = ~n16743 & ~n17241;
  assign n17243 = pi0215 & ~n17242;
  assign n17244 = n2926 & n17168;
  assign n17245 = n16825 & n17244;
  assign n17246 = n16684 & n17168;
  assign n17247 = n6195 & n17246;
  assign n17248 = ~n17167 & n17235;
  assign n17249 = n17167 & n17246;
  assign n17250 = ~n17248 & ~n17249;
  assign n17251 = ~n6195 & ~n17250;
  assign n17252 = ~n17247 & ~n17251;
  assign n17253 = n6242 & n17252;
  assign n17254 = n17143 & n17168;
  assign n17255 = ~n6242 & ~n17254;
  assign n17256 = ~n3448 & ~n17253;
  assign n17257 = ~n17255 & n17256;
  assign n17258 = ~pi0215 & ~n17245;
  assign n17259 = ~n17257 & n17258;
  assign n17260 = pi0299 & ~n17243;
  assign n17261 = ~n17259 & n17260;
  assign n17262 = ~n16724 & ~n17241;
  assign n17263 = pi0223 & ~n17262;
  assign n17264 = n6205 & n17252;
  assign n17265 = ~n6205 & ~n17254;
  assign n17266 = ~n2603 & ~n17264;
  assign n17267 = ~n17265 & n17266;
  assign n17268 = n16654 & n17168;
  assign n17269 = ~pi0223 & ~n17268;
  assign n17270 = ~n17267 & n17269;
  assign n17271 = ~pi0299 & ~n17263;
  assign n17272 = ~n17270 & n17271;
  assign n17273 = ~n17261 & ~n17272;
  assign n17274 = pi0039 & n17273;
  assign n17275 = ~n17234 & ~n17274;
  assign n17276 = pi0140 & ~pi0761;
  assign n17277 = n17275 & n17276;
  assign n17278 = ~n17225 & ~n17277;
  assign n17279 = ~pi0038 & ~n17278;
  assign n17280 = n6284 & n17244;
  assign n17281 = ~pi0761 & n17280;
  assign n17282 = ~n16642 & ~n17281;
  assign n17283 = pi0038 & ~n17282;
  assign n17284 = ~n17279 & ~n17283;
  assign n17285 = n2571 & n17284;
  assign n17286 = ~n16640 & ~n17285;
  assign n17287 = ~n17117 & ~n17286;
  assign n17288 = ~n17060 & n17117;
  assign n17289 = ~n17287 & ~n17288;
  assign n17290 = ~pi0785 & ~n17289;
  assign n17291 = pi0609 & ~n17117;
  assign n17292 = ~n17060 & ~n17291;
  assign n17293 = pi0609 & n17287;
  assign n17294 = ~n17292 & ~n17293;
  assign n17295 = pi1155 & ~n17294;
  assign n17296 = ~pi0609 & ~n17117;
  assign n17297 = ~n17060 & ~n17296;
  assign n17298 = ~pi0609 & n17287;
  assign n17299 = ~n17297 & ~n17298;
  assign n17300 = ~pi1155 & ~n17299;
  assign n17301 = ~n17295 & ~n17300;
  assign n17302 = pi0785 & ~n17301;
  assign n17303 = ~n17290 & ~n17302;
  assign n17304 = ~pi0781 & ~n17303;
  assign n17305 = ~pi0618 & n17060;
  assign n17306 = pi0618 & n17303;
  assign n17307 = pi1154 & ~n17305;
  assign n17308 = ~n17306 & n17307;
  assign n17309 = ~pi0618 & n17303;
  assign n17310 = pi0618 & n17060;
  assign n17311 = ~pi1154 & ~n17310;
  assign n17312 = ~n17309 & n17311;
  assign n17313 = ~n17308 & ~n17312;
  assign n17314 = pi0781 & ~n17313;
  assign n17315 = ~n17304 & ~n17314;
  assign n17316 = pi0619 & n17315;
  assign n17317 = pi1159 & ~n17113;
  assign n17318 = ~n17316 & n17317;
  assign n17319 = pi0738 & ~n17284;
  assign n17320 = ~n16721 & n17235;
  assign n17321 = ~n16805 & ~n17320;
  assign n17322 = n6195 & n17321;
  assign n17323 = pi0680 & ~n16657;
  assign n17324 = ~n16756 & ~n16805;
  assign n17325 = ~n17237 & n17324;
  assign n17326 = ~n17167 & n17325;
  assign n17327 = ~pi0603 & n16756;
  assign n17328 = n17321 & ~n17327;
  assign n17329 = n17167 & n17328;
  assign n17330 = ~n17326 & ~n17329;
  assign n17331 = n17323 & ~n17330;
  assign n17332 = ~n17322 & ~n17331;
  assign n17333 = ~n16815 & n17332;
  assign n17334 = ~n6205 & ~n17333;
  assign n17335 = n16808 & ~n17236;
  assign n17336 = ~n16643 & ~n17168;
  assign n17337 = n16653 & ~n17336;
  assign n17338 = pi0616 & ~n17337;
  assign n17339 = pi0614 & ~n17337;
  assign n17340 = pi0642 & ~n17337;
  assign n17341 = ~pi0642 & ~n16807;
  assign n17342 = ~n17236 & n17341;
  assign n17343 = n17328 & n17342;
  assign n17344 = ~n17340 & ~n17343;
  assign n17345 = ~pi0614 & ~n17344;
  assign n17346 = ~n17339 & ~n17345;
  assign n17347 = ~pi0616 & ~n17346;
  assign n17348 = ~n17338 & ~n17347;
  assign n17349 = n17323 & ~n17348;
  assign n17350 = ~n16804 & ~n17335;
  assign n17351 = ~n17349 & n17350;
  assign n17352 = n6205 & ~n17351;
  assign n17353 = pi0223 & ~n17334;
  assign n17354 = ~n17352 & n17353;
  assign n17355 = pi0680 & n17336;
  assign n17356 = n16653 & ~n17355;
  assign n17357 = n2603 & ~n17356;
  assign n17358 = n16769 & ~n17336;
  assign n17359 = ~pi0642 & ~n17358;
  assign n17360 = ~n17340 & ~n17359;
  assign n17361 = ~pi0614 & ~n17360;
  assign n17362 = ~n17339 & ~n17361;
  assign n17363 = ~pi0616 & ~n17362;
  assign n17364 = ~n17338 & ~n17363;
  assign n17365 = n17323 & ~n17364;
  assign n17366 = ~pi0603 & ~n16781;
  assign n17367 = pi0603 & ~pi0665;
  assign n17368 = n17144 & n17367;
  assign n17369 = ~n16768 & ~n17368;
  assign n17370 = ~n17366 & n17369;
  assign n17371 = n6195 & ~n17370;
  assign n17372 = ~n16777 & ~n17371;
  assign n17373 = ~n17365 & n17372;
  assign n17374 = n6205 & n17373;
  assign n17375 = pi0603 & n17147;
  assign n17376 = pi0603 & ~pi0621;
  assign n17377 = n16754 & ~n17376;
  assign n17378 = n6195 & ~n17377;
  assign n17379 = ~n17375 & n17378;
  assign n17380 = n16702 & ~n17336;
  assign n17381 = n17323 & ~n17380;
  assign n17382 = ~n16753 & ~n17379;
  assign n17383 = ~n17381 & n17382;
  assign n17384 = ~n6205 & n17383;
  assign n17385 = ~n2603 & ~n17384;
  assign n17386 = ~n17374 & n17385;
  assign n17387 = ~pi0223 & ~n17357;
  assign n17388 = ~n17386 & n17387;
  assign n17389 = ~n17354 & ~n17388;
  assign n17390 = ~pi0299 & ~n17389;
  assign n17391 = n3448 & ~n17356;
  assign n17392 = ~n6242 & ~n17383;
  assign n17393 = n6242 & ~n17373;
  assign n17394 = ~n17392 & ~n17393;
  assign n17395 = ~n3448 & ~n17394;
  assign n17396 = ~pi0215 & ~n17391;
  assign n17397 = ~n17395 & n17396;
  assign n17398 = n6242 & ~n17351;
  assign n17399 = ~n6242 & ~n17333;
  assign n17400 = pi0215 & ~n17399;
  assign n17401 = ~n17398 & n17400;
  assign n17402 = ~n17397 & ~n17401;
  assign n17403 = pi0299 & ~n17402;
  assign n17404 = ~n17390 & ~n17403;
  assign n17405 = ~pi0140 & n17404;
  assign n17406 = n17026 & n17355;
  assign n17407 = ~n16643 & n17169;
  assign n17408 = pi0616 & ~n17407;
  assign n17409 = n17323 & ~n17408;
  assign n17410 = ~n17166 & n17407;
  assign n17411 = pi0603 & pi0665;
  assign n17412 = ~pi0603 & ~n16658;
  assign n17413 = ~n17411 & ~n17412;
  assign n17414 = ~n17163 & n17413;
  assign n17415 = n17166 & n17414;
  assign n17416 = ~pi0616 & ~n17410;
  assign n17417 = ~n17415 & n17416;
  assign n17418 = n17409 & ~n17417;
  assign n17419 = n16684 & n17371;
  assign n17420 = ~n17418 & ~n17419;
  assign n17421 = n6242 & n17420;
  assign n17422 = ~n16687 & n17154;
  assign n17423 = pi0616 & ~n17422;
  assign n17424 = ~pi0665 & n17145;
  assign n17425 = pi0603 & ~n17424;
  assign n17426 = ~n16687 & ~n16699;
  assign n17427 = ~pi0603 & ~n17426;
  assign n17428 = ~n17425 & ~n17427;
  assign n17429 = n17166 & n17428;
  assign n17430 = n17167 & ~n17428;
  assign n17431 = n17422 & ~n17430;
  assign n17432 = ~pi0616 & ~n17429;
  assign n17433 = ~n17431 & n17432;
  assign n17434 = ~n17423 & ~n17433;
  assign n17435 = ~n16657 & ~n17434;
  assign n17436 = n16696 & ~n17425;
  assign n17437 = ~n17323 & ~n17436;
  assign n17438 = ~n17435 & ~n17437;
  assign n17439 = ~n6242 & ~n17438;
  assign n17440 = ~n3448 & ~n17421;
  assign n17441 = ~n17439 & n17440;
  assign n17442 = ~pi0215 & ~n17406;
  assign n17443 = ~n17441 & n17442;
  assign n17444 = ~n16643 & ~n17196;
  assign n17445 = ~pi0616 & ~n17444;
  assign n17446 = n17409 & ~n17445;
  assign n17447 = n17199 & n17413;
  assign n17448 = ~n17446 & ~n17447;
  assign n17449 = n6242 & ~n17448;
  assign n17450 = n17183 & n17413;
  assign n17451 = pi0616 & ~n17450;
  assign n17452 = pi0614 & ~pi0616;
  assign n17453 = ~n17450 & n17452;
  assign n17454 = ~n17194 & n17413;
  assign n17455 = ~pi0642 & ~n17454;
  assign n17456 = n17450 & ~n17455;
  assign n17457 = n6191 & ~n17456;
  assign n17458 = ~n17453 & ~n17457;
  assign n17459 = ~n17451 & n17458;
  assign n17460 = ~n16657 & ~n17459;
  assign n17461 = ~n16721 & n17355;
  assign n17462 = ~n17323 & ~n17461;
  assign n17463 = ~n17460 & ~n17462;
  assign n17464 = ~n6242 & n17463;
  assign n17465 = pi0215 & ~n17449;
  assign n17466 = ~n17464 & n17465;
  assign n17467 = ~n17443 & ~n17466;
  assign n17468 = pi0299 & ~n17467;
  assign n17469 = n16645 & ~n17168;
  assign n17470 = ~n17244 & ~n17469;
  assign n17471 = n16653 & ~n17470;
  assign n17472 = n2603 & ~n17471;
  assign n17473 = ~n6205 & n17438;
  assign n17474 = n6205 & ~n17420;
  assign n17475 = ~n2603 & ~n17474;
  assign n17476 = ~n17473 & n17475;
  assign n17477 = n17269 & ~n17472;
  assign n17478 = ~n17476 & n17477;
  assign n17479 = n6205 & n17448;
  assign n17480 = ~n6205 & ~n17463;
  assign n17481 = pi0223 & ~n17479;
  assign n17482 = ~n17480 & n17481;
  assign n17483 = ~pi0299 & ~n17482;
  assign n17484 = ~n17478 & n17483;
  assign n17485 = ~n17468 & ~n17484;
  assign n17486 = pi0140 & n17485;
  assign n17487 = pi0761 & ~n17486;
  assign n17488 = ~n17405 & n17487;
  assign n17489 = ~n16644 & ~n17168;
  assign n17490 = n16667 & n17489;
  assign n17491 = ~n16650 & n17490;
  assign n17492 = n2603 & n17491;
  assign n17493 = n16643 & ~n17376;
  assign n17494 = ~n16758 & n17493;
  assign n17495 = n17323 & ~n17494;
  assign n17496 = n16702 & ~n17168;
  assign n17497 = ~pi0680 & ~n17496;
  assign n17498 = ~n17378 & ~n17495;
  assign n17499 = ~n17497 & n17498;
  assign n17500 = ~n6205 & n17499;
  assign n17501 = ~pi0680 & n17173;
  assign n17502 = n16781 & n17493;
  assign n17503 = n6195 & ~n17502;
  assign n17504 = n16778 & ~n17376;
  assign n17505 = ~n17167 & n17504;
  assign n17506 = n16643 & n17172;
  assign n17507 = n17323 & ~n17505;
  assign n17508 = ~n17506 & n17507;
  assign n17509 = ~n17501 & ~n17503;
  assign n17510 = ~n17508 & n17509;
  assign n17511 = n6205 & n17510;
  assign n17512 = ~n17500 & ~n17511;
  assign n17513 = ~n2603 & ~n17512;
  assign n17514 = ~pi0223 & ~n17492;
  assign n17515 = ~n17513 & n17514;
  assign n17516 = ~n16644 & n17197;
  assign n17517 = n6195 & ~n17376;
  assign n17518 = n16807 & n17517;
  assign n17519 = ~n17516 & ~n17518;
  assign n17520 = n6205 & ~n17519;
  assign n17521 = ~pi0680 & ~n17185;
  assign n17522 = ~n16816 & ~n17376;
  assign n17523 = n6195 & ~n17522;
  assign n17524 = ~n17196 & ~n17324;
  assign n17525 = n17323 & ~n17524;
  assign n17526 = ~n17521 & ~n17523;
  assign n17527 = ~n17525 & n17526;
  assign n17528 = ~n6205 & n17527;
  assign n17529 = pi0223 & ~n17520;
  assign n17530 = ~n17528 & n17529;
  assign n17531 = ~n17515 & ~n17530;
  assign n17532 = ~pi0299 & ~n17531;
  assign n17533 = n3448 & n17491;
  assign n17534 = ~n6242 & n17499;
  assign n17535 = n6242 & n17510;
  assign n17536 = ~n17534 & ~n17535;
  assign n17537 = ~n3448 & ~n17536;
  assign n17538 = ~pi0215 & ~n17533;
  assign n17539 = ~n17537 & n17538;
  assign n17540 = n6242 & ~n17519;
  assign n17541 = ~n6242 & n17527;
  assign n17542 = pi0215 & ~n17540;
  assign n17543 = ~n17541 & n17542;
  assign n17544 = ~n17539 & ~n17543;
  assign n17545 = pi0299 & ~n17544;
  assign n17546 = ~n17532 & ~n17545;
  assign n17547 = ~pi0140 & ~n17546;
  assign n17548 = n16653 & ~n17493;
  assign n17549 = ~n17167 & n17548;
  assign n17550 = n17323 & ~n17549;
  assign n17551 = n16727 & ~n17236;
  assign n17552 = n17167 & ~n17551;
  assign n17553 = n17550 & ~n17552;
  assign n17554 = pi0680 & ~n16730;
  assign n17555 = n17241 & ~n17554;
  assign n17556 = ~n17553 & ~n17555;
  assign n17557 = n6205 & ~n17556;
  assign n17558 = ~n17240 & ~n17320;
  assign n17559 = n16658 & ~n16723;
  assign n17560 = ~n16727 & n17554;
  assign n17561 = n17559 & n17560;
  assign n17562 = n17558 & ~n17561;
  assign n17563 = ~n6205 & n17562;
  assign n17564 = pi0223 & ~n17563;
  assign n17565 = ~n17557 & n17564;
  assign n17566 = ~pi0680 & n17250;
  assign n17567 = ~n17246 & ~n17414;
  assign n17568 = n17167 & ~n17567;
  assign n17569 = n17550 & ~n17568;
  assign n17570 = n6195 & ~n16688;
  assign n17571 = ~n17246 & n17570;
  assign n17572 = ~n17566 & ~n17571;
  assign n17573 = ~n17569 & n17572;
  assign n17574 = n6205 & n17573;
  assign n17575 = ~n17375 & ~n17428;
  assign n17576 = n17167 & ~n17575;
  assign n17577 = ~n16699 & n17168;
  assign n17578 = ~n17426 & ~n17577;
  assign n17579 = ~n17167 & ~n17578;
  assign n17580 = n17323 & ~n17579;
  assign n17581 = ~n17576 & n17580;
  assign n17582 = ~n16696 & ~n17323;
  assign n17583 = ~n17254 & n17582;
  assign n17584 = ~n17581 & ~n17583;
  assign n17585 = ~n6205 & n17584;
  assign n17586 = ~n2603 & ~n17574;
  assign n17587 = ~n17585 & n17586;
  assign n17588 = ~pi0223 & ~n17472;
  assign n17589 = ~n17587 & n17588;
  assign n17590 = ~pi0299 & ~n17565;
  assign n17591 = ~n17589 & n17590;
  assign n17592 = n3448 & n17471;
  assign n17593 = ~n6242 & n17584;
  assign n17594 = n6242 & n17573;
  assign n17595 = ~n17593 & ~n17594;
  assign n17596 = ~n3448 & ~n17595;
  assign n17597 = ~pi0215 & ~n17592;
  assign n17598 = ~n17596 & n17597;
  assign n17599 = ~n6242 & ~n17562;
  assign n17600 = n6242 & n17556;
  assign n17601 = pi0215 & ~n17599;
  assign n17602 = ~n17600 & n17601;
  assign n17603 = ~n17598 & ~n17602;
  assign n17604 = pi0299 & ~n17603;
  assign n17605 = ~n17591 & ~n17604;
  assign n17606 = pi0140 & n17605;
  assign n17607 = ~pi0761 & ~n17547;
  assign n17608 = ~n17606 & n17607;
  assign n17609 = ~n17488 & ~n17608;
  assign n17610 = pi0039 & ~n17609;
  assign n17611 = pi0680 & n17233;
  assign n17612 = ~n16948 & ~n17611;
  assign n17613 = ~pi0140 & ~n17612;
  assign n17614 = pi0603 & ~n17128;
  assign n17615 = ~pi0603 & ~n16918;
  assign n17616 = ~n17411 & ~n17614;
  assign n17617 = ~n17615 & n17616;
  assign n17618 = pi0680 & n17617;
  assign n17619 = ~pi0299 & ~n17618;
  assign n17620 = ~pi0603 & ~n16923;
  assign n17621 = ~n17123 & ~n17411;
  assign n17622 = ~n17620 & n17621;
  assign n17623 = pi0680 & n17622;
  assign n17624 = pi0299 & ~n17623;
  assign n17625 = ~n17619 & ~n17624;
  assign n17626 = pi0140 & ~n17625;
  assign n17627 = pi0761 & ~n17613;
  assign n17628 = ~n17626 & n17627;
  assign n17629 = n16948 & n17139;
  assign n17630 = ~pi0140 & n17629;
  assign n17631 = ~n16926 & ~n17233;
  assign n17632 = pi0140 & n17631;
  assign n17633 = ~pi0761 & ~n17632;
  assign n17634 = ~n17630 & n17633;
  assign n17635 = ~pi0039 & ~n17634;
  assign n17636 = ~n17628 & n17635;
  assign n17637 = ~pi0038 & ~n17636;
  assign n17638 = ~n17610 & n17637;
  assign n17639 = pi0140 & ~n17470;
  assign n17640 = n2521 & n17639;
  assign n17641 = ~pi0140 & ~n17490;
  assign n17642 = ~pi0761 & ~n17640;
  assign n17643 = ~n17641 & n17642;
  assign n17644 = ~pi0140 & ~n16667;
  assign n17645 = n16667 & n17355;
  assign n17646 = pi0761 & ~n17644;
  assign n17647 = ~n17645 & n17646;
  assign n17648 = ~n17643 & ~n17647;
  assign n17649 = ~pi0039 & ~n17648;
  assign n17650 = pi0038 & ~n16751;
  assign n17651 = ~n17649 & n17650;
  assign n17652 = ~n17638 & ~n17651;
  assign n17653 = ~pi0738 & ~n17652;
  assign n17654 = n2571 & ~n17319;
  assign n17655 = ~n17653 & n17654;
  assign n17656 = ~n16640 & ~n17655;
  assign n17657 = ~pi0625 & n17656;
  assign n17658 = pi0625 & n17286;
  assign n17659 = ~pi1153 & ~n17658;
  assign n17660 = ~n17657 & n17659;
  assign n17661 = ~pi0608 & ~n17064;
  assign n17662 = ~n17660 & n17661;
  assign n17663 = ~pi0625 & n17286;
  assign n17664 = pi0625 & n17656;
  assign n17665 = pi1153 & ~n17663;
  assign n17666 = ~n17664 & n17665;
  assign n17667 = pi0608 & ~n17068;
  assign n17668 = ~n17666 & n17667;
  assign n17669 = ~n17662 & ~n17668;
  assign n17670 = pi0778 & ~n17669;
  assign n17671 = ~pi0778 & n17656;
  assign n17672 = ~n17670 & ~n17671;
  assign n17673 = ~pi0609 & ~n17672;
  assign n17674 = pi0609 & n17071;
  assign n17675 = ~pi1155 & ~n17674;
  assign n17676 = ~n17673 & n17675;
  assign n17677 = ~pi0660 & ~n17295;
  assign n17678 = ~n17676 & n17677;
  assign n17679 = ~pi0609 & n17071;
  assign n17680 = pi0609 & ~n17672;
  assign n17681 = pi1155 & ~n17679;
  assign n17682 = ~n17680 & n17681;
  assign n17683 = pi0660 & ~n17300;
  assign n17684 = ~n17682 & n17683;
  assign n17685 = ~n17678 & ~n17684;
  assign n17686 = pi0785 & ~n17685;
  assign n17687 = ~pi0785 & ~n17672;
  assign n17688 = ~n17686 & ~n17687;
  assign n17689 = ~pi0618 & ~n17688;
  assign n17690 = pi0618 & n17078;
  assign n17691 = ~pi1154 & ~n17690;
  assign n17692 = ~n17689 & n17691;
  assign n17693 = ~pi0627 & ~n17308;
  assign n17694 = ~n17692 & n17693;
  assign n17695 = ~pi0618 & n17078;
  assign n17696 = pi0618 & ~n17688;
  assign n17697 = pi1154 & ~n17695;
  assign n17698 = ~n17696 & n17697;
  assign n17699 = pi0627 & ~n17312;
  assign n17700 = ~n17698 & n17699;
  assign n17701 = ~n17694 & ~n17700;
  assign n17702 = pi0781 & ~n17701;
  assign n17703 = ~pi0781 & ~n17688;
  assign n17704 = ~n17702 & ~n17703;
  assign n17705 = ~pi0619 & ~n17704;
  assign n17706 = pi0619 & ~n17081;
  assign n17707 = ~pi1159 & ~n17706;
  assign n17708 = ~n17705 & n17707;
  assign n17709 = ~pi0648 & ~n17318;
  assign n17710 = ~n17708 & n17709;
  assign n17711 = ~pi0619 & n17315;
  assign n17712 = pi0619 & n17060;
  assign n17713 = ~pi1159 & ~n17712;
  assign n17714 = ~n17711 & n17713;
  assign n17715 = pi0619 & ~n17704;
  assign n17716 = ~pi0619 & ~n17081;
  assign n17717 = pi1159 & ~n17716;
  assign n17718 = ~n17715 & n17717;
  assign n17719 = pi0648 & ~n17714;
  assign n17720 = ~n17718 & n17719;
  assign n17721 = ~n17710 & ~n17720;
  assign n17722 = pi0789 & ~n17721;
  assign n17723 = ~pi0789 & ~n17704;
  assign n17724 = ~n17722 & ~n17723;
  assign n17725 = ~pi0788 & n17724;
  assign n17726 = ~pi0626 & n17724;
  assign n17727 = pi0626 & ~n17084;
  assign n17728 = ~pi0641 & ~n17727;
  assign n17729 = ~n17726 & n17728;
  assign n17730 = ~pi0641 & ~pi1158;
  assign n17731 = ~pi0789 & ~n17315;
  assign n17732 = ~n17318 & ~n17714;
  assign n17733 = pi0789 & ~n17732;
  assign n17734 = ~n17731 & ~n17733;
  assign n17735 = ~pi0626 & n17734;
  assign n17736 = pi0626 & n17060;
  assign n17737 = ~pi1158 & ~n17736;
  assign n17738 = ~n17735 & n17737;
  assign n17739 = ~n17730 & ~n17738;
  assign n17740 = ~n17729 & ~n17739;
  assign n17741 = pi0626 & n17724;
  assign n17742 = ~pi0626 & ~n17084;
  assign n17743 = pi0641 & ~n17742;
  assign n17744 = ~n17741 & n17743;
  assign n17745 = pi0641 & pi1158;
  assign n17746 = ~pi0626 & n17060;
  assign n17747 = pi0626 & n17734;
  assign n17748 = pi1158 & ~n17746;
  assign n17749 = ~n17747 & n17748;
  assign n17750 = ~n17745 & ~n17749;
  assign n17751 = ~n17744 & ~n17750;
  assign n17752 = ~n17740 & ~n17751;
  assign n17753 = pi0788 & ~n17752;
  assign n17754 = ~n17725 & ~n17753;
  assign n17755 = ~pi0628 & n17754;
  assign n17756 = ~n17738 & ~n17749;
  assign n17757 = pi0788 & ~n17756;
  assign n17758 = ~pi0788 & ~n17734;
  assign n17759 = ~n17757 & ~n17758;
  assign n17760 = pi0628 & n17759;
  assign n17761 = ~pi1156 & ~n17760;
  assign n17762 = ~n17755 & n17761;
  assign n17763 = ~pi0629 & ~n17092;
  assign n17764 = ~n17762 & n17763;
  assign n17765 = pi0628 & n17754;
  assign n17766 = ~pi0628 & n17759;
  assign n17767 = pi1156 & ~n17766;
  assign n17768 = ~n17765 & n17767;
  assign n17769 = pi0629 & ~n17096;
  assign n17770 = ~n17768 & n17769;
  assign n17771 = ~n17764 & ~n17770;
  assign n17772 = pi0792 & ~n17771;
  assign n17773 = ~pi0792 & n17754;
  assign n17774 = ~n17772 & ~n17773;
  assign n17775 = ~pi0647 & ~n17774;
  assign n17776 = ~pi0629 & pi1156;
  assign n17777 = pi0629 & ~pi1156;
  assign n17778 = ~n17776 & ~n17777;
  assign n17779 = pi0792 & ~n17778;
  assign n17780 = n17759 & ~n17779;
  assign n17781 = n17060 & n17779;
  assign n17782 = ~n17780 & ~n17781;
  assign n17783 = pi0647 & ~n17782;
  assign n17784 = ~pi1157 & ~n17783;
  assign n17785 = ~n17775 & n17784;
  assign n17786 = ~pi0630 & ~n17104;
  assign n17787 = ~n17785 & n17786;
  assign n17788 = pi0647 & ~n17774;
  assign n17789 = ~pi0647 & ~n17782;
  assign n17790 = pi1157 & ~n17789;
  assign n17791 = ~n17788 & n17790;
  assign n17792 = pi0630 & ~n17108;
  assign n17793 = ~n17791 & n17792;
  assign n17794 = ~n17787 & ~n17793;
  assign n17795 = pi0787 & ~n17794;
  assign n17796 = ~pi0787 & ~n17774;
  assign n17797 = ~n17795 & ~n17796;
  assign n17798 = pi0644 & ~n17797;
  assign n17799 = pi0715 & ~n17112;
  assign n17800 = ~n17798 & n17799;
  assign n17801 = ~pi0630 & pi1157;
  assign n17802 = pi0630 & ~pi1157;
  assign n17803 = ~n17801 & ~n17802;
  assign n17804 = pi0787 & ~n17803;
  assign n17805 = n17782 & ~n17804;
  assign n17806 = ~n17060 & n17804;
  assign n17807 = ~n17805 & ~n17806;
  assign n17808 = pi0644 & n17807;
  assign n17809 = ~pi0644 & n17060;
  assign n17810 = ~pi0715 & ~n17809;
  assign n17811 = ~n17808 & n17810;
  assign n17812 = pi1160 & ~n17811;
  assign n17813 = ~n17800 & n17812;
  assign n17814 = ~pi0644 & ~n17797;
  assign n17815 = pi0644 & n17111;
  assign n17816 = ~pi0715 & ~n17815;
  assign n17817 = ~n17814 & n17816;
  assign n17818 = ~pi0644 & n17807;
  assign n17819 = pi0644 & n17060;
  assign n17820 = pi0715 & ~n17819;
  assign n17821 = ~n17818 & n17820;
  assign n17822 = ~pi1160 & ~n17821;
  assign n17823 = ~n17817 & n17822;
  assign n17824 = pi0790 & ~n17813;
  assign n17825 = ~n17823 & n17824;
  assign n17826 = ~pi0790 & n17797;
  assign n17827 = ~po1038 & ~n17826;
  assign n17828 = ~n17825 & n17827;
  assign n17829 = ~pi0140 & po1038;
  assign n17830 = ~pi0832 & ~n17829;
  assign n17831 = ~n17828 & n17830;
  assign n17832 = ~pi0140 & ~n2926;
  assign n17833 = ~pi0647 & n17832;
  assign n17834 = ~pi0738 & n16645;
  assign n17835 = ~n17832 & ~n17834;
  assign n17836 = ~pi0778 & n17835;
  assign n17837 = ~pi0625 & n17834;
  assign n17838 = ~n17835 & ~n17837;
  assign n17839 = pi1153 & ~n17838;
  assign n17840 = ~pi1153 & ~n17832;
  assign n17841 = ~n17837 & n17840;
  assign n17842 = ~n17839 & ~n17841;
  assign n17843 = pi0778 & ~n17842;
  assign n17844 = ~n17836 & ~n17843;
  assign n17845 = n2926 & n17075;
  assign n17846 = n17844 & ~n17845;
  assign n17847 = n2926 & n16639;
  assign n17848 = n17846 & ~n17847;
  assign n17849 = n2926 & n16635;
  assign n17850 = n17848 & ~n17849;
  assign n17851 = n2926 & n16631;
  assign n17852 = n17850 & ~n17851;
  assign n17853 = ~pi0628 & pi1156;
  assign n17854 = pi0628 & ~pi1156;
  assign n17855 = ~n17853 & ~n17854;
  assign n17856 = pi0792 & ~n17855;
  assign n17857 = n2926 & n17856;
  assign n17858 = n17852 & ~n17857;
  assign n17859 = pi0647 & n17858;
  assign n17860 = pi1157 & ~n17833;
  assign n17861 = ~n17859 & n17860;
  assign n17862 = ~pi0628 & n2926;
  assign n17863 = n17852 & ~n17862;
  assign n17864 = pi1156 & ~n17863;
  assign n17865 = ~pi0626 & pi1158;
  assign n17866 = pi0626 & ~pi1158;
  assign n17867 = ~n17865 & ~n17866;
  assign n17868 = ~pi0626 & pi0641;
  assign n17869 = pi0626 & ~pi0641;
  assign n17870 = ~n17868 & ~n17869;
  assign n17871 = ~n17867 & ~n17870;
  assign n17872 = n17850 & n17871;
  assign n17873 = ~pi0626 & n17832;
  assign n17874 = n2926 & n17117;
  assign n17875 = ~pi0761 & n17244;
  assign n17876 = ~n17832 & ~n17875;
  assign n17877 = ~n17874 & ~n17876;
  assign n17878 = ~pi0785 & ~n17877;
  assign n17879 = n2926 & ~n17291;
  assign n17880 = ~n17876 & ~n17879;
  assign n17881 = pi1155 & ~n17880;
  assign n17882 = pi0609 & n2926;
  assign n17883 = n17877 & ~n17882;
  assign n17884 = ~pi1155 & ~n17883;
  assign n17885 = ~n17881 & ~n17884;
  assign n17886 = pi0785 & ~n17885;
  assign n17887 = ~n17878 & ~n17886;
  assign n17888 = ~pi0781 & ~n17887;
  assign n17889 = ~pi0618 & n2926;
  assign n17890 = n17887 & ~n17889;
  assign n17891 = pi1154 & ~n17890;
  assign n17892 = pi0618 & n2926;
  assign n17893 = n17887 & ~n17892;
  assign n17894 = ~pi1154 & ~n17893;
  assign n17895 = ~n17891 & ~n17894;
  assign n17896 = pi0781 & ~n17895;
  assign n17897 = ~n17888 & ~n17896;
  assign n17898 = ~pi0789 & ~n17897;
  assign n17899 = ~pi0619 & n17832;
  assign n17900 = pi0619 & n17897;
  assign n17901 = pi1159 & ~n17899;
  assign n17902 = ~n17900 & n17901;
  assign n17903 = ~pi0619 & n17897;
  assign n17904 = pi0619 & n17832;
  assign n17905 = ~pi1159 & ~n17904;
  assign n17906 = ~n17903 & n17905;
  assign n17907 = ~n17902 & ~n17906;
  assign n17908 = pi0789 & ~n17907;
  assign n17909 = ~n17898 & ~n17908;
  assign n17910 = pi0626 & n17909;
  assign n17911 = pi1158 & ~n17873;
  assign n17912 = ~n17910 & n17911;
  assign n17913 = ~pi0626 & n17909;
  assign n17914 = pi0626 & n17832;
  assign n17915 = ~pi1158 & ~n17914;
  assign n17916 = ~n17913 & n17915;
  assign n17917 = ~n17912 & ~n17916;
  assign n17918 = ~n16630 & n17917;
  assign n17919 = ~n17872 & ~n17918;
  assign n17920 = pi0788 & ~n17919;
  assign n17921 = pi0618 & n17846;
  assign n17922 = pi0609 & n17844;
  assign n17923 = ~n17168 & ~n17835;
  assign n17924 = pi0625 & n17923;
  assign n17925 = n17876 & ~n17923;
  assign n17926 = ~n17924 & ~n17925;
  assign n17927 = n17840 & ~n17926;
  assign n17928 = ~pi0608 & ~n17839;
  assign n17929 = ~n17927 & n17928;
  assign n17930 = pi1153 & n17876;
  assign n17931 = ~n17924 & n17930;
  assign n17932 = pi0608 & ~n17841;
  assign n17933 = ~n17931 & n17932;
  assign n17934 = ~n17929 & ~n17933;
  assign n17935 = pi0778 & ~n17934;
  assign n17936 = ~pi0778 & ~n17925;
  assign n17937 = ~n17935 & ~n17936;
  assign n17938 = ~pi0609 & ~n17937;
  assign n17939 = ~pi1155 & ~n17922;
  assign n17940 = ~n17938 & n17939;
  assign n17941 = ~pi0660 & ~n17881;
  assign n17942 = ~n17940 & n17941;
  assign n17943 = ~pi0609 & n17844;
  assign n17944 = pi0609 & ~n17937;
  assign n17945 = pi1155 & ~n17943;
  assign n17946 = ~n17944 & n17945;
  assign n17947 = pi0660 & ~n17884;
  assign n17948 = ~n17946 & n17947;
  assign n17949 = ~n17942 & ~n17948;
  assign n17950 = pi0785 & ~n17949;
  assign n17951 = ~pi0785 & ~n17937;
  assign n17952 = ~n17950 & ~n17951;
  assign n17953 = ~pi0618 & ~n17952;
  assign n17954 = ~pi1154 & ~n17921;
  assign n17955 = ~n17953 & n17954;
  assign n17956 = ~pi0627 & ~n17891;
  assign n17957 = ~n17955 & n17956;
  assign n17958 = ~pi0618 & n17846;
  assign n17959 = pi0618 & ~n17952;
  assign n17960 = pi1154 & ~n17958;
  assign n17961 = ~n17959 & n17960;
  assign n17962 = pi0627 & ~n17894;
  assign n17963 = ~n17961 & n17962;
  assign n17964 = ~n17957 & ~n17963;
  assign n17965 = pi0781 & ~n17964;
  assign n17966 = ~pi0781 & ~n17952;
  assign n17967 = ~n17965 & ~n17966;
  assign n17968 = ~pi0789 & n17967;
  assign n17969 = pi0788 & ~n17867;
  assign n17970 = ~n16631 & ~n17969;
  assign n17971 = ~pi0619 & ~n17967;
  assign n17972 = pi0619 & n17848;
  assign n17973 = ~pi1159 & ~n17972;
  assign n17974 = ~n17971 & n17973;
  assign n17975 = ~pi0648 & ~n17902;
  assign n17976 = ~n17974 & n17975;
  assign n17977 = ~pi0619 & n17848;
  assign n17978 = pi0619 & ~n17967;
  assign n17979 = pi1159 & ~n17977;
  assign n17980 = ~n17978 & n17979;
  assign n17981 = pi0648 & ~n17906;
  assign n17982 = ~n17980 & n17981;
  assign n17983 = pi0789 & ~n17976;
  assign n17984 = ~n17982 & n17983;
  assign n17985 = ~n17968 & n17970;
  assign n17986 = ~n17984 & n17985;
  assign n17987 = ~n17920 & ~n17986;
  assign n17988 = ~pi0628 & ~n17987;
  assign n17989 = ~pi0788 & ~n17909;
  assign n17990 = pi0788 & ~n17917;
  assign n17991 = ~n17989 & ~n17990;
  assign n17992 = pi0628 & n17991;
  assign n17993 = ~pi1156 & ~n17992;
  assign n17994 = ~n17988 & n17993;
  assign n17995 = ~pi0629 & ~n17864;
  assign n17996 = ~n17994 & n17995;
  assign n17997 = pi0628 & n2926;
  assign n17998 = n17852 & ~n17997;
  assign n17999 = ~pi1156 & ~n17998;
  assign n18000 = ~pi0628 & n17991;
  assign n18001 = pi0628 & ~n17987;
  assign n18002 = pi1156 & ~n18000;
  assign n18003 = ~n18001 & n18002;
  assign n18004 = pi0629 & ~n17999;
  assign n18005 = ~n18003 & n18004;
  assign n18006 = ~n17996 & ~n18005;
  assign n18007 = pi0792 & ~n18006;
  assign n18008 = ~pi0792 & ~n17987;
  assign n18009 = ~n18007 & ~n18008;
  assign n18010 = ~pi0647 & ~n18009;
  assign n18011 = ~n17779 & n17991;
  assign n18012 = n17779 & n17832;
  assign n18013 = ~n18011 & ~n18012;
  assign n18014 = pi0647 & ~n18013;
  assign n18015 = ~pi1157 & ~n18014;
  assign n18016 = ~n18010 & n18015;
  assign n18017 = ~pi0630 & ~n17861;
  assign n18018 = ~n18016 & n18017;
  assign n18019 = ~pi0647 & n17858;
  assign n18020 = pi0647 & n17832;
  assign n18021 = ~pi1157 & ~n18020;
  assign n18022 = ~n18019 & n18021;
  assign n18023 = pi0647 & ~n18009;
  assign n18024 = ~pi0647 & ~n18013;
  assign n18025 = pi1157 & ~n18024;
  assign n18026 = ~n18023 & n18025;
  assign n18027 = pi0630 & ~n18022;
  assign n18028 = ~n18026 & n18027;
  assign n18029 = ~n18018 & ~n18028;
  assign n18030 = pi0787 & ~n18029;
  assign n18031 = ~pi0787 & ~n18009;
  assign n18032 = ~n18030 & ~n18031;
  assign n18033 = ~pi0790 & ~n18032;
  assign n18034 = ~pi0787 & ~n17858;
  assign n18035 = ~n17861 & ~n18022;
  assign n18036 = pi0787 & ~n18035;
  assign n18037 = ~n18034 & ~n18036;
  assign n18038 = ~pi0644 & n18037;
  assign n18039 = pi0644 & ~n18032;
  assign n18040 = pi0715 & ~n18038;
  assign n18041 = ~n18039 & n18040;
  assign n18042 = n17804 & ~n17832;
  assign n18043 = ~n17804 & n18013;
  assign n18044 = ~n18042 & ~n18043;
  assign n18045 = pi0644 & n18044;
  assign n18046 = ~pi0644 & n17832;
  assign n18047 = ~pi0715 & ~n18046;
  assign n18048 = ~n18045 & n18047;
  assign n18049 = pi1160 & ~n18048;
  assign n18050 = ~n18041 & n18049;
  assign n18051 = ~pi0644 & n18044;
  assign n18052 = pi0644 & n17832;
  assign n18053 = pi0715 & ~n18052;
  assign n18054 = ~n18051 & n18053;
  assign n18055 = pi0644 & n18037;
  assign n18056 = ~pi0644 & ~n18032;
  assign n18057 = ~pi0715 & ~n18055;
  assign n18058 = ~n18056 & n18057;
  assign n18059 = ~pi1160 & ~n18054;
  assign n18060 = ~n18058 & n18059;
  assign n18061 = ~n18050 & ~n18060;
  assign n18062 = pi0790 & ~n18061;
  assign n18063 = pi0832 & ~n18033;
  assign n18064 = ~n18062 & n18063;
  assign po0297 = ~n17831 & ~n18064;
  assign n18066 = ~pi0141 & ~n17059;
  assign n18067 = n16635 & ~n18066;
  assign n18068 = pi0141 & ~n2571;
  assign n18069 = ~pi0141 & ~n16641;
  assign n18070 = n16647 & ~n18069;
  assign n18071 = ~pi0039 & n16948;
  assign n18072 = ~n16841 & ~n18071;
  assign n18073 = ~pi0141 & n18072;
  assign n18074 = pi0039 & ~n16749;
  assign n18075 = ~pi0039 & n16926;
  assign n18076 = ~n18074 & ~n18075;
  assign n18077 = pi0141 & ~n18076;
  assign n18078 = ~pi0038 & ~n18077;
  assign n18079 = ~n18073 & n18078;
  assign n18080 = pi0706 & ~n18070;
  assign n18081 = ~n18079 & n18080;
  assign n18082 = ~pi0141 & ~pi0706;
  assign n18083 = ~n17052 & n18082;
  assign n18084 = n2571 & ~n18083;
  assign n18085 = ~n18081 & n18084;
  assign n18086 = ~n18068 & ~n18085;
  assign n18087 = ~pi0778 & ~n18086;
  assign n18088 = ~pi0625 & n18066;
  assign n18089 = pi0625 & n18086;
  assign n18090 = pi1153 & ~n18088;
  assign n18091 = ~n18089 & n18090;
  assign n18092 = ~pi0625 & n18086;
  assign n18093 = pi0625 & n18066;
  assign n18094 = ~pi1153 & ~n18093;
  assign n18095 = ~n18092 & n18094;
  assign n18096 = ~n18091 & ~n18095;
  assign n18097 = pi0778 & ~n18096;
  assign n18098 = ~n18087 & ~n18097;
  assign n18099 = ~n17075 & ~n18098;
  assign n18100 = n17075 & ~n18066;
  assign n18101 = ~n18099 & ~n18100;
  assign n18102 = ~n16639 & n18101;
  assign n18103 = n16639 & n18066;
  assign n18104 = ~n18102 & ~n18103;
  assign n18105 = ~n16635 & n18104;
  assign n18106 = ~n18067 & ~n18105;
  assign n18107 = ~n16631 & n18106;
  assign n18108 = n16631 & n18066;
  assign n18109 = ~n18107 & ~n18108;
  assign n18110 = ~pi0792 & n18109;
  assign n18111 = ~pi0628 & n18066;
  assign n18112 = pi0628 & ~n18109;
  assign n18113 = pi1156 & ~n18111;
  assign n18114 = ~n18112 & n18113;
  assign n18115 = pi0628 & n18066;
  assign n18116 = ~pi0628 & ~n18109;
  assign n18117 = ~pi1156 & ~n18115;
  assign n18118 = ~n18116 & n18117;
  assign n18119 = ~n18114 & ~n18118;
  assign n18120 = pi0792 & ~n18119;
  assign n18121 = ~n18110 & ~n18120;
  assign n18122 = ~pi0787 & ~n18121;
  assign n18123 = ~pi0647 & n18066;
  assign n18124 = pi0647 & n18121;
  assign n18125 = pi1157 & ~n18123;
  assign n18126 = ~n18124 & n18125;
  assign n18127 = ~pi0647 & n18121;
  assign n18128 = pi0647 & n18066;
  assign n18129 = ~pi1157 & ~n18128;
  assign n18130 = ~n18127 & n18129;
  assign n18131 = ~n18126 & ~n18130;
  assign n18132 = pi0787 & ~n18131;
  assign n18133 = ~n18122 & ~n18132;
  assign n18134 = ~pi0644 & n18133;
  assign n18135 = ~pi0618 & n18066;
  assign n18136 = pi0749 & n17280;
  assign n18137 = ~n18069 & ~n18136;
  assign n18138 = pi0038 & ~n18137;
  assign n18139 = ~pi0749 & n17046;
  assign n18140 = pi0141 & n17273;
  assign n18141 = ~n18139 & ~n18140;
  assign n18142 = pi0039 & ~n18141;
  assign n18143 = ~pi0141 & n17221;
  assign n18144 = pi0141 & n17234;
  assign n18145 = pi0749 & ~n18144;
  assign n18146 = ~n18143 & n18145;
  assign n18147 = ~pi0039 & n16958;
  assign n18148 = ~pi0141 & ~pi0749;
  assign n18149 = ~n18147 & n18148;
  assign n18150 = ~n18146 & ~n18149;
  assign n18151 = ~pi0038 & ~n18150;
  assign n18152 = ~n18142 & n18151;
  assign n18153 = ~n18138 & ~n18152;
  assign n18154 = n2571 & n18153;
  assign n18155 = ~n18068 & ~n18154;
  assign n18156 = ~n17117 & ~n18155;
  assign n18157 = n17117 & ~n18066;
  assign n18158 = ~n18156 & ~n18157;
  assign n18159 = ~pi0785 & ~n18158;
  assign n18160 = ~n17291 & ~n18066;
  assign n18161 = pi0609 & n18156;
  assign n18162 = ~n18160 & ~n18161;
  assign n18163 = pi1155 & ~n18162;
  assign n18164 = ~n17296 & ~n18066;
  assign n18165 = ~pi0609 & n18156;
  assign n18166 = ~n18164 & ~n18165;
  assign n18167 = ~pi1155 & ~n18166;
  assign n18168 = ~n18163 & ~n18167;
  assign n18169 = pi0785 & ~n18168;
  assign n18170 = ~n18159 & ~n18169;
  assign n18171 = pi0618 & n18170;
  assign n18172 = pi1154 & ~n18135;
  assign n18173 = ~n18171 & n18172;
  assign n18174 = ~pi0706 & ~n18153;
  assign n18175 = ~pi0039 & n17645;
  assign n18176 = pi0038 & ~n18175;
  assign n18177 = n18137 & n18176;
  assign n18178 = ~pi0141 & ~n17629;
  assign n18179 = pi0141 & ~n17631;
  assign n18180 = pi0749 & ~n18179;
  assign n18181 = ~n18178 & n18180;
  assign n18182 = ~pi0141 & n17612;
  assign n18183 = pi0141 & n17625;
  assign n18184 = ~pi0749 & ~n18182;
  assign n18185 = ~n18183 & n18184;
  assign n18186 = ~pi0039 & ~n18181;
  assign n18187 = ~n18185 & n18186;
  assign n18188 = pi0141 & n17605;
  assign n18189 = ~pi0141 & ~n17546;
  assign n18190 = pi0749 & ~n18189;
  assign n18191 = ~n18188 & n18190;
  assign n18192 = ~pi0141 & n17404;
  assign n18193 = pi0141 & n17485;
  assign n18194 = ~pi0749 & ~n18193;
  assign n18195 = ~n18192 & n18194;
  assign n18196 = pi0039 & ~n18191;
  assign n18197 = ~n18195 & n18196;
  assign n18198 = ~pi0038 & ~n18187;
  assign n18199 = ~n18197 & n18198;
  assign n18200 = pi0706 & ~n18177;
  assign n18201 = ~n18199 & n18200;
  assign n18202 = n2571 & ~n18174;
  assign n18203 = ~n18201 & n18202;
  assign n18204 = ~n18068 & ~n18203;
  assign n18205 = ~pi0625 & n18204;
  assign n18206 = pi0625 & n18155;
  assign n18207 = ~pi1153 & ~n18206;
  assign n18208 = ~n18205 & n18207;
  assign n18209 = ~pi0608 & ~n18091;
  assign n18210 = ~n18208 & n18209;
  assign n18211 = ~pi0625 & n18155;
  assign n18212 = pi0625 & n18204;
  assign n18213 = pi1153 & ~n18211;
  assign n18214 = ~n18212 & n18213;
  assign n18215 = pi0608 & ~n18095;
  assign n18216 = ~n18214 & n18215;
  assign n18217 = ~n18210 & ~n18216;
  assign n18218 = pi0778 & ~n18217;
  assign n18219 = ~pi0778 & n18204;
  assign n18220 = ~n18218 & ~n18219;
  assign n18221 = ~pi0609 & ~n18220;
  assign n18222 = pi0609 & n18098;
  assign n18223 = ~pi1155 & ~n18222;
  assign n18224 = ~n18221 & n18223;
  assign n18225 = ~pi0660 & ~n18163;
  assign n18226 = ~n18224 & n18225;
  assign n18227 = ~pi0609 & n18098;
  assign n18228 = pi0609 & ~n18220;
  assign n18229 = pi1155 & ~n18227;
  assign n18230 = ~n18228 & n18229;
  assign n18231 = pi0660 & ~n18167;
  assign n18232 = ~n18230 & n18231;
  assign n18233 = ~n18226 & ~n18232;
  assign n18234 = pi0785 & ~n18233;
  assign n18235 = ~pi0785 & ~n18220;
  assign n18236 = ~n18234 & ~n18235;
  assign n18237 = ~pi0618 & ~n18236;
  assign n18238 = pi0618 & n18101;
  assign n18239 = ~pi1154 & ~n18238;
  assign n18240 = ~n18237 & n18239;
  assign n18241 = ~pi0627 & ~n18173;
  assign n18242 = ~n18240 & n18241;
  assign n18243 = ~pi0618 & n18170;
  assign n18244 = pi0618 & n18066;
  assign n18245 = ~pi1154 & ~n18244;
  assign n18246 = ~n18243 & n18245;
  assign n18247 = ~pi0618 & n18101;
  assign n18248 = pi0618 & ~n18236;
  assign n18249 = pi1154 & ~n18247;
  assign n18250 = ~n18248 & n18249;
  assign n18251 = pi0627 & ~n18246;
  assign n18252 = ~n18250 & n18251;
  assign n18253 = ~n18242 & ~n18252;
  assign n18254 = pi0781 & ~n18253;
  assign n18255 = ~pi0781 & ~n18236;
  assign n18256 = ~n18254 & ~n18255;
  assign n18257 = ~pi0619 & ~n18256;
  assign n18258 = pi0619 & ~n18104;
  assign n18259 = ~pi1159 & ~n18258;
  assign n18260 = ~n18257 & n18259;
  assign n18261 = ~pi0619 & n18066;
  assign n18262 = ~pi0781 & ~n18170;
  assign n18263 = ~n18173 & ~n18246;
  assign n18264 = pi0781 & ~n18263;
  assign n18265 = ~n18262 & ~n18264;
  assign n18266 = pi0619 & n18265;
  assign n18267 = pi1159 & ~n18261;
  assign n18268 = ~n18266 & n18267;
  assign n18269 = ~pi0648 & ~n18268;
  assign n18270 = ~n18260 & n18269;
  assign n18271 = pi0619 & ~n18256;
  assign n18272 = ~pi0619 & ~n18104;
  assign n18273 = pi1159 & ~n18272;
  assign n18274 = ~n18271 & n18273;
  assign n18275 = ~pi0619 & n18265;
  assign n18276 = pi0619 & n18066;
  assign n18277 = ~pi1159 & ~n18276;
  assign n18278 = ~n18275 & n18277;
  assign n18279 = pi0648 & ~n18278;
  assign n18280 = ~n18274 & n18279;
  assign n18281 = ~n18270 & ~n18280;
  assign n18282 = pi0789 & ~n18281;
  assign n18283 = ~pi0789 & ~n18256;
  assign n18284 = ~n18282 & ~n18283;
  assign n18285 = ~pi0788 & n18284;
  assign n18286 = ~pi0626 & n18284;
  assign n18287 = pi0626 & ~n18106;
  assign n18288 = ~pi0641 & ~n18287;
  assign n18289 = ~n18286 & n18288;
  assign n18290 = ~pi0789 & ~n18265;
  assign n18291 = ~n18268 & ~n18278;
  assign n18292 = pi0789 & ~n18291;
  assign n18293 = ~n18290 & ~n18292;
  assign n18294 = ~pi0626 & n18293;
  assign n18295 = pi0626 & n18066;
  assign n18296 = ~pi1158 & ~n18295;
  assign n18297 = ~n18294 & n18296;
  assign n18298 = ~n17730 & ~n18297;
  assign n18299 = ~n18289 & ~n18298;
  assign n18300 = pi0626 & n18284;
  assign n18301 = ~pi0626 & ~n18106;
  assign n18302 = pi0641 & ~n18301;
  assign n18303 = ~n18300 & n18302;
  assign n18304 = ~pi0626 & n18066;
  assign n18305 = pi0626 & n18293;
  assign n18306 = pi1158 & ~n18304;
  assign n18307 = ~n18305 & n18306;
  assign n18308 = ~n17745 & ~n18307;
  assign n18309 = ~n18303 & ~n18308;
  assign n18310 = ~n18299 & ~n18309;
  assign n18311 = pi0788 & ~n18310;
  assign n18312 = ~n18285 & ~n18311;
  assign n18313 = ~pi0628 & n18312;
  assign n18314 = ~n18297 & ~n18307;
  assign n18315 = pi0788 & ~n18314;
  assign n18316 = ~pi0788 & ~n18293;
  assign n18317 = ~n18315 & ~n18316;
  assign n18318 = pi0628 & n18317;
  assign n18319 = ~pi1156 & ~n18318;
  assign n18320 = ~n18313 & n18319;
  assign n18321 = ~pi0629 & ~n18114;
  assign n18322 = ~n18320 & n18321;
  assign n18323 = pi0628 & n18312;
  assign n18324 = ~pi0628 & n18317;
  assign n18325 = pi1156 & ~n18324;
  assign n18326 = ~n18323 & n18325;
  assign n18327 = pi0629 & ~n18118;
  assign n18328 = ~n18326 & n18327;
  assign n18329 = ~n18322 & ~n18328;
  assign n18330 = pi0792 & ~n18329;
  assign n18331 = ~pi0792 & n18312;
  assign n18332 = ~n18330 & ~n18331;
  assign n18333 = ~pi0647 & ~n18332;
  assign n18334 = ~n17779 & n18317;
  assign n18335 = n17779 & n18066;
  assign n18336 = ~n18334 & ~n18335;
  assign n18337 = pi0647 & ~n18336;
  assign n18338 = ~pi1157 & ~n18337;
  assign n18339 = ~n18333 & n18338;
  assign n18340 = ~pi0630 & ~n18126;
  assign n18341 = ~n18339 & n18340;
  assign n18342 = pi0647 & ~n18332;
  assign n18343 = ~pi0647 & ~n18336;
  assign n18344 = pi1157 & ~n18343;
  assign n18345 = ~n18342 & n18344;
  assign n18346 = pi0630 & ~n18130;
  assign n18347 = ~n18345 & n18346;
  assign n18348 = ~n18341 & ~n18347;
  assign n18349 = pi0787 & ~n18348;
  assign n18350 = ~pi0787 & ~n18332;
  assign n18351 = ~n18349 & ~n18350;
  assign n18352 = pi0644 & ~n18351;
  assign n18353 = pi0715 & ~n18134;
  assign n18354 = ~n18352 & n18353;
  assign n18355 = n17804 & ~n18066;
  assign n18356 = ~n17804 & n18336;
  assign n18357 = ~n18355 & ~n18356;
  assign n18358 = pi0644 & n18357;
  assign n18359 = ~pi0644 & n18066;
  assign n18360 = ~pi0715 & ~n18359;
  assign n18361 = ~n18358 & n18360;
  assign n18362 = pi1160 & ~n18361;
  assign n18363 = ~n18354 & n18362;
  assign n18364 = ~pi0644 & ~n18351;
  assign n18365 = pi0644 & n18133;
  assign n18366 = ~pi0715 & ~n18365;
  assign n18367 = ~n18364 & n18366;
  assign n18368 = ~pi0644 & n18357;
  assign n18369 = pi0644 & n18066;
  assign n18370 = pi0715 & ~n18369;
  assign n18371 = ~n18368 & n18370;
  assign n18372 = ~pi1160 & ~n18371;
  assign n18373 = ~n18367 & n18372;
  assign n18374 = pi0790 & ~n18363;
  assign n18375 = ~n18373 & n18374;
  assign n18376 = ~pi0790 & n18351;
  assign n18377 = ~po1038 & ~n18376;
  assign n18378 = ~n18375 & n18377;
  assign n18379 = ~pi0141 & po1038;
  assign n18380 = ~pi0832 & ~n18379;
  assign n18381 = ~n18378 & n18380;
  assign n18382 = ~pi0141 & ~n2926;
  assign n18383 = ~pi0647 & n18382;
  assign n18384 = pi0706 & n16645;
  assign n18385 = ~n18382 & ~n18384;
  assign n18386 = ~pi0778 & n18385;
  assign n18387 = ~pi0625 & n18384;
  assign n18388 = ~n18385 & ~n18387;
  assign n18389 = pi1153 & ~n18388;
  assign n18390 = ~pi1153 & ~n18382;
  assign n18391 = ~n18387 & n18390;
  assign n18392 = ~n18389 & ~n18391;
  assign n18393 = pi0778 & ~n18392;
  assign n18394 = ~n18386 & ~n18393;
  assign n18395 = ~n17845 & n18394;
  assign n18396 = ~n17847 & n18395;
  assign n18397 = ~n17849 & n18396;
  assign n18398 = ~n17851 & n18397;
  assign n18399 = ~n17857 & n18398;
  assign n18400 = pi0647 & n18399;
  assign n18401 = pi1157 & ~n18383;
  assign n18402 = ~n18400 & n18401;
  assign n18403 = ~n17862 & n18398;
  assign n18404 = pi1156 & ~n18403;
  assign n18405 = n17871 & n18397;
  assign n18406 = ~pi0626 & n18382;
  assign n18407 = pi0749 & n17244;
  assign n18408 = ~n18382 & ~n18407;
  assign n18409 = ~n17874 & ~n18408;
  assign n18410 = ~pi0785 & ~n18409;
  assign n18411 = ~n17879 & ~n18408;
  assign n18412 = pi1155 & ~n18411;
  assign n18413 = ~n17882 & n18409;
  assign n18414 = ~pi1155 & ~n18413;
  assign n18415 = ~n18412 & ~n18414;
  assign n18416 = pi0785 & ~n18415;
  assign n18417 = ~n18410 & ~n18416;
  assign n18418 = ~pi0781 & ~n18417;
  assign n18419 = ~n17889 & n18417;
  assign n18420 = pi1154 & ~n18419;
  assign n18421 = ~n17892 & n18417;
  assign n18422 = ~pi1154 & ~n18421;
  assign n18423 = ~n18420 & ~n18422;
  assign n18424 = pi0781 & ~n18423;
  assign n18425 = ~n18418 & ~n18424;
  assign n18426 = ~pi0789 & ~n18425;
  assign n18427 = ~pi0619 & n18382;
  assign n18428 = pi0619 & n18425;
  assign n18429 = pi1159 & ~n18427;
  assign n18430 = ~n18428 & n18429;
  assign n18431 = ~pi0619 & n18425;
  assign n18432 = pi0619 & n18382;
  assign n18433 = ~pi1159 & ~n18432;
  assign n18434 = ~n18431 & n18433;
  assign n18435 = ~n18430 & ~n18434;
  assign n18436 = pi0789 & ~n18435;
  assign n18437 = ~n18426 & ~n18436;
  assign n18438 = pi0626 & n18437;
  assign n18439 = pi1158 & ~n18406;
  assign n18440 = ~n18438 & n18439;
  assign n18441 = ~pi0626 & n18437;
  assign n18442 = pi0626 & n18382;
  assign n18443 = ~pi1158 & ~n18442;
  assign n18444 = ~n18441 & n18443;
  assign n18445 = ~n18440 & ~n18444;
  assign n18446 = ~n16630 & n18445;
  assign n18447 = ~n18405 & ~n18446;
  assign n18448 = pi0788 & ~n18447;
  assign n18449 = pi0618 & n18395;
  assign n18450 = pi0609 & n18394;
  assign n18451 = ~n17168 & ~n18385;
  assign n18452 = pi0625 & n18451;
  assign n18453 = n18408 & ~n18451;
  assign n18454 = ~n18452 & ~n18453;
  assign n18455 = n18390 & ~n18454;
  assign n18456 = ~pi0608 & ~n18389;
  assign n18457 = ~n18455 & n18456;
  assign n18458 = pi1153 & n18408;
  assign n18459 = ~n18452 & n18458;
  assign n18460 = pi0608 & ~n18391;
  assign n18461 = ~n18459 & n18460;
  assign n18462 = ~n18457 & ~n18461;
  assign n18463 = pi0778 & ~n18462;
  assign n18464 = ~pi0778 & ~n18453;
  assign n18465 = ~n18463 & ~n18464;
  assign n18466 = ~pi0609 & ~n18465;
  assign n18467 = ~pi1155 & ~n18450;
  assign n18468 = ~n18466 & n18467;
  assign n18469 = ~pi0660 & ~n18412;
  assign n18470 = ~n18468 & n18469;
  assign n18471 = ~pi0609 & n18394;
  assign n18472 = pi0609 & ~n18465;
  assign n18473 = pi1155 & ~n18471;
  assign n18474 = ~n18472 & n18473;
  assign n18475 = pi0660 & ~n18414;
  assign n18476 = ~n18474 & n18475;
  assign n18477 = ~n18470 & ~n18476;
  assign n18478 = pi0785 & ~n18477;
  assign n18479 = ~pi0785 & ~n18465;
  assign n18480 = ~n18478 & ~n18479;
  assign n18481 = ~pi0618 & ~n18480;
  assign n18482 = ~pi1154 & ~n18449;
  assign n18483 = ~n18481 & n18482;
  assign n18484 = ~pi0627 & ~n18420;
  assign n18485 = ~n18483 & n18484;
  assign n18486 = ~pi0618 & n18395;
  assign n18487 = pi0618 & ~n18480;
  assign n18488 = pi1154 & ~n18486;
  assign n18489 = ~n18487 & n18488;
  assign n18490 = pi0627 & ~n18422;
  assign n18491 = ~n18489 & n18490;
  assign n18492 = ~n18485 & ~n18491;
  assign n18493 = pi0781 & ~n18492;
  assign n18494 = ~pi0781 & ~n18480;
  assign n18495 = ~n18493 & ~n18494;
  assign n18496 = ~pi0789 & n18495;
  assign n18497 = ~pi0619 & ~n18495;
  assign n18498 = pi0619 & n18396;
  assign n18499 = ~pi1159 & ~n18498;
  assign n18500 = ~n18497 & n18499;
  assign n18501 = ~pi0648 & ~n18430;
  assign n18502 = ~n18500 & n18501;
  assign n18503 = ~pi0619 & n18396;
  assign n18504 = pi0619 & ~n18495;
  assign n18505 = pi1159 & ~n18503;
  assign n18506 = ~n18504 & n18505;
  assign n18507 = pi0648 & ~n18434;
  assign n18508 = ~n18506 & n18507;
  assign n18509 = pi0789 & ~n18502;
  assign n18510 = ~n18508 & n18509;
  assign n18511 = n17970 & ~n18496;
  assign n18512 = ~n18510 & n18511;
  assign n18513 = ~n18448 & ~n18512;
  assign n18514 = ~pi0628 & ~n18513;
  assign n18515 = ~pi0788 & ~n18437;
  assign n18516 = pi0788 & ~n18445;
  assign n18517 = ~n18515 & ~n18516;
  assign n18518 = pi0628 & n18517;
  assign n18519 = ~pi1156 & ~n18518;
  assign n18520 = ~n18514 & n18519;
  assign n18521 = ~pi0629 & ~n18404;
  assign n18522 = ~n18520 & n18521;
  assign n18523 = ~n17997 & n18398;
  assign n18524 = ~pi1156 & ~n18523;
  assign n18525 = ~pi0628 & n18517;
  assign n18526 = pi0628 & ~n18513;
  assign n18527 = pi1156 & ~n18525;
  assign n18528 = ~n18526 & n18527;
  assign n18529 = pi0629 & ~n18524;
  assign n18530 = ~n18528 & n18529;
  assign n18531 = ~n18522 & ~n18530;
  assign n18532 = pi0792 & ~n18531;
  assign n18533 = ~pi0792 & ~n18513;
  assign n18534 = ~n18532 & ~n18533;
  assign n18535 = ~pi0647 & ~n18534;
  assign n18536 = ~n17779 & n18517;
  assign n18537 = n17779 & n18382;
  assign n18538 = ~n18536 & ~n18537;
  assign n18539 = pi0647 & ~n18538;
  assign n18540 = ~pi1157 & ~n18539;
  assign n18541 = ~n18535 & n18540;
  assign n18542 = ~pi0630 & ~n18402;
  assign n18543 = ~n18541 & n18542;
  assign n18544 = ~pi0647 & n18399;
  assign n18545 = pi0647 & n18382;
  assign n18546 = ~pi1157 & ~n18545;
  assign n18547 = ~n18544 & n18546;
  assign n18548 = pi0647 & ~n18534;
  assign n18549 = ~pi0647 & ~n18538;
  assign n18550 = pi1157 & ~n18549;
  assign n18551 = ~n18548 & n18550;
  assign n18552 = pi0630 & ~n18547;
  assign n18553 = ~n18551 & n18552;
  assign n18554 = ~n18543 & ~n18553;
  assign n18555 = pi0787 & ~n18554;
  assign n18556 = ~pi0787 & ~n18534;
  assign n18557 = ~n18555 & ~n18556;
  assign n18558 = ~pi0790 & ~n18557;
  assign n18559 = ~pi0787 & ~n18399;
  assign n18560 = ~n18402 & ~n18547;
  assign n18561 = pi0787 & ~n18560;
  assign n18562 = ~n18559 & ~n18561;
  assign n18563 = ~pi0644 & n18562;
  assign n18564 = pi0644 & ~n18557;
  assign n18565 = pi0715 & ~n18563;
  assign n18566 = ~n18564 & n18565;
  assign n18567 = n17804 & ~n18382;
  assign n18568 = ~n17804 & n18538;
  assign n18569 = ~n18567 & ~n18568;
  assign n18570 = pi0644 & n18569;
  assign n18571 = ~pi0644 & n18382;
  assign n18572 = ~pi0715 & ~n18571;
  assign n18573 = ~n18570 & n18572;
  assign n18574 = pi1160 & ~n18573;
  assign n18575 = ~n18566 & n18574;
  assign n18576 = ~pi0644 & n18569;
  assign n18577 = pi0644 & n18382;
  assign n18578 = pi0715 & ~n18577;
  assign n18579 = ~n18576 & n18578;
  assign n18580 = pi0644 & n18562;
  assign n18581 = ~pi0644 & ~n18557;
  assign n18582 = ~pi0715 & ~n18580;
  assign n18583 = ~n18581 & n18582;
  assign n18584 = ~pi1160 & ~n18579;
  assign n18585 = ~n18583 & n18584;
  assign n18586 = ~n18575 & ~n18585;
  assign n18587 = pi0790 & ~n18586;
  assign n18588 = pi0832 & ~n18558;
  assign n18589 = ~n18587 & n18588;
  assign po0298 = ~n18381 & ~n18589;
  assign n18591 = n2571 & ~n17051;
  assign n18592 = pi0142 & ~n18591;
  assign n18593 = pi0039 & ~n17025;
  assign n18594 = pi0142 & ~n18147;
  assign n18595 = ~n18593 & n18594;
  assign n18596 = pi0142 & ~n16970;
  assign n18597 = ~n6242 & ~n18596;
  assign n18598 = pi0142 & ~n16990;
  assign n18599 = n6242 & ~n18598;
  assign n18600 = pi0215 & ~n18599;
  assign n18601 = ~n18597 & n18600;
  assign n18602 = pi0142 & ~n16653;
  assign n18603 = n3448 & ~n18602;
  assign n18604 = pi0142 & ~n17018;
  assign n18605 = ~n6242 & ~n18604;
  assign n18606 = pi0142 & ~n17011;
  assign n18607 = n6242 & ~n18606;
  assign n18608 = ~n18605 & ~n18607;
  assign n18609 = ~n3448 & ~n18608;
  assign n18610 = ~pi0215 & ~n18603;
  assign n18611 = ~n18609 & n18610;
  assign n18612 = ~n18601 & ~n18611;
  assign n18613 = pi0039 & pi0299;
  assign n18614 = ~n18612 & n18613;
  assign n18615 = ~n18595 & ~n18614;
  assign n18616 = n14873 & ~n18615;
  assign n18617 = ~n18592 & ~n18616;
  assign n18618 = n16639 & ~n18617;
  assign n18619 = pi0142 & ~n2571;
  assign n18620 = pi0039 & pi0142;
  assign n18621 = pi0038 & ~n18620;
  assign n18622 = pi0142 & ~n16667;
  assign n18623 = pi0735 & n16645;
  assign n18624 = n2521 & n18623;
  assign n18625 = ~n18622 & ~n18624;
  assign n18626 = ~pi0039 & ~n18625;
  assign n18627 = n18621 & ~n18626;
  assign n18628 = ~pi0142 & ~n16926;
  assign n18629 = pi0142 & n16948;
  assign n18630 = pi0735 & ~n18628;
  assign n18631 = ~n18629 & n18630;
  assign n18632 = pi0142 & ~pi0735;
  assign n18633 = ~n16958 & n18632;
  assign n18634 = ~n18631 & ~n18633;
  assign n18635 = ~pi0039 & ~n18634;
  assign n18636 = n16652 & n18623;
  assign n18637 = ~n18602 & ~n18636;
  assign n18638 = n3448 & n18637;
  assign n18639 = ~pi0142 & ~n16694;
  assign n18640 = pi0142 & ~n16791;
  assign n18641 = ~n18639 & ~n18640;
  assign n18642 = pi0735 & ~n18641;
  assign n18643 = ~pi0735 & ~n18606;
  assign n18644 = ~n18642 & ~n18643;
  assign n18645 = n6242 & n18644;
  assign n18646 = ~pi0142 & n16705;
  assign n18647 = pi0142 & n16763;
  assign n18648 = ~n18646 & ~n18647;
  assign n18649 = pi0735 & ~n18648;
  assign n18650 = ~pi0735 & ~n18604;
  assign n18651 = ~n18649 & ~n18650;
  assign n18652 = ~n6242 & n18651;
  assign n18653 = ~n3448 & ~n18652;
  assign n18654 = ~n18645 & n18653;
  assign n18655 = ~pi0215 & ~n18638;
  assign n18656 = ~n18654 & n18655;
  assign n18657 = ~pi0735 & ~n18598;
  assign n18658 = ~pi0142 & n17560;
  assign n18659 = pi0142 & ~n16811;
  assign n18660 = pi0735 & ~n18658;
  assign n18661 = ~n18659 & n18660;
  assign n18662 = ~n18657 & ~n18661;
  assign n18663 = n6242 & ~n18662;
  assign n18664 = ~pi0735 & ~n18596;
  assign n18665 = pi0142 & ~n16819;
  assign n18666 = n17559 & n18658;
  assign n18667 = pi0735 & ~n18666;
  assign n18668 = ~n18665 & n18667;
  assign n18669 = ~n18664 & ~n18668;
  assign n18670 = ~n6242 & ~n18669;
  assign n18671 = pi0215 & ~n18663;
  assign n18672 = ~n18670 & n18671;
  assign n18673 = pi0299 & ~n18672;
  assign n18674 = ~n18656 & n18673;
  assign n18675 = n6205 & ~n18662;
  assign n18676 = ~n6205 & ~n18669;
  assign n18677 = pi0223 & ~n18675;
  assign n18678 = ~n18676 & n18677;
  assign n18679 = n2603 & n18637;
  assign n18680 = n6205 & n18644;
  assign n18681 = ~n6205 & n18651;
  assign n18682 = ~n2603 & ~n18681;
  assign n18683 = ~n18680 & n18682;
  assign n18684 = ~pi0223 & ~n18679;
  assign n18685 = ~n18683 & n18684;
  assign n18686 = ~pi0299 & ~n18678;
  assign n18687 = ~n18685 & n18686;
  assign n18688 = pi0039 & ~n18674;
  assign n18689 = ~n18687 & n18688;
  assign n18690 = ~pi0038 & ~n18635;
  assign n18691 = ~n18689 & n18690;
  assign n18692 = n2571 & ~n18627;
  assign n18693 = ~n18691 & n18692;
  assign n18694 = ~n18619 & ~n18693;
  assign n18695 = ~pi0778 & ~n18694;
  assign n18696 = ~pi0625 & n18694;
  assign n18697 = pi0625 & n18617;
  assign n18698 = ~pi1153 & ~n18697;
  assign n18699 = ~n18696 & n18698;
  assign n18700 = ~pi0625 & n18617;
  assign n18701 = pi0625 & n18694;
  assign n18702 = pi1153 & ~n18700;
  assign n18703 = ~n18701 & n18702;
  assign n18704 = ~n18699 & ~n18703;
  assign n18705 = pi0778 & ~n18704;
  assign n18706 = ~n18695 & ~n18705;
  assign n18707 = ~n17075 & n18706;
  assign n18708 = n17075 & n18617;
  assign n18709 = ~n18707 & ~n18708;
  assign n18710 = ~n16639 & n18709;
  assign n18711 = ~n18618 & ~n18710;
  assign n18712 = ~n16635 & n18711;
  assign n18713 = n16635 & n18617;
  assign n18714 = ~n18712 & ~n18713;
  assign n18715 = ~n16631 & ~n18714;
  assign n18716 = n16631 & n18617;
  assign n18717 = ~n18715 & ~n18716;
  assign n18718 = ~pi0792 & n18717;
  assign n18719 = ~pi0628 & n18617;
  assign n18720 = pi0628 & ~n18717;
  assign n18721 = pi1156 & ~n18719;
  assign n18722 = ~n18720 & n18721;
  assign n18723 = pi0628 & n18617;
  assign n18724 = ~pi0628 & ~n18717;
  assign n18725 = ~pi1156 & ~n18723;
  assign n18726 = ~n18724 & n18725;
  assign n18727 = ~n18722 & ~n18726;
  assign n18728 = pi0792 & ~n18727;
  assign n18729 = ~n18718 & ~n18728;
  assign n18730 = ~pi0787 & ~n18729;
  assign n18731 = ~pi0647 & n18617;
  assign n18732 = pi0647 & n18729;
  assign n18733 = pi1157 & ~n18731;
  assign n18734 = ~n18732 & n18733;
  assign n18735 = ~pi0647 & n18729;
  assign n18736 = pi0647 & n18617;
  assign n18737 = ~pi1157 & ~n18736;
  assign n18738 = ~n18735 & n18737;
  assign n18739 = ~n18734 & ~n18738;
  assign n18740 = pi0787 & ~n18739;
  assign n18741 = ~n18730 & ~n18740;
  assign n18742 = ~pi0644 & n18741;
  assign n18743 = ~pi0618 & n18617;
  assign n18744 = pi0743 & n17244;
  assign n18745 = n2521 & n18744;
  assign n18746 = ~n18622 & ~n18745;
  assign n18747 = ~pi0039 & ~n18746;
  assign n18748 = n18621 & ~n18747;
  assign n18749 = pi0142 & ~pi0743;
  assign n18750 = ~n16930 & n18749;
  assign n18751 = ~pi0142 & ~n17226;
  assign n18752 = pi0142 & ~n17137;
  assign n18753 = pi0743 & ~n18751;
  assign n18754 = ~n18752 & n18753;
  assign n18755 = ~pi0299 & ~n18750;
  assign n18756 = ~n18754 & n18755;
  assign n18757 = ~pi0142 & ~n17231;
  assign n18758 = pi0142 & ~n16941;
  assign n18759 = ~pi0743 & ~n18758;
  assign n18760 = pi0142 & n17124;
  assign n18761 = ~n18757 & ~n18759;
  assign n18762 = ~n18760 & n18761;
  assign n18763 = pi0299 & ~n18762;
  assign n18764 = ~n18756 & ~n18763;
  assign n18765 = ~pi0039 & n18764;
  assign n18766 = ~pi0743 & ~n18596;
  assign n18767 = pi0142 & ~n17189;
  assign n18768 = pi0743 & n17558;
  assign n18769 = ~n18767 & n18768;
  assign n18770 = ~n18766 & ~n18769;
  assign n18771 = ~n6205 & ~n18770;
  assign n18772 = ~pi0743 & ~n18598;
  assign n18773 = pi0142 & n17200;
  assign n18774 = pi0743 & n17241;
  assign n18775 = ~n18773 & n18774;
  assign n18776 = ~n18772 & ~n18775;
  assign n18777 = n6205 & ~n18776;
  assign n18778 = pi0223 & ~n18777;
  assign n18779 = ~n18771 & n18778;
  assign n18780 = ~pi0743 & ~n18604;
  assign n18781 = pi0142 & ~n17157;
  assign n18782 = pi0743 & ~n17254;
  assign n18783 = ~n18781 & n18782;
  assign n18784 = ~n18780 & ~n18783;
  assign n18785 = ~n6205 & n18784;
  assign n18786 = ~pi0142 & n17252;
  assign n18787 = pi0142 & n17175;
  assign n18788 = ~n18786 & ~n18787;
  assign n18789 = pi0743 & ~n18788;
  assign n18790 = ~pi0743 & ~n18606;
  assign n18791 = ~n18789 & ~n18790;
  assign n18792 = n6205 & n18791;
  assign n18793 = ~n2603 & ~n18785;
  assign n18794 = ~n18792 & n18793;
  assign n18795 = pi0743 & n17235;
  assign n18796 = ~n18602 & ~n18795;
  assign n18797 = n2603 & n18796;
  assign n18798 = ~pi0223 & ~n18797;
  assign n18799 = ~n18794 & n18798;
  assign n18800 = ~pi0299 & ~n18779;
  assign n18801 = ~n18799 & n18800;
  assign n18802 = n3448 & ~n18796;
  assign n18803 = ~n6242 & n18784;
  assign n18804 = n6242 & n18791;
  assign n18805 = ~n18803 & ~n18804;
  assign n18806 = ~n3448 & ~n18805;
  assign n18807 = ~pi0215 & ~n18802;
  assign n18808 = ~n18806 & n18807;
  assign n18809 = ~n6242 & n18770;
  assign n18810 = n6242 & n18776;
  assign n18811 = pi0215 & ~n18810;
  assign n18812 = ~n18809 & n18811;
  assign n18813 = ~n18808 & ~n18812;
  assign n18814 = pi0299 & ~n18813;
  assign n18815 = pi0039 & ~n18801;
  assign n18816 = ~n18814 & n18815;
  assign n18817 = ~pi0038 & ~n18765;
  assign n18818 = ~n18816 & n18817;
  assign n18819 = n2571 & ~n18748;
  assign n18820 = ~n18818 & n18819;
  assign n18821 = ~n18619 & ~n18820;
  assign n18822 = ~n17117 & ~n18821;
  assign n18823 = n17117 & ~n18617;
  assign n18824 = ~n18822 & ~n18823;
  assign n18825 = ~pi0785 & ~n18824;
  assign n18826 = ~n17291 & ~n18617;
  assign n18827 = pi0609 & n18822;
  assign n18828 = ~n18826 & ~n18827;
  assign n18829 = pi1155 & ~n18828;
  assign n18830 = ~n17296 & ~n18617;
  assign n18831 = ~pi0609 & n18822;
  assign n18832 = ~n18830 & ~n18831;
  assign n18833 = ~pi1155 & ~n18832;
  assign n18834 = ~n18829 & ~n18833;
  assign n18835 = pi0785 & ~n18834;
  assign n18836 = ~n18825 & ~n18835;
  assign n18837 = pi0618 & n18836;
  assign n18838 = pi1154 & ~n18743;
  assign n18839 = ~n18837 & n18838;
  assign n18840 = pi0609 & n18706;
  assign n18841 = ~pi0625 & n18821;
  assign n18842 = ~pi0735 & n18764;
  assign n18843 = n16937 & n18752;
  assign n18844 = ~n16919 & n18751;
  assign n18845 = ~n18843 & ~n18844;
  assign n18846 = pi0743 & ~n18845;
  assign n18847 = pi0142 & ~n16937;
  assign n18848 = ~n17226 & n18847;
  assign n18849 = ~pi0142 & n17618;
  assign n18850 = ~pi0743 & ~n18848;
  assign n18851 = ~n18849 & n18850;
  assign n18852 = ~pi0299 & ~n18851;
  assign n18853 = ~n18846 & n18852;
  assign n18854 = ~n16924 & n18757;
  assign n18855 = ~n16945 & n18760;
  assign n18856 = ~n18854 & ~n18855;
  assign n18857 = pi0743 & ~n18856;
  assign n18858 = ~pi0142 & n17623;
  assign n18859 = pi0142 & ~n16946;
  assign n18860 = ~n17231 & n18859;
  assign n18861 = ~pi0743 & ~n18860;
  assign n18862 = ~n18858 & n18861;
  assign n18863 = pi0299 & ~n18857;
  assign n18864 = ~n18862 & n18863;
  assign n18865 = ~n18853 & ~n18864;
  assign n18866 = pi0735 & ~n18865;
  assign n18867 = ~pi0039 & ~n18842;
  assign n18868 = ~n18866 & n18867;
  assign n18869 = ~pi0142 & ~n17556;
  assign n18870 = pi0142 & ~n17519;
  assign n18871 = pi0743 & ~n18869;
  assign n18872 = ~n18870 & n18871;
  assign n18873 = ~pi0142 & n17448;
  assign n18874 = pi0142 & n17351;
  assign n18875 = ~pi0743 & ~n18873;
  assign n18876 = ~n18874 & n18875;
  assign n18877 = ~n18872 & ~n18876;
  assign n18878 = pi0735 & ~n18877;
  assign n18879 = ~pi0735 & n18776;
  assign n18880 = ~n18878 & ~n18879;
  assign n18881 = n6205 & n18880;
  assign n18882 = ~pi0142 & n17562;
  assign n18883 = pi0142 & n17527;
  assign n18884 = pi0743 & ~n18882;
  assign n18885 = ~n18883 & n18884;
  assign n18886 = ~pi0142 & ~n17463;
  assign n18887 = pi0142 & n17333;
  assign n18888 = ~pi0743 & ~n18887;
  assign n18889 = ~n18886 & n18888;
  assign n18890 = ~n18885 & ~n18889;
  assign n18891 = pi0735 & ~n18890;
  assign n18892 = ~pi0735 & n18770;
  assign n18893 = ~n18891 & ~n18892;
  assign n18894 = ~n6205 & n18893;
  assign n18895 = pi0223 & ~n18881;
  assign n18896 = ~n18894 & n18895;
  assign n18897 = ~pi0735 & n18796;
  assign n18898 = ~n17645 & n18746;
  assign n18899 = ~n16650 & ~n18898;
  assign n18900 = pi0735 & ~n18899;
  assign n18901 = ~n18602 & n18900;
  assign n18902 = ~n18897 & ~n18901;
  assign n18903 = n2603 & ~n18902;
  assign n18904 = pi0142 & n17510;
  assign n18905 = ~pi0142 & ~n17573;
  assign n18906 = pi0743 & ~n18904;
  assign n18907 = ~n18905 & n18906;
  assign n18908 = ~pi0142 & n17420;
  assign n18909 = pi0142 & n17373;
  assign n18910 = ~pi0743 & ~n18908;
  assign n18911 = ~n18909 & n18910;
  assign n18912 = ~n18907 & ~n18911;
  assign n18913 = pi0735 & ~n18912;
  assign n18914 = ~pi0735 & n18791;
  assign n18915 = ~n18913 & ~n18914;
  assign n18916 = n6205 & ~n18915;
  assign n18917 = ~pi0142 & ~n17584;
  assign n18918 = pi0142 & n17499;
  assign n18919 = pi0743 & ~n18918;
  assign n18920 = ~n18917 & n18919;
  assign n18921 = ~pi0142 & ~n17438;
  assign n18922 = pi0142 & n17383;
  assign n18923 = ~pi0743 & ~n18922;
  assign n18924 = ~n18921 & n18923;
  assign n18925 = ~n18920 & ~n18924;
  assign n18926 = pi0735 & ~n18925;
  assign n18927 = ~pi0735 & n18784;
  assign n18928 = ~n18926 & ~n18927;
  assign n18929 = ~n6205 & ~n18928;
  assign n18930 = ~n2603 & ~n18929;
  assign n18931 = ~n18916 & n18930;
  assign n18932 = ~pi0223 & ~n18903;
  assign n18933 = ~n18931 & n18932;
  assign n18934 = ~n18896 & ~n18933;
  assign n18935 = ~pi0299 & ~n18934;
  assign n18936 = n6242 & n18880;
  assign n18937 = ~n6242 & n18893;
  assign n18938 = pi0215 & ~n18936;
  assign n18939 = ~n18937 & n18938;
  assign n18940 = n3448 & ~n18902;
  assign n18941 = ~n6242 & ~n18928;
  assign n18942 = n6242 & ~n18915;
  assign n18943 = ~n3448 & ~n18941;
  assign n18944 = ~n18942 & n18943;
  assign n18945 = ~pi0215 & ~n18940;
  assign n18946 = ~n18944 & n18945;
  assign n18947 = ~n18939 & ~n18946;
  assign n18948 = pi0299 & ~n18947;
  assign n18949 = pi0039 & ~n18935;
  assign n18950 = ~n18948 & n18949;
  assign n18951 = ~n18868 & ~n18950;
  assign n18952 = ~pi0038 & ~n18951;
  assign n18953 = pi0735 & n17645;
  assign n18954 = n18746 & ~n18953;
  assign n18955 = ~pi0039 & ~n18954;
  assign n18956 = n18621 & ~n18955;
  assign n18957 = n2571 & ~n18956;
  assign n18958 = ~n18952 & n18957;
  assign n18959 = ~n18619 & ~n18958;
  assign n18960 = pi0625 & n18959;
  assign n18961 = pi1153 & ~n18841;
  assign n18962 = ~n18960 & n18961;
  assign n18963 = pi0608 & ~n18699;
  assign n18964 = ~n18962 & n18963;
  assign n18965 = ~pi0625 & n18959;
  assign n18966 = pi0625 & n18821;
  assign n18967 = ~pi1153 & ~n18966;
  assign n18968 = ~n18965 & n18967;
  assign n18969 = ~pi0608 & ~n18703;
  assign n18970 = ~n18968 & n18969;
  assign n18971 = ~n18964 & ~n18970;
  assign n18972 = pi0778 & ~n18971;
  assign n18973 = ~pi0778 & n18959;
  assign n18974 = ~n18972 & ~n18973;
  assign n18975 = ~pi0609 & ~n18974;
  assign n18976 = ~pi1155 & ~n18840;
  assign n18977 = ~n18975 & n18976;
  assign n18978 = ~pi0660 & ~n18829;
  assign n18979 = ~n18977 & n18978;
  assign n18980 = ~pi0609 & n18706;
  assign n18981 = pi0609 & ~n18974;
  assign n18982 = pi1155 & ~n18980;
  assign n18983 = ~n18981 & n18982;
  assign n18984 = pi0660 & ~n18833;
  assign n18985 = ~n18983 & n18984;
  assign n18986 = ~n18979 & ~n18985;
  assign n18987 = pi0785 & ~n18986;
  assign n18988 = ~pi0785 & ~n18974;
  assign n18989 = ~n18987 & ~n18988;
  assign n18990 = ~pi0618 & ~n18989;
  assign n18991 = pi0618 & ~n18709;
  assign n18992 = ~pi1154 & ~n18991;
  assign n18993 = ~n18990 & n18992;
  assign n18994 = ~pi0627 & ~n18839;
  assign n18995 = ~n18993 & n18994;
  assign n18996 = ~pi0618 & n18836;
  assign n18997 = pi0618 & n18617;
  assign n18998 = ~pi1154 & ~n18997;
  assign n18999 = ~n18996 & n18998;
  assign n19000 = pi0618 & ~n18989;
  assign n19001 = ~pi0618 & ~n18709;
  assign n19002 = pi1154 & ~n19001;
  assign n19003 = ~n19000 & n19002;
  assign n19004 = pi0627 & ~n18999;
  assign n19005 = ~n19003 & n19004;
  assign n19006 = ~n18995 & ~n19005;
  assign n19007 = pi0781 & ~n19006;
  assign n19008 = ~pi0781 & ~n18989;
  assign n19009 = ~n19007 & ~n19008;
  assign n19010 = ~pi0619 & ~n19009;
  assign n19011 = pi0619 & n18711;
  assign n19012 = ~pi1159 & ~n19011;
  assign n19013 = ~n19010 & n19012;
  assign n19014 = ~pi0619 & n18617;
  assign n19015 = ~pi0781 & ~n18836;
  assign n19016 = ~n18839 & ~n18999;
  assign n19017 = pi0781 & ~n19016;
  assign n19018 = ~n19015 & ~n19017;
  assign n19019 = pi0619 & n19018;
  assign n19020 = pi1159 & ~n19014;
  assign n19021 = ~n19019 & n19020;
  assign n19022 = ~pi0648 & ~n19021;
  assign n19023 = ~n19013 & n19022;
  assign n19024 = pi0619 & ~n19009;
  assign n19025 = ~pi0619 & n18711;
  assign n19026 = pi1159 & ~n19025;
  assign n19027 = ~n19024 & n19026;
  assign n19028 = ~pi0619 & n19018;
  assign n19029 = pi0619 & n18617;
  assign n19030 = ~pi1159 & ~n19029;
  assign n19031 = ~n19028 & n19030;
  assign n19032 = pi0648 & ~n19031;
  assign n19033 = ~n19027 & n19032;
  assign n19034 = ~n19023 & ~n19033;
  assign n19035 = pi0789 & ~n19034;
  assign n19036 = ~pi0789 & ~n19009;
  assign n19037 = ~n19035 & ~n19036;
  assign n19038 = ~pi0788 & n19037;
  assign n19039 = ~pi0626 & n19037;
  assign n19040 = pi0626 & n18714;
  assign n19041 = ~pi0641 & ~n19040;
  assign n19042 = ~n19039 & n19041;
  assign n19043 = ~pi0789 & ~n19018;
  assign n19044 = ~n19021 & ~n19031;
  assign n19045 = pi0789 & ~n19044;
  assign n19046 = ~n19043 & ~n19045;
  assign n19047 = ~pi0626 & n19046;
  assign n19048 = pi0626 & n18617;
  assign n19049 = ~pi1158 & ~n19048;
  assign n19050 = ~n19047 & n19049;
  assign n19051 = ~n17730 & ~n19050;
  assign n19052 = ~n19042 & ~n19051;
  assign n19053 = pi0626 & n19037;
  assign n19054 = ~pi0626 & n18714;
  assign n19055 = pi0641 & ~n19054;
  assign n19056 = ~n19053 & n19055;
  assign n19057 = ~pi0626 & n18617;
  assign n19058 = pi0626 & n19046;
  assign n19059 = pi1158 & ~n19057;
  assign n19060 = ~n19058 & n19059;
  assign n19061 = ~n17745 & ~n19060;
  assign n19062 = ~n19056 & ~n19061;
  assign n19063 = ~n19052 & ~n19062;
  assign n19064 = pi0788 & ~n19063;
  assign n19065 = ~n19038 & ~n19064;
  assign n19066 = ~pi0628 & n19065;
  assign n19067 = ~n19050 & ~n19060;
  assign n19068 = pi0788 & ~n19067;
  assign n19069 = ~pi0788 & ~n19046;
  assign n19070 = ~n19068 & ~n19069;
  assign n19071 = pi0628 & n19070;
  assign n19072 = ~pi1156 & ~n19071;
  assign n19073 = ~n19066 & n19072;
  assign n19074 = ~pi0629 & ~n18722;
  assign n19075 = ~n19073 & n19074;
  assign n19076 = pi0628 & n19065;
  assign n19077 = ~pi0628 & n19070;
  assign n19078 = pi1156 & ~n19077;
  assign n19079 = ~n19076 & n19078;
  assign n19080 = pi0629 & ~n18726;
  assign n19081 = ~n19079 & n19080;
  assign n19082 = ~n19075 & ~n19081;
  assign n19083 = pi0792 & ~n19082;
  assign n19084 = ~pi0792 & n19065;
  assign n19085 = ~n19083 & ~n19084;
  assign n19086 = ~pi0647 & ~n19085;
  assign n19087 = ~n17779 & n19070;
  assign n19088 = n17779 & n18617;
  assign n19089 = ~n19087 & ~n19088;
  assign n19090 = pi0647 & ~n19089;
  assign n19091 = ~pi1157 & ~n19090;
  assign n19092 = ~n19086 & n19091;
  assign n19093 = ~pi0630 & ~n18734;
  assign n19094 = ~n19092 & n19093;
  assign n19095 = pi0647 & ~n19085;
  assign n19096 = ~pi0647 & ~n19089;
  assign n19097 = pi1157 & ~n19096;
  assign n19098 = ~n19095 & n19097;
  assign n19099 = pi0630 & ~n18738;
  assign n19100 = ~n19098 & n19099;
  assign n19101 = ~n19094 & ~n19100;
  assign n19102 = pi0787 & ~n19101;
  assign n19103 = ~pi0787 & ~n19085;
  assign n19104 = ~n19102 & ~n19103;
  assign n19105 = pi0644 & ~n19104;
  assign n19106 = pi0715 & ~n18742;
  assign n19107 = ~n19105 & n19106;
  assign n19108 = n17804 & ~n18617;
  assign n19109 = ~n17804 & n19089;
  assign n19110 = ~n19108 & ~n19109;
  assign n19111 = pi0644 & n19110;
  assign n19112 = ~pi0644 & n18617;
  assign n19113 = ~pi0715 & ~n19112;
  assign n19114 = ~n19111 & n19113;
  assign n19115 = pi1160 & ~n19114;
  assign n19116 = ~n19107 & n19115;
  assign n19117 = ~pi0644 & ~n19104;
  assign n19118 = pi0644 & n18741;
  assign n19119 = ~pi0715 & ~n19118;
  assign n19120 = ~n19117 & n19119;
  assign n19121 = ~pi0644 & n19110;
  assign n19122 = pi0644 & n18617;
  assign n19123 = pi0715 & ~n19122;
  assign n19124 = ~n19121 & n19123;
  assign n19125 = ~pi1160 & ~n19124;
  assign n19126 = ~n19120 & n19125;
  assign n19127 = pi0790 & ~n19116;
  assign n19128 = ~n19126 & n19127;
  assign n19129 = ~pi0790 & n19104;
  assign n19130 = n6305 & ~n19129;
  assign n19131 = ~n19128 & n19130;
  assign n19132 = ~pi0142 & ~n6305;
  assign n19133 = ~pi0057 & ~n19132;
  assign n19134 = ~n19131 & n19133;
  assign n19135 = pi0057 & pi0142;
  assign n19136 = ~pi0832 & ~n19135;
  assign n19137 = ~n19134 & n19136;
  assign n19138 = pi0142 & ~n2926;
  assign n19139 = pi0628 & pi1156;
  assign n19140 = ~pi0628 & ~pi1156;
  assign n19141 = pi0792 & ~n19139;
  assign n19142 = ~n19140 & n19141;
  assign n19143 = ~pi0625 & pi1153;
  assign n19144 = pi0625 & ~pi1153;
  assign n19145 = ~n19143 & ~n19144;
  assign n19146 = pi0778 & ~n19145;
  assign n19147 = n18623 & ~n19146;
  assign n19148 = ~n19138 & ~n19147;
  assign n19149 = ~n16631 & ~n16635;
  assign n19150 = ~n16639 & ~n17075;
  assign n19151 = n19149 & n19150;
  assign n19152 = ~n19148 & n19151;
  assign n19153 = ~n19142 & n19152;
  assign n19154 = pi0647 & n19153;
  assign n19155 = pi1157 & ~n19138;
  assign n19156 = ~n19154 & n19155;
  assign n19157 = pi0628 & n19152;
  assign n19158 = ~n19138 & ~n19157;
  assign n19159 = pi1156 & ~n19158;
  assign n19160 = ~pi0626 & n19138;
  assign n19161 = ~n17117 & n18744;
  assign n19162 = pi0609 & n19161;
  assign n19163 = pi1155 & ~n19138;
  assign n19164 = ~n19162 & n19163;
  assign n19165 = ~pi0609 & n19161;
  assign n19166 = ~pi1155 & ~n19138;
  assign n19167 = ~n19165 & n19166;
  assign n19168 = ~n19164 & ~n19167;
  assign n19169 = pi0785 & ~n19168;
  assign n19170 = ~pi0785 & ~n19138;
  assign n19171 = ~n19161 & n19170;
  assign n19172 = ~n19169 & ~n19171;
  assign n19173 = ~pi0781 & ~n19172;
  assign n19174 = ~pi0618 & n19138;
  assign n19175 = pi0618 & n19172;
  assign n19176 = pi1154 & ~n19174;
  assign n19177 = ~n19175 & n19176;
  assign n19178 = ~pi0618 & n19172;
  assign n19179 = pi0618 & n19138;
  assign n19180 = ~pi1154 & ~n19179;
  assign n19181 = ~n19178 & n19180;
  assign n19182 = ~n19177 & ~n19181;
  assign n19183 = pi0781 & ~n19182;
  assign n19184 = ~n19173 & ~n19183;
  assign n19185 = ~pi0789 & ~n19184;
  assign n19186 = ~pi0619 & n19138;
  assign n19187 = pi0619 & n19184;
  assign n19188 = pi1159 & ~n19186;
  assign n19189 = ~n19187 & n19188;
  assign n19190 = ~pi0619 & n19184;
  assign n19191 = pi0619 & n19138;
  assign n19192 = ~pi1159 & ~n19191;
  assign n19193 = ~n19190 & n19192;
  assign n19194 = ~n19189 & ~n19193;
  assign n19195 = pi0789 & ~n19194;
  assign n19196 = ~n19185 & ~n19195;
  assign n19197 = pi0626 & n19196;
  assign n19198 = pi1158 & ~n19160;
  assign n19199 = ~n19197 & n19198;
  assign n19200 = ~pi0626 & n19196;
  assign n19201 = pi0626 & n19138;
  assign n19202 = ~pi1158 & ~n19201;
  assign n19203 = ~n19200 & n19202;
  assign n19204 = ~n19199 & ~n19203;
  assign n19205 = ~n16630 & n19204;
  assign n19206 = n16635 & ~n19138;
  assign n19207 = ~n17075 & ~n19148;
  assign n19208 = ~n16639 & n19207;
  assign n19209 = ~n19138 & ~n19208;
  assign n19210 = n17871 & ~n19206;
  assign n19211 = ~n19209 & n19210;
  assign n19212 = ~n19205 & ~n19211;
  assign n19213 = pi0788 & ~n19212;
  assign n19214 = ~n19138 & ~n19207;
  assign n19215 = pi0618 & ~n19214;
  assign n19216 = pi0625 & n18623;
  assign n19217 = pi1153 & ~n19138;
  assign n19218 = ~n19216 & n19217;
  assign n19219 = pi0735 & n17469;
  assign n19220 = pi0625 & n19219;
  assign n19221 = ~n18744 & ~n19138;
  assign n19222 = ~n19219 & n19221;
  assign n19223 = ~n19220 & ~n19222;
  assign n19224 = ~pi1153 & ~n19223;
  assign n19225 = ~pi0608 & ~n19218;
  assign n19226 = ~n19224 & n19225;
  assign n19227 = ~n18744 & ~n19220;
  assign n19228 = pi1153 & ~n19227;
  assign n19229 = ~pi0625 & ~pi1153;
  assign n19230 = n18623 & n19229;
  assign n19231 = ~n19138 & ~n19230;
  assign n19232 = ~n19228 & n19231;
  assign n19233 = pi0608 & ~n19232;
  assign n19234 = ~n19226 & ~n19233;
  assign n19235 = pi0778 & ~n19234;
  assign n19236 = ~pi0778 & ~n19222;
  assign n19237 = ~n19235 & ~n19236;
  assign n19238 = ~pi0609 & ~n19237;
  assign n19239 = pi0609 & ~n19148;
  assign n19240 = ~pi1155 & ~n19239;
  assign n19241 = ~n19238 & n19240;
  assign n19242 = ~pi0660 & ~n19164;
  assign n19243 = ~n19241 & n19242;
  assign n19244 = pi0609 & ~n19237;
  assign n19245 = ~pi0609 & ~n19148;
  assign n19246 = pi1155 & ~n19245;
  assign n19247 = ~n19244 & n19246;
  assign n19248 = pi0660 & ~n19167;
  assign n19249 = ~n19247 & n19248;
  assign n19250 = ~n19243 & ~n19249;
  assign n19251 = pi0785 & ~n19250;
  assign n19252 = ~pi0785 & ~n19237;
  assign n19253 = ~n19251 & ~n19252;
  assign n19254 = ~pi0618 & ~n19253;
  assign n19255 = ~pi1154 & ~n19215;
  assign n19256 = ~n19254 & n19255;
  assign n19257 = ~pi0627 & ~n19177;
  assign n19258 = ~n19256 & n19257;
  assign n19259 = ~pi0618 & ~n19214;
  assign n19260 = pi0618 & ~n19253;
  assign n19261 = pi1154 & ~n19259;
  assign n19262 = ~n19260 & n19261;
  assign n19263 = pi0627 & ~n19181;
  assign n19264 = ~n19262 & n19263;
  assign n19265 = ~n19258 & ~n19264;
  assign n19266 = pi0781 & ~n19265;
  assign n19267 = ~pi0781 & ~n19253;
  assign n19268 = ~n19266 & ~n19267;
  assign n19269 = ~pi0789 & n19268;
  assign n19270 = ~pi0619 & ~n19268;
  assign n19271 = pi0619 & ~n19209;
  assign n19272 = ~pi1159 & ~n19271;
  assign n19273 = ~n19270 & n19272;
  assign n19274 = ~pi0648 & ~n19189;
  assign n19275 = ~n19273 & n19274;
  assign n19276 = pi0619 & ~n19268;
  assign n19277 = ~pi0619 & ~n19209;
  assign n19278 = pi1159 & ~n19277;
  assign n19279 = ~n19276 & n19278;
  assign n19280 = pi0648 & ~n19193;
  assign n19281 = ~n19279 & n19280;
  assign n19282 = pi0789 & ~n19275;
  assign n19283 = ~n19281 & n19282;
  assign n19284 = n17970 & ~n19269;
  assign n19285 = ~n19283 & n19284;
  assign n19286 = ~n19213 & ~n19285;
  assign n19287 = ~pi0628 & n19286;
  assign n19288 = ~pi0788 & ~n19196;
  assign n19289 = pi0788 & ~n19204;
  assign n19290 = ~n19288 & ~n19289;
  assign n19291 = pi0628 & ~n19290;
  assign n19292 = ~pi1156 & ~n19291;
  assign n19293 = ~n19287 & n19292;
  assign n19294 = ~pi0629 & ~n19159;
  assign n19295 = ~n19293 & n19294;
  assign n19296 = ~pi0628 & n19152;
  assign n19297 = ~n19138 & ~n19296;
  assign n19298 = ~pi1156 & ~n19297;
  assign n19299 = pi0628 & n19286;
  assign n19300 = ~pi0628 & ~n19290;
  assign n19301 = pi1156 & ~n19300;
  assign n19302 = ~n19299 & n19301;
  assign n19303 = pi0629 & ~n19298;
  assign n19304 = ~n19302 & n19303;
  assign n19305 = ~n19295 & ~n19304;
  assign n19306 = pi0792 & ~n19305;
  assign n19307 = ~pi0792 & n19286;
  assign n19308 = ~n19306 & ~n19307;
  assign n19309 = ~pi0647 & n19308;
  assign n19310 = ~n17779 & n19290;
  assign n19311 = n17779 & n19138;
  assign n19312 = ~n19310 & ~n19311;
  assign n19313 = pi0647 & ~n19312;
  assign n19314 = ~pi1157 & ~n19313;
  assign n19315 = ~n19309 & n19314;
  assign n19316 = ~pi0630 & ~n19156;
  assign n19317 = ~n19315 & n19316;
  assign n19318 = ~pi0647 & n19153;
  assign n19319 = ~pi1157 & ~n19138;
  assign n19320 = ~n19318 & n19319;
  assign n19321 = ~pi0647 & ~n19312;
  assign n19322 = pi0647 & n19308;
  assign n19323 = pi1157 & ~n19321;
  assign n19324 = ~n19322 & n19323;
  assign n19325 = pi0630 & ~n19320;
  assign n19326 = ~n19324 & n19325;
  assign n19327 = ~n19317 & ~n19326;
  assign n19328 = pi0787 & ~n19327;
  assign n19329 = ~pi0787 & n19308;
  assign n19330 = ~n19328 & ~n19329;
  assign n19331 = ~pi0790 & ~n19330;
  assign n19332 = n17804 & ~n19138;
  assign n19333 = ~n17804 & n19312;
  assign n19334 = ~n19332 & ~n19333;
  assign n19335 = pi0644 & n19334;
  assign n19336 = ~pi0644 & n19138;
  assign n19337 = ~pi0715 & ~n19336;
  assign n19338 = ~n19335 & n19337;
  assign n19339 = ~pi0647 & pi1157;
  assign n19340 = pi0647 & ~pi1157;
  assign n19341 = ~n19339 & ~n19340;
  assign n19342 = pi0787 & ~n19341;
  assign n19343 = n19153 & ~n19342;
  assign n19344 = ~n19138 & ~n19343;
  assign n19345 = ~pi0644 & ~n19344;
  assign n19346 = pi0644 & ~n19330;
  assign n19347 = pi0715 & ~n19345;
  assign n19348 = ~n19346 & n19347;
  assign n19349 = pi1160 & ~n19338;
  assign n19350 = ~n19348 & n19349;
  assign n19351 = ~pi0644 & n19334;
  assign n19352 = pi0644 & n19138;
  assign n19353 = pi0715 & ~n19352;
  assign n19354 = ~n19351 & n19353;
  assign n19355 = pi0644 & ~n19344;
  assign n19356 = ~pi0644 & ~n19330;
  assign n19357 = ~pi0715 & ~n19355;
  assign n19358 = ~n19356 & n19357;
  assign n19359 = ~pi1160 & ~n19354;
  assign n19360 = ~n19358 & n19359;
  assign n19361 = ~n19350 & ~n19360;
  assign n19362 = pi0790 & ~n19361;
  assign n19363 = pi0832 & ~n19331;
  assign n19364 = ~n19362 & n19363;
  assign po0299 = ~n19137 & ~n19364;
  assign n19366 = ~pi0143 & ~n17059;
  assign n19367 = n16635 & ~n19366;
  assign n19368 = pi0143 & ~n2571;
  assign n19369 = ~pi0143 & ~n17052;
  assign n19370 = ~pi0687 & n19369;
  assign n19371 = ~pi0143 & ~n16641;
  assign n19372 = n16647 & ~n19371;
  assign n19373 = ~pi0143 & n18072;
  assign n19374 = pi0143 & ~n18076;
  assign n19375 = ~pi0038 & ~n19374;
  assign n19376 = ~n19373 & n19375;
  assign n19377 = pi0687 & ~n19372;
  assign n19378 = ~n19376 & n19377;
  assign n19379 = n2571 & ~n19370;
  assign n19380 = ~n19378 & n19379;
  assign n19381 = ~n19368 & ~n19380;
  assign n19382 = ~pi0778 & ~n19381;
  assign n19383 = ~pi0625 & n19366;
  assign n19384 = pi0625 & n19381;
  assign n19385 = pi1153 & ~n19383;
  assign n19386 = ~n19384 & n19385;
  assign n19387 = ~pi0625 & n19381;
  assign n19388 = pi0625 & n19366;
  assign n19389 = ~pi1153 & ~n19388;
  assign n19390 = ~n19387 & n19389;
  assign n19391 = ~n19386 & ~n19390;
  assign n19392 = pi0778 & ~n19391;
  assign n19393 = ~n19382 & ~n19392;
  assign n19394 = ~n17075 & ~n19393;
  assign n19395 = n17075 & ~n19366;
  assign n19396 = ~n19394 & ~n19395;
  assign n19397 = ~n16639 & n19396;
  assign n19398 = n16639 & n19366;
  assign n19399 = ~n19397 & ~n19398;
  assign n19400 = ~n16635 & n19399;
  assign n19401 = ~n19367 & ~n19400;
  assign n19402 = ~n16631 & n19401;
  assign n19403 = n16631 & n19366;
  assign n19404 = ~n19402 & ~n19403;
  assign n19405 = ~pi0792 & n19404;
  assign n19406 = ~pi0628 & n19366;
  assign n19407 = pi0628 & ~n19404;
  assign n19408 = pi1156 & ~n19406;
  assign n19409 = ~n19407 & n19408;
  assign n19410 = pi0628 & n19366;
  assign n19411 = ~pi0628 & ~n19404;
  assign n19412 = ~pi1156 & ~n19410;
  assign n19413 = ~n19411 & n19412;
  assign n19414 = ~n19409 & ~n19413;
  assign n19415 = pi0792 & ~n19414;
  assign n19416 = ~n19405 & ~n19415;
  assign n19417 = ~pi0787 & ~n19416;
  assign n19418 = ~pi0647 & n19366;
  assign n19419 = pi0647 & n19416;
  assign n19420 = pi1157 & ~n19418;
  assign n19421 = ~n19419 & n19420;
  assign n19422 = ~pi0647 & n19416;
  assign n19423 = pi0647 & n19366;
  assign n19424 = ~pi1157 & ~n19423;
  assign n19425 = ~n19422 & n19424;
  assign n19426 = ~n19421 & ~n19425;
  assign n19427 = pi0787 & ~n19426;
  assign n19428 = ~n19417 & ~n19427;
  assign n19429 = ~pi0644 & n19428;
  assign n19430 = ~pi0618 & n19366;
  assign n19431 = pi0774 & ~n19369;
  assign n19432 = n6135 & n17244;
  assign n19433 = pi0038 & n19432;
  assign n19434 = ~pi0038 & n17275;
  assign n19435 = pi0143 & ~n19434;
  assign n19436 = ~pi0038 & ~n17221;
  assign n19437 = n6284 & n17182;
  assign n19438 = pi0038 & ~n19437;
  assign n19439 = ~n19436 & ~n19438;
  assign n19440 = ~pi0143 & ~pi0774;
  assign n19441 = n19439 & n19440;
  assign n19442 = ~n19435 & ~n19441;
  assign n19443 = ~n19433 & ~n19442;
  assign n19444 = ~n19431 & ~n19443;
  assign n19445 = n2571 & ~n19444;
  assign n19446 = ~n19368 & ~n19445;
  assign n19447 = ~n17117 & ~n19446;
  assign n19448 = n17117 & ~n19366;
  assign n19449 = ~n19447 & ~n19448;
  assign n19450 = ~pi0785 & ~n19449;
  assign n19451 = ~n17291 & ~n19366;
  assign n19452 = pi0609 & n19447;
  assign n19453 = ~n19451 & ~n19452;
  assign n19454 = pi1155 & ~n19453;
  assign n19455 = ~n17296 & ~n19366;
  assign n19456 = ~pi0609 & n19447;
  assign n19457 = ~n19455 & ~n19456;
  assign n19458 = ~pi1155 & ~n19457;
  assign n19459 = ~n19454 & ~n19458;
  assign n19460 = pi0785 & ~n19459;
  assign n19461 = ~n19450 & ~n19460;
  assign n19462 = pi0618 & n19461;
  assign n19463 = pi1154 & ~n19430;
  assign n19464 = ~n19462 & n19463;
  assign n19465 = ~pi0039 & ~n17625;
  assign n19466 = pi0039 & ~n17485;
  assign n19467 = ~n19465 & ~n19466;
  assign n19468 = ~pi0038 & n19467;
  assign n19469 = pi0143 & n19468;
  assign n19470 = pi0038 & n18175;
  assign n19471 = n16641 & ~n17355;
  assign n19472 = pi0038 & n19471;
  assign n19473 = pi0039 & ~n17404;
  assign n19474 = ~pi0039 & ~n17612;
  assign n19475 = ~n19473 & ~n19474;
  assign n19476 = ~pi0038 & ~n19475;
  assign n19477 = ~n19472 & ~n19476;
  assign n19478 = ~pi0143 & n19477;
  assign n19479 = pi0774 & ~n19470;
  assign n19480 = ~n19469 & n19479;
  assign n19481 = ~n19478 & n19480;
  assign n19482 = ~pi0039 & ~n17629;
  assign n19483 = ~pi0038 & n19482;
  assign n19484 = pi0039 & ~n17546;
  assign n19485 = ~pi0039 & n17490;
  assign n19486 = pi0038 & ~n19485;
  assign n19487 = ~n19483 & ~n19486;
  assign n19488 = ~n19484 & n19487;
  assign n19489 = ~pi0143 & ~n19488;
  assign n19490 = n6284 & ~n17470;
  assign n19491 = pi0038 & ~n19490;
  assign n19492 = pi0039 & ~n17605;
  assign n19493 = ~n16926 & n17234;
  assign n19494 = ~n19492 & ~n19493;
  assign n19495 = ~pi0038 & ~n19494;
  assign n19496 = ~n19491 & ~n19495;
  assign n19497 = pi0143 & n19496;
  assign n19498 = ~pi0774 & ~n19489;
  assign n19499 = ~n19497 & n19498;
  assign n19500 = pi0687 & ~n19499;
  assign n19501 = ~n19481 & n19500;
  assign n19502 = ~pi0687 & n19444;
  assign n19503 = n2571 & ~n19501;
  assign n19504 = ~n19502 & n19503;
  assign n19505 = ~n19368 & ~n19504;
  assign n19506 = ~pi0625 & n19505;
  assign n19507 = pi0625 & n19446;
  assign n19508 = ~pi1153 & ~n19507;
  assign n19509 = ~n19506 & n19508;
  assign n19510 = ~pi0608 & ~n19386;
  assign n19511 = ~n19509 & n19510;
  assign n19512 = ~pi0625 & n19446;
  assign n19513 = pi0625 & n19505;
  assign n19514 = pi1153 & ~n19512;
  assign n19515 = ~n19513 & n19514;
  assign n19516 = pi0608 & ~n19390;
  assign n19517 = ~n19515 & n19516;
  assign n19518 = ~n19511 & ~n19517;
  assign n19519 = pi0778 & ~n19518;
  assign n19520 = ~pi0778 & n19505;
  assign n19521 = ~n19519 & ~n19520;
  assign n19522 = ~pi0609 & ~n19521;
  assign n19523 = pi0609 & n19393;
  assign n19524 = ~pi1155 & ~n19523;
  assign n19525 = ~n19522 & n19524;
  assign n19526 = ~pi0660 & ~n19454;
  assign n19527 = ~n19525 & n19526;
  assign n19528 = ~pi0609 & n19393;
  assign n19529 = pi0609 & ~n19521;
  assign n19530 = pi1155 & ~n19528;
  assign n19531 = ~n19529 & n19530;
  assign n19532 = pi0660 & ~n19458;
  assign n19533 = ~n19531 & n19532;
  assign n19534 = ~n19527 & ~n19533;
  assign n19535 = pi0785 & ~n19534;
  assign n19536 = ~pi0785 & ~n19521;
  assign n19537 = ~n19535 & ~n19536;
  assign n19538 = ~pi0618 & ~n19537;
  assign n19539 = pi0618 & n19396;
  assign n19540 = ~pi1154 & ~n19539;
  assign n19541 = ~n19538 & n19540;
  assign n19542 = ~pi0627 & ~n19464;
  assign n19543 = ~n19541 & n19542;
  assign n19544 = ~pi0618 & n19461;
  assign n19545 = pi0618 & n19366;
  assign n19546 = ~pi1154 & ~n19545;
  assign n19547 = ~n19544 & n19546;
  assign n19548 = ~pi0618 & n19396;
  assign n19549 = pi0618 & ~n19537;
  assign n19550 = pi1154 & ~n19548;
  assign n19551 = ~n19549 & n19550;
  assign n19552 = pi0627 & ~n19547;
  assign n19553 = ~n19551 & n19552;
  assign n19554 = ~n19543 & ~n19553;
  assign n19555 = pi0781 & ~n19554;
  assign n19556 = ~pi0781 & ~n19537;
  assign n19557 = ~n19555 & ~n19556;
  assign n19558 = ~pi0619 & ~n19557;
  assign n19559 = pi0619 & ~n19399;
  assign n19560 = ~pi1159 & ~n19559;
  assign n19561 = ~n19558 & n19560;
  assign n19562 = ~pi0619 & n19366;
  assign n19563 = ~pi0781 & ~n19461;
  assign n19564 = ~n19464 & ~n19547;
  assign n19565 = pi0781 & ~n19564;
  assign n19566 = ~n19563 & ~n19565;
  assign n19567 = pi0619 & n19566;
  assign n19568 = pi1159 & ~n19562;
  assign n19569 = ~n19567 & n19568;
  assign n19570 = ~pi0648 & ~n19569;
  assign n19571 = ~n19561 & n19570;
  assign n19572 = pi0619 & ~n19557;
  assign n19573 = ~pi0619 & ~n19399;
  assign n19574 = pi1159 & ~n19573;
  assign n19575 = ~n19572 & n19574;
  assign n19576 = ~pi0619 & n19566;
  assign n19577 = pi0619 & n19366;
  assign n19578 = ~pi1159 & ~n19577;
  assign n19579 = ~n19576 & n19578;
  assign n19580 = pi0648 & ~n19579;
  assign n19581 = ~n19575 & n19580;
  assign n19582 = ~n19571 & ~n19581;
  assign n19583 = pi0789 & ~n19582;
  assign n19584 = ~pi0789 & ~n19557;
  assign n19585 = ~n19583 & ~n19584;
  assign n19586 = ~pi0788 & n19585;
  assign n19587 = ~pi0626 & n19585;
  assign n19588 = pi0626 & ~n19401;
  assign n19589 = ~pi0641 & ~n19588;
  assign n19590 = ~n19587 & n19589;
  assign n19591 = ~pi0789 & ~n19566;
  assign n19592 = ~n19569 & ~n19579;
  assign n19593 = pi0789 & ~n19592;
  assign n19594 = ~n19591 & ~n19593;
  assign n19595 = ~pi0626 & n19594;
  assign n19596 = pi0626 & n19366;
  assign n19597 = ~pi1158 & ~n19596;
  assign n19598 = ~n19595 & n19597;
  assign n19599 = ~n17730 & ~n19598;
  assign n19600 = ~n19590 & ~n19599;
  assign n19601 = pi0626 & n19585;
  assign n19602 = ~pi0626 & ~n19401;
  assign n19603 = pi0641 & ~n19602;
  assign n19604 = ~n19601 & n19603;
  assign n19605 = ~pi0626 & n19366;
  assign n19606 = pi0626 & n19594;
  assign n19607 = pi1158 & ~n19605;
  assign n19608 = ~n19606 & n19607;
  assign n19609 = ~n17745 & ~n19608;
  assign n19610 = ~n19604 & ~n19609;
  assign n19611 = ~n19600 & ~n19610;
  assign n19612 = pi0788 & ~n19611;
  assign n19613 = ~n19586 & ~n19612;
  assign n19614 = ~pi0628 & n19613;
  assign n19615 = ~n19598 & ~n19608;
  assign n19616 = pi0788 & ~n19615;
  assign n19617 = ~pi0788 & ~n19594;
  assign n19618 = ~n19616 & ~n19617;
  assign n19619 = pi0628 & n19618;
  assign n19620 = ~pi1156 & ~n19619;
  assign n19621 = ~n19614 & n19620;
  assign n19622 = ~pi0629 & ~n19409;
  assign n19623 = ~n19621 & n19622;
  assign n19624 = pi0628 & n19613;
  assign n19625 = ~pi0628 & n19618;
  assign n19626 = pi1156 & ~n19625;
  assign n19627 = ~n19624 & n19626;
  assign n19628 = pi0629 & ~n19413;
  assign n19629 = ~n19627 & n19628;
  assign n19630 = ~n19623 & ~n19629;
  assign n19631 = pi0792 & ~n19630;
  assign n19632 = ~pi0792 & n19613;
  assign n19633 = ~n19631 & ~n19632;
  assign n19634 = ~pi0647 & ~n19633;
  assign n19635 = ~n17779 & n19618;
  assign n19636 = n17779 & n19366;
  assign n19637 = ~n19635 & ~n19636;
  assign n19638 = pi0647 & ~n19637;
  assign n19639 = ~pi1157 & ~n19638;
  assign n19640 = ~n19634 & n19639;
  assign n19641 = ~pi0630 & ~n19421;
  assign n19642 = ~n19640 & n19641;
  assign n19643 = pi0647 & ~n19633;
  assign n19644 = ~pi0647 & ~n19637;
  assign n19645 = pi1157 & ~n19644;
  assign n19646 = ~n19643 & n19645;
  assign n19647 = pi0630 & ~n19425;
  assign n19648 = ~n19646 & n19647;
  assign n19649 = ~n19642 & ~n19648;
  assign n19650 = pi0787 & ~n19649;
  assign n19651 = ~pi0787 & ~n19633;
  assign n19652 = ~n19650 & ~n19651;
  assign n19653 = pi0644 & ~n19652;
  assign n19654 = pi0715 & ~n19429;
  assign n19655 = ~n19653 & n19654;
  assign n19656 = n17804 & ~n19366;
  assign n19657 = ~n17804 & n19637;
  assign n19658 = ~n19656 & ~n19657;
  assign n19659 = pi0644 & n19658;
  assign n19660 = ~pi0644 & n19366;
  assign n19661 = ~pi0715 & ~n19660;
  assign n19662 = ~n19659 & n19661;
  assign n19663 = pi1160 & ~n19662;
  assign n19664 = ~n19655 & n19663;
  assign n19665 = ~pi0644 & ~n19652;
  assign n19666 = pi0644 & n19428;
  assign n19667 = ~pi0715 & ~n19666;
  assign n19668 = ~n19665 & n19667;
  assign n19669 = ~pi0644 & n19658;
  assign n19670 = pi0644 & n19366;
  assign n19671 = pi0715 & ~n19670;
  assign n19672 = ~n19669 & n19671;
  assign n19673 = ~pi1160 & ~n19672;
  assign n19674 = ~n19668 & n19673;
  assign n19675 = pi0790 & ~n19664;
  assign n19676 = ~n19674 & n19675;
  assign n19677 = ~pi0790 & n19652;
  assign n19678 = ~po1038 & ~n19677;
  assign n19679 = ~n19676 & n19678;
  assign n19680 = ~pi0143 & po1038;
  assign n19681 = ~pi0832 & ~n19680;
  assign n19682 = ~n19679 & n19681;
  assign n19683 = ~pi0143 & ~n2926;
  assign n19684 = ~pi0647 & n19683;
  assign n19685 = pi0687 & n16645;
  assign n19686 = ~n19683 & ~n19685;
  assign n19687 = ~pi0778 & n19686;
  assign n19688 = ~pi0625 & n19685;
  assign n19689 = ~n19686 & ~n19688;
  assign n19690 = pi1153 & ~n19689;
  assign n19691 = ~pi1153 & ~n19683;
  assign n19692 = ~n19688 & n19691;
  assign n19693 = ~n19690 & ~n19692;
  assign n19694 = pi0778 & ~n19693;
  assign n19695 = ~n19687 & ~n19694;
  assign n19696 = ~n17845 & n19695;
  assign n19697 = ~n17847 & n19696;
  assign n19698 = ~n17849 & n19697;
  assign n19699 = ~n17851 & n19698;
  assign n19700 = ~n17857 & n19699;
  assign n19701 = pi0647 & n19700;
  assign n19702 = pi1157 & ~n19684;
  assign n19703 = ~n19701 & n19702;
  assign n19704 = ~n17862 & n19699;
  assign n19705 = pi1156 & ~n19704;
  assign n19706 = n17871 & n19698;
  assign n19707 = ~pi0626 & n19683;
  assign n19708 = ~pi0774 & n17244;
  assign n19709 = ~n19683 & ~n19708;
  assign n19710 = ~n17874 & ~n19709;
  assign n19711 = ~pi0785 & ~n19710;
  assign n19712 = ~n17879 & ~n19709;
  assign n19713 = pi1155 & ~n19712;
  assign n19714 = ~n17882 & n19710;
  assign n19715 = ~pi1155 & ~n19714;
  assign n19716 = ~n19713 & ~n19715;
  assign n19717 = pi0785 & ~n19716;
  assign n19718 = ~n19711 & ~n19717;
  assign n19719 = ~pi0781 & ~n19718;
  assign n19720 = ~n17889 & n19718;
  assign n19721 = pi1154 & ~n19720;
  assign n19722 = ~n17892 & n19718;
  assign n19723 = ~pi1154 & ~n19722;
  assign n19724 = ~n19721 & ~n19723;
  assign n19725 = pi0781 & ~n19724;
  assign n19726 = ~n19719 & ~n19725;
  assign n19727 = ~pi0789 & ~n19726;
  assign n19728 = ~pi0619 & n19683;
  assign n19729 = pi0619 & n19726;
  assign n19730 = pi1159 & ~n19728;
  assign n19731 = ~n19729 & n19730;
  assign n19732 = ~pi0619 & n19726;
  assign n19733 = pi0619 & n19683;
  assign n19734 = ~pi1159 & ~n19733;
  assign n19735 = ~n19732 & n19734;
  assign n19736 = ~n19731 & ~n19735;
  assign n19737 = pi0789 & ~n19736;
  assign n19738 = ~n19727 & ~n19737;
  assign n19739 = pi0626 & n19738;
  assign n19740 = pi1158 & ~n19707;
  assign n19741 = ~n19739 & n19740;
  assign n19742 = ~pi0626 & n19738;
  assign n19743 = pi0626 & n19683;
  assign n19744 = ~pi1158 & ~n19743;
  assign n19745 = ~n19742 & n19744;
  assign n19746 = ~n19741 & ~n19745;
  assign n19747 = ~n16630 & n19746;
  assign n19748 = ~n19706 & ~n19747;
  assign n19749 = pi0788 & ~n19748;
  assign n19750 = pi0618 & n19696;
  assign n19751 = pi0609 & n19695;
  assign n19752 = ~n17168 & ~n19686;
  assign n19753 = pi0625 & n19752;
  assign n19754 = n19709 & ~n19752;
  assign n19755 = ~n19753 & ~n19754;
  assign n19756 = n19691 & ~n19755;
  assign n19757 = ~pi0608 & ~n19690;
  assign n19758 = ~n19756 & n19757;
  assign n19759 = pi1153 & n19709;
  assign n19760 = ~n19753 & n19759;
  assign n19761 = pi0608 & ~n19692;
  assign n19762 = ~n19760 & n19761;
  assign n19763 = ~n19758 & ~n19762;
  assign n19764 = pi0778 & ~n19763;
  assign n19765 = ~pi0778 & ~n19754;
  assign n19766 = ~n19764 & ~n19765;
  assign n19767 = ~pi0609 & ~n19766;
  assign n19768 = ~pi1155 & ~n19751;
  assign n19769 = ~n19767 & n19768;
  assign n19770 = ~pi0660 & ~n19713;
  assign n19771 = ~n19769 & n19770;
  assign n19772 = ~pi0609 & n19695;
  assign n19773 = pi0609 & ~n19766;
  assign n19774 = pi1155 & ~n19772;
  assign n19775 = ~n19773 & n19774;
  assign n19776 = pi0660 & ~n19715;
  assign n19777 = ~n19775 & n19776;
  assign n19778 = ~n19771 & ~n19777;
  assign n19779 = pi0785 & ~n19778;
  assign n19780 = ~pi0785 & ~n19766;
  assign n19781 = ~n19779 & ~n19780;
  assign n19782 = ~pi0618 & ~n19781;
  assign n19783 = ~pi1154 & ~n19750;
  assign n19784 = ~n19782 & n19783;
  assign n19785 = ~pi0627 & ~n19721;
  assign n19786 = ~n19784 & n19785;
  assign n19787 = ~pi0618 & n19696;
  assign n19788 = pi0618 & ~n19781;
  assign n19789 = pi1154 & ~n19787;
  assign n19790 = ~n19788 & n19789;
  assign n19791 = pi0627 & ~n19723;
  assign n19792 = ~n19790 & n19791;
  assign n19793 = ~n19786 & ~n19792;
  assign n19794 = pi0781 & ~n19793;
  assign n19795 = ~pi0781 & ~n19781;
  assign n19796 = ~n19794 & ~n19795;
  assign n19797 = ~pi0789 & n19796;
  assign n19798 = ~pi0619 & ~n19796;
  assign n19799 = pi0619 & n19697;
  assign n19800 = ~pi1159 & ~n19799;
  assign n19801 = ~n19798 & n19800;
  assign n19802 = ~pi0648 & ~n19731;
  assign n19803 = ~n19801 & n19802;
  assign n19804 = ~pi0619 & n19697;
  assign n19805 = pi0619 & ~n19796;
  assign n19806 = pi1159 & ~n19804;
  assign n19807 = ~n19805 & n19806;
  assign n19808 = pi0648 & ~n19735;
  assign n19809 = ~n19807 & n19808;
  assign n19810 = pi0789 & ~n19803;
  assign n19811 = ~n19809 & n19810;
  assign n19812 = n17970 & ~n19797;
  assign n19813 = ~n19811 & n19812;
  assign n19814 = ~n19749 & ~n19813;
  assign n19815 = ~pi0628 & ~n19814;
  assign n19816 = ~pi0788 & ~n19738;
  assign n19817 = pi0788 & ~n19746;
  assign n19818 = ~n19816 & ~n19817;
  assign n19819 = pi0628 & n19818;
  assign n19820 = ~pi1156 & ~n19819;
  assign n19821 = ~n19815 & n19820;
  assign n19822 = ~pi0629 & ~n19705;
  assign n19823 = ~n19821 & n19822;
  assign n19824 = ~n17997 & n19699;
  assign n19825 = ~pi1156 & ~n19824;
  assign n19826 = ~pi0628 & n19818;
  assign n19827 = pi0628 & ~n19814;
  assign n19828 = pi1156 & ~n19826;
  assign n19829 = ~n19827 & n19828;
  assign n19830 = pi0629 & ~n19825;
  assign n19831 = ~n19829 & n19830;
  assign n19832 = ~n19823 & ~n19831;
  assign n19833 = pi0792 & ~n19832;
  assign n19834 = ~pi0792 & ~n19814;
  assign n19835 = ~n19833 & ~n19834;
  assign n19836 = ~pi0647 & ~n19835;
  assign n19837 = ~n17779 & n19818;
  assign n19838 = n17779 & n19683;
  assign n19839 = ~n19837 & ~n19838;
  assign n19840 = pi0647 & ~n19839;
  assign n19841 = ~pi1157 & ~n19840;
  assign n19842 = ~n19836 & n19841;
  assign n19843 = ~pi0630 & ~n19703;
  assign n19844 = ~n19842 & n19843;
  assign n19845 = ~pi0647 & n19700;
  assign n19846 = pi0647 & n19683;
  assign n19847 = ~pi1157 & ~n19846;
  assign n19848 = ~n19845 & n19847;
  assign n19849 = pi0647 & ~n19835;
  assign n19850 = ~pi0647 & ~n19839;
  assign n19851 = pi1157 & ~n19850;
  assign n19852 = ~n19849 & n19851;
  assign n19853 = pi0630 & ~n19848;
  assign n19854 = ~n19852 & n19853;
  assign n19855 = ~n19844 & ~n19854;
  assign n19856 = pi0787 & ~n19855;
  assign n19857 = ~pi0787 & ~n19835;
  assign n19858 = ~n19856 & ~n19857;
  assign n19859 = ~pi0790 & ~n19858;
  assign n19860 = ~pi0787 & ~n19700;
  assign n19861 = ~n19703 & ~n19848;
  assign n19862 = pi0787 & ~n19861;
  assign n19863 = ~n19860 & ~n19862;
  assign n19864 = ~pi0644 & n19863;
  assign n19865 = pi0644 & ~n19858;
  assign n19866 = pi0715 & ~n19864;
  assign n19867 = ~n19865 & n19866;
  assign n19868 = n17804 & ~n19683;
  assign n19869 = ~n17804 & n19839;
  assign n19870 = ~n19868 & ~n19869;
  assign n19871 = pi0644 & n19870;
  assign n19872 = ~pi0644 & n19683;
  assign n19873 = ~pi0715 & ~n19872;
  assign n19874 = ~n19871 & n19873;
  assign n19875 = pi1160 & ~n19874;
  assign n19876 = ~n19867 & n19875;
  assign n19877 = ~pi0644 & n19870;
  assign n19878 = pi0644 & n19683;
  assign n19879 = pi0715 & ~n19878;
  assign n19880 = ~n19877 & n19879;
  assign n19881 = pi0644 & n19863;
  assign n19882 = ~pi0644 & ~n19858;
  assign n19883 = ~pi0715 & ~n19881;
  assign n19884 = ~n19882 & n19883;
  assign n19885 = ~pi1160 & ~n19880;
  assign n19886 = ~n19884 & n19885;
  assign n19887 = ~n19876 & ~n19886;
  assign n19888 = pi0790 & ~n19887;
  assign n19889 = pi0832 & ~n19859;
  assign n19890 = ~n19888 & n19889;
  assign po0300 = ~n19682 & ~n19890;
  assign n19892 = pi0144 & ~n17059;
  assign n19893 = n16635 & ~n19892;
  assign n19894 = n17075 & ~n19892;
  assign n19895 = pi0736 & n2571;
  assign n19896 = ~n19892 & ~n19895;
  assign n19897 = ~pi0144 & ~n16641;
  assign n19898 = n16641 & ~n16644;
  assign n19899 = pi0038 & ~n19898;
  assign n19900 = ~n19897 & n19899;
  assign n19901 = ~pi0144 & n18076;
  assign n19902 = pi0144 & ~n18072;
  assign n19903 = ~pi0038 & ~n19901;
  assign n19904 = ~n19902 & n19903;
  assign n19905 = n19895 & ~n19900;
  assign n19906 = ~n19904 & n19905;
  assign n19907 = ~n19896 & ~n19906;
  assign n19908 = ~pi0778 & n19907;
  assign n19909 = ~pi0625 & ~n19892;
  assign n19910 = pi0625 & ~n19907;
  assign n19911 = pi1153 & ~n19909;
  assign n19912 = ~n19910 & n19911;
  assign n19913 = ~pi0625 & ~n19907;
  assign n19914 = pi0625 & ~n19892;
  assign n19915 = ~pi1153 & ~n19914;
  assign n19916 = ~n19913 & n19915;
  assign n19917 = ~n19912 & ~n19916;
  assign n19918 = pi0778 & ~n19917;
  assign n19919 = ~n19908 & ~n19918;
  assign n19920 = ~n17075 & n19919;
  assign n19921 = ~n19894 & ~n19920;
  assign n19922 = ~n16639 & n19921;
  assign n19923 = n16639 & n19892;
  assign n19924 = ~n19922 & ~n19923;
  assign n19925 = ~n16635 & n19924;
  assign n19926 = ~n19893 & ~n19925;
  assign n19927 = ~n16631 & n19926;
  assign n19928 = n16631 & n19892;
  assign n19929 = ~n19927 & ~n19928;
  assign n19930 = ~pi0792 & ~n19929;
  assign n19931 = ~pi0628 & ~n19892;
  assign n19932 = pi0628 & n19929;
  assign n19933 = pi1156 & ~n19931;
  assign n19934 = ~n19932 & n19933;
  assign n19935 = pi0628 & ~n19892;
  assign n19936 = ~pi0628 & n19929;
  assign n19937 = ~pi1156 & ~n19935;
  assign n19938 = ~n19936 & n19937;
  assign n19939 = ~n19934 & ~n19938;
  assign n19940 = pi0792 & ~n19939;
  assign n19941 = ~n19930 & ~n19940;
  assign n19942 = ~pi0787 & ~n19941;
  assign n19943 = ~pi0647 & ~n19892;
  assign n19944 = pi0647 & n19941;
  assign n19945 = pi1157 & ~n19943;
  assign n19946 = ~n19944 & n19945;
  assign n19947 = pi0647 & ~n19892;
  assign n19948 = ~pi0647 & n19941;
  assign n19949 = ~pi1157 & ~n19947;
  assign n19950 = ~n19948 & n19949;
  assign n19951 = ~n19946 & ~n19950;
  assign n19952 = pi0787 & ~n19951;
  assign n19953 = ~n19942 & ~n19952;
  assign n19954 = ~pi0644 & n19953;
  assign n19955 = ~pi0619 & ~n19892;
  assign n19956 = n17117 & ~n19892;
  assign n19957 = pi0144 & ~n2571;
  assign n19958 = ~pi0758 & ~n17046;
  assign n19959 = pi0758 & n17219;
  assign n19960 = ~n19958 & ~n19959;
  assign n19961 = pi0039 & ~n19960;
  assign n19962 = ~pi0758 & n16958;
  assign n19963 = pi0758 & n17139;
  assign n19964 = ~pi0039 & ~n19962;
  assign n19965 = ~n19963 & n19964;
  assign n19966 = ~n19961 & ~n19965;
  assign n19967 = pi0144 & ~n19966;
  assign n19968 = ~pi0144 & pi0758;
  assign n19969 = n17275 & n19968;
  assign n19970 = ~n19967 & ~n19969;
  assign n19971 = ~pi0038 & ~n19970;
  assign n19972 = pi0758 & n17168;
  assign n19973 = n16641 & ~n19972;
  assign n19974 = pi0038 & ~n19897;
  assign n19975 = ~n19973 & n19974;
  assign n19976 = ~n19971 & ~n19975;
  assign n19977 = n2571 & ~n19976;
  assign n19978 = ~n19957 & ~n19977;
  assign n19979 = ~n17117 & n19978;
  assign n19980 = ~n19956 & ~n19979;
  assign n19981 = ~pi0785 & n19980;
  assign n19982 = ~pi0609 & ~n19892;
  assign n19983 = pi0609 & ~n19980;
  assign n19984 = pi1155 & ~n19982;
  assign n19985 = ~n19983 & n19984;
  assign n19986 = ~pi0609 & ~n19980;
  assign n19987 = pi0609 & ~n19892;
  assign n19988 = ~pi1155 & ~n19987;
  assign n19989 = ~n19986 & n19988;
  assign n19990 = ~n19985 & ~n19989;
  assign n19991 = pi0785 & ~n19990;
  assign n19992 = ~n19981 & ~n19991;
  assign n19993 = ~pi0781 & ~n19992;
  assign n19994 = ~pi0618 & ~n19892;
  assign n19995 = pi0618 & n19992;
  assign n19996 = pi1154 & ~n19994;
  assign n19997 = ~n19995 & n19996;
  assign n19998 = pi0618 & ~n19892;
  assign n19999 = ~pi0618 & n19992;
  assign n20000 = ~pi1154 & ~n19998;
  assign n20001 = ~n19999 & n20000;
  assign n20002 = ~n19997 & ~n20001;
  assign n20003 = pi0781 & ~n20002;
  assign n20004 = ~n19993 & ~n20003;
  assign n20005 = pi0619 & n20004;
  assign n20006 = pi1159 & ~n19955;
  assign n20007 = ~n20005 & n20006;
  assign n20008 = ~pi0736 & n19976;
  assign n20009 = ~pi0144 & ~n17605;
  assign n20010 = pi0144 & n17546;
  assign n20011 = pi0758 & ~n20010;
  assign n20012 = ~n20009 & n20011;
  assign n20013 = pi0144 & ~n17404;
  assign n20014 = ~pi0144 & ~n17485;
  assign n20015 = ~pi0758 & ~n20014;
  assign n20016 = ~n20013 & n20015;
  assign n20017 = pi0039 & ~n20012;
  assign n20018 = ~n20016 & n20017;
  assign n20019 = ~pi0144 & n17631;
  assign n20020 = pi0144 & n17629;
  assign n20021 = pi0758 & ~n20019;
  assign n20022 = ~n20020 & n20021;
  assign n20023 = ~pi0144 & ~n17625;
  assign n20024 = pi0144 & ~n17612;
  assign n20025 = ~pi0758 & ~n20023;
  assign n20026 = ~n20024 & n20025;
  assign n20027 = ~pi0039 & ~n20022;
  assign n20028 = ~n20026 & n20027;
  assign n20029 = ~pi0038 & ~n20028;
  assign n20030 = ~n20018 & n20029;
  assign n20031 = pi0736 & ~n19470;
  assign n20032 = ~n19975 & n20031;
  assign n20033 = ~n20030 & n20032;
  assign n20034 = n2571 & ~n20033;
  assign n20035 = ~n20008 & n20034;
  assign n20036 = ~n19957 & ~n20035;
  assign n20037 = ~pi0625 & n20036;
  assign n20038 = pi0625 & n19978;
  assign n20039 = ~pi1153 & ~n20038;
  assign n20040 = ~n20037 & n20039;
  assign n20041 = ~pi0608 & ~n19912;
  assign n20042 = ~n20040 & n20041;
  assign n20043 = ~pi0625 & n19978;
  assign n20044 = pi0625 & n20036;
  assign n20045 = pi1153 & ~n20043;
  assign n20046 = ~n20044 & n20045;
  assign n20047 = pi0608 & ~n19916;
  assign n20048 = ~n20046 & n20047;
  assign n20049 = ~n20042 & ~n20048;
  assign n20050 = pi0778 & ~n20049;
  assign n20051 = ~pi0778 & n20036;
  assign n20052 = ~n20050 & ~n20051;
  assign n20053 = ~pi0609 & ~n20052;
  assign n20054 = pi0609 & n19919;
  assign n20055 = ~pi1155 & ~n20054;
  assign n20056 = ~n20053 & n20055;
  assign n20057 = ~pi0660 & ~n19985;
  assign n20058 = ~n20056 & n20057;
  assign n20059 = ~pi0609 & n19919;
  assign n20060 = pi0609 & ~n20052;
  assign n20061 = pi1155 & ~n20059;
  assign n20062 = ~n20060 & n20061;
  assign n20063 = pi0660 & ~n19989;
  assign n20064 = ~n20062 & n20063;
  assign n20065 = ~n20058 & ~n20064;
  assign n20066 = pi0785 & ~n20065;
  assign n20067 = ~pi0785 & ~n20052;
  assign n20068 = ~n20066 & ~n20067;
  assign n20069 = ~pi0618 & ~n20068;
  assign n20070 = pi0618 & ~n19921;
  assign n20071 = ~pi1154 & ~n20070;
  assign n20072 = ~n20069 & n20071;
  assign n20073 = ~pi0627 & ~n19997;
  assign n20074 = ~n20072 & n20073;
  assign n20075 = pi0618 & ~n20068;
  assign n20076 = ~pi0618 & ~n19921;
  assign n20077 = pi1154 & ~n20076;
  assign n20078 = ~n20075 & n20077;
  assign n20079 = pi0627 & ~n20001;
  assign n20080 = ~n20078 & n20079;
  assign n20081 = ~n20074 & ~n20080;
  assign n20082 = pi0781 & ~n20081;
  assign n20083 = ~pi0781 & ~n20068;
  assign n20084 = ~n20082 & ~n20083;
  assign n20085 = ~pi0619 & ~n20084;
  assign n20086 = pi0619 & n19924;
  assign n20087 = ~pi1159 & ~n20086;
  assign n20088 = ~n20085 & n20087;
  assign n20089 = ~pi0648 & ~n20007;
  assign n20090 = ~n20088 & n20089;
  assign n20091 = pi0619 & ~n19892;
  assign n20092 = ~pi0619 & n20004;
  assign n20093 = ~pi1159 & ~n20091;
  assign n20094 = ~n20092 & n20093;
  assign n20095 = ~pi0619 & n19924;
  assign n20096 = pi0619 & ~n20084;
  assign n20097 = pi1159 & ~n20095;
  assign n20098 = ~n20096 & n20097;
  assign n20099 = pi0648 & ~n20094;
  assign n20100 = ~n20098 & n20099;
  assign n20101 = ~n20090 & ~n20100;
  assign n20102 = pi0789 & ~n20101;
  assign n20103 = ~pi0789 & ~n20084;
  assign n20104 = ~n20102 & ~n20103;
  assign n20105 = ~pi0788 & n20104;
  assign n20106 = ~pi0626 & n20104;
  assign n20107 = pi0626 & n19926;
  assign n20108 = ~pi0641 & ~n20107;
  assign n20109 = ~n20106 & n20108;
  assign n20110 = ~pi0789 & ~n20004;
  assign n20111 = ~n20007 & ~n20094;
  assign n20112 = pi0789 & ~n20111;
  assign n20113 = ~n20110 & ~n20112;
  assign n20114 = ~pi0626 & n20113;
  assign n20115 = pi0626 & ~n19892;
  assign n20116 = ~pi1158 & ~n20115;
  assign n20117 = ~n20114 & n20116;
  assign n20118 = ~n17730 & ~n20117;
  assign n20119 = ~n20109 & ~n20118;
  assign n20120 = pi0626 & n20104;
  assign n20121 = ~pi0626 & n19926;
  assign n20122 = pi0641 & ~n20121;
  assign n20123 = ~n20120 & n20122;
  assign n20124 = pi0626 & n20113;
  assign n20125 = ~pi0626 & ~n19892;
  assign n20126 = pi1158 & ~n20125;
  assign n20127 = ~n20124 & n20126;
  assign n20128 = ~n17745 & ~n20127;
  assign n20129 = ~n20123 & ~n20128;
  assign n20130 = ~n20119 & ~n20129;
  assign n20131 = pi0788 & ~n20130;
  assign n20132 = ~n20105 & ~n20131;
  assign n20133 = ~pi0628 & n20132;
  assign n20134 = ~n20117 & ~n20127;
  assign n20135 = pi0788 & ~n20134;
  assign n20136 = ~pi0788 & ~n20113;
  assign n20137 = ~n20135 & ~n20136;
  assign n20138 = pi0628 & n20137;
  assign n20139 = ~pi1156 & ~n20138;
  assign n20140 = ~n20133 & n20139;
  assign n20141 = ~pi0629 & ~n19934;
  assign n20142 = ~n20140 & n20141;
  assign n20143 = pi0628 & n20132;
  assign n20144 = ~pi0628 & n20137;
  assign n20145 = pi1156 & ~n20144;
  assign n20146 = ~n20143 & n20145;
  assign n20147 = pi0629 & ~n19938;
  assign n20148 = ~n20146 & n20147;
  assign n20149 = ~n20142 & ~n20148;
  assign n20150 = pi0792 & ~n20149;
  assign n20151 = ~pi0792 & n20132;
  assign n20152 = ~n20150 & ~n20151;
  assign n20153 = ~pi0647 & ~n20152;
  assign n20154 = ~n17779 & ~n20137;
  assign n20155 = n17779 & n19892;
  assign n20156 = ~n20154 & ~n20155;
  assign n20157 = pi0647 & n20156;
  assign n20158 = ~pi1157 & ~n20157;
  assign n20159 = ~n20153 & n20158;
  assign n20160 = ~pi0630 & ~n19946;
  assign n20161 = ~n20159 & n20160;
  assign n20162 = pi0647 & ~n20152;
  assign n20163 = ~pi0647 & n20156;
  assign n20164 = pi1157 & ~n20163;
  assign n20165 = ~n20162 & n20164;
  assign n20166 = pi0630 & ~n19950;
  assign n20167 = ~n20165 & n20166;
  assign n20168 = ~n20161 & ~n20167;
  assign n20169 = pi0787 & ~n20168;
  assign n20170 = ~pi0787 & ~n20152;
  assign n20171 = ~n20169 & ~n20170;
  assign n20172 = pi0644 & ~n20171;
  assign n20173 = pi0715 & ~n19954;
  assign n20174 = ~n20172 & n20173;
  assign n20175 = n17804 & ~n19892;
  assign n20176 = ~n17804 & n20156;
  assign n20177 = ~n20175 & ~n20176;
  assign n20178 = pi0644 & ~n20177;
  assign n20179 = ~pi0644 & ~n19892;
  assign n20180 = ~pi0715 & ~n20179;
  assign n20181 = ~n20178 & n20180;
  assign n20182 = pi1160 & ~n20181;
  assign n20183 = ~n20174 & n20182;
  assign n20184 = ~pi0644 & ~n20171;
  assign n20185 = pi0644 & n19953;
  assign n20186 = ~pi0715 & ~n20185;
  assign n20187 = ~n20184 & n20186;
  assign n20188 = ~pi0644 & ~n20177;
  assign n20189 = pi0644 & ~n19892;
  assign n20190 = pi0715 & ~n20189;
  assign n20191 = ~n20188 & n20190;
  assign n20192 = ~pi1160 & ~n20191;
  assign n20193 = ~n20187 & n20192;
  assign n20194 = pi0790 & ~n20183;
  assign n20195 = ~n20193 & n20194;
  assign n20196 = ~pi0790 & n20171;
  assign n20197 = n6305 & ~n20196;
  assign n20198 = ~n20195 & n20197;
  assign n20199 = ~pi0144 & ~n6305;
  assign n20200 = ~pi0057 & ~n20199;
  assign n20201 = ~n20198 & n20200;
  assign n20202 = pi0057 & pi0144;
  assign n20203 = ~pi0832 & ~n20202;
  assign n20204 = ~n20201 & n20203;
  assign n20205 = n17803 & n19341;
  assign n20206 = pi0787 & ~n20205;
  assign n20207 = pi0144 & ~n2926;
  assign n20208 = pi0736 & n16645;
  assign n20209 = ~n20207 & ~n20208;
  assign n20210 = ~pi0778 & n20209;
  assign n20211 = pi0625 & n20208;
  assign n20212 = ~n20209 & ~n20211;
  assign n20213 = ~pi1153 & ~n20212;
  assign n20214 = pi1153 & ~n20207;
  assign n20215 = ~n20211 & n20214;
  assign n20216 = ~n20213 & ~n20215;
  assign n20217 = pi0778 & ~n20216;
  assign n20218 = ~n20210 & ~n20217;
  assign n20219 = n19151 & n20218;
  assign n20220 = ~pi0628 & n20219;
  assign n20221 = pi0629 & ~n20220;
  assign n20222 = ~pi0609 & ~pi1155;
  assign n20223 = pi0609 & pi1155;
  assign n20224 = pi0785 & ~n20222;
  assign n20225 = ~n20223 & n20224;
  assign n20226 = pi0758 & n17244;
  assign n20227 = ~n20225 & n20226;
  assign n20228 = ~pi0619 & pi1159;
  assign n20229 = pi0619 & ~pi1159;
  assign n20230 = ~n20228 & ~n20229;
  assign n20231 = pi0789 & ~n20230;
  assign n20232 = ~pi0618 & ~pi1154;
  assign n20233 = pi0618 & pi1154;
  assign n20234 = pi0781 & ~n20232;
  assign n20235 = ~n20233 & n20234;
  assign n20236 = ~n17117 & ~n20231;
  assign n20237 = ~n20235 & n20236;
  assign n20238 = n20227 & n20237;
  assign n20239 = ~n17969 & n20238;
  assign n20240 = pi0628 & ~n20239;
  assign n20241 = ~n20221 & ~n20240;
  assign n20242 = ~pi1156 & ~n20241;
  assign n20243 = pi0628 & n20219;
  assign n20244 = ~pi0628 & ~n20239;
  assign n20245 = pi0629 & ~n20244;
  assign n20246 = pi1156 & ~n20245;
  assign n20247 = ~n20243 & n20246;
  assign n20248 = ~n20242 & ~n20247;
  assign n20249 = ~n20207 & ~n20248;
  assign n20250 = pi0792 & n20249;
  assign n20251 = n16635 & ~n20207;
  assign n20252 = ~n17075 & n20218;
  assign n20253 = ~n16639 & n20252;
  assign n20254 = ~n20207 & ~n20253;
  assign n20255 = ~n20251 & ~n20254;
  assign n20256 = n17865 & n20255;
  assign n20257 = ~pi0626 & n20238;
  assign n20258 = ~n20207 & ~n20257;
  assign n20259 = ~pi1158 & ~n20258;
  assign n20260 = pi0641 & ~n20259;
  assign n20261 = ~n20256 & n20260;
  assign n20262 = pi0626 & n20238;
  assign n20263 = ~n20207 & ~n20262;
  assign n20264 = pi1158 & ~n20263;
  assign n20265 = n17866 & n20255;
  assign n20266 = ~pi0641 & ~n20264;
  assign n20267 = ~n20265 & n20266;
  assign n20268 = pi0788 & ~n20261;
  assign n20269 = ~n20267 & n20268;
  assign n20270 = pi0618 & ~n17117;
  assign n20271 = n20227 & n20270;
  assign n20272 = pi1154 & ~n20207;
  assign n20273 = ~n20271 & n20272;
  assign n20274 = ~n20207 & ~n20252;
  assign n20275 = pi0618 & ~n20274;
  assign n20276 = n17291 & n20226;
  assign n20277 = pi1155 & ~n20207;
  assign n20278 = ~n20276 & n20277;
  assign n20279 = pi0609 & n20218;
  assign n20280 = ~n20207 & ~n20226;
  assign n20281 = pi0736 & n17469;
  assign n20282 = n20280 & ~n20281;
  assign n20283 = pi0625 & n20281;
  assign n20284 = ~n20282 & ~n20283;
  assign n20285 = ~pi1153 & ~n20284;
  assign n20286 = ~pi0608 & ~n20215;
  assign n20287 = ~n20285 & n20286;
  assign n20288 = pi1153 & n20280;
  assign n20289 = ~n20283 & n20288;
  assign n20290 = pi0608 & ~n20213;
  assign n20291 = ~n20289 & n20290;
  assign n20292 = ~n20287 & ~n20291;
  assign n20293 = pi0778 & ~n20292;
  assign n20294 = ~pi0778 & ~n20282;
  assign n20295 = ~n20293 & ~n20294;
  assign n20296 = ~pi0609 & ~n20295;
  assign n20297 = ~pi1155 & ~n20279;
  assign n20298 = ~n20296 & n20297;
  assign n20299 = ~pi0660 & ~n20278;
  assign n20300 = ~n20298 & n20299;
  assign n20301 = n17296 & n20226;
  assign n20302 = ~pi1155 & ~n20207;
  assign n20303 = ~n20301 & n20302;
  assign n20304 = ~pi0609 & n20218;
  assign n20305 = pi0609 & ~n20295;
  assign n20306 = pi1155 & ~n20304;
  assign n20307 = ~n20305 & n20306;
  assign n20308 = pi0660 & ~n20303;
  assign n20309 = ~n20307 & n20308;
  assign n20310 = ~n20300 & ~n20309;
  assign n20311 = pi0785 & ~n20310;
  assign n20312 = ~pi0785 & ~n20295;
  assign n20313 = ~n20311 & ~n20312;
  assign n20314 = ~pi0618 & ~n20313;
  assign n20315 = ~pi1154 & ~n20275;
  assign n20316 = ~n20314 & n20315;
  assign n20317 = ~pi0627 & ~n20273;
  assign n20318 = ~n20316 & n20317;
  assign n20319 = ~pi0618 & ~n17117;
  assign n20320 = n20227 & n20319;
  assign n20321 = ~pi1154 & ~n20207;
  assign n20322 = ~n20320 & n20321;
  assign n20323 = ~pi0618 & ~n20274;
  assign n20324 = pi0618 & ~n20313;
  assign n20325 = pi1154 & ~n20323;
  assign n20326 = ~n20324 & n20325;
  assign n20327 = pi0627 & ~n20322;
  assign n20328 = ~n20326 & n20327;
  assign n20329 = ~n20318 & ~n20328;
  assign n20330 = pi0781 & ~n20329;
  assign n20331 = ~pi0781 & ~n20313;
  assign n20332 = ~n20330 & ~n20331;
  assign n20333 = ~pi0789 & n20332;
  assign n20334 = n20227 & ~n20235;
  assign n20335 = pi0619 & ~n17117;
  assign n20336 = n20334 & n20335;
  assign n20337 = pi1159 & ~n20207;
  assign n20338 = ~n20336 & n20337;
  assign n20339 = pi0619 & ~n20254;
  assign n20340 = ~pi0619 & ~n20332;
  assign n20341 = ~pi1159 & ~n20339;
  assign n20342 = ~n20340 & n20341;
  assign n20343 = ~pi0648 & ~n20338;
  assign n20344 = ~n20342 & n20343;
  assign n20345 = ~pi0619 & ~n17117;
  assign n20346 = n20334 & n20345;
  assign n20347 = ~pi1159 & ~n20207;
  assign n20348 = ~n20346 & n20347;
  assign n20349 = ~pi0619 & ~n20254;
  assign n20350 = pi0619 & ~n20332;
  assign n20351 = pi1159 & ~n20349;
  assign n20352 = ~n20350 & n20351;
  assign n20353 = pi0648 & ~n20348;
  assign n20354 = ~n20352 & n20353;
  assign n20355 = pi0789 & ~n20344;
  assign n20356 = ~n20354 & n20355;
  assign n20357 = n17970 & ~n20333;
  assign n20358 = ~n20356 & n20357;
  assign n20359 = ~n20269 & ~n20358;
  assign n20360 = ~n20250 & ~n20359;
  assign n20361 = pi0629 & n19139;
  assign n20362 = ~pi0629 & n19140;
  assign n20363 = pi0792 & ~n20361;
  assign n20364 = ~n20362 & n20363;
  assign n20365 = ~n20249 & n20364;
  assign n20366 = ~n20206 & ~n20365;
  assign n20367 = ~n20360 & n20366;
  assign n20368 = ~n17779 & n20239;
  assign n20369 = ~pi0630 & n20368;
  assign n20370 = pi0647 & ~n20369;
  assign n20371 = ~n19142 & n20219;
  assign n20372 = pi0630 & ~n20371;
  assign n20373 = ~n20370 & ~n20372;
  assign n20374 = ~pi1157 & ~n20373;
  assign n20375 = pi0630 & n20368;
  assign n20376 = ~pi0630 & ~n20371;
  assign n20377 = pi0647 & ~n20376;
  assign n20378 = pi1157 & ~n20375;
  assign n20379 = ~n20377 & n20378;
  assign n20380 = ~n20374 & ~n20379;
  assign n20381 = pi0787 & ~n20207;
  assign n20382 = ~n20380 & n20381;
  assign n20383 = ~n20367 & ~n20382;
  assign n20384 = ~pi0790 & n20383;
  assign n20385 = ~n17804 & n20368;
  assign n20386 = pi0644 & n20385;
  assign n20387 = ~pi0715 & ~n20207;
  assign n20388 = ~n20386 & n20387;
  assign n20389 = ~n19342 & n20371;
  assign n20390 = ~n20207 & ~n20389;
  assign n20391 = ~pi0644 & ~n20390;
  assign n20392 = pi0644 & n20383;
  assign n20393 = pi0715 & ~n20391;
  assign n20394 = ~n20392 & n20393;
  assign n20395 = pi1160 & ~n20388;
  assign n20396 = ~n20394 & n20395;
  assign n20397 = ~pi0644 & n20385;
  assign n20398 = pi0715 & ~n20207;
  assign n20399 = ~n20397 & n20398;
  assign n20400 = ~pi0644 & n20383;
  assign n20401 = pi0644 & ~n20390;
  assign n20402 = ~pi0715 & ~n20401;
  assign n20403 = ~n20400 & n20402;
  assign n20404 = ~pi1160 & ~n20399;
  assign n20405 = ~n20403 & n20404;
  assign n20406 = ~n20396 & ~n20405;
  assign n20407 = pi0790 & ~n20406;
  assign n20408 = pi0832 & ~n20384;
  assign n20409 = ~n20407 & n20408;
  assign po0301 = ~n20204 & ~n20409;
  assign n20411 = ~pi0145 & po1038;
  assign n20412 = ~pi0145 & ~n17059;
  assign n20413 = n16635 & ~n20412;
  assign n20414 = ~pi0698 & n2571;
  assign n20415 = n20412 & ~n20414;
  assign n20416 = ~pi0145 & ~n16641;
  assign n20417 = n16647 & ~n20416;
  assign n20418 = pi0145 & ~n18076;
  assign n20419 = ~pi0038 & ~n20418;
  assign n20420 = n2571 & ~n20419;
  assign n20421 = ~pi0145 & n18072;
  assign n20422 = ~n20420 & ~n20421;
  assign n20423 = ~pi0698 & ~n20417;
  assign n20424 = ~n20422 & n20423;
  assign n20425 = ~n20415 & ~n20424;
  assign n20426 = ~pi0778 & n20425;
  assign n20427 = ~pi0625 & n20412;
  assign n20428 = pi0625 & ~n20425;
  assign n20429 = pi1153 & ~n20427;
  assign n20430 = ~n20428 & n20429;
  assign n20431 = pi0625 & n20412;
  assign n20432 = ~pi0625 & ~n20425;
  assign n20433 = ~pi1153 & ~n20431;
  assign n20434 = ~n20432 & n20433;
  assign n20435 = ~n20430 & ~n20434;
  assign n20436 = pi0778 & ~n20435;
  assign n20437 = ~n20426 & ~n20436;
  assign n20438 = ~n17075 & ~n20437;
  assign n20439 = n17075 & ~n20412;
  assign n20440 = ~n20438 & ~n20439;
  assign n20441 = ~n16639 & n20440;
  assign n20442 = n16639 & n20412;
  assign n20443 = ~n20441 & ~n20442;
  assign n20444 = ~n16635 & n20443;
  assign n20445 = ~n20413 & ~n20444;
  assign n20446 = ~n16631 & n20445;
  assign n20447 = n16631 & n20412;
  assign n20448 = ~n20446 & ~n20447;
  assign n20449 = ~pi0792 & n20448;
  assign n20450 = pi0628 & ~n20448;
  assign n20451 = ~pi0628 & n20412;
  assign n20452 = pi1156 & ~n20451;
  assign n20453 = ~n20450 & n20452;
  assign n20454 = pi0628 & n20412;
  assign n20455 = ~pi0628 & ~n20448;
  assign n20456 = ~pi1156 & ~n20454;
  assign n20457 = ~n20455 & n20456;
  assign n20458 = ~n20453 & ~n20457;
  assign n20459 = pi0792 & ~n20458;
  assign n20460 = ~n20449 & ~n20459;
  assign n20461 = ~pi0647 & ~n20460;
  assign n20462 = pi0647 & ~n20412;
  assign n20463 = ~n20461 & ~n20462;
  assign n20464 = ~pi1157 & n20463;
  assign n20465 = pi0647 & ~n20460;
  assign n20466 = ~pi0647 & ~n20412;
  assign n20467 = ~n20465 & ~n20466;
  assign n20468 = pi1157 & n20467;
  assign n20469 = ~n20464 & ~n20468;
  assign n20470 = pi0787 & ~n20469;
  assign n20471 = ~pi0787 & n20460;
  assign n20472 = ~n20470 & ~n20471;
  assign n20473 = ~pi0644 & ~n20472;
  assign n20474 = pi0715 & ~n20473;
  assign n20475 = pi0145 & ~n2571;
  assign n20476 = pi0145 & ~n17275;
  assign n20477 = ~pi0145 & ~n17048;
  assign n20478 = pi0767 & ~n20477;
  assign n20479 = ~pi0145 & ~pi0767;
  assign n20480 = n17221 & n20479;
  assign n20481 = ~n20476 & ~n20480;
  assign n20482 = ~n20478 & n20481;
  assign n20483 = ~pi0038 & ~n20482;
  assign n20484 = ~pi0767 & n17280;
  assign n20485 = pi0038 & ~n20416;
  assign n20486 = ~n20484 & n20485;
  assign n20487 = ~n20483 & ~n20486;
  assign n20488 = n2571 & ~n20487;
  assign n20489 = ~n20475 & ~n20488;
  assign n20490 = ~n17117 & ~n20489;
  assign n20491 = n17117 & ~n20412;
  assign n20492 = ~n20490 & ~n20491;
  assign n20493 = ~pi0785 & ~n20492;
  assign n20494 = ~n17291 & ~n20412;
  assign n20495 = pi0609 & n20490;
  assign n20496 = ~n20494 & ~n20495;
  assign n20497 = pi1155 & ~n20496;
  assign n20498 = ~n17296 & ~n20412;
  assign n20499 = ~pi0609 & n20490;
  assign n20500 = ~n20498 & ~n20499;
  assign n20501 = ~pi1155 & ~n20500;
  assign n20502 = ~n20497 & ~n20501;
  assign n20503 = pi0785 & ~n20502;
  assign n20504 = ~n20493 & ~n20503;
  assign n20505 = ~pi0781 & ~n20504;
  assign n20506 = ~pi0618 & n20412;
  assign n20507 = pi0618 & n20504;
  assign n20508 = pi1154 & ~n20506;
  assign n20509 = ~n20507 & n20508;
  assign n20510 = ~pi0618 & n20504;
  assign n20511 = pi0618 & n20412;
  assign n20512 = ~pi1154 & ~n20511;
  assign n20513 = ~n20510 & n20512;
  assign n20514 = ~n20509 & ~n20513;
  assign n20515 = pi0781 & ~n20514;
  assign n20516 = ~n20505 & ~n20515;
  assign n20517 = ~pi0789 & ~n20516;
  assign n20518 = ~pi0619 & n20412;
  assign n20519 = pi0619 & n20516;
  assign n20520 = pi1159 & ~n20518;
  assign n20521 = ~n20519 & n20520;
  assign n20522 = ~pi0619 & n20516;
  assign n20523 = pi0619 & n20412;
  assign n20524 = ~pi1159 & ~n20523;
  assign n20525 = ~n20522 & n20524;
  assign n20526 = ~n20521 & ~n20525;
  assign n20527 = pi0789 & ~n20526;
  assign n20528 = ~n20517 & ~n20527;
  assign n20529 = ~pi0788 & ~n20528;
  assign n20530 = ~pi0626 & n20412;
  assign n20531 = pi0626 & n20528;
  assign n20532 = pi1158 & ~n20530;
  assign n20533 = ~n20531 & n20532;
  assign n20534 = ~pi0626 & n20528;
  assign n20535 = pi0626 & n20412;
  assign n20536 = ~pi1158 & ~n20535;
  assign n20537 = ~n20534 & n20536;
  assign n20538 = ~n20533 & ~n20537;
  assign n20539 = pi0788 & ~n20538;
  assign n20540 = ~n20529 & ~n20539;
  assign n20541 = ~n17779 & n20540;
  assign n20542 = n17779 & n20412;
  assign n20543 = ~n20541 & ~n20542;
  assign n20544 = ~n17804 & ~n20543;
  assign n20545 = n17804 & n20412;
  assign n20546 = ~n20544 & ~n20545;
  assign n20547 = pi0644 & ~n20546;
  assign n20548 = ~pi0644 & n20412;
  assign n20549 = ~pi0715 & ~n20548;
  assign n20550 = ~n20547 & n20549;
  assign n20551 = pi1160 & ~n20550;
  assign n20552 = ~n20474 & n20551;
  assign n20553 = pi0644 & ~n20472;
  assign n20554 = n17802 & ~n20463;
  assign n20555 = pi0630 & ~pi0647;
  assign n20556 = pi1157 & n20555;
  assign n20557 = ~pi0630 & pi0647;
  assign n20558 = ~pi1157 & n20557;
  assign n20559 = ~n20556 & ~n20558;
  assign n20560 = n20543 & ~n20559;
  assign n20561 = n17801 & ~n20467;
  assign n20562 = ~n20554 & ~n20561;
  assign n20563 = ~n20560 & n20562;
  assign n20564 = pi0787 & ~n20563;
  assign n20565 = ~pi0629 & n20453;
  assign n20566 = ~pi0628 & pi0629;
  assign n20567 = pi1156 & n20566;
  assign n20568 = pi0628 & ~pi0629;
  assign n20569 = ~pi1156 & n20568;
  assign n20570 = ~n20567 & ~n20569;
  assign n20571 = ~n20540 & ~n20570;
  assign n20572 = pi0629 & n20457;
  assign n20573 = ~n20565 & ~n20572;
  assign n20574 = ~n20571 & n20573;
  assign n20575 = pi0792 & ~n20574;
  assign n20576 = pi0609 & n20437;
  assign n20577 = pi0145 & ~n17625;
  assign n20578 = ~pi0145 & ~n17612;
  assign n20579 = pi0767 & ~n20577;
  assign n20580 = ~n20578 & n20579;
  assign n20581 = ~pi0145 & n17629;
  assign n20582 = pi0145 & n17631;
  assign n20583 = ~pi0767 & ~n20582;
  assign n20584 = ~n20581 & n20583;
  assign n20585 = ~n20580 & ~n20584;
  assign n20586 = ~pi0039 & ~n20585;
  assign n20587 = pi0145 & n17605;
  assign n20588 = ~pi0145 & ~n17546;
  assign n20589 = ~pi0767 & ~n20588;
  assign n20590 = ~n20587 & n20589;
  assign n20591 = ~pi0145 & n17404;
  assign n20592 = pi0145 & n17485;
  assign n20593 = pi0767 & ~n20592;
  assign n20594 = ~n20591 & n20593;
  assign n20595 = pi0039 & ~n20590;
  assign n20596 = ~n20594 & n20595;
  assign n20597 = ~pi0038 & ~n20586;
  assign n20598 = ~n20596 & n20597;
  assign n20599 = ~pi0767 & ~n17490;
  assign n20600 = n19471 & ~n20599;
  assign n20601 = ~pi0145 & ~n20600;
  assign n20602 = ~pi0767 & n17244;
  assign n20603 = ~n17469 & ~n20602;
  assign n20604 = pi0145 & ~n20603;
  assign n20605 = n6284 & n20604;
  assign n20606 = pi0038 & ~n20605;
  assign n20607 = ~n20601 & n20606;
  assign n20608 = ~pi0698 & ~n20607;
  assign n20609 = ~n20598 & n20608;
  assign n20610 = pi0698 & n20487;
  assign n20611 = n2571 & ~n20609;
  assign n20612 = ~n20610 & n20611;
  assign n20613 = ~n20475 & ~n20612;
  assign n20614 = ~pi0625 & n20613;
  assign n20615 = pi0625 & n20489;
  assign n20616 = ~pi1153 & ~n20615;
  assign n20617 = ~n20614 & n20616;
  assign n20618 = ~pi0608 & ~n20430;
  assign n20619 = ~n20617 & n20618;
  assign n20620 = ~pi0625 & n20489;
  assign n20621 = pi0625 & n20613;
  assign n20622 = pi1153 & ~n20620;
  assign n20623 = ~n20621 & n20622;
  assign n20624 = pi0608 & ~n20434;
  assign n20625 = ~n20623 & n20624;
  assign n20626 = ~n20619 & ~n20625;
  assign n20627 = pi0778 & ~n20626;
  assign n20628 = ~pi0778 & n20613;
  assign n20629 = ~n20627 & ~n20628;
  assign n20630 = ~pi0609 & ~n20629;
  assign n20631 = ~pi1155 & ~n20576;
  assign n20632 = ~n20630 & n20631;
  assign n20633 = ~pi0660 & ~n20497;
  assign n20634 = ~n20632 & n20633;
  assign n20635 = ~pi0609 & n20437;
  assign n20636 = pi0609 & ~n20629;
  assign n20637 = pi1155 & ~n20635;
  assign n20638 = ~n20636 & n20637;
  assign n20639 = pi0660 & ~n20501;
  assign n20640 = ~n20638 & n20639;
  assign n20641 = ~n20634 & ~n20640;
  assign n20642 = pi0785 & ~n20641;
  assign n20643 = ~pi0785 & ~n20629;
  assign n20644 = ~n20642 & ~n20643;
  assign n20645 = ~pi0618 & ~n20644;
  assign n20646 = pi0618 & n20440;
  assign n20647 = ~pi1154 & ~n20646;
  assign n20648 = ~n20645 & n20647;
  assign n20649 = ~pi0627 & ~n20509;
  assign n20650 = ~n20648 & n20649;
  assign n20651 = ~pi0618 & n20440;
  assign n20652 = pi0618 & ~n20644;
  assign n20653 = pi1154 & ~n20651;
  assign n20654 = ~n20652 & n20653;
  assign n20655 = pi0627 & ~n20513;
  assign n20656 = ~n20654 & n20655;
  assign n20657 = ~n20650 & ~n20656;
  assign n20658 = pi0781 & ~n20657;
  assign n20659 = ~pi0781 & ~n20644;
  assign n20660 = ~n20658 & ~n20659;
  assign n20661 = ~pi0789 & n20660;
  assign n20662 = pi0619 & ~n20443;
  assign n20663 = ~pi0619 & ~n20660;
  assign n20664 = ~pi1159 & ~n20662;
  assign n20665 = ~n20663 & n20664;
  assign n20666 = ~pi0648 & ~n20521;
  assign n20667 = ~n20665 & n20666;
  assign n20668 = pi0619 & ~n20660;
  assign n20669 = ~pi0619 & ~n20443;
  assign n20670 = pi1159 & ~n20669;
  assign n20671 = ~n20668 & n20670;
  assign n20672 = pi0648 & ~n20525;
  assign n20673 = ~n20671 & n20672;
  assign n20674 = pi0789 & ~n20667;
  assign n20675 = ~n20673 & n20674;
  assign n20676 = n17970 & ~n20661;
  assign n20677 = ~n20675 & n20676;
  assign n20678 = n17871 & n20445;
  assign n20679 = ~n16630 & n20538;
  assign n20680 = ~n20678 & ~n20679;
  assign n20681 = pi0788 & ~n20680;
  assign n20682 = ~n20364 & ~n20681;
  assign n20683 = ~n20677 & n20682;
  assign n20684 = ~n20575 & ~n20683;
  assign n20685 = ~n20206 & ~n20684;
  assign n20686 = ~n20564 & ~n20685;
  assign n20687 = ~pi0644 & n20686;
  assign n20688 = ~pi0715 & ~n20553;
  assign n20689 = ~n20687 & n20688;
  assign n20690 = pi0644 & n20412;
  assign n20691 = ~pi0644 & ~n20546;
  assign n20692 = pi0715 & ~n20690;
  assign n20693 = ~n20691 & n20692;
  assign n20694 = ~pi1160 & ~n20693;
  assign n20695 = ~n20689 & n20694;
  assign n20696 = ~n20552 & ~n20695;
  assign n20697 = pi0790 & ~n20696;
  assign n20698 = pi0644 & n20551;
  assign n20699 = pi0790 & ~n20698;
  assign n20700 = n20686 & ~n20699;
  assign n20701 = ~n20697 & ~n20700;
  assign n20702 = ~po1038 & ~n20701;
  assign n20703 = ~pi0832 & ~n20411;
  assign n20704 = ~n20702 & n20703;
  assign n20705 = ~pi0145 & ~n2926;
  assign n20706 = ~pi0698 & n16645;
  assign n20707 = ~n20705 & ~n20706;
  assign n20708 = ~pi0778 & n20707;
  assign n20709 = ~pi0625 & n20706;
  assign n20710 = ~n20707 & ~n20709;
  assign n20711 = pi1153 & ~n20710;
  assign n20712 = ~pi1153 & ~n20705;
  assign n20713 = ~n20709 & n20712;
  assign n20714 = ~n20711 & ~n20713;
  assign n20715 = pi0778 & ~n20714;
  assign n20716 = ~n20708 & ~n20715;
  assign n20717 = ~n17845 & n20716;
  assign n20718 = ~n17847 & n20717;
  assign n20719 = ~n17849 & n20718;
  assign n20720 = ~n17851 & n20719;
  assign n20721 = ~n17857 & n20720;
  assign n20722 = ~pi0647 & n20721;
  assign n20723 = pi0647 & n20705;
  assign n20724 = ~pi1157 & ~n20723;
  assign n20725 = ~n20722 & n20724;
  assign n20726 = pi0630 & n20725;
  assign n20727 = ~n20602 & ~n20705;
  assign n20728 = ~n17874 & ~n20727;
  assign n20729 = ~pi0785 & ~n20728;
  assign n20730 = ~n17879 & ~n20727;
  assign n20731 = pi1155 & ~n20730;
  assign n20732 = ~n17882 & n20728;
  assign n20733 = ~pi1155 & ~n20732;
  assign n20734 = ~n20731 & ~n20733;
  assign n20735 = pi0785 & ~n20734;
  assign n20736 = ~n20729 & ~n20735;
  assign n20737 = ~pi0781 & ~n20736;
  assign n20738 = ~n17889 & n20736;
  assign n20739 = pi1154 & ~n20738;
  assign n20740 = ~n17892 & n20736;
  assign n20741 = ~pi1154 & ~n20740;
  assign n20742 = ~n20739 & ~n20741;
  assign n20743 = pi0781 & ~n20742;
  assign n20744 = ~n20737 & ~n20743;
  assign n20745 = ~pi0789 & ~n20744;
  assign n20746 = ~pi0619 & n20705;
  assign n20747 = pi0619 & n20744;
  assign n20748 = pi1159 & ~n20746;
  assign n20749 = ~n20747 & n20748;
  assign n20750 = ~pi0619 & n20744;
  assign n20751 = pi0619 & n20705;
  assign n20752 = ~pi1159 & ~n20751;
  assign n20753 = ~n20750 & n20752;
  assign n20754 = ~n20749 & ~n20753;
  assign n20755 = pi0789 & ~n20754;
  assign n20756 = ~n20745 & ~n20755;
  assign n20757 = ~pi0788 & ~n20756;
  assign n20758 = ~pi0626 & n20705;
  assign n20759 = pi0626 & n20756;
  assign n20760 = pi1158 & ~n20758;
  assign n20761 = ~n20759 & n20760;
  assign n20762 = ~pi0626 & n20756;
  assign n20763 = pi0626 & n20705;
  assign n20764 = ~pi1158 & ~n20763;
  assign n20765 = ~n20762 & n20764;
  assign n20766 = ~n20761 & ~n20765;
  assign n20767 = pi0788 & ~n20766;
  assign n20768 = ~n20757 & ~n20767;
  assign n20769 = ~n17779 & n20768;
  assign n20770 = n17779 & n20705;
  assign n20771 = ~n20769 & ~n20770;
  assign n20772 = ~n20559 & n20771;
  assign n20773 = pi0647 & ~n20721;
  assign n20774 = ~pi0647 & ~n20705;
  assign n20775 = ~n20773 & ~n20774;
  assign n20776 = n17801 & ~n20775;
  assign n20777 = ~n20726 & ~n20776;
  assign n20778 = ~n20772 & n20777;
  assign n20779 = pi0787 & ~n20778;
  assign n20780 = n17871 & n20719;
  assign n20781 = ~n16630 & n20766;
  assign n20782 = ~n20780 & ~n20781;
  assign n20783 = pi0788 & ~n20782;
  assign n20784 = pi0618 & n20717;
  assign n20785 = pi0609 & n20716;
  assign n20786 = ~n17168 & ~n20707;
  assign n20787 = pi0625 & n20786;
  assign n20788 = n20727 & ~n20786;
  assign n20789 = ~n20787 & ~n20788;
  assign n20790 = n20712 & ~n20789;
  assign n20791 = ~pi0608 & ~n20711;
  assign n20792 = ~n20790 & n20791;
  assign n20793 = pi1153 & n20727;
  assign n20794 = ~n20787 & n20793;
  assign n20795 = pi0608 & ~n20713;
  assign n20796 = ~n20794 & n20795;
  assign n20797 = ~n20792 & ~n20796;
  assign n20798 = pi0778 & ~n20797;
  assign n20799 = ~pi0778 & ~n20788;
  assign n20800 = ~n20798 & ~n20799;
  assign n20801 = ~pi0609 & ~n20800;
  assign n20802 = ~pi1155 & ~n20785;
  assign n20803 = ~n20801 & n20802;
  assign n20804 = ~pi0660 & ~n20731;
  assign n20805 = ~n20803 & n20804;
  assign n20806 = ~pi0609 & n20716;
  assign n20807 = pi0609 & ~n20800;
  assign n20808 = pi1155 & ~n20806;
  assign n20809 = ~n20807 & n20808;
  assign n20810 = pi0660 & ~n20733;
  assign n20811 = ~n20809 & n20810;
  assign n20812 = ~n20805 & ~n20811;
  assign n20813 = pi0785 & ~n20812;
  assign n20814 = ~pi0785 & ~n20800;
  assign n20815 = ~n20813 & ~n20814;
  assign n20816 = ~pi0618 & ~n20815;
  assign n20817 = ~pi1154 & ~n20784;
  assign n20818 = ~n20816 & n20817;
  assign n20819 = ~pi0627 & ~n20739;
  assign n20820 = ~n20818 & n20819;
  assign n20821 = ~pi0618 & n20717;
  assign n20822 = pi0618 & ~n20815;
  assign n20823 = pi1154 & ~n20821;
  assign n20824 = ~n20822 & n20823;
  assign n20825 = pi0627 & ~n20741;
  assign n20826 = ~n20824 & n20825;
  assign n20827 = ~n20820 & ~n20826;
  assign n20828 = pi0781 & ~n20827;
  assign n20829 = ~pi0781 & ~n20815;
  assign n20830 = ~n20828 & ~n20829;
  assign n20831 = ~pi0789 & n20830;
  assign n20832 = ~pi0619 & ~n20830;
  assign n20833 = pi0619 & n20718;
  assign n20834 = ~pi1159 & ~n20833;
  assign n20835 = ~n20832 & n20834;
  assign n20836 = ~pi0648 & ~n20749;
  assign n20837 = ~n20835 & n20836;
  assign n20838 = ~pi0619 & n20718;
  assign n20839 = pi0619 & ~n20830;
  assign n20840 = pi1159 & ~n20838;
  assign n20841 = ~n20839 & n20840;
  assign n20842 = pi0648 & ~n20753;
  assign n20843 = ~n20841 & n20842;
  assign n20844 = pi0789 & ~n20837;
  assign n20845 = ~n20843 & n20844;
  assign n20846 = n17970 & ~n20831;
  assign n20847 = ~n20845 & n20846;
  assign n20848 = ~n20783 & ~n20847;
  assign n20849 = ~n20364 & ~n20848;
  assign n20850 = n17854 & n20768;
  assign n20851 = pi1156 & ~n17862;
  assign n20852 = n20720 & n20851;
  assign n20853 = ~n20850 & ~n20852;
  assign n20854 = ~pi0629 & ~n20853;
  assign n20855 = ~pi1156 & ~n17997;
  assign n20856 = n20720 & n20855;
  assign n20857 = n17853 & n20768;
  assign n20858 = ~n20856 & ~n20857;
  assign n20859 = pi0629 & ~n20858;
  assign n20860 = ~n20854 & ~n20859;
  assign n20861 = pi0792 & ~n20860;
  assign n20862 = ~n20206 & ~n20861;
  assign n20863 = ~n20849 & n20862;
  assign n20864 = ~n20779 & ~n20863;
  assign n20865 = ~pi0790 & n20864;
  assign n20866 = ~pi0787 & ~n20721;
  assign n20867 = pi1157 & ~n20775;
  assign n20868 = ~n20725 & ~n20867;
  assign n20869 = pi0787 & ~n20868;
  assign n20870 = ~n20866 & ~n20869;
  assign n20871 = ~pi0644 & n20870;
  assign n20872 = pi0644 & n20864;
  assign n20873 = pi0715 & ~n20871;
  assign n20874 = ~n20872 & n20873;
  assign n20875 = ~n17804 & ~n20771;
  assign n20876 = n17804 & n20705;
  assign n20877 = ~n20875 & ~n20876;
  assign n20878 = pi0644 & ~n20877;
  assign n20879 = ~pi0644 & n20705;
  assign n20880 = ~pi0715 & ~n20879;
  assign n20881 = ~n20878 & n20880;
  assign n20882 = pi1160 & ~n20881;
  assign n20883 = ~n20874 & n20882;
  assign n20884 = ~pi0644 & ~n20877;
  assign n20885 = pi0644 & n20705;
  assign n20886 = pi0715 & ~n20885;
  assign n20887 = ~n20884 & n20886;
  assign n20888 = pi0644 & n20870;
  assign n20889 = ~pi0644 & n20864;
  assign n20890 = ~pi0715 & ~n20888;
  assign n20891 = ~n20889 & n20890;
  assign n20892 = ~pi1160 & ~n20887;
  assign n20893 = ~n20891 & n20892;
  assign n20894 = ~n20883 & ~n20893;
  assign n20895 = pi0790 & ~n20894;
  assign n20896 = pi0832 & ~n20865;
  assign n20897 = ~n20895 & n20896;
  assign po0302 = ~n20704 & ~n20897;
  assign n20899 = ~pi0146 & ~n10197;
  assign n20900 = ~pi0146 & ~n16641;
  assign n20901 = pi0743 & pi0947;
  assign n20902 = pi0907 & ~pi0947;
  assign n20903 = pi0735 & n20902;
  assign n20904 = ~n20901 & ~n20903;
  assign n20905 = n2926 & n20904;
  assign n20906 = n6284 & n20905;
  assign n20907 = pi0038 & ~n20906;
  assign n20908 = ~n20900 & n20907;
  assign n20909 = ~pi0146 & ~n16941;
  assign n20910 = n16941 & n20904;
  assign n20911 = pi0299 & ~n20909;
  assign n20912 = ~n20910 & n20911;
  assign n20913 = ~pi0146 & ~n16930;
  assign n20914 = n16930 & n20904;
  assign n20915 = ~pi0299 & ~n20913;
  assign n20916 = ~n20914 & n20915;
  assign n20917 = ~pi0039 & ~n20912;
  assign n20918 = ~n20916 & n20917;
  assign n20919 = n16653 & ~n20904;
  assign n20920 = pi0146 & ~n16653;
  assign n20921 = ~n20919 & ~n20920;
  assign n20922 = n3448 & ~n20921;
  assign n20923 = ~pi0907 & n6241;
  assign n20924 = pi0146 & ~n17018;
  assign n20925 = ~n20923 & n20924;
  assign n20926 = pi0735 & pi0907;
  assign n20927 = n17018 & n20926;
  assign n20928 = pi0146 & ~n17011;
  assign n20929 = n20923 & n20928;
  assign n20930 = ~pi0947 & ~n20927;
  assign n20931 = ~n20929 & n20930;
  assign n20932 = pi0743 & n17018;
  assign n20933 = pi0947 & ~n20924;
  assign n20934 = ~n20932 & n20933;
  assign n20935 = ~n20931 & ~n20934;
  assign n20936 = ~n20925 & ~n20935;
  assign n20937 = ~n3448 & ~n20936;
  assign n20938 = ~pi0215 & ~n20922;
  assign n20939 = ~n20937 & n20938;
  assign n20940 = n16970 & ~n20904;
  assign n20941 = pi0146 & n17042;
  assign n20942 = pi0215 & ~n20940;
  assign n20943 = ~n20941 & n20942;
  assign n20944 = ~n20939 & ~n20943;
  assign n20945 = pi0299 & ~n20944;
  assign n20946 = pi0146 & ~n16970;
  assign n20947 = ~n20940 & ~n20946;
  assign n20948 = ~n6205 & ~n20947;
  assign n20949 = ~pi0146 & ~n16990;
  assign n20950 = n16990 & n20904;
  assign n20951 = n6205 & ~n20949;
  assign n20952 = ~n20950 & n20951;
  assign n20953 = ~n20948 & ~n20952;
  assign n20954 = pi0223 & ~n20953;
  assign n20955 = n2603 & n20921;
  assign n20956 = n17018 & ~n20904;
  assign n20957 = ~n6205 & ~n20924;
  assign n20958 = ~n20956 & n20957;
  assign n20959 = n17011 & ~n20904;
  assign n20960 = n6205 & ~n20928;
  assign n20961 = ~n20959 & n20960;
  assign n20962 = ~n20958 & ~n20961;
  assign n20963 = ~n2603 & ~n20962;
  assign n20964 = ~pi0223 & ~n20955;
  assign n20965 = ~n20963 & n20964;
  assign n20966 = ~pi0299 & ~n20954;
  assign n20967 = ~n20965 & n20966;
  assign n20968 = ~n20945 & ~n20967;
  assign n20969 = pi0039 & ~n20968;
  assign n20970 = ~pi0038 & ~n20918;
  assign n20971 = ~n20969 & n20970;
  assign n20972 = n10197 & ~n20908;
  assign n20973 = ~n20971 & n20972;
  assign n20974 = ~pi0832 & ~n20899;
  assign n20975 = ~n20973 & n20974;
  assign n20976 = ~pi0146 & ~n2926;
  assign n20977 = pi0832 & ~n20976;
  assign n20978 = ~n20905 & n20977;
  assign po0303 = n20975 | n20978;
  assign n20980 = ~pi0147 & ~n2926;
  assign n20981 = ~pi0770 & pi0947;
  assign n20982 = pi0726 & n20902;
  assign n20983 = ~n20981 & ~n20982;
  assign n20984 = n2926 & ~n20983;
  assign n20985 = pi0832 & ~n20980;
  assign n20986 = ~n20984 & n20985;
  assign n20987 = ~pi0147 & ~n10197;
  assign n20988 = ~pi0947 & n16958;
  assign n20989 = ~pi0039 & ~n20988;
  assign n20990 = ~pi0299 & n17024;
  assign n20991 = pi0947 & n20990;
  assign n20992 = ~pi0947 & n17026;
  assign n20993 = n17018 & n20902;
  assign n20994 = ~n17030 & ~n20993;
  assign n20995 = ~n3448 & ~n20994;
  assign n20996 = ~pi0215 & ~n20995;
  assign n20997 = ~n20992 & n20996;
  assign n20998 = pi0215 & ~n17041;
  assign n20999 = n16970 & n20902;
  assign n21000 = n20998 & ~n20999;
  assign n21001 = ~n20997 & ~n21000;
  assign n21002 = pi0299 & ~n21001;
  assign n21003 = ~n17025 & ~n21002;
  assign n21004 = ~n20991 & n21003;
  assign n21005 = pi0039 & ~n21004;
  assign n21006 = ~n20989 & ~n21005;
  assign n21007 = ~pi0038 & n21006;
  assign n21008 = pi0038 & ~pi0947;
  assign n21009 = n17050 & n21008;
  assign n21010 = ~n21007 & ~n21009;
  assign n21011 = ~pi0770 & n21010;
  assign n21012 = pi0770 & ~n17052;
  assign n21013 = ~n21011 & ~n21012;
  assign n21014 = ~pi0147 & ~n21013;
  assign n21015 = ~n17051 & ~n21009;
  assign n21016 = pi0947 & n16958;
  assign n21017 = ~pi0039 & ~n21016;
  assign n21018 = pi0947 & n17024;
  assign n21019 = ~pi0299 & ~n21018;
  assign n21020 = pi0215 & pi0947;
  assign n21021 = n16970 & n21020;
  assign n21022 = pi0299 & ~n21021;
  assign n21023 = pi0947 & n17018;
  assign n21024 = ~n3448 & ~n21023;
  assign n21025 = pi0947 & n16653;
  assign n21026 = n3448 & ~n21025;
  assign n21027 = ~pi0215 & ~n21026;
  assign n21028 = ~n21024 & n21027;
  assign n21029 = n21022 & ~n21028;
  assign n21030 = ~n21019 & ~n21029;
  assign n21031 = pi0039 & ~n21030;
  assign n21032 = ~n21017 & ~n21031;
  assign n21033 = ~pi0038 & ~n21032;
  assign n21034 = n21015 & ~n21033;
  assign n21035 = pi0147 & ~pi0770;
  assign n21036 = n21034 & n21035;
  assign n21037 = ~pi0726 & ~n21036;
  assign n21038 = ~n21014 & n21037;
  assign n21039 = n6236 & n17050;
  assign n21040 = ~pi0147 & ~n21039;
  assign n21041 = ~n6236 & n16641;
  assign n21042 = pi0038 & ~n21041;
  assign n21043 = ~n21040 & n21042;
  assign n21044 = pi0299 & pi0947;
  assign n21045 = n17026 & ~n20902;
  assign n21046 = ~n17030 & ~n21023;
  assign n21047 = ~n3448 & ~n21046;
  assign n21048 = ~pi0215 & ~n21047;
  assign n21049 = ~n21045 & n21048;
  assign n21050 = ~n20998 & ~n21049;
  assign n21051 = pi0299 & ~n21050;
  assign n21052 = ~pi0947 & n16992;
  assign n21053 = pi0223 & ~n21052;
  assign n21054 = n16992 & ~n20902;
  assign n21055 = pi0223 & ~n21054;
  assign n21056 = n2521 & n16654;
  assign n21057 = ~n17021 & ~n21056;
  assign n21058 = n6236 & ~n21057;
  assign n21059 = ~pi0223 & ~n21058;
  assign n21060 = ~n21053 & ~n21055;
  assign n21061 = ~n21059 & n21060;
  assign n21062 = ~pi0299 & ~n21061;
  assign n21063 = ~n21044 & ~n21051;
  assign n21064 = ~n21062 & n21063;
  assign n21065 = pi0039 & n21064;
  assign n21066 = ~n6236 & n16958;
  assign n21067 = ~pi0039 & ~n21066;
  assign n21068 = n16958 & n21067;
  assign n21069 = ~n21065 & ~n21068;
  assign n21070 = ~pi0147 & n21069;
  assign n21071 = ~n6236 & n17024;
  assign n21072 = ~pi0299 & n21071;
  assign n21073 = pi0215 & ~n17037;
  assign n21074 = ~n6236 & n16653;
  assign n21075 = n3448 & n21074;
  assign n21076 = ~pi0215 & ~n21075;
  assign n21077 = ~n17033 & n21076;
  assign n21078 = pi0299 & ~n21073;
  assign n21079 = ~n21077 & n21078;
  assign n21080 = ~n21072 & ~n21079;
  assign n21081 = pi0039 & n21080;
  assign n21082 = ~n21067 & ~n21081;
  assign n21083 = pi0147 & n21082;
  assign n21084 = ~pi0038 & ~n21083;
  assign n21085 = ~n21070 & n21084;
  assign n21086 = ~pi0770 & ~n21043;
  assign n21087 = ~n21085 & n21086;
  assign n21088 = ~pi0147 & ~n16641;
  assign n21089 = n16641 & n20902;
  assign n21090 = pi0038 & ~n21089;
  assign n21091 = ~n21088 & n21090;
  assign n21092 = ~n21021 & ~n21050;
  assign n21093 = pi0299 & ~n21092;
  assign n21094 = ~n20902 & n20990;
  assign n21095 = ~n21093 & ~n21094;
  assign n21096 = pi0039 & ~n21095;
  assign n21097 = n16958 & ~n20902;
  assign n21098 = ~pi0039 & n21097;
  assign n21099 = ~n21096 & ~n21098;
  assign n21100 = ~pi0147 & n21099;
  assign n21101 = pi0215 & ~n20999;
  assign n21102 = ~n3448 & ~n20993;
  assign n21103 = pi0907 & n16653;
  assign n21104 = ~pi0947 & n21103;
  assign n21105 = n3448 & ~n21104;
  assign n21106 = ~n21102 & ~n21105;
  assign n21107 = ~pi0215 & ~n21106;
  assign n21108 = ~n21101 & ~n21107;
  assign n21109 = pi0299 & ~n21108;
  assign n21110 = n17024 & n20902;
  assign n21111 = ~pi0299 & ~n21110;
  assign n21112 = ~n21109 & ~n21111;
  assign n21113 = pi0039 & ~n21112;
  assign n21114 = n16958 & n20902;
  assign n21115 = ~pi0039 & ~n21114;
  assign n21116 = ~n21113 & ~n21115;
  assign n21117 = pi0147 & n21116;
  assign n21118 = ~pi0038 & ~n21117;
  assign n21119 = ~n21100 & n21118;
  assign n21120 = pi0770 & ~n21091;
  assign n21121 = ~n21119 & n21120;
  assign n21122 = pi0726 & ~n21087;
  assign n21123 = ~n21121 & n21122;
  assign n21124 = n10197 & ~n21123;
  assign n21125 = ~n21038 & n21124;
  assign n21126 = ~pi0832 & ~n20987;
  assign n21127 = ~n21125 & n21126;
  assign po0304 = ~n20986 & ~n21127;
  assign n21129 = pi0057 & pi0148;
  assign n21130 = n2571 & n6305;
  assign n21131 = ~pi0148 & ~n21130;
  assign n21132 = ~pi0749 & pi0947;
  assign n21133 = n21041 & ~n21132;
  assign n21134 = ~pi0148 & ~n16641;
  assign n21135 = ~n21133 & ~n21134;
  assign n21136 = pi0038 & ~n21135;
  assign n21137 = ~n17025 & ~n21109;
  assign n21138 = pi0148 & ~n21137;
  assign n21139 = ~n9737 & ~n21095;
  assign n21140 = ~pi0749 & ~n21138;
  assign n21141 = ~n21139 & n21140;
  assign n21142 = ~pi0148 & n21064;
  assign n21143 = pi0148 & n21080;
  assign n21144 = pi0749 & ~n21143;
  assign n21145 = ~n21142 & n21144;
  assign n21146 = pi0039 & ~n21141;
  assign n21147 = ~n21145 & n21146;
  assign n21148 = ~pi0148 & ~n16958;
  assign n21149 = ~pi0039 & ~n21148;
  assign n21150 = n21066 & ~n21132;
  assign n21151 = n21149 & ~n21150;
  assign n21152 = ~pi0038 & ~n21151;
  assign n21153 = ~n21147 & n21152;
  assign n21154 = pi0706 & ~n21136;
  assign n21155 = ~n21153 & n21154;
  assign n21156 = pi0749 & pi0947;
  assign n21157 = n16958 & n21156;
  assign n21158 = n21149 & ~n21157;
  assign n21159 = ~pi0148 & ~pi0749;
  assign n21160 = ~n17046 & n21159;
  assign n21161 = ~pi0148 & ~n21001;
  assign n21162 = ~n21021 & ~n21028;
  assign n21163 = pi0148 & ~n21162;
  assign n21164 = pi0299 & ~n21163;
  assign n21165 = ~n21161 & n21164;
  assign n21166 = ~pi0148 & ~n17024;
  assign n21167 = n21019 & ~n21166;
  assign n21168 = pi0749 & ~n21167;
  assign n21169 = ~n21165 & n21168;
  assign n21170 = pi0039 & ~n21160;
  assign n21171 = ~n21169 & n21170;
  assign n21172 = ~pi0038 & ~n21158;
  assign n21173 = ~n21171 & n21172;
  assign n21174 = n16641 & ~n21156;
  assign n21175 = pi0148 & ~n17050;
  assign n21176 = pi0038 & ~n21174;
  assign n21177 = ~n21175 & n21176;
  assign n21178 = ~pi0706 & ~n21177;
  assign n21179 = ~n21173 & n21178;
  assign n21180 = n21130 & ~n21179;
  assign n21181 = ~n21155 & n21180;
  assign n21182 = ~pi0057 & ~n21131;
  assign n21183 = ~n21181 & n21182;
  assign n21184 = ~pi0832 & ~n21129;
  assign n21185 = ~n21183 & n21184;
  assign n21186 = pi0706 & n20902;
  assign n21187 = n2926 & ~n21156;
  assign n21188 = ~n21186 & n21187;
  assign n21189 = pi0148 & ~n2926;
  assign n21190 = pi0832 & ~n21189;
  assign n21191 = ~n21188 & n21190;
  assign po0305 = n21185 | n21191;
  assign n21193 = ~pi0149 & ~n2926;
  assign n21194 = ~pi0755 & pi0947;
  assign n21195 = ~pi0725 & n20902;
  assign n21196 = ~n21194 & ~n21195;
  assign n21197 = n2926 & ~n21196;
  assign n21198 = pi0832 & ~n21193;
  assign n21199 = ~n21197 & n21198;
  assign n21200 = ~pi0149 & ~n10197;
  assign n21201 = n16641 & ~n21194;
  assign n21202 = pi0149 & ~n17050;
  assign n21203 = pi0038 & ~n21201;
  assign n21204 = ~n21202 & n21203;
  assign n21205 = ~pi0149 & ~n16958;
  assign n21206 = n16958 & n21194;
  assign n21207 = ~pi0039 & ~n21205;
  assign n21208 = ~n21206 & n21207;
  assign n21209 = ~pi0149 & ~n17024;
  assign n21210 = n21019 & ~n21209;
  assign n21211 = ~pi0149 & ~n21001;
  assign n21212 = ~n16116 & ~n21029;
  assign n21213 = ~n21211 & ~n21212;
  assign n21214 = ~pi0755 & ~n21210;
  assign n21215 = ~n21213 & n21214;
  assign n21216 = ~pi0149 & pi0755;
  assign n21217 = ~n17046 & n21216;
  assign n21218 = pi0039 & ~n21217;
  assign n21219 = ~n21215 & n21218;
  assign n21220 = ~pi0038 & ~n21208;
  assign n21221 = ~n21219 & n21220;
  assign n21222 = ~n21204 & ~n21221;
  assign n21223 = pi0725 & ~n21222;
  assign n21224 = ~n21114 & n21208;
  assign n21225 = ~pi0149 & n21064;
  assign n21226 = pi0149 & n21080;
  assign n21227 = ~pi0755 & ~n21226;
  assign n21228 = ~n21225 & n21227;
  assign n21229 = ~pi0149 & n21093;
  assign n21230 = pi0149 & ~n21137;
  assign n21231 = pi0755 & ~n21094;
  assign n21232 = ~n21230 & n21231;
  assign n21233 = ~n21229 & n21232;
  assign n21234 = pi0039 & ~n21233;
  assign n21235 = ~n21228 & n21234;
  assign n21236 = ~n21224 & ~n21235;
  assign n21237 = ~pi0038 & ~n21236;
  assign n21238 = ~pi0149 & ~n16641;
  assign n21239 = ~n6236 & n16667;
  assign n21240 = pi0755 & pi0947;
  assign n21241 = ~pi0039 & ~n21240;
  assign n21242 = n21239 & n21241;
  assign n21243 = pi0038 & ~n21238;
  assign n21244 = ~n21242 & n21243;
  assign n21245 = ~pi0725 & ~n21244;
  assign n21246 = ~n21237 & n21245;
  assign n21247 = ~n21223 & ~n21246;
  assign n21248 = n10197 & ~n21247;
  assign n21249 = ~pi0832 & ~n21200;
  assign n21250 = ~n21248 & n21249;
  assign po0306 = ~n21199 & ~n21250;
  assign n21252 = ~pi0150 & ~n10197;
  assign n21253 = pi0150 & ~n17050;
  assign n21254 = ~pi0751 & pi0947;
  assign n21255 = n16641 & ~n21254;
  assign n21256 = ~n21253 & ~n21255;
  assign n21257 = pi0038 & ~n21256;
  assign n21258 = pi0150 & ~n16958;
  assign n21259 = pi0751 & n16958;
  assign n21260 = ~n21258 & ~n21259;
  assign n21261 = n20989 & n21260;
  assign n21262 = ~pi0150 & n21004;
  assign n21263 = pi0150 & ~n21030;
  assign n21264 = ~pi0751 & ~n21263;
  assign n21265 = ~n21262 & n21264;
  assign n21266 = ~pi0150 & pi0751;
  assign n21267 = ~n17046 & n21266;
  assign n21268 = ~n21265 & ~n21267;
  assign n21269 = pi0039 & ~n21268;
  assign n21270 = ~pi0038 & ~n21261;
  assign n21271 = ~n21269 & n21270;
  assign n21272 = pi0701 & ~n21257;
  assign n21273 = ~n21271 & n21272;
  assign n21274 = ~pi0150 & ~n16641;
  assign n21275 = pi0751 & pi0947;
  assign n21276 = ~pi0039 & ~n21275;
  assign n21277 = n21239 & n21276;
  assign n21278 = pi0038 & ~n21274;
  assign n21279 = ~n21277 & n21278;
  assign n21280 = n21097 & ~n21254;
  assign n21281 = ~pi0039 & ~n21258;
  assign n21282 = ~n21280 & n21281;
  assign n21283 = ~pi0150 & ~n21095;
  assign n21284 = pi0150 & ~n21112;
  assign n21285 = pi0751 & ~n21284;
  assign n21286 = ~n21283 & n21285;
  assign n21287 = ~pi0150 & n21064;
  assign n21288 = pi0150 & n21080;
  assign n21289 = ~pi0751 & ~n21288;
  assign n21290 = ~n21287 & n21289;
  assign n21291 = ~n21286 & ~n21290;
  assign n21292 = pi0039 & ~n21291;
  assign n21293 = ~pi0038 & ~n21282;
  assign n21294 = ~n21292 & n21293;
  assign n21295 = ~pi0701 & ~n21279;
  assign n21296 = ~n21294 & n21295;
  assign n21297 = ~n21273 & ~n21296;
  assign n21298 = n10197 & ~n21297;
  assign n21299 = ~pi0832 & ~n21252;
  assign n21300 = ~n21298 & n21299;
  assign n21301 = ~pi0150 & ~n2926;
  assign n21302 = ~pi0701 & n20902;
  assign n21303 = ~n21254 & ~n21302;
  assign n21304 = n2926 & ~n21303;
  assign n21305 = pi0832 & ~n21301;
  assign n21306 = ~n21304 & n21305;
  assign po0307 = ~n21300 & ~n21306;
  assign n21308 = ~pi0151 & ~n2926;
  assign n21309 = ~pi0745 & pi0947;
  assign n21310 = ~pi0723 & n20902;
  assign n21311 = ~n21309 & ~n21310;
  assign n21312 = n2926 & ~n21311;
  assign n21313 = pi0832 & ~n21308;
  assign n21314 = ~n21312 & n21313;
  assign n21315 = ~pi0151 & ~n10197;
  assign n21316 = ~pi0151 & ~n16641;
  assign n21317 = pi0745 & pi0947;
  assign n21318 = ~pi0039 & ~n21317;
  assign n21319 = n21239 & n21318;
  assign n21320 = pi0038 & ~n21316;
  assign n21321 = ~n21319 & n21320;
  assign n21322 = ~pi0151 & ~n16958;
  assign n21323 = ~pi0745 & n21016;
  assign n21324 = ~n21322 & ~n21323;
  assign n21325 = n21115 & n21324;
  assign n21326 = ~n17041 & ~n20999;
  assign n21327 = ~pi0151 & n21326;
  assign n21328 = ~n17037 & ~n21327;
  assign n21329 = pi0215 & ~n21328;
  assign n21330 = pi0151 & ~n3448;
  assign n21331 = ~n17032 & n21330;
  assign n21332 = ~n17031 & ~n21331;
  assign n21333 = ~pi0151 & ~n16653;
  assign n21334 = n21105 & ~n21333;
  assign n21335 = ~n21074 & n21334;
  assign n21336 = ~pi0215 & ~n21335;
  assign n21337 = n21332 & n21336;
  assign n21338 = ~n21329 & ~n21337;
  assign n21339 = pi0299 & ~n21338;
  assign n21340 = pi0151 & ~n21071;
  assign n21341 = n21062 & ~n21340;
  assign n21342 = ~n21339 & ~n21341;
  assign n21343 = ~pi0745 & ~n21342;
  assign n21344 = n21332 & ~n21334;
  assign n21345 = n21048 & n21344;
  assign n21346 = ~n21329 & ~n21345;
  assign n21347 = ~n21021 & ~n21346;
  assign n21348 = pi0299 & ~n21347;
  assign n21349 = ~pi0151 & ~n17024;
  assign n21350 = n21111 & ~n21349;
  assign n21351 = pi0745 & ~n21350;
  assign n21352 = ~n21348 & n21351;
  assign n21353 = pi0039 & ~n21352;
  assign n21354 = ~n21343 & n21353;
  assign n21355 = ~n21325 & ~n21354;
  assign n21356 = ~pi0038 & ~n21355;
  assign n21357 = ~pi0723 & ~n21321;
  assign n21358 = ~n21356 & n21357;
  assign n21359 = pi0151 & ~n17050;
  assign n21360 = n16641 & ~n21309;
  assign n21361 = ~n21359 & ~n21360;
  assign n21362 = pi0038 & ~n21361;
  assign n21363 = ~pi0039 & ~n21324;
  assign n21364 = ~pi0745 & ~n17025;
  assign n21365 = ~pi0151 & ~n17046;
  assign n21366 = ~n21364 & n21365;
  assign n21367 = n21026 & ~n21333;
  assign n21368 = n21332 & ~n21367;
  assign n21369 = n20996 & n21368;
  assign n21370 = n21101 & ~n21328;
  assign n21371 = pi0299 & ~n21370;
  assign n21372 = ~n21369 & n21371;
  assign n21373 = ~pi0745 & ~n21019;
  assign n21374 = ~n21372 & n21373;
  assign n21375 = ~n21366 & ~n21374;
  assign n21376 = pi0039 & ~n21375;
  assign n21377 = ~pi0038 & ~n21363;
  assign n21378 = ~n21376 & n21377;
  assign n21379 = pi0723 & ~n21362;
  assign n21380 = ~n21378 & n21379;
  assign n21381 = ~n21358 & ~n21380;
  assign n21382 = n10197 & ~n21381;
  assign n21383 = ~pi0832 & ~n21315;
  assign n21384 = ~n21382 & n21383;
  assign po0308 = ~n21314 & ~n21384;
  assign n21386 = ~pi0152 & ~n10197;
  assign n21387 = ~pi0152 & ~n16641;
  assign n21388 = pi0759 & pi0947;
  assign n21389 = ~pi0039 & ~n21388;
  assign n21390 = n16667 & ~n20902;
  assign n21391 = n21389 & n21390;
  assign n21392 = pi0038 & ~n21387;
  assign n21393 = ~n21391 & n21392;
  assign n21394 = pi0152 & ~n16958;
  assign n21395 = ~n16959 & ~n21389;
  assign n21396 = ~n21394 & ~n21395;
  assign n21397 = ~n21114 & n21396;
  assign n21398 = ~pi0152 & ~n17037;
  assign n21399 = n20998 & ~n21398;
  assign n21400 = ~n20902 & ~n21073;
  assign n21401 = n21399 & ~n21400;
  assign n21402 = pi0152 & n21046;
  assign n21403 = n21102 & ~n21402;
  assign n21404 = pi0152 & ~n16653;
  assign n21405 = ~n21074 & ~n21404;
  assign n21406 = n3448 & n21405;
  assign n21407 = ~pi0215 & ~n21406;
  assign n21408 = ~n21045 & n21407;
  assign n21409 = ~n21403 & n21408;
  assign n21410 = pi0299 & ~n21401;
  assign n21411 = ~n21409 & n21410;
  assign n21412 = ~n21104 & ~n21404;
  assign n21413 = n2603 & ~n21412;
  assign n21414 = ~pi0152 & ~n17020;
  assign n21415 = n17020 & ~n20902;
  assign n21416 = ~n2603 & ~n21415;
  assign n21417 = ~n21414 & n21416;
  assign n21418 = ~n21413 & ~n21417;
  assign n21419 = ~pi0223 & ~n21418;
  assign n21420 = ~pi0152 & ~n16992;
  assign n21421 = n21055 & ~n21420;
  assign n21422 = ~pi0299 & ~n21421;
  assign n21423 = ~n21419 & n21422;
  assign n21424 = ~pi0759 & ~n21411;
  assign n21425 = ~n21423 & n21424;
  assign n21426 = ~n17032 & n21403;
  assign n21427 = n21407 & ~n21426;
  assign n21428 = pi0299 & ~n21399;
  assign n21429 = ~n21427 & n21428;
  assign n21430 = n2603 & n21405;
  assign n21431 = ~pi0947 & n17020;
  assign n21432 = ~n2603 & ~n21431;
  assign n21433 = ~n21414 & n21432;
  assign n21434 = ~n6236 & n17020;
  assign n21435 = ~n2603 & ~n21434;
  assign n21436 = ~n21433 & n21435;
  assign n21437 = ~pi0223 & ~n21430;
  assign n21438 = ~n21436 & n21437;
  assign n21439 = n21053 & ~n21420;
  assign n21440 = ~pi0299 & ~n21439;
  assign n21441 = ~n21421 & n21440;
  assign n21442 = ~n21438 & n21441;
  assign n21443 = pi0759 & ~n21429;
  assign n21444 = ~n21442 & n21443;
  assign n21445 = pi0039 & ~n21425;
  assign n21446 = ~n21444 & n21445;
  assign n21447 = ~pi0038 & ~n21397;
  assign n21448 = ~n21446 & n21447;
  assign n21449 = pi0696 & ~n21393;
  assign n21450 = ~n21448 & n21449;
  assign n21451 = ~pi0152 & ~n17050;
  assign n21452 = n16641 & ~n21388;
  assign n21453 = pi0038 & ~n21452;
  assign n21454 = ~n21451 & n21453;
  assign n21455 = ~n21025 & ~n21404;
  assign n21456 = n2603 & ~n21455;
  assign n21457 = ~n21433 & ~n21456;
  assign n21458 = ~pi0223 & ~n21457;
  assign n21459 = n21440 & ~n21458;
  assign n21460 = pi0152 & n21000;
  assign n21461 = n3448 & n21455;
  assign n21462 = ~n20995 & ~n21403;
  assign n21463 = ~n21023 & ~n21462;
  assign n21464 = ~pi0215 & ~n21461;
  assign n21465 = ~n21463 & n21464;
  assign n21466 = n21022 & ~n21460;
  assign n21467 = ~n21465 & n21466;
  assign n21468 = pi0759 & ~n21459;
  assign n21469 = ~n21467 & n21468;
  assign n21470 = ~pi0759 & ~n17046;
  assign n21471 = pi0152 & n21470;
  assign n21472 = pi0039 & ~n21471;
  assign n21473 = ~n21469 & n21472;
  assign n21474 = ~pi0038 & ~n21396;
  assign n21475 = ~n21473 & n21474;
  assign n21476 = ~pi0696 & ~n21454;
  assign n21477 = ~n21475 & n21476;
  assign n21478 = ~n21450 & ~n21477;
  assign n21479 = n10197 & ~n21478;
  assign n21480 = ~pi0832 & ~n21386;
  assign n21481 = ~n21479 & n21480;
  assign n21482 = ~pi0152 & ~n2926;
  assign n21483 = pi0696 & n20902;
  assign n21484 = n2926 & ~n21388;
  assign n21485 = ~n21483 & n21484;
  assign n21486 = pi0832 & ~n21482;
  assign n21487 = ~n21485 & n21486;
  assign po0309 = n21481 | n21487;
  assign n21489 = pi0153 & ~n2926;
  assign n21490 = pi0766 & pi0947;
  assign n21491 = n2926 & ~n21490;
  assign n21492 = pi0700 & n20902;
  assign n21493 = n21491 & ~n21492;
  assign n21494 = pi0832 & ~n21489;
  assign n21495 = ~n21493 & n21494;
  assign n21496 = pi0057 & pi0153;
  assign n21497 = ~pi0153 & ~n21130;
  assign n21498 = ~pi0153 & ~n16958;
  assign n21499 = ~pi0766 & n18147;
  assign n21500 = ~n21017 & ~n21499;
  assign n21501 = ~n21498 & ~n21500;
  assign n21502 = ~n21114 & n21501;
  assign n21503 = ~pi0153 & ~n17024;
  assign n21504 = n21111 & ~n21503;
  assign n21505 = pi0153 & ~n17037;
  assign n21506 = n20998 & ~n21505;
  assign n21507 = n21073 & ~n21506;
  assign n21508 = pi0153 & ~n3448;
  assign n21509 = ~n17032 & n21508;
  assign n21510 = ~n17031 & ~n21509;
  assign n21511 = ~pi0153 & ~n16653;
  assign n21512 = n21105 & ~n21511;
  assign n21513 = ~n21047 & ~n21512;
  assign n21514 = n21510 & n21513;
  assign n21515 = ~pi0215 & ~n21514;
  assign n21516 = ~n21021 & ~n21507;
  assign n21517 = ~n21515 & n21516;
  assign n21518 = pi0299 & ~n21517;
  assign n21519 = ~pi0766 & ~n21504;
  assign n21520 = ~n21518 & n21519;
  assign n21521 = n21026 & ~n21511;
  assign n21522 = ~n21103 & n21521;
  assign n21523 = ~pi0215 & ~n21522;
  assign n21524 = n21510 & n21523;
  assign n21525 = ~n21506 & ~n21524;
  assign n21526 = pi0299 & ~n21525;
  assign n21527 = pi0153 & ~n21071;
  assign n21528 = n21062 & ~n21527;
  assign n21529 = ~n21526 & ~n21528;
  assign n21530 = pi0766 & ~n21529;
  assign n21531 = pi0039 & ~n21520;
  assign n21532 = ~n21530 & n21531;
  assign n21533 = ~n21502 & ~n21532;
  assign n21534 = ~pi0038 & ~n21533;
  assign n21535 = ~pi0153 & ~n16641;
  assign n21536 = ~pi0766 & pi0947;
  assign n21537 = ~pi0039 & ~n21536;
  assign n21538 = n21239 & n21537;
  assign n21539 = pi0038 & ~n21535;
  assign n21540 = ~n21538 & n21539;
  assign n21541 = ~n21534 & ~n21540;
  assign n21542 = pi0700 & ~n21541;
  assign n21543 = n6284 & n21491;
  assign n21544 = pi0153 & ~n17050;
  assign n21545 = pi0038 & ~n21543;
  assign n21546 = ~n21544 & n21545;
  assign n21547 = n21019 & ~n21503;
  assign n21548 = n21000 & ~n21505;
  assign n21549 = n21510 & ~n21521;
  assign n21550 = n20996 & n21549;
  assign n21551 = pi0299 & ~n21548;
  assign n21552 = ~n21550 & n21551;
  assign n21553 = pi0766 & ~n21552;
  assign n21554 = ~n21547 & n21553;
  assign n21555 = ~pi0153 & ~pi0766;
  assign n21556 = ~n17046 & n21555;
  assign n21557 = pi0039 & ~n21556;
  assign n21558 = ~n21554 & n21557;
  assign n21559 = ~pi0038 & ~n21501;
  assign n21560 = ~n21558 & n21559;
  assign n21561 = ~pi0700 & ~n21546;
  assign n21562 = ~n21560 & n21561;
  assign n21563 = n21130 & ~n21562;
  assign n21564 = ~n21542 & n21563;
  assign n21565 = ~pi0057 & ~n21497;
  assign n21566 = ~n21564 & n21565;
  assign n21567 = ~pi0832 & ~n21496;
  assign n21568 = ~n21566 & n21567;
  assign po0310 = n21495 | n21568;
  assign n21570 = ~pi0154 & ~n2926;
  assign n21571 = ~pi0742 & pi0947;
  assign n21572 = ~pi0704 & n20902;
  assign n21573 = ~n21571 & ~n21572;
  assign n21574 = n2926 & ~n21573;
  assign n21575 = pi0832 & ~n21570;
  assign n21576 = ~n21574 & n21575;
  assign n21577 = ~pi0154 & ~n10197;
  assign n21578 = ~pi0154 & ~n16641;
  assign n21579 = n21090 & ~n21578;
  assign n21580 = ~pi0154 & ~n16958;
  assign n21581 = n21115 & ~n21580;
  assign n21582 = ~pi0154 & n21095;
  assign n21583 = pi0154 & n21112;
  assign n21584 = pi0039 & ~n21583;
  assign n21585 = ~n21582 & n21584;
  assign n21586 = ~n21581 & ~n21585;
  assign n21587 = ~pi0038 & ~n21586;
  assign n21588 = pi0742 & ~n21579;
  assign n21589 = ~n21587 & n21588;
  assign n21590 = n21042 & ~n21578;
  assign n21591 = ~n21066 & n21581;
  assign n21592 = ~pi0154 & ~n21064;
  assign n21593 = pi0154 & ~n21080;
  assign n21594 = pi0039 & ~n21593;
  assign n21595 = ~n21592 & n21594;
  assign n21596 = ~n21591 & ~n21595;
  assign n21597 = ~pi0038 & ~n21596;
  assign n21598 = ~pi0742 & ~n21590;
  assign n21599 = ~n21597 & n21598;
  assign n21600 = ~pi0704 & ~n21589;
  assign n21601 = ~n21599 & n21600;
  assign n21602 = ~pi0154 & ~n17050;
  assign n21603 = ~n21015 & ~n21602;
  assign n21604 = n21017 & ~n21580;
  assign n21605 = pi0154 & n21030;
  assign n21606 = ~pi0154 & ~n21004;
  assign n21607 = pi0039 & ~n21605;
  assign n21608 = ~n21606 & n21607;
  assign n21609 = ~n21604 & ~n21608;
  assign n21610 = ~pi0038 & ~n21609;
  assign n21611 = ~pi0742 & ~n21603;
  assign n21612 = ~n21610 & n21611;
  assign n21613 = ~pi0154 & pi0742;
  assign n21614 = ~n17052 & n21613;
  assign n21615 = pi0704 & ~n21614;
  assign n21616 = ~n21612 & n21615;
  assign n21617 = n10197 & ~n21616;
  assign n21618 = ~n21601 & n21617;
  assign n21619 = ~pi0832 & ~n21577;
  assign n21620 = ~n21618 & n21619;
  assign po0311 = ~n21576 & ~n21620;
  assign n21622 = ~pi0757 & n21034;
  assign n21623 = pi0686 & ~n21622;
  assign n21624 = ~pi0038 & ~n21082;
  assign n21625 = ~n21042 & ~n21624;
  assign n21626 = ~pi0757 & n21625;
  assign n21627 = ~pi0038 & ~n21116;
  assign n21628 = ~n21090 & ~n21627;
  assign n21629 = pi0757 & n21628;
  assign n21630 = ~pi0686 & ~n21626;
  assign n21631 = ~n21629 & n21630;
  assign n21632 = n10197 & ~n21623;
  assign n21633 = ~n21631 & n21632;
  assign n21634 = pi0155 & ~n21633;
  assign n21635 = ~pi0038 & ~n21069;
  assign n21636 = pi0038 & n21039;
  assign n21637 = ~n21635 & ~n21636;
  assign n21638 = ~pi0757 & n21637;
  assign n21639 = ~pi0038 & ~n21099;
  assign n21640 = n16641 & n21090;
  assign n21641 = ~n21639 & ~n21640;
  assign n21642 = pi0757 & n21641;
  assign n21643 = ~pi0686 & ~n21638;
  assign n21644 = ~n21642 & n21643;
  assign n21645 = ~pi0757 & n21010;
  assign n21646 = pi0757 & ~n17052;
  assign n21647 = pi0686 & ~n21646;
  assign n21648 = ~n21645 & n21647;
  assign n21649 = ~n21644 & ~n21648;
  assign n21650 = ~pi0155 & n10197;
  assign n21651 = ~n21649 & n21650;
  assign n21652 = ~n21634 & ~n21651;
  assign n21653 = ~pi0832 & ~n21652;
  assign n21654 = ~pi0155 & ~n2926;
  assign n21655 = ~pi0757 & pi0947;
  assign n21656 = ~pi0686 & n20902;
  assign n21657 = ~n21655 & ~n21656;
  assign n21658 = n2926 & ~n21657;
  assign n21659 = pi0832 & ~n21654;
  assign n21660 = ~n21658 & n21659;
  assign po0312 = ~n21653 & ~n21660;
  assign n21662 = ~pi0156 & ~n2926;
  assign n21663 = ~pi0741 & pi0947;
  assign n21664 = ~pi0724 & n20902;
  assign n21665 = ~n21663 & ~n21664;
  assign n21666 = n2926 & ~n21665;
  assign n21667 = pi0832 & ~n21662;
  assign n21668 = ~n21666 & n21667;
  assign n21669 = ~pi0741 & ~n21637;
  assign n21670 = pi0741 & ~n21641;
  assign n21671 = ~pi0724 & ~n21669;
  assign n21672 = ~n21670 & n21671;
  assign n21673 = ~pi0741 & ~n21010;
  assign n21674 = pi0741 & n17052;
  assign n21675 = pi0724 & ~n21674;
  assign n21676 = ~n21673 & n21675;
  assign n21677 = n10197 & ~n21676;
  assign n21678 = ~n21672 & n21677;
  assign n21679 = ~pi0156 & ~n21678;
  assign n21680 = ~pi0741 & ~n21625;
  assign n21681 = pi0741 & ~n21628;
  assign n21682 = ~pi0724 & ~n21680;
  assign n21683 = ~n21681 & n21682;
  assign n21684 = pi0724 & ~pi0741;
  assign n21685 = n21034 & n21684;
  assign n21686 = ~n21683 & ~n21685;
  assign n21687 = pi0156 & n10197;
  assign n21688 = ~n21686 & n21687;
  assign n21689 = ~pi0832 & ~n21688;
  assign n21690 = ~n21679 & n21689;
  assign po0313 = ~n21668 & ~n21690;
  assign n21692 = ~pi0157 & ~n2926;
  assign n21693 = ~pi0760 & pi0947;
  assign n21694 = ~pi0688 & n20902;
  assign n21695 = ~n21693 & ~n21694;
  assign n21696 = n2926 & ~n21695;
  assign n21697 = pi0832 & ~n21692;
  assign n21698 = ~n21696 & n21697;
  assign n21699 = ~pi0157 & ~n10197;
  assign n21700 = n16641 & ~n21693;
  assign n21701 = pi0157 & ~n17050;
  assign n21702 = pi0038 & ~n21700;
  assign n21703 = ~n21701 & n21702;
  assign n21704 = ~pi0157 & pi0760;
  assign n21705 = ~n17046 & n21704;
  assign n21706 = ~pi0157 & ~n17024;
  assign n21707 = n21019 & ~n21706;
  assign n21708 = ~pi0157 & ~n21001;
  assign n21709 = ~n13717 & ~n21029;
  assign n21710 = ~n21708 & ~n21709;
  assign n21711 = ~pi0760 & ~n21707;
  assign n21712 = ~n21710 & n21711;
  assign n21713 = pi0039 & ~n21705;
  assign n21714 = ~n21712 & n21713;
  assign n21715 = ~pi0157 & ~n16958;
  assign n21716 = n16958 & n21693;
  assign n21717 = ~pi0039 & ~n21715;
  assign n21718 = ~n21716 & n21717;
  assign n21719 = ~pi0038 & ~n21718;
  assign n21720 = ~n21714 & n21719;
  assign n21721 = ~n21703 & ~n21720;
  assign n21722 = pi0688 & ~n21721;
  assign n21723 = ~n21114 & n21718;
  assign n21724 = ~pi0760 & n21080;
  assign n21725 = pi0760 & ~n21112;
  assign n21726 = pi0157 & ~n21724;
  assign n21727 = ~n21725 & n21726;
  assign n21728 = pi0760 & ~n21095;
  assign n21729 = ~pi0760 & n21064;
  assign n21730 = ~pi0157 & ~n21728;
  assign n21731 = ~n21729 & n21730;
  assign n21732 = pi0039 & ~n21727;
  assign n21733 = ~n21731 & n21732;
  assign n21734 = ~n21723 & ~n21733;
  assign n21735 = ~pi0038 & ~n21734;
  assign n21736 = ~pi0157 & ~n16641;
  assign n21737 = pi0760 & pi0947;
  assign n21738 = ~pi0039 & ~n21737;
  assign n21739 = n21239 & n21738;
  assign n21740 = pi0038 & ~n21736;
  assign n21741 = ~n21739 & n21740;
  assign n21742 = ~pi0688 & ~n21741;
  assign n21743 = ~n21735 & n21742;
  assign n21744 = ~n21722 & ~n21743;
  assign n21745 = n10197 & ~n21744;
  assign n21746 = ~pi0832 & ~n21699;
  assign n21747 = ~n21745 & n21746;
  assign po0314 = ~n21698 & ~n21747;
  assign n21749 = ~pi0158 & ~n10197;
  assign n21750 = pi0158 & ~n17050;
  assign n21751 = ~pi0753 & pi0947;
  assign n21752 = n16641 & ~n21751;
  assign n21753 = ~n21750 & ~n21752;
  assign n21754 = pi0038 & ~n21753;
  assign n21755 = pi0158 & ~n16958;
  assign n21756 = pi0753 & n16958;
  assign n21757 = ~n21755 & ~n21756;
  assign n21758 = n20989 & n21757;
  assign n21759 = ~pi0158 & n21004;
  assign n21760 = pi0158 & ~n21030;
  assign n21761 = ~pi0753 & ~n21760;
  assign n21762 = ~n21759 & n21761;
  assign n21763 = ~pi0158 & pi0753;
  assign n21764 = ~n17046 & n21763;
  assign n21765 = ~n21762 & ~n21764;
  assign n21766 = pi0039 & ~n21765;
  assign n21767 = ~pi0038 & ~n21758;
  assign n21768 = ~n21766 & n21767;
  assign n21769 = pi0702 & ~n21754;
  assign n21770 = ~n21768 & n21769;
  assign n21771 = ~pi0158 & ~n16641;
  assign n21772 = pi0753 & pi0947;
  assign n21773 = ~pi0039 & ~n21772;
  assign n21774 = n21239 & n21773;
  assign n21775 = pi0038 & ~n21771;
  assign n21776 = ~n21774 & n21775;
  assign n21777 = n21097 & ~n21751;
  assign n21778 = ~pi0039 & ~n21755;
  assign n21779 = ~n21777 & n21778;
  assign n21780 = ~pi0158 & ~n21095;
  assign n21781 = pi0158 & ~n21112;
  assign n21782 = pi0753 & ~n21781;
  assign n21783 = ~n21780 & n21782;
  assign n21784 = ~pi0158 & n21064;
  assign n21785 = pi0158 & n21080;
  assign n21786 = ~pi0753 & ~n21785;
  assign n21787 = ~n21784 & n21786;
  assign n21788 = ~n21783 & ~n21787;
  assign n21789 = pi0039 & ~n21788;
  assign n21790 = ~pi0038 & ~n21779;
  assign n21791 = ~n21789 & n21790;
  assign n21792 = ~pi0702 & ~n21776;
  assign n21793 = ~n21791 & n21792;
  assign n21794 = ~n21770 & ~n21793;
  assign n21795 = n10197 & ~n21794;
  assign n21796 = ~pi0832 & ~n21749;
  assign n21797 = ~n21795 & n21796;
  assign n21798 = ~pi0158 & ~n2926;
  assign n21799 = ~pi0702 & n20902;
  assign n21800 = ~n21751 & ~n21799;
  assign n21801 = n2926 & ~n21800;
  assign n21802 = pi0832 & ~n21798;
  assign n21803 = ~n21801 & n21802;
  assign po0315 = ~n21797 & ~n21803;
  assign n21805 = ~pi0159 & ~n10197;
  assign n21806 = pi0159 & ~n17050;
  assign n21807 = ~pi0754 & pi0947;
  assign n21808 = n16641 & ~n21807;
  assign n21809 = ~n21806 & ~n21808;
  assign n21810 = pi0038 & ~n21809;
  assign n21811 = pi0159 & ~n16958;
  assign n21812 = pi0754 & n16958;
  assign n21813 = ~n21811 & ~n21812;
  assign n21814 = n20989 & n21813;
  assign n21815 = ~pi0159 & n21004;
  assign n21816 = pi0159 & ~n21030;
  assign n21817 = ~pi0754 & ~n21816;
  assign n21818 = ~n21815 & n21817;
  assign n21819 = ~pi0159 & pi0754;
  assign n21820 = ~n17046 & n21819;
  assign n21821 = ~n21818 & ~n21820;
  assign n21822 = pi0039 & ~n21821;
  assign n21823 = ~pi0038 & ~n21814;
  assign n21824 = ~n21822 & n21823;
  assign n21825 = pi0709 & ~n21810;
  assign n21826 = ~n21824 & n21825;
  assign n21827 = ~pi0159 & ~n16641;
  assign n21828 = pi0754 & pi0947;
  assign n21829 = ~pi0039 & ~n21828;
  assign n21830 = n21239 & n21829;
  assign n21831 = pi0038 & ~n21827;
  assign n21832 = ~n21830 & n21831;
  assign n21833 = n21097 & ~n21807;
  assign n21834 = ~pi0039 & ~n21811;
  assign n21835 = ~n21833 & n21834;
  assign n21836 = ~pi0159 & ~n21095;
  assign n21837 = pi0159 & ~n21112;
  assign n21838 = pi0754 & ~n21837;
  assign n21839 = ~n21836 & n21838;
  assign n21840 = ~pi0159 & n21064;
  assign n21841 = pi0159 & n21080;
  assign n21842 = ~pi0754 & ~n21841;
  assign n21843 = ~n21840 & n21842;
  assign n21844 = ~n21839 & ~n21843;
  assign n21845 = pi0039 & ~n21844;
  assign n21846 = ~pi0038 & ~n21835;
  assign n21847 = ~n21845 & n21846;
  assign n21848 = ~pi0709 & ~n21832;
  assign n21849 = ~n21847 & n21848;
  assign n21850 = ~n21826 & ~n21849;
  assign n21851 = n10197 & ~n21850;
  assign n21852 = ~pi0832 & ~n21805;
  assign n21853 = ~n21851 & n21852;
  assign n21854 = ~pi0159 & ~n2926;
  assign n21855 = ~pi0709 & n20902;
  assign n21856 = ~n21807 & ~n21855;
  assign n21857 = n2926 & ~n21856;
  assign n21858 = pi0832 & ~n21854;
  assign n21859 = ~n21857 & n21858;
  assign po0316 = ~n21853 & ~n21859;
  assign n21861 = ~pi0160 & ~n2926;
  assign n21862 = ~pi0756 & pi0947;
  assign n21863 = ~pi0734 & n20902;
  assign n21864 = ~n21862 & ~n21863;
  assign n21865 = n2926 & ~n21864;
  assign n21866 = pi0832 & ~n21861;
  assign n21867 = ~n21865 & n21866;
  assign n21868 = ~pi0160 & ~n10197;
  assign n21869 = n16641 & ~n21862;
  assign n21870 = pi0160 & ~n17050;
  assign n21871 = pi0038 & ~n21869;
  assign n21872 = ~n21870 & n21871;
  assign n21873 = ~pi0160 & ~n16958;
  assign n21874 = n16958 & n21862;
  assign n21875 = ~pi0039 & ~n21873;
  assign n21876 = ~n21874 & n21875;
  assign n21877 = ~pi0160 & ~n21001;
  assign n21878 = pi0160 & ~n21162;
  assign n21879 = pi0299 & ~n21878;
  assign n21880 = ~n21877 & n21879;
  assign n21881 = ~pi0160 & ~n17024;
  assign n21882 = n21019 & ~n21881;
  assign n21883 = ~pi0756 & ~n21882;
  assign n21884 = ~n21880 & n21883;
  assign n21885 = ~pi0160 & pi0756;
  assign n21886 = ~n17046 & n21885;
  assign n21887 = pi0039 & ~n21886;
  assign n21888 = ~n21884 & n21887;
  assign n21889 = ~pi0038 & ~n21876;
  assign n21890 = ~n21888 & n21889;
  assign n21891 = ~n21872 & ~n21890;
  assign n21892 = pi0734 & ~n21891;
  assign n21893 = ~n21114 & n21876;
  assign n21894 = ~pi0160 & n21064;
  assign n21895 = pi0160 & n21080;
  assign n21896 = ~pi0756 & ~n21895;
  assign n21897 = ~n21894 & n21896;
  assign n21898 = pi0160 & ~n21137;
  assign n21899 = ~pi0160 & n21093;
  assign n21900 = pi0756 & ~n21094;
  assign n21901 = ~n21898 & n21900;
  assign n21902 = ~n21899 & n21901;
  assign n21903 = pi0039 & ~n21902;
  assign n21904 = ~n21897 & n21903;
  assign n21905 = ~n21893 & ~n21904;
  assign n21906 = ~pi0038 & ~n21905;
  assign n21907 = ~pi0160 & ~n16641;
  assign n21908 = pi0756 & pi0947;
  assign n21909 = ~pi0039 & ~n21908;
  assign n21910 = n21239 & n21909;
  assign n21911 = pi0038 & ~n21907;
  assign n21912 = ~n21910 & n21911;
  assign n21913 = ~pi0734 & ~n21912;
  assign n21914 = ~n21906 & n21913;
  assign n21915 = ~n21892 & ~n21914;
  assign n21916 = n10197 & ~n21915;
  assign n21917 = ~pi0832 & ~n21868;
  assign n21918 = ~n21916 & n21917;
  assign po0317 = ~n21867 & ~n21918;
  assign n21920 = ~pi0161 & ~n10197;
  assign n21921 = ~pi0161 & ~n16641;
  assign n21922 = pi0758 & pi0947;
  assign n21923 = ~pi0039 & ~n21922;
  assign n21924 = n21390 & n21923;
  assign n21925 = pi0038 & ~n21921;
  assign n21926 = ~n21924 & n21925;
  assign n21927 = n16958 & n21922;
  assign n21928 = pi0161 & ~n16958;
  assign n21929 = ~pi0039 & ~n21927;
  assign n21930 = ~n21928 & n21929;
  assign n21931 = ~n21114 & n21930;
  assign n21932 = ~pi0161 & ~n17037;
  assign n21933 = n20998 & ~n21932;
  assign n21934 = ~n21400 & n21933;
  assign n21935 = pi0161 & n21046;
  assign n21936 = n21102 & ~n21935;
  assign n21937 = pi0161 & ~n16653;
  assign n21938 = ~n21074 & ~n21937;
  assign n21939 = n3448 & n21938;
  assign n21940 = ~pi0215 & ~n21939;
  assign n21941 = ~n21045 & n21940;
  assign n21942 = ~n21936 & n21941;
  assign n21943 = pi0299 & ~n21934;
  assign n21944 = ~n21942 & n21943;
  assign n21945 = ~n21104 & ~n21937;
  assign n21946 = n2603 & ~n21945;
  assign n21947 = ~pi0161 & ~n17020;
  assign n21948 = n21416 & ~n21947;
  assign n21949 = ~n21946 & ~n21948;
  assign n21950 = ~pi0223 & ~n21949;
  assign n21951 = ~pi0161 & ~n16992;
  assign n21952 = n21055 & ~n21951;
  assign n21953 = ~pi0299 & ~n21952;
  assign n21954 = ~n21950 & n21953;
  assign n21955 = ~pi0758 & ~n21944;
  assign n21956 = ~n21954 & n21955;
  assign n21957 = ~n17032 & n21936;
  assign n21958 = n21940 & ~n21957;
  assign n21959 = pi0299 & ~n21933;
  assign n21960 = ~n21958 & n21959;
  assign n21961 = n2603 & n21938;
  assign n21962 = n21432 & ~n21947;
  assign n21963 = n21435 & ~n21962;
  assign n21964 = ~pi0223 & ~n21961;
  assign n21965 = ~n21963 & n21964;
  assign n21966 = n21053 & ~n21951;
  assign n21967 = ~pi0299 & ~n21966;
  assign n21968 = ~n21952 & n21967;
  assign n21969 = ~n21965 & n21968;
  assign n21970 = pi0758 & ~n21960;
  assign n21971 = ~n21969 & n21970;
  assign n21972 = pi0039 & ~n21956;
  assign n21973 = ~n21971 & n21972;
  assign n21974 = ~pi0038 & ~n21931;
  assign n21975 = ~n21973 & n21974;
  assign n21976 = pi0736 & ~n21926;
  assign n21977 = ~n21975 & n21976;
  assign n21978 = ~pi0161 & ~n17050;
  assign n21979 = n16641 & ~n21922;
  assign n21980 = pi0038 & ~n21979;
  assign n21981 = ~n21978 & n21980;
  assign n21982 = ~n21025 & ~n21937;
  assign n21983 = n2603 & ~n21982;
  assign n21984 = ~n21962 & ~n21983;
  assign n21985 = ~pi0223 & ~n21984;
  assign n21986 = n21967 & ~n21985;
  assign n21987 = pi0161 & n21000;
  assign n21988 = n3448 & n21982;
  assign n21989 = ~n20995 & ~n21936;
  assign n21990 = ~n21023 & ~n21989;
  assign n21991 = ~pi0215 & ~n21988;
  assign n21992 = ~n21990 & n21991;
  assign n21993 = n21022 & ~n21987;
  assign n21994 = ~n21992 & n21993;
  assign n21995 = pi0758 & ~n21986;
  assign n21996 = ~n21994 & n21995;
  assign n21997 = pi0161 & n19958;
  assign n21998 = pi0039 & ~n21997;
  assign n21999 = ~n21996 & n21998;
  assign n22000 = ~pi0038 & ~n21930;
  assign n22001 = ~n21999 & n22000;
  assign n22002 = ~pi0736 & ~n21981;
  assign n22003 = ~n22001 & n22002;
  assign n22004 = ~n21977 & ~n22003;
  assign n22005 = n10197 & ~n22004;
  assign n22006 = ~pi0832 & ~n21920;
  assign n22007 = ~n22005 & n22006;
  assign n22008 = ~pi0161 & ~n2926;
  assign n22009 = pi0736 & n20902;
  assign n22010 = n2926 & ~n21922;
  assign n22011 = ~n22009 & n22010;
  assign n22012 = pi0832 & ~n22008;
  assign n22013 = ~n22011 & n22012;
  assign po0318 = n22007 | n22013;
  assign n22015 = ~pi0162 & ~n10197;
  assign n22016 = ~pi0761 & pi0947;
  assign n22017 = n16641 & ~n22016;
  assign n22018 = pi0162 & ~n17050;
  assign n22019 = pi0038 & ~n22017;
  assign n22020 = ~n22018 & n22019;
  assign n22021 = ~pi0162 & ~n16958;
  assign n22022 = n16958 & n22016;
  assign n22023 = ~pi0039 & ~n22021;
  assign n22024 = ~n22022 & n22023;
  assign n22025 = n14933 & ~n21162;
  assign n22026 = ~n20991 & ~n22025;
  assign n22027 = ~pi0761 & ~n22026;
  assign n22028 = ~pi0761 & n21003;
  assign n22029 = pi0761 & n17046;
  assign n22030 = ~pi0162 & ~n22029;
  assign n22031 = ~n22028 & n22030;
  assign n22032 = pi0039 & ~n22027;
  assign n22033 = ~n22031 & n22032;
  assign n22034 = ~pi0038 & ~n22024;
  assign n22035 = ~n22033 & n22034;
  assign n22036 = ~n22020 & ~n22035;
  assign n22037 = pi0738 & ~n22036;
  assign n22038 = ~n21114 & n22024;
  assign n22039 = pi0162 & ~n21137;
  assign n22040 = ~n14933 & ~n21095;
  assign n22041 = pi0761 & ~n22039;
  assign n22042 = ~n22040 & n22041;
  assign n22043 = ~pi0162 & n21064;
  assign n22044 = pi0162 & n21080;
  assign n22045 = ~pi0761 & ~n22044;
  assign n22046 = ~n22043 & n22045;
  assign n22047 = pi0039 & ~n22042;
  assign n22048 = ~n22046 & n22047;
  assign n22049 = ~n22038 & ~n22048;
  assign n22050 = ~pi0038 & ~n22049;
  assign n22051 = ~pi0162 & ~n16641;
  assign n22052 = pi0761 & pi0947;
  assign n22053 = ~pi0039 & ~n22052;
  assign n22054 = n21239 & n22053;
  assign n22055 = pi0038 & ~n22051;
  assign n22056 = ~n22054 & n22055;
  assign n22057 = ~pi0738 & ~n22056;
  assign n22058 = ~n22050 & n22057;
  assign n22059 = ~n22037 & ~n22058;
  assign n22060 = n10197 & ~n22059;
  assign n22061 = ~pi0832 & ~n22015;
  assign n22062 = ~n22060 & n22061;
  assign n22063 = ~pi0162 & ~n2926;
  assign n22064 = ~pi0738 & n20902;
  assign n22065 = ~n22016 & ~n22064;
  assign n22066 = n2926 & ~n22065;
  assign n22067 = pi0832 & ~n22063;
  assign n22068 = ~n22066 & n22067;
  assign po0319 = ~n22062 & ~n22068;
  assign n22070 = ~pi0163 & ~n2926;
  assign n22071 = ~pi0777 & pi0947;
  assign n22072 = ~pi0737 & n20902;
  assign n22073 = ~n22071 & ~n22072;
  assign n22074 = n2926 & ~n22073;
  assign n22075 = pi0832 & ~n22070;
  assign n22076 = ~n22074 & n22075;
  assign n22077 = ~pi0163 & ~n10197;
  assign n22078 = n16641 & ~n22071;
  assign n22079 = pi0163 & ~n17050;
  assign n22080 = pi0038 & ~n22078;
  assign n22081 = ~n22079 & n22080;
  assign n22082 = ~pi0163 & ~n16958;
  assign n22083 = n16958 & n22071;
  assign n22084 = ~pi0039 & ~n22082;
  assign n22085 = ~n22083 & n22084;
  assign n22086 = ~pi0163 & ~n17024;
  assign n22087 = n21019 & ~n22086;
  assign n22088 = ~pi0163 & ~n21001;
  assign n22089 = ~n14735 & ~n21029;
  assign n22090 = ~n22088 & ~n22089;
  assign n22091 = ~pi0777 & ~n22087;
  assign n22092 = ~n22090 & n22091;
  assign n22093 = ~pi0163 & pi0777;
  assign n22094 = ~n17046 & n22093;
  assign n22095 = pi0039 & ~n22094;
  assign n22096 = ~n22092 & n22095;
  assign n22097 = ~pi0038 & ~n22085;
  assign n22098 = ~n22096 & n22097;
  assign n22099 = ~n22081 & ~n22098;
  assign n22100 = pi0737 & ~n22099;
  assign n22101 = ~n21114 & n22085;
  assign n22102 = ~pi0163 & n21064;
  assign n22103 = pi0163 & n21080;
  assign n22104 = ~pi0777 & ~n22103;
  assign n22105 = ~n22102 & n22104;
  assign n22106 = ~pi0163 & n21093;
  assign n22107 = pi0163 & ~n21137;
  assign n22108 = pi0777 & ~n21094;
  assign n22109 = ~n22107 & n22108;
  assign n22110 = ~n22106 & n22109;
  assign n22111 = pi0039 & ~n22110;
  assign n22112 = ~n22105 & n22111;
  assign n22113 = ~n22101 & ~n22112;
  assign n22114 = ~pi0038 & ~n22113;
  assign n22115 = ~pi0163 & ~n16641;
  assign n22116 = pi0777 & pi0947;
  assign n22117 = ~pi0039 & ~n22116;
  assign n22118 = n21239 & n22117;
  assign n22119 = pi0038 & ~n22115;
  assign n22120 = ~n22118 & n22119;
  assign n22121 = ~pi0737 & ~n22120;
  assign n22122 = ~n22114 & n22121;
  assign n22123 = ~n22100 & ~n22122;
  assign n22124 = n10197 & ~n22123;
  assign n22125 = ~pi0832 & ~n22077;
  assign n22126 = ~n22124 & n22125;
  assign po0320 = ~n22076 & ~n22126;
  assign n22128 = ~pi0164 & ~n2926;
  assign n22129 = ~pi0752 & pi0947;
  assign n22130 = pi0703 & n20902;
  assign n22131 = ~n22129 & ~n22130;
  assign n22132 = n2926 & ~n22131;
  assign n22133 = pi0832 & ~n22128;
  assign n22134 = ~n22132 & n22133;
  assign n22135 = ~pi0164 & ~n10197;
  assign n22136 = ~pi0164 & ~n21039;
  assign n22137 = n21042 & ~n22136;
  assign n22138 = ~pi0164 & n21069;
  assign n22139 = pi0164 & n21082;
  assign n22140 = ~pi0038 & ~n22139;
  assign n22141 = ~n22138 & n22140;
  assign n22142 = ~pi0752 & ~n22137;
  assign n22143 = ~n22141 & n22142;
  assign n22144 = ~pi0164 & ~n16641;
  assign n22145 = n21090 & ~n22144;
  assign n22146 = ~pi0164 & n21099;
  assign n22147 = pi0164 & n21116;
  assign n22148 = ~pi0038 & ~n22147;
  assign n22149 = ~n22146 & n22148;
  assign n22150 = pi0752 & ~n22145;
  assign n22151 = ~n22149 & n22150;
  assign n22152 = ~n22143 & ~n22151;
  assign n22153 = pi0703 & ~n22152;
  assign n22154 = pi0752 & n17052;
  assign n22155 = ~pi0752 & n21034;
  assign n22156 = pi0164 & ~n22155;
  assign n22157 = pi0164 & ~n21009;
  assign n22158 = ~pi0752 & ~n22157;
  assign n22159 = ~n21010 & n22158;
  assign n22160 = ~pi0703 & ~n22154;
  assign n22161 = ~n22156 & n22160;
  assign n22162 = ~n22159 & n22161;
  assign n22163 = ~n22153 & ~n22162;
  assign n22164 = n10197 & ~n22163;
  assign n22165 = ~pi0832 & ~n22135;
  assign n22166 = ~n22164 & n22165;
  assign po0321 = ~n22134 & ~n22166;
  assign n22168 = ~pi0165 & ~n2926;
  assign n22169 = ~pi0774 & pi0947;
  assign n22170 = pi0687 & n20902;
  assign n22171 = ~n22169 & ~n22170;
  assign n22172 = n2926 & ~n22171;
  assign n22173 = pi0832 & ~n22168;
  assign n22174 = ~n22172 & n22173;
  assign n22175 = ~pi0165 & ~n10197;
  assign n22176 = ~pi0165 & ~n21039;
  assign n22177 = n21042 & ~n22176;
  assign n22178 = ~pi0165 & n21069;
  assign n22179 = pi0165 & n21082;
  assign n22180 = ~pi0038 & ~n22179;
  assign n22181 = ~n22178 & n22180;
  assign n22182 = ~pi0774 & ~n22177;
  assign n22183 = ~n22181 & n22182;
  assign n22184 = ~pi0165 & ~n16641;
  assign n22185 = n21090 & ~n22184;
  assign n22186 = ~pi0165 & n21099;
  assign n22187 = pi0165 & n21116;
  assign n22188 = ~pi0038 & ~n22187;
  assign n22189 = ~n22186 & n22188;
  assign n22190 = pi0774 & ~n22185;
  assign n22191 = ~n22189 & n22190;
  assign n22192 = ~n22183 & ~n22191;
  assign n22193 = pi0687 & ~n22192;
  assign n22194 = pi0774 & n17052;
  assign n22195 = ~pi0774 & n21034;
  assign n22196 = pi0165 & ~n22195;
  assign n22197 = pi0165 & ~n21009;
  assign n22198 = ~pi0774 & ~n22197;
  assign n22199 = ~n21010 & n22198;
  assign n22200 = ~pi0687 & ~n22194;
  assign n22201 = ~n22196 & n22200;
  assign n22202 = ~n22199 & n22201;
  assign n22203 = ~n22193 & ~n22202;
  assign n22204 = n10197 & ~n22203;
  assign n22205 = ~pi0832 & ~n22175;
  assign n22206 = ~n22204 & n22205;
  assign po0322 = ~n22174 & ~n22206;
  assign n22208 = ~pi0166 & ~n10197;
  assign n22209 = ~pi0166 & ~n17050;
  assign n22210 = pi0772 & pi0947;
  assign n22211 = n16641 & ~n22210;
  assign n22212 = pi0038 & ~n22211;
  assign n22213 = ~n22209 & n22212;
  assign n22214 = pi0166 & ~n16958;
  assign n22215 = ~pi0039 & ~n22210;
  assign n22216 = ~n16959 & ~n22215;
  assign n22217 = ~n22214 & ~n22216;
  assign n22218 = ~pi0166 & ~n16992;
  assign n22219 = n21053 & ~n22218;
  assign n22220 = ~pi0299 & ~n22219;
  assign n22221 = pi0166 & ~n16653;
  assign n22222 = ~n21025 & ~n22221;
  assign n22223 = n2603 & ~n22222;
  assign n22224 = ~pi0166 & ~n17020;
  assign n22225 = n21432 & ~n22224;
  assign n22226 = ~n22223 & ~n22225;
  assign n22227 = ~pi0223 & ~n22226;
  assign n22228 = n22220 & ~n22227;
  assign n22229 = pi0166 & n21000;
  assign n22230 = n3448 & n22222;
  assign n22231 = pi0166 & n21046;
  assign n22232 = n21102 & ~n22231;
  assign n22233 = ~n20995 & ~n22232;
  assign n22234 = ~n21023 & ~n22233;
  assign n22235 = ~pi0215 & ~n22230;
  assign n22236 = ~n22234 & n22235;
  assign n22237 = n21022 & ~n22229;
  assign n22238 = ~n22236 & n22237;
  assign n22239 = pi0772 & ~n22228;
  assign n22240 = ~n22238 & n22239;
  assign n22241 = ~pi0772 & ~n17046;
  assign n22242 = pi0166 & n22241;
  assign n22243 = pi0039 & ~n22242;
  assign n22244 = ~n22240 & n22243;
  assign n22245 = ~pi0038 & ~n22217;
  assign n22246 = ~n22244 & n22245;
  assign n22247 = ~pi0727 & ~n22213;
  assign n22248 = ~n22246 & n22247;
  assign n22249 = n21390 & n22215;
  assign n22250 = ~pi0166 & ~n16641;
  assign n22251 = pi0038 & ~n22249;
  assign n22252 = ~n22250 & n22251;
  assign n22253 = ~n21114 & n22217;
  assign n22254 = ~n6236 & n16992;
  assign n22255 = ~pi0166 & ~n22254;
  assign n22256 = n21055 & ~n22255;
  assign n22257 = ~n21074 & ~n22221;
  assign n22258 = n2603 & n22257;
  assign n22259 = ~pi0223 & ~n22258;
  assign n22260 = ~n21415 & ~n22224;
  assign n22261 = n21435 & ~n22260;
  assign n22262 = n22259 & ~n22261;
  assign n22263 = n22220 & ~n22256;
  assign n22264 = ~n22262 & n22263;
  assign n22265 = ~pi0166 & ~n17037;
  assign n22266 = n20998 & ~n22265;
  assign n22267 = n3448 & n22257;
  assign n22268 = ~pi0215 & ~n22267;
  assign n22269 = ~n17032 & n22232;
  assign n22270 = n22268 & ~n22269;
  assign n22271 = pi0299 & ~n22266;
  assign n22272 = ~n22270 & n22271;
  assign n22273 = pi0772 & ~n22264;
  assign n22274 = ~n22272 & n22273;
  assign n22275 = ~n2603 & ~n22260;
  assign n22276 = n2603 & n21025;
  assign n22277 = n22259 & ~n22276;
  assign n22278 = ~n22275 & n22277;
  assign n22279 = ~pi0299 & ~n22256;
  assign n22280 = ~n22278 & n22279;
  assign n22281 = ~n21045 & n22268;
  assign n22282 = ~n22232 & n22281;
  assign n22283 = ~n21400 & n22266;
  assign n22284 = pi0299 & ~n22283;
  assign n22285 = ~n22282 & n22284;
  assign n22286 = ~pi0772 & ~n22280;
  assign n22287 = ~n22285 & n22286;
  assign n22288 = pi0039 & ~n22274;
  assign n22289 = ~n22287 & n22288;
  assign n22290 = ~pi0038 & ~n22253;
  assign n22291 = ~n22289 & n22290;
  assign n22292 = pi0727 & ~n22252;
  assign n22293 = ~n22291 & n22292;
  assign n22294 = ~n22248 & ~n22293;
  assign n22295 = n10197 & ~n22294;
  assign n22296 = ~pi0832 & ~n22208;
  assign n22297 = ~n22295 & n22296;
  assign n22298 = ~pi0166 & ~n2926;
  assign n22299 = pi0727 & n20902;
  assign n22300 = n2926 & ~n22210;
  assign n22301 = ~n22299 & n22300;
  assign n22302 = pi0832 & ~n22298;
  assign n22303 = ~n22301 & n22302;
  assign po0323 = n22297 | n22303;
  assign n22305 = ~pi0167 & ~n2926;
  assign n22306 = ~pi0768 & pi0947;
  assign n22307 = pi0705 & n20902;
  assign n22308 = ~n22306 & ~n22307;
  assign n22309 = n2926 & ~n22308;
  assign n22310 = pi0832 & ~n22305;
  assign n22311 = ~n22309 & n22310;
  assign n22312 = ~pi0167 & ~n10197;
  assign n22313 = pi0768 & ~n17052;
  assign n22314 = ~pi0167 & n22313;
  assign n22315 = ~pi0167 & ~n17050;
  assign n22316 = ~n21015 & ~n22315;
  assign n22317 = pi0167 & n21032;
  assign n22318 = ~pi0167 & ~n21006;
  assign n22319 = ~pi0038 & ~n22317;
  assign n22320 = ~n22318 & n22319;
  assign n22321 = ~pi0768 & ~n22316;
  assign n22322 = ~n22320 & n22321;
  assign n22323 = ~pi0705 & ~n22314;
  assign n22324 = ~n22322 & n22323;
  assign n22325 = ~pi0167 & ~n16641;
  assign n22326 = n21090 & ~n22325;
  assign n22327 = ~pi0167 & n21099;
  assign n22328 = pi0167 & n21116;
  assign n22329 = ~pi0038 & ~n22328;
  assign n22330 = ~n22327 & n22329;
  assign n22331 = pi0768 & ~n22326;
  assign n22332 = ~n22330 & n22331;
  assign n22333 = ~pi0167 & ~n21039;
  assign n22334 = n21042 & ~n22333;
  assign n22335 = ~pi0167 & n21069;
  assign n22336 = pi0167 & n21082;
  assign n22337 = ~pi0038 & ~n22336;
  assign n22338 = ~n22335 & n22337;
  assign n22339 = ~pi0768 & ~n22334;
  assign n22340 = ~n22338 & n22339;
  assign n22341 = pi0705 & ~n22332;
  assign n22342 = ~n22340 & n22341;
  assign n22343 = n10197 & ~n22324;
  assign n22344 = ~n22342 & n22343;
  assign n22345 = ~pi0832 & ~n22312;
  assign n22346 = ~n22344 & n22345;
  assign po0324 = ~n22311 & ~n22346;
  assign n22348 = pi0168 & ~n2926;
  assign n22349 = pi0763 & pi0947;
  assign n22350 = n2926 & ~n22349;
  assign n22351 = pi0699 & n20902;
  assign n22352 = n22350 & ~n22351;
  assign n22353 = pi0832 & ~n22348;
  assign n22354 = ~n22352 & n22353;
  assign n22355 = pi0057 & pi0168;
  assign n22356 = ~pi0168 & ~n21130;
  assign n22357 = ~pi0168 & ~n16958;
  assign n22358 = ~pi0763 & n18147;
  assign n22359 = ~n21017 & ~n22358;
  assign n22360 = ~n22357 & ~n22359;
  assign n22361 = ~n21114 & n22360;
  assign n22362 = ~pi0168 & ~n17024;
  assign n22363 = n21111 & ~n22362;
  assign n22364 = pi0168 & ~n17037;
  assign n22365 = n20998 & ~n22364;
  assign n22366 = n21073 & ~n22365;
  assign n22367 = pi0168 & ~n3448;
  assign n22368 = ~n17032 & n22367;
  assign n22369 = ~n17031 & ~n22368;
  assign n22370 = ~pi0168 & ~n16653;
  assign n22371 = n21105 & ~n22370;
  assign n22372 = ~n21047 & ~n22371;
  assign n22373 = n22369 & n22372;
  assign n22374 = ~pi0215 & ~n22373;
  assign n22375 = ~n21021 & ~n22366;
  assign n22376 = ~n22374 & n22375;
  assign n22377 = pi0299 & ~n22376;
  assign n22378 = ~pi0763 & ~n22363;
  assign n22379 = ~n22377 & n22378;
  assign n22380 = n21026 & ~n22370;
  assign n22381 = ~n21103 & n22380;
  assign n22382 = ~pi0215 & ~n22381;
  assign n22383 = n22369 & n22382;
  assign n22384 = ~n22365 & ~n22383;
  assign n22385 = pi0299 & ~n22384;
  assign n22386 = pi0168 & ~n21071;
  assign n22387 = n21062 & ~n22386;
  assign n22388 = ~n22385 & ~n22387;
  assign n22389 = pi0763 & ~n22388;
  assign n22390 = pi0039 & ~n22379;
  assign n22391 = ~n22389 & n22390;
  assign n22392 = ~n22361 & ~n22391;
  assign n22393 = ~pi0038 & ~n22392;
  assign n22394 = ~pi0168 & ~n16641;
  assign n22395 = ~pi0763 & pi0947;
  assign n22396 = ~pi0039 & ~n22395;
  assign n22397 = n21239 & n22396;
  assign n22398 = pi0038 & ~n22394;
  assign n22399 = ~n22397 & n22398;
  assign n22400 = ~n22393 & ~n22399;
  assign n22401 = pi0699 & ~n22400;
  assign n22402 = n6284 & n22350;
  assign n22403 = pi0168 & ~n17050;
  assign n22404 = pi0038 & ~n22402;
  assign n22405 = ~n22403 & n22404;
  assign n22406 = n21019 & ~n22362;
  assign n22407 = n21000 & ~n22364;
  assign n22408 = n22369 & ~n22380;
  assign n22409 = n20996 & n22408;
  assign n22410 = pi0299 & ~n22407;
  assign n22411 = ~n22409 & n22410;
  assign n22412 = pi0763 & ~n22411;
  assign n22413 = ~n22406 & n22412;
  assign n22414 = ~pi0168 & ~pi0763;
  assign n22415 = ~n17046 & n22414;
  assign n22416 = pi0039 & ~n22415;
  assign n22417 = ~n22413 & n22416;
  assign n22418 = ~pi0038 & ~n22360;
  assign n22419 = ~n22417 & n22418;
  assign n22420 = ~pi0699 & ~n22405;
  assign n22421 = ~n22419 & n22420;
  assign n22422 = n21130 & ~n22421;
  assign n22423 = ~n22401 & n22422;
  assign n22424 = ~pi0057 & ~n22356;
  assign n22425 = ~n22423 & n22424;
  assign n22426 = ~pi0832 & ~n22355;
  assign n22427 = ~n22425 & n22426;
  assign po0325 = n22354 | n22427;
  assign n22429 = pi0169 & ~n2926;
  assign n22430 = pi0746 & pi0947;
  assign n22431 = n2926 & ~n22430;
  assign n22432 = pi0729 & n20902;
  assign n22433 = n22431 & ~n22432;
  assign n22434 = pi0832 & ~n22429;
  assign n22435 = ~n22433 & n22434;
  assign n22436 = pi0057 & pi0169;
  assign n22437 = ~pi0169 & ~n21130;
  assign n22438 = ~pi0169 & ~n16958;
  assign n22439 = ~pi0746 & n18147;
  assign n22440 = ~n21017 & ~n22439;
  assign n22441 = ~n22438 & ~n22440;
  assign n22442 = ~n21114 & n22441;
  assign n22443 = ~pi0169 & ~n17024;
  assign n22444 = n21111 & ~n22443;
  assign n22445 = pi0169 & ~n17037;
  assign n22446 = n20998 & ~n22445;
  assign n22447 = n21073 & ~n22446;
  assign n22448 = pi0169 & ~n3448;
  assign n22449 = ~n17032 & n22448;
  assign n22450 = ~n17031 & ~n22449;
  assign n22451 = ~pi0169 & ~n16653;
  assign n22452 = n21105 & ~n22451;
  assign n22453 = ~n21047 & ~n22452;
  assign n22454 = n22450 & n22453;
  assign n22455 = ~pi0215 & ~n22454;
  assign n22456 = ~n21021 & ~n22447;
  assign n22457 = ~n22455 & n22456;
  assign n22458 = pi0299 & ~n22457;
  assign n22459 = ~pi0746 & ~n22444;
  assign n22460 = ~n22458 & n22459;
  assign n22461 = n21026 & ~n22451;
  assign n22462 = ~n21103 & n22461;
  assign n22463 = ~pi0215 & ~n22462;
  assign n22464 = n22450 & n22463;
  assign n22465 = ~n22446 & ~n22464;
  assign n22466 = pi0299 & ~n22465;
  assign n22467 = pi0169 & ~n21071;
  assign n22468 = n21062 & ~n22467;
  assign n22469 = ~n22466 & ~n22468;
  assign n22470 = pi0746 & ~n22469;
  assign n22471 = pi0039 & ~n22460;
  assign n22472 = ~n22470 & n22471;
  assign n22473 = ~n22442 & ~n22472;
  assign n22474 = ~pi0038 & ~n22473;
  assign n22475 = ~pi0169 & ~n16641;
  assign n22476 = ~pi0746 & pi0947;
  assign n22477 = ~pi0039 & ~n22476;
  assign n22478 = n21239 & n22477;
  assign n22479 = pi0038 & ~n22475;
  assign n22480 = ~n22478 & n22479;
  assign n22481 = ~n22474 & ~n22480;
  assign n22482 = pi0729 & ~n22481;
  assign n22483 = n6284 & n22431;
  assign n22484 = pi0169 & ~n17050;
  assign n22485 = pi0038 & ~n22483;
  assign n22486 = ~n22484 & n22485;
  assign n22487 = n21019 & ~n22443;
  assign n22488 = n21000 & ~n22445;
  assign n22489 = n22450 & ~n22461;
  assign n22490 = n20996 & n22489;
  assign n22491 = pi0299 & ~n22488;
  assign n22492 = ~n22490 & n22491;
  assign n22493 = pi0746 & ~n22492;
  assign n22494 = ~n22487 & n22493;
  assign n22495 = ~pi0169 & ~pi0746;
  assign n22496 = ~n17046 & n22495;
  assign n22497 = pi0039 & ~n22496;
  assign n22498 = ~n22494 & n22497;
  assign n22499 = ~pi0038 & ~n22441;
  assign n22500 = ~n22498 & n22499;
  assign n22501 = ~pi0729 & ~n22486;
  assign n22502 = ~n22500 & n22501;
  assign n22503 = n21130 & ~n22502;
  assign n22504 = ~n22482 & n22503;
  assign n22505 = ~pi0057 & ~n22437;
  assign n22506 = ~n22504 & n22505;
  assign n22507 = ~pi0832 & ~n22436;
  assign n22508 = ~n22506 & n22507;
  assign po0326 = n22435 | n22508;
  assign n22510 = pi0730 & n20902;
  assign n22511 = pi0748 & pi0947;
  assign n22512 = n2926 & ~n22511;
  assign n22513 = ~n22510 & n22512;
  assign n22514 = pi0170 & ~n2926;
  assign n22515 = pi0832 & ~n22514;
  assign n22516 = ~n22513 & n22515;
  assign n22517 = pi0057 & pi0170;
  assign n22518 = ~pi0170 & ~n21130;
  assign n22519 = ~pi0170 & ~n16641;
  assign n22520 = n21090 & ~n22519;
  assign n22521 = pi0170 & ~n17037;
  assign n22522 = n20998 & ~n22521;
  assign n22523 = n21073 & ~n22522;
  assign n22524 = pi0170 & ~n3448;
  assign n22525 = ~n17032 & n22524;
  assign n22526 = ~n17031 & ~n22525;
  assign n22527 = ~pi0170 & ~n16653;
  assign n22528 = n21105 & ~n22527;
  assign n22529 = ~n21047 & ~n22528;
  assign n22530 = n22526 & n22529;
  assign n22531 = ~pi0215 & ~n22530;
  assign n22532 = ~n21021 & ~n22523;
  assign n22533 = ~n22531 & n22532;
  assign n22534 = pi0299 & ~n22533;
  assign n22535 = ~pi0170 & ~n17024;
  assign n22536 = ~pi0299 & ~n22535;
  assign n22537 = ~n21110 & n22536;
  assign n22538 = ~n22534 & ~n22537;
  assign n22539 = pi0039 & ~n22538;
  assign n22540 = ~pi0170 & ~n16958;
  assign n22541 = n21115 & ~n22540;
  assign n22542 = ~n22539 & ~n22541;
  assign n22543 = ~pi0038 & ~n22542;
  assign n22544 = ~pi0748 & ~n22520;
  assign n22545 = ~n22543 & n22544;
  assign n22546 = n21042 & ~n22519;
  assign n22547 = n21067 & ~n22540;
  assign n22548 = n21026 & ~n22527;
  assign n22549 = ~n21103 & n22548;
  assign n22550 = ~pi0215 & ~n22549;
  assign n22551 = n22526 & n22550;
  assign n22552 = ~n22522 & ~n22551;
  assign n22553 = pi0299 & ~n22552;
  assign n22554 = pi0170 & ~n21071;
  assign n22555 = n21062 & ~n22554;
  assign n22556 = pi0039 & ~n22553;
  assign n22557 = ~n22555 & n22556;
  assign n22558 = ~n22547 & ~n22557;
  assign n22559 = ~pi0038 & ~n22558;
  assign n22560 = pi0748 & ~n22546;
  assign n22561 = ~n22559 & n22560;
  assign n22562 = pi0730 & ~n22561;
  assign n22563 = ~n22545 & n22562;
  assign n22564 = ~pi0170 & ~n17050;
  assign n22565 = ~n21015 & ~n22564;
  assign n22566 = n21017 & ~n22540;
  assign n22567 = n21000 & ~n22521;
  assign n22568 = n22526 & ~n22548;
  assign n22569 = n20996 & n22568;
  assign n22570 = pi0299 & ~n22567;
  assign n22571 = ~n22569 & n22570;
  assign n22572 = ~n21018 & n22536;
  assign n22573 = ~n22571 & ~n22572;
  assign n22574 = pi0039 & ~n22573;
  assign n22575 = ~n22566 & ~n22574;
  assign n22576 = ~pi0038 & ~n22575;
  assign n22577 = pi0748 & ~n22565;
  assign n22578 = ~n22576 & n22577;
  assign n22579 = ~pi0170 & ~pi0748;
  assign n22580 = ~n17052 & n22579;
  assign n22581 = ~pi0730 & ~n22580;
  assign n22582 = ~n22578 & n22581;
  assign n22583 = n21130 & ~n22582;
  assign n22584 = ~n22563 & n22583;
  assign n22585 = ~pi0057 & ~n22518;
  assign n22586 = ~n22584 & n22585;
  assign n22587 = ~pi0832 & ~n22517;
  assign n22588 = ~n22586 & n22587;
  assign po0327 = n22516 | n22588;
  assign n22590 = pi0171 & ~n2926;
  assign n22591 = pi0764 & pi0947;
  assign n22592 = n2926 & ~n22591;
  assign n22593 = pi0691 & n20902;
  assign n22594 = n22592 & ~n22593;
  assign n22595 = pi0832 & ~n22590;
  assign n22596 = ~n22594 & n22595;
  assign n22597 = pi0057 & pi0171;
  assign n22598 = ~pi0171 & ~n21130;
  assign n22599 = ~pi0171 & ~n16958;
  assign n22600 = ~pi0764 & n18147;
  assign n22601 = ~n21017 & ~n22600;
  assign n22602 = ~n22599 & ~n22601;
  assign n22603 = ~n21114 & n22602;
  assign n22604 = ~pi0171 & ~n17024;
  assign n22605 = n21111 & ~n22604;
  assign n22606 = pi0171 & ~n17037;
  assign n22607 = n20998 & ~n22606;
  assign n22608 = n21073 & ~n22607;
  assign n22609 = pi0171 & ~n3448;
  assign n22610 = ~n17032 & n22609;
  assign n22611 = ~n17031 & ~n22610;
  assign n22612 = ~pi0171 & ~n16653;
  assign n22613 = n21105 & ~n22612;
  assign n22614 = ~n21047 & ~n22613;
  assign n22615 = n22611 & n22614;
  assign n22616 = ~pi0215 & ~n22615;
  assign n22617 = ~n21021 & ~n22608;
  assign n22618 = ~n22616 & n22617;
  assign n22619 = pi0299 & ~n22618;
  assign n22620 = ~pi0764 & ~n22605;
  assign n22621 = ~n22619 & n22620;
  assign n22622 = n21026 & ~n22612;
  assign n22623 = ~n21103 & n22622;
  assign n22624 = ~pi0215 & ~n22623;
  assign n22625 = n22611 & n22624;
  assign n22626 = ~n22607 & ~n22625;
  assign n22627 = pi0299 & ~n22626;
  assign n22628 = pi0171 & ~n21071;
  assign n22629 = n21062 & ~n22628;
  assign n22630 = ~n22627 & ~n22629;
  assign n22631 = pi0764 & ~n22630;
  assign n22632 = pi0039 & ~n22621;
  assign n22633 = ~n22631 & n22632;
  assign n22634 = ~n22603 & ~n22633;
  assign n22635 = ~pi0038 & ~n22634;
  assign n22636 = ~pi0171 & ~n16641;
  assign n22637 = ~pi0764 & pi0947;
  assign n22638 = ~pi0039 & ~n22637;
  assign n22639 = n21239 & n22638;
  assign n22640 = pi0038 & ~n22636;
  assign n22641 = ~n22639 & n22640;
  assign n22642 = ~n22635 & ~n22641;
  assign n22643 = pi0691 & ~n22642;
  assign n22644 = n6284 & n22592;
  assign n22645 = pi0171 & ~n17050;
  assign n22646 = pi0038 & ~n22644;
  assign n22647 = ~n22645 & n22646;
  assign n22648 = n21019 & ~n22604;
  assign n22649 = n21000 & ~n22606;
  assign n22650 = n22611 & ~n22622;
  assign n22651 = n20996 & n22650;
  assign n22652 = pi0299 & ~n22649;
  assign n22653 = ~n22651 & n22652;
  assign n22654 = pi0764 & ~n22653;
  assign n22655 = ~n22648 & n22654;
  assign n22656 = ~pi0171 & ~pi0764;
  assign n22657 = ~n17046 & n22656;
  assign n22658 = pi0039 & ~n22657;
  assign n22659 = ~n22655 & n22658;
  assign n22660 = ~pi0038 & ~n22602;
  assign n22661 = ~n22659 & n22660;
  assign n22662 = ~pi0691 & ~n22647;
  assign n22663 = ~n22661 & n22662;
  assign n22664 = n21130 & ~n22663;
  assign n22665 = ~n22643 & n22664;
  assign n22666 = ~pi0057 & ~n22598;
  assign n22667 = ~n22665 & n22666;
  assign n22668 = ~pi0832 & ~n22597;
  assign n22669 = ~n22667 & n22668;
  assign po0328 = n22596 | n22669;
  assign n22671 = pi0172 & ~n2926;
  assign n22672 = pi0739 & pi0947;
  assign n22673 = n2926 & ~n22672;
  assign n22674 = pi0690 & n20902;
  assign n22675 = n22673 & ~n22674;
  assign n22676 = pi0832 & ~n22671;
  assign n22677 = ~n22675 & n22676;
  assign n22678 = pi0057 & pi0172;
  assign n22679 = ~pi0172 & ~n21130;
  assign n22680 = ~pi0172 & ~n16958;
  assign n22681 = n16958 & n22672;
  assign n22682 = ~pi0039 & ~n22680;
  assign n22683 = ~n22681 & n22682;
  assign n22684 = ~n21114 & n22683;
  assign n22685 = ~pi0172 & ~n17024;
  assign n22686 = n21111 & ~n22685;
  assign n22687 = pi0172 & ~n17037;
  assign n22688 = n20998 & ~n22687;
  assign n22689 = n21073 & ~n22688;
  assign n22690 = pi0172 & ~n3448;
  assign n22691 = ~n17032 & n22690;
  assign n22692 = ~n17031 & ~n22691;
  assign n22693 = ~pi0172 & ~n16653;
  assign n22694 = n21105 & ~n22693;
  assign n22695 = ~n21047 & ~n22694;
  assign n22696 = n22692 & n22695;
  assign n22697 = ~pi0215 & ~n22696;
  assign n22698 = ~n21021 & ~n22689;
  assign n22699 = ~n22697 & n22698;
  assign n22700 = pi0299 & ~n22699;
  assign n22701 = ~pi0739 & ~n22686;
  assign n22702 = ~n22700 & n22701;
  assign n22703 = n21026 & ~n22693;
  assign n22704 = ~n21103 & n22703;
  assign n22705 = ~pi0215 & ~n22704;
  assign n22706 = n22692 & n22705;
  assign n22707 = ~n22688 & ~n22706;
  assign n22708 = pi0299 & ~n22707;
  assign n22709 = pi0172 & ~n21071;
  assign n22710 = n21062 & ~n22709;
  assign n22711 = ~n22708 & ~n22710;
  assign n22712 = pi0739 & ~n22711;
  assign n22713 = pi0039 & ~n22702;
  assign n22714 = ~n22712 & n22713;
  assign n22715 = ~n22684 & ~n22714;
  assign n22716 = ~pi0038 & ~n22715;
  assign n22717 = ~pi0172 & ~n16641;
  assign n22718 = ~pi0739 & pi0947;
  assign n22719 = ~pi0039 & ~n22718;
  assign n22720 = n21239 & n22719;
  assign n22721 = pi0038 & ~n22717;
  assign n22722 = ~n22720 & n22721;
  assign n22723 = ~n22716 & ~n22722;
  assign n22724 = pi0690 & ~n22723;
  assign n22725 = n6284 & n22673;
  assign n22726 = pi0172 & ~n17050;
  assign n22727 = pi0038 & ~n22725;
  assign n22728 = ~n22726 & n22727;
  assign n22729 = n21019 & ~n22685;
  assign n22730 = n21000 & ~n22687;
  assign n22731 = n22692 & ~n22703;
  assign n22732 = n20996 & n22731;
  assign n22733 = pi0299 & ~n22730;
  assign n22734 = ~n22732 & n22733;
  assign n22735 = pi0739 & ~n22734;
  assign n22736 = ~n22729 & n22735;
  assign n22737 = ~pi0172 & ~pi0739;
  assign n22738 = ~n17046 & n22737;
  assign n22739 = pi0039 & ~n22738;
  assign n22740 = ~n22736 & n22739;
  assign n22741 = ~pi0038 & ~n22683;
  assign n22742 = ~n22740 & n22741;
  assign n22743 = ~pi0690 & ~n22728;
  assign n22744 = ~n22742 & n22743;
  assign n22745 = n21130 & ~n22744;
  assign n22746 = ~n22724 & n22745;
  assign n22747 = ~pi0057 & ~n22679;
  assign n22748 = ~n22746 & n22747;
  assign n22749 = ~pi0832 & ~n22678;
  assign n22750 = ~n22748 & n22749;
  assign po0329 = n22677 | n22750;
  assign n22752 = ~pi0173 & po1038;
  assign n22753 = ~pi0173 & ~n17059;
  assign n22754 = n16635 & ~n22753;
  assign n22755 = ~pi0723 & n2571;
  assign n22756 = n22753 & ~n22755;
  assign n22757 = ~pi0173 & ~n16641;
  assign n22758 = n16647 & ~n22757;
  assign n22759 = pi0173 & ~n18076;
  assign n22760 = ~pi0038 & ~n22759;
  assign n22761 = n2571 & ~n22760;
  assign n22762 = ~pi0173 & n18072;
  assign n22763 = ~n22761 & ~n22762;
  assign n22764 = ~pi0723 & ~n22758;
  assign n22765 = ~n22763 & n22764;
  assign n22766 = ~n22756 & ~n22765;
  assign n22767 = ~pi0778 & n22766;
  assign n22768 = ~pi0625 & n22753;
  assign n22769 = pi0625 & ~n22766;
  assign n22770 = pi1153 & ~n22768;
  assign n22771 = ~n22769 & n22770;
  assign n22772 = pi0625 & n22753;
  assign n22773 = ~pi0625 & ~n22766;
  assign n22774 = ~pi1153 & ~n22772;
  assign n22775 = ~n22773 & n22774;
  assign n22776 = ~n22771 & ~n22775;
  assign n22777 = pi0778 & ~n22776;
  assign n22778 = ~n22767 & ~n22777;
  assign n22779 = ~n17075 & ~n22778;
  assign n22780 = n17075 & ~n22753;
  assign n22781 = ~n22779 & ~n22780;
  assign n22782 = ~n16639 & n22781;
  assign n22783 = n16639 & n22753;
  assign n22784 = ~n22782 & ~n22783;
  assign n22785 = ~n16635 & n22784;
  assign n22786 = ~n22754 & ~n22785;
  assign n22787 = ~n16631 & n22786;
  assign n22788 = n16631 & n22753;
  assign n22789 = ~n22787 & ~n22788;
  assign n22790 = ~pi0792 & n22789;
  assign n22791 = pi0628 & ~n22789;
  assign n22792 = ~pi0628 & n22753;
  assign n22793 = pi1156 & ~n22792;
  assign n22794 = ~n22791 & n22793;
  assign n22795 = pi0628 & n22753;
  assign n22796 = ~pi0628 & ~n22789;
  assign n22797 = ~pi1156 & ~n22795;
  assign n22798 = ~n22796 & n22797;
  assign n22799 = ~n22794 & ~n22798;
  assign n22800 = pi0792 & ~n22799;
  assign n22801 = ~n22790 & ~n22800;
  assign n22802 = ~pi0647 & ~n22801;
  assign n22803 = pi0647 & ~n22753;
  assign n22804 = ~n22802 & ~n22803;
  assign n22805 = ~pi1157 & n22804;
  assign n22806 = pi0647 & ~n22801;
  assign n22807 = ~pi0647 & ~n22753;
  assign n22808 = ~n22806 & ~n22807;
  assign n22809 = pi1157 & n22808;
  assign n22810 = ~n22805 & ~n22809;
  assign n22811 = pi0787 & ~n22810;
  assign n22812 = ~pi0787 & n22801;
  assign n22813 = ~n22811 & ~n22812;
  assign n22814 = ~pi0644 & ~n22813;
  assign n22815 = pi0715 & ~n22814;
  assign n22816 = pi0173 & ~n2571;
  assign n22817 = pi0173 & ~n17275;
  assign n22818 = ~pi0173 & ~n17048;
  assign n22819 = pi0745 & ~n22818;
  assign n22820 = ~pi0173 & ~pi0745;
  assign n22821 = n17221 & n22820;
  assign n22822 = ~n22817 & ~n22821;
  assign n22823 = ~n22819 & n22822;
  assign n22824 = ~pi0038 & ~n22823;
  assign n22825 = ~pi0745 & n17280;
  assign n22826 = pi0038 & ~n22757;
  assign n22827 = ~n22825 & n22826;
  assign n22828 = ~n22824 & ~n22827;
  assign n22829 = n2571 & ~n22828;
  assign n22830 = ~n22816 & ~n22829;
  assign n22831 = ~n17117 & ~n22830;
  assign n22832 = n17117 & ~n22753;
  assign n22833 = ~n22831 & ~n22832;
  assign n22834 = ~pi0785 & ~n22833;
  assign n22835 = ~n17291 & ~n22753;
  assign n22836 = pi0609 & n22831;
  assign n22837 = ~n22835 & ~n22836;
  assign n22838 = pi1155 & ~n22837;
  assign n22839 = ~n17296 & ~n22753;
  assign n22840 = ~pi0609 & n22831;
  assign n22841 = ~n22839 & ~n22840;
  assign n22842 = ~pi1155 & ~n22841;
  assign n22843 = ~n22838 & ~n22842;
  assign n22844 = pi0785 & ~n22843;
  assign n22845 = ~n22834 & ~n22844;
  assign n22846 = ~pi0781 & ~n22845;
  assign n22847 = ~pi0618 & n22753;
  assign n22848 = pi0618 & n22845;
  assign n22849 = pi1154 & ~n22847;
  assign n22850 = ~n22848 & n22849;
  assign n22851 = ~pi0618 & n22845;
  assign n22852 = pi0618 & n22753;
  assign n22853 = ~pi1154 & ~n22852;
  assign n22854 = ~n22851 & n22853;
  assign n22855 = ~n22850 & ~n22854;
  assign n22856 = pi0781 & ~n22855;
  assign n22857 = ~n22846 & ~n22856;
  assign n22858 = ~pi0789 & ~n22857;
  assign n22859 = ~pi0619 & n22753;
  assign n22860 = pi0619 & n22857;
  assign n22861 = pi1159 & ~n22859;
  assign n22862 = ~n22860 & n22861;
  assign n22863 = ~pi0619 & n22857;
  assign n22864 = pi0619 & n22753;
  assign n22865 = ~pi1159 & ~n22864;
  assign n22866 = ~n22863 & n22865;
  assign n22867 = ~n22862 & ~n22866;
  assign n22868 = pi0789 & ~n22867;
  assign n22869 = ~n22858 & ~n22868;
  assign n22870 = ~pi0788 & ~n22869;
  assign n22871 = ~pi0626 & n22753;
  assign n22872 = pi0626 & n22869;
  assign n22873 = pi1158 & ~n22871;
  assign n22874 = ~n22872 & n22873;
  assign n22875 = ~pi0626 & n22869;
  assign n22876 = pi0626 & n22753;
  assign n22877 = ~pi1158 & ~n22876;
  assign n22878 = ~n22875 & n22877;
  assign n22879 = ~n22874 & ~n22878;
  assign n22880 = pi0788 & ~n22879;
  assign n22881 = ~n22870 & ~n22880;
  assign n22882 = ~n17779 & n22881;
  assign n22883 = n17779 & n22753;
  assign n22884 = ~n22882 & ~n22883;
  assign n22885 = ~n17804 & ~n22884;
  assign n22886 = n17804 & n22753;
  assign n22887 = ~n22885 & ~n22886;
  assign n22888 = pi0644 & ~n22887;
  assign n22889 = ~pi0644 & n22753;
  assign n22890 = ~pi0715 & ~n22889;
  assign n22891 = ~n22888 & n22890;
  assign n22892 = pi1160 & ~n22891;
  assign n22893 = ~n22815 & n22892;
  assign n22894 = pi0644 & ~n22813;
  assign n22895 = n17802 & ~n22804;
  assign n22896 = ~n20559 & n22884;
  assign n22897 = n17801 & ~n22808;
  assign n22898 = ~n22895 & ~n22897;
  assign n22899 = ~n22896 & n22898;
  assign n22900 = pi0787 & ~n22899;
  assign n22901 = ~pi0629 & n22794;
  assign n22902 = ~n20570 & ~n22881;
  assign n22903 = pi0629 & n22798;
  assign n22904 = ~n22901 & ~n22903;
  assign n22905 = ~n22902 & n22904;
  assign n22906 = pi0792 & ~n22905;
  assign n22907 = pi0609 & n22778;
  assign n22908 = pi0173 & ~n17625;
  assign n22909 = ~pi0173 & ~n17612;
  assign n22910 = pi0745 & ~n22908;
  assign n22911 = ~n22909 & n22910;
  assign n22912 = ~pi0173 & n17629;
  assign n22913 = pi0173 & n17631;
  assign n22914 = ~pi0745 & ~n22913;
  assign n22915 = ~n22912 & n22914;
  assign n22916 = ~n22911 & ~n22915;
  assign n22917 = ~pi0039 & ~n22916;
  assign n22918 = pi0173 & n17605;
  assign n22919 = ~pi0173 & ~n17546;
  assign n22920 = ~pi0745 & ~n22919;
  assign n22921 = ~n22918 & n22920;
  assign n22922 = ~pi0173 & n17404;
  assign n22923 = pi0173 & n17485;
  assign n22924 = pi0745 & ~n22923;
  assign n22925 = ~n22922 & n22924;
  assign n22926 = pi0039 & ~n22921;
  assign n22927 = ~n22925 & n22926;
  assign n22928 = ~pi0038 & ~n22917;
  assign n22929 = ~n22927 & n22928;
  assign n22930 = ~pi0745 & ~n17490;
  assign n22931 = n19471 & ~n22930;
  assign n22932 = ~pi0173 & ~n22931;
  assign n22933 = ~pi0745 & n17244;
  assign n22934 = ~n17469 & ~n22933;
  assign n22935 = pi0173 & ~n22934;
  assign n22936 = n6284 & n22935;
  assign n22937 = pi0038 & ~n22936;
  assign n22938 = ~n22932 & n22937;
  assign n22939 = ~pi0723 & ~n22938;
  assign n22940 = ~n22929 & n22939;
  assign n22941 = pi0723 & n22828;
  assign n22942 = n2571 & ~n22940;
  assign n22943 = ~n22941 & n22942;
  assign n22944 = ~n22816 & ~n22943;
  assign n22945 = ~pi0625 & n22944;
  assign n22946 = pi0625 & n22830;
  assign n22947 = ~pi1153 & ~n22946;
  assign n22948 = ~n22945 & n22947;
  assign n22949 = ~pi0608 & ~n22771;
  assign n22950 = ~n22948 & n22949;
  assign n22951 = ~pi0625 & n22830;
  assign n22952 = pi0625 & n22944;
  assign n22953 = pi1153 & ~n22951;
  assign n22954 = ~n22952 & n22953;
  assign n22955 = pi0608 & ~n22775;
  assign n22956 = ~n22954 & n22955;
  assign n22957 = ~n22950 & ~n22956;
  assign n22958 = pi0778 & ~n22957;
  assign n22959 = ~pi0778 & n22944;
  assign n22960 = ~n22958 & ~n22959;
  assign n22961 = ~pi0609 & ~n22960;
  assign n22962 = ~pi1155 & ~n22907;
  assign n22963 = ~n22961 & n22962;
  assign n22964 = ~pi0660 & ~n22838;
  assign n22965 = ~n22963 & n22964;
  assign n22966 = ~pi0609 & n22778;
  assign n22967 = pi0609 & ~n22960;
  assign n22968 = pi1155 & ~n22966;
  assign n22969 = ~n22967 & n22968;
  assign n22970 = pi0660 & ~n22842;
  assign n22971 = ~n22969 & n22970;
  assign n22972 = ~n22965 & ~n22971;
  assign n22973 = pi0785 & ~n22972;
  assign n22974 = ~pi0785 & ~n22960;
  assign n22975 = ~n22973 & ~n22974;
  assign n22976 = ~pi0618 & ~n22975;
  assign n22977 = pi0618 & n22781;
  assign n22978 = ~pi1154 & ~n22977;
  assign n22979 = ~n22976 & n22978;
  assign n22980 = ~pi0627 & ~n22850;
  assign n22981 = ~n22979 & n22980;
  assign n22982 = ~pi0618 & n22781;
  assign n22983 = pi0618 & ~n22975;
  assign n22984 = pi1154 & ~n22982;
  assign n22985 = ~n22983 & n22984;
  assign n22986 = pi0627 & ~n22854;
  assign n22987 = ~n22985 & n22986;
  assign n22988 = ~n22981 & ~n22987;
  assign n22989 = pi0781 & ~n22988;
  assign n22990 = ~pi0781 & ~n22975;
  assign n22991 = ~n22989 & ~n22990;
  assign n22992 = ~pi0789 & n22991;
  assign n22993 = pi0619 & ~n22784;
  assign n22994 = ~pi0619 & ~n22991;
  assign n22995 = ~pi1159 & ~n22993;
  assign n22996 = ~n22994 & n22995;
  assign n22997 = ~pi0648 & ~n22862;
  assign n22998 = ~n22996 & n22997;
  assign n22999 = pi0619 & ~n22991;
  assign n23000 = ~pi0619 & ~n22784;
  assign n23001 = pi1159 & ~n23000;
  assign n23002 = ~n22999 & n23001;
  assign n23003 = pi0648 & ~n22866;
  assign n23004 = ~n23002 & n23003;
  assign n23005 = pi0789 & ~n22998;
  assign n23006 = ~n23004 & n23005;
  assign n23007 = n17970 & ~n22992;
  assign n23008 = ~n23006 & n23007;
  assign n23009 = n17871 & n22786;
  assign n23010 = ~n16630 & n22879;
  assign n23011 = ~n23009 & ~n23010;
  assign n23012 = pi0788 & ~n23011;
  assign n23013 = ~n20364 & ~n23012;
  assign n23014 = ~n23008 & n23013;
  assign n23015 = ~n22906 & ~n23014;
  assign n23016 = ~n20206 & ~n23015;
  assign n23017 = ~n22900 & ~n23016;
  assign n23018 = ~pi0644 & n23017;
  assign n23019 = ~pi0715 & ~n22894;
  assign n23020 = ~n23018 & n23019;
  assign n23021 = pi0644 & n22753;
  assign n23022 = ~pi0644 & ~n22887;
  assign n23023 = pi0715 & ~n23021;
  assign n23024 = ~n23022 & n23023;
  assign n23025 = ~pi1160 & ~n23024;
  assign n23026 = ~n23020 & n23025;
  assign n23027 = ~n22893 & ~n23026;
  assign n23028 = pi0790 & ~n23027;
  assign n23029 = pi0644 & n22892;
  assign n23030 = pi0790 & ~n23029;
  assign n23031 = n23017 & ~n23030;
  assign n23032 = ~n23028 & ~n23031;
  assign n23033 = ~po1038 & ~n23032;
  assign n23034 = ~pi0832 & ~n22752;
  assign n23035 = ~n23033 & n23034;
  assign n23036 = ~pi0173 & ~n2926;
  assign n23037 = ~pi0723 & n16645;
  assign n23038 = ~n23036 & ~n23037;
  assign n23039 = ~pi0778 & ~n23038;
  assign n23040 = ~pi0625 & n23037;
  assign n23041 = ~n23038 & ~n23040;
  assign n23042 = pi1153 & ~n23041;
  assign n23043 = ~pi1153 & ~n23036;
  assign n23044 = ~n23040 & n23043;
  assign n23045 = pi0778 & ~n23044;
  assign n23046 = ~n23042 & n23045;
  assign n23047 = ~n23039 & ~n23046;
  assign n23048 = ~n17845 & ~n23047;
  assign n23049 = ~n17847 & n23048;
  assign n23050 = ~n17849 & n23049;
  assign n23051 = ~n17851 & n23050;
  assign n23052 = ~n17857 & n23051;
  assign n23053 = ~pi0647 & n23052;
  assign n23054 = pi0647 & n23036;
  assign n23055 = ~pi1157 & ~n23054;
  assign n23056 = ~n23053 & n23055;
  assign n23057 = pi0630 & n23056;
  assign n23058 = ~n22933 & ~n23036;
  assign n23059 = ~n17874 & ~n23058;
  assign n23060 = ~pi0785 & ~n23059;
  assign n23061 = n17296 & n22933;
  assign n23062 = n23059 & ~n23061;
  assign n23063 = pi1155 & ~n23062;
  assign n23064 = ~pi1155 & ~n23036;
  assign n23065 = ~n23061 & n23064;
  assign n23066 = ~n23063 & ~n23065;
  assign n23067 = pi0785 & ~n23066;
  assign n23068 = ~n23060 & ~n23067;
  assign n23069 = ~pi0781 & ~n23068;
  assign n23070 = ~n17889 & n23068;
  assign n23071 = pi1154 & ~n23070;
  assign n23072 = ~n17892 & n23068;
  assign n23073 = ~pi1154 & ~n23072;
  assign n23074 = ~n23071 & ~n23073;
  assign n23075 = pi0781 & ~n23074;
  assign n23076 = ~n23069 & ~n23075;
  assign n23077 = ~pi0789 & ~n23076;
  assign n23078 = ~pi0619 & n2926;
  assign n23079 = n23076 & ~n23078;
  assign n23080 = pi1159 & ~n23079;
  assign n23081 = pi0619 & n2926;
  assign n23082 = n23076 & ~n23081;
  assign n23083 = ~pi1159 & ~n23082;
  assign n23084 = ~n23080 & ~n23083;
  assign n23085 = pi0789 & ~n23084;
  assign n23086 = ~n23077 & ~n23085;
  assign n23087 = ~pi0788 & ~n23086;
  assign n23088 = ~pi0626 & n23036;
  assign n23089 = pi0626 & n23086;
  assign n23090 = pi1158 & ~n23088;
  assign n23091 = ~n23089 & n23090;
  assign n23092 = ~pi0626 & n23086;
  assign n23093 = pi0626 & n23036;
  assign n23094 = ~pi1158 & ~n23093;
  assign n23095 = ~n23092 & n23094;
  assign n23096 = ~n23091 & ~n23095;
  assign n23097 = pi0788 & ~n23096;
  assign n23098 = ~n23087 & ~n23097;
  assign n23099 = ~n17779 & n23098;
  assign n23100 = n17779 & n23036;
  assign n23101 = ~n23099 & ~n23100;
  assign n23102 = ~n20559 & n23101;
  assign n23103 = pi0647 & ~n23052;
  assign n23104 = ~pi0647 & ~n23036;
  assign n23105 = ~n23103 & ~n23104;
  assign n23106 = n17801 & ~n23105;
  assign n23107 = ~n23057 & ~n23106;
  assign n23108 = ~n23102 & n23107;
  assign n23109 = pi0787 & ~n23108;
  assign n23110 = n17871 & n23050;
  assign n23111 = ~n16630 & n23096;
  assign n23112 = ~n23110 & ~n23111;
  assign n23113 = pi0788 & ~n23112;
  assign n23114 = pi0618 & n23048;
  assign n23115 = ~n17168 & ~n23038;
  assign n23116 = pi0625 & n23115;
  assign n23117 = n23058 & ~n23115;
  assign n23118 = ~n23116 & ~n23117;
  assign n23119 = n23043 & ~n23118;
  assign n23120 = ~pi0608 & ~n23042;
  assign n23121 = ~n23119 & n23120;
  assign n23122 = pi1153 & n23058;
  assign n23123 = ~n23116 & n23122;
  assign n23124 = pi0608 & ~n23044;
  assign n23125 = ~n23123 & n23124;
  assign n23126 = ~n23121 & ~n23125;
  assign n23127 = pi0778 & ~n23126;
  assign n23128 = ~pi0778 & ~n23117;
  assign n23129 = ~n23127 & ~n23128;
  assign n23130 = ~pi0609 & ~n23129;
  assign n23131 = pi0609 & ~n23047;
  assign n23132 = ~pi1155 & ~n23131;
  assign n23133 = ~n23130 & n23132;
  assign n23134 = ~pi0660 & ~n23063;
  assign n23135 = ~n23133 & n23134;
  assign n23136 = pi0609 & ~n23129;
  assign n23137 = ~pi0609 & ~n23047;
  assign n23138 = pi1155 & ~n23137;
  assign n23139 = ~n23136 & n23138;
  assign n23140 = pi0660 & ~n23065;
  assign n23141 = ~n23139 & n23140;
  assign n23142 = ~n23135 & ~n23141;
  assign n23143 = pi0785 & ~n23142;
  assign n23144 = ~pi0785 & ~n23129;
  assign n23145 = ~n23143 & ~n23144;
  assign n23146 = ~pi0618 & ~n23145;
  assign n23147 = ~pi1154 & ~n23114;
  assign n23148 = ~n23146 & n23147;
  assign n23149 = ~pi0627 & ~n23071;
  assign n23150 = ~n23148 & n23149;
  assign n23151 = ~pi0618 & n23048;
  assign n23152 = pi0618 & ~n23145;
  assign n23153 = pi1154 & ~n23151;
  assign n23154 = ~n23152 & n23153;
  assign n23155 = pi0627 & ~n23073;
  assign n23156 = ~n23154 & n23155;
  assign n23157 = ~n23150 & ~n23156;
  assign n23158 = pi0781 & ~n23157;
  assign n23159 = ~pi0781 & ~n23145;
  assign n23160 = ~n23158 & ~n23159;
  assign n23161 = ~pi0789 & n23160;
  assign n23162 = ~pi0619 & ~n23160;
  assign n23163 = pi0619 & n23049;
  assign n23164 = ~pi1159 & ~n23163;
  assign n23165 = ~n23162 & n23164;
  assign n23166 = ~pi0648 & ~n23080;
  assign n23167 = ~n23165 & n23166;
  assign n23168 = ~pi0619 & n23049;
  assign n23169 = pi0619 & ~n23160;
  assign n23170 = pi1159 & ~n23168;
  assign n23171 = ~n23169 & n23170;
  assign n23172 = pi0648 & ~n23083;
  assign n23173 = ~n23171 & n23172;
  assign n23174 = pi0789 & ~n23167;
  assign n23175 = ~n23173 & n23174;
  assign n23176 = n17970 & ~n23161;
  assign n23177 = ~n23175 & n23176;
  assign n23178 = ~n23113 & ~n23177;
  assign n23179 = ~n20364 & ~n23178;
  assign n23180 = n17854 & n23098;
  assign n23181 = n20851 & n23051;
  assign n23182 = ~n23180 & ~n23181;
  assign n23183 = ~pi0629 & ~n23182;
  assign n23184 = n20855 & n23051;
  assign n23185 = n17853 & n23098;
  assign n23186 = ~n23184 & ~n23185;
  assign n23187 = pi0629 & ~n23186;
  assign n23188 = ~n23183 & ~n23187;
  assign n23189 = pi0792 & ~n23188;
  assign n23190 = ~n20206 & ~n23189;
  assign n23191 = ~n23179 & n23190;
  assign n23192 = ~n23109 & ~n23191;
  assign n23193 = ~pi0790 & n23192;
  assign n23194 = ~pi0787 & ~n23052;
  assign n23195 = pi1157 & ~n23105;
  assign n23196 = ~n23056 & ~n23195;
  assign n23197 = pi0787 & ~n23196;
  assign n23198 = ~n23194 & ~n23197;
  assign n23199 = ~pi0644 & n23198;
  assign n23200 = pi0644 & n23192;
  assign n23201 = pi0715 & ~n23199;
  assign n23202 = ~n23200 & n23201;
  assign n23203 = ~n17804 & ~n23101;
  assign n23204 = n17804 & n23036;
  assign n23205 = ~n23203 & ~n23204;
  assign n23206 = pi0644 & ~n23205;
  assign n23207 = ~pi0644 & n23036;
  assign n23208 = ~pi0715 & ~n23207;
  assign n23209 = ~n23206 & n23208;
  assign n23210 = pi1160 & ~n23209;
  assign n23211 = ~n23202 & n23210;
  assign n23212 = ~pi0644 & ~n23205;
  assign n23213 = pi0644 & n23036;
  assign n23214 = pi0715 & ~n23213;
  assign n23215 = ~n23212 & n23214;
  assign n23216 = pi0644 & n23198;
  assign n23217 = ~pi0644 & n23192;
  assign n23218 = ~pi0715 & ~n23216;
  assign n23219 = ~n23217 & n23218;
  assign n23220 = ~pi1160 & ~n23215;
  assign n23221 = ~n23219 & n23220;
  assign n23222 = ~n23211 & ~n23221;
  assign n23223 = pi0790 & ~n23222;
  assign n23224 = pi0832 & ~n23193;
  assign n23225 = ~n23223 & n23224;
  assign po0330 = ~n23035 & ~n23225;
  assign n23227 = pi0174 & ~n17059;
  assign n23228 = n16635 & ~n23227;
  assign n23229 = n17075 & ~n23227;
  assign n23230 = pi0696 & n2571;
  assign n23231 = ~n23227 & ~n23230;
  assign n23232 = ~pi0174 & ~n16641;
  assign n23233 = n19899 & ~n23232;
  assign n23234 = ~pi0174 & n18076;
  assign n23235 = pi0174 & ~n18072;
  assign n23236 = ~pi0038 & ~n23234;
  assign n23237 = ~n23235 & n23236;
  assign n23238 = n23230 & ~n23233;
  assign n23239 = ~n23237 & n23238;
  assign n23240 = ~n23231 & ~n23239;
  assign n23241 = ~pi0778 & n23240;
  assign n23242 = ~pi0625 & ~n23227;
  assign n23243 = pi0625 & ~n23240;
  assign n23244 = pi1153 & ~n23242;
  assign n23245 = ~n23243 & n23244;
  assign n23246 = ~pi0625 & ~n23240;
  assign n23247 = pi0625 & ~n23227;
  assign n23248 = ~pi1153 & ~n23247;
  assign n23249 = ~n23246 & n23248;
  assign n23250 = ~n23245 & ~n23249;
  assign n23251 = pi0778 & ~n23250;
  assign n23252 = ~n23241 & ~n23251;
  assign n23253 = ~n17075 & n23252;
  assign n23254 = ~n23229 & ~n23253;
  assign n23255 = ~n16639 & n23254;
  assign n23256 = n16639 & n23227;
  assign n23257 = ~n23255 & ~n23256;
  assign n23258 = ~n16635 & n23257;
  assign n23259 = ~n23228 & ~n23258;
  assign n23260 = ~n16631 & n23259;
  assign n23261 = n16631 & n23227;
  assign n23262 = ~n23260 & ~n23261;
  assign n23263 = ~pi0792 & ~n23262;
  assign n23264 = ~pi0628 & ~n23227;
  assign n23265 = pi0628 & n23262;
  assign n23266 = pi1156 & ~n23264;
  assign n23267 = ~n23265 & n23266;
  assign n23268 = pi0628 & ~n23227;
  assign n23269 = ~pi0628 & n23262;
  assign n23270 = ~pi1156 & ~n23268;
  assign n23271 = ~n23269 & n23270;
  assign n23272 = ~n23267 & ~n23271;
  assign n23273 = pi0792 & ~n23272;
  assign n23274 = ~n23263 & ~n23273;
  assign n23275 = ~pi0787 & ~n23274;
  assign n23276 = ~pi0647 & ~n23227;
  assign n23277 = pi0647 & n23274;
  assign n23278 = pi1157 & ~n23276;
  assign n23279 = ~n23277 & n23278;
  assign n23280 = pi0647 & ~n23227;
  assign n23281 = ~pi0647 & n23274;
  assign n23282 = ~pi1157 & ~n23280;
  assign n23283 = ~n23281 & n23282;
  assign n23284 = ~n23279 & ~n23283;
  assign n23285 = pi0787 & ~n23284;
  assign n23286 = ~n23275 & ~n23285;
  assign n23287 = ~pi0644 & n23286;
  assign n23288 = ~pi0619 & ~n23227;
  assign n23289 = n17117 & ~n23227;
  assign n23290 = pi0174 & ~n2571;
  assign n23291 = pi0759 & n17219;
  assign n23292 = ~n21470 & ~n23291;
  assign n23293 = pi0039 & ~n23292;
  assign n23294 = ~pi0759 & n16958;
  assign n23295 = pi0759 & n17139;
  assign n23296 = ~pi0039 & ~n23294;
  assign n23297 = ~n23295 & n23296;
  assign n23298 = ~n23293 & ~n23297;
  assign n23299 = pi0174 & ~n23298;
  assign n23300 = ~pi0174 & pi0759;
  assign n23301 = n17275 & n23300;
  assign n23302 = ~n23299 & ~n23301;
  assign n23303 = ~pi0038 & ~n23302;
  assign n23304 = pi0759 & n17168;
  assign n23305 = n16641 & ~n23304;
  assign n23306 = pi0038 & ~n23232;
  assign n23307 = ~n23305 & n23306;
  assign n23308 = ~n23303 & ~n23307;
  assign n23309 = n2571 & ~n23308;
  assign n23310 = ~n23290 & ~n23309;
  assign n23311 = ~n17117 & n23310;
  assign n23312 = ~n23289 & ~n23311;
  assign n23313 = ~pi0785 & n23312;
  assign n23314 = ~pi0609 & ~n23227;
  assign n23315 = pi0609 & ~n23312;
  assign n23316 = pi1155 & ~n23314;
  assign n23317 = ~n23315 & n23316;
  assign n23318 = ~pi0609 & ~n23312;
  assign n23319 = pi0609 & ~n23227;
  assign n23320 = ~pi1155 & ~n23319;
  assign n23321 = ~n23318 & n23320;
  assign n23322 = ~n23317 & ~n23321;
  assign n23323 = pi0785 & ~n23322;
  assign n23324 = ~n23313 & ~n23323;
  assign n23325 = ~pi0781 & ~n23324;
  assign n23326 = ~pi0618 & ~n23227;
  assign n23327 = pi0618 & n23324;
  assign n23328 = pi1154 & ~n23326;
  assign n23329 = ~n23327 & n23328;
  assign n23330 = pi0618 & ~n23227;
  assign n23331 = ~pi0618 & n23324;
  assign n23332 = ~pi1154 & ~n23330;
  assign n23333 = ~n23331 & n23332;
  assign n23334 = ~n23329 & ~n23333;
  assign n23335 = pi0781 & ~n23334;
  assign n23336 = ~n23325 & ~n23335;
  assign n23337 = pi0619 & n23336;
  assign n23338 = pi1159 & ~n23288;
  assign n23339 = ~n23337 & n23338;
  assign n23340 = ~pi0696 & n23308;
  assign n23341 = ~pi0174 & ~n17605;
  assign n23342 = pi0174 & n17546;
  assign n23343 = pi0759 & ~n23342;
  assign n23344 = ~n23341 & n23343;
  assign n23345 = pi0174 & ~n17404;
  assign n23346 = ~pi0174 & ~n17485;
  assign n23347 = ~pi0759 & ~n23346;
  assign n23348 = ~n23345 & n23347;
  assign n23349 = pi0039 & ~n23344;
  assign n23350 = ~n23348 & n23349;
  assign n23351 = ~pi0174 & n17631;
  assign n23352 = pi0174 & n17629;
  assign n23353 = pi0759 & ~n23351;
  assign n23354 = ~n23352 & n23353;
  assign n23355 = ~pi0174 & ~n17625;
  assign n23356 = pi0174 & ~n17612;
  assign n23357 = ~pi0759 & ~n23355;
  assign n23358 = ~n23356 & n23357;
  assign n23359 = ~pi0039 & ~n23354;
  assign n23360 = ~n23358 & n23359;
  assign n23361 = ~pi0038 & ~n23360;
  assign n23362 = ~n23350 & n23361;
  assign n23363 = pi0696 & ~n19470;
  assign n23364 = ~n23307 & n23363;
  assign n23365 = ~n23362 & n23364;
  assign n23366 = n2571 & ~n23365;
  assign n23367 = ~n23340 & n23366;
  assign n23368 = ~n23290 & ~n23367;
  assign n23369 = ~pi0625 & n23368;
  assign n23370 = pi0625 & n23310;
  assign n23371 = ~pi1153 & ~n23370;
  assign n23372 = ~n23369 & n23371;
  assign n23373 = ~pi0608 & ~n23245;
  assign n23374 = ~n23372 & n23373;
  assign n23375 = ~pi0625 & n23310;
  assign n23376 = pi0625 & n23368;
  assign n23377 = pi1153 & ~n23375;
  assign n23378 = ~n23376 & n23377;
  assign n23379 = pi0608 & ~n23249;
  assign n23380 = ~n23378 & n23379;
  assign n23381 = ~n23374 & ~n23380;
  assign n23382 = pi0778 & ~n23381;
  assign n23383 = ~pi0778 & n23368;
  assign n23384 = ~n23382 & ~n23383;
  assign n23385 = ~pi0609 & ~n23384;
  assign n23386 = pi0609 & n23252;
  assign n23387 = ~pi1155 & ~n23386;
  assign n23388 = ~n23385 & n23387;
  assign n23389 = ~pi0660 & ~n23317;
  assign n23390 = ~n23388 & n23389;
  assign n23391 = ~pi0609 & n23252;
  assign n23392 = pi0609 & ~n23384;
  assign n23393 = pi1155 & ~n23391;
  assign n23394 = ~n23392 & n23393;
  assign n23395 = pi0660 & ~n23321;
  assign n23396 = ~n23394 & n23395;
  assign n23397 = ~n23390 & ~n23396;
  assign n23398 = pi0785 & ~n23397;
  assign n23399 = ~pi0785 & ~n23384;
  assign n23400 = ~n23398 & ~n23399;
  assign n23401 = ~pi0618 & ~n23400;
  assign n23402 = pi0618 & ~n23254;
  assign n23403 = ~pi1154 & ~n23402;
  assign n23404 = ~n23401 & n23403;
  assign n23405 = ~pi0627 & ~n23329;
  assign n23406 = ~n23404 & n23405;
  assign n23407 = pi0618 & ~n23400;
  assign n23408 = ~pi0618 & ~n23254;
  assign n23409 = pi1154 & ~n23408;
  assign n23410 = ~n23407 & n23409;
  assign n23411 = pi0627 & ~n23333;
  assign n23412 = ~n23410 & n23411;
  assign n23413 = ~n23406 & ~n23412;
  assign n23414 = pi0781 & ~n23413;
  assign n23415 = ~pi0781 & ~n23400;
  assign n23416 = ~n23414 & ~n23415;
  assign n23417 = ~pi0619 & ~n23416;
  assign n23418 = pi0619 & n23257;
  assign n23419 = ~pi1159 & ~n23418;
  assign n23420 = ~n23417 & n23419;
  assign n23421 = ~pi0648 & ~n23339;
  assign n23422 = ~n23420 & n23421;
  assign n23423 = pi0619 & ~n23227;
  assign n23424 = ~pi0619 & n23336;
  assign n23425 = ~pi1159 & ~n23423;
  assign n23426 = ~n23424 & n23425;
  assign n23427 = ~pi0619 & n23257;
  assign n23428 = pi0619 & ~n23416;
  assign n23429 = pi1159 & ~n23427;
  assign n23430 = ~n23428 & n23429;
  assign n23431 = pi0648 & ~n23426;
  assign n23432 = ~n23430 & n23431;
  assign n23433 = ~n23422 & ~n23432;
  assign n23434 = pi0789 & ~n23433;
  assign n23435 = ~pi0789 & ~n23416;
  assign n23436 = ~n23434 & ~n23435;
  assign n23437 = ~pi0788 & n23436;
  assign n23438 = ~pi0626 & n23436;
  assign n23439 = pi0626 & n23259;
  assign n23440 = ~pi0641 & ~n23439;
  assign n23441 = ~n23438 & n23440;
  assign n23442 = ~pi0789 & ~n23336;
  assign n23443 = ~n23339 & ~n23426;
  assign n23444 = pi0789 & ~n23443;
  assign n23445 = ~n23442 & ~n23444;
  assign n23446 = ~pi0626 & ~n23445;
  assign n23447 = pi0626 & n23227;
  assign n23448 = pi0641 & ~n23447;
  assign n23449 = ~n23446 & n23448;
  assign n23450 = ~pi1158 & ~n23449;
  assign n23451 = ~n23441 & n23450;
  assign n23452 = pi0626 & n23436;
  assign n23453 = ~pi0626 & n23259;
  assign n23454 = pi0641 & ~n23453;
  assign n23455 = ~n23452 & n23454;
  assign n23456 = pi0626 & ~n23445;
  assign n23457 = ~pi0626 & n23227;
  assign n23458 = ~pi0641 & ~n23457;
  assign n23459 = ~n23456 & n23458;
  assign n23460 = pi1158 & ~n23459;
  assign n23461 = ~n23455 & n23460;
  assign n23462 = ~n23451 & ~n23461;
  assign n23463 = pi0788 & ~n23462;
  assign n23464 = ~n23437 & ~n23463;
  assign n23465 = ~pi0628 & n23464;
  assign n23466 = ~n17969 & ~n23445;
  assign n23467 = n17969 & n23227;
  assign n23468 = ~n23466 & ~n23467;
  assign n23469 = pi0628 & n23468;
  assign n23470 = ~pi1156 & ~n23469;
  assign n23471 = ~n23465 & n23470;
  assign n23472 = ~pi0629 & ~n23267;
  assign n23473 = ~n23471 & n23472;
  assign n23474 = pi0628 & n23464;
  assign n23475 = ~pi0628 & n23468;
  assign n23476 = pi1156 & ~n23475;
  assign n23477 = ~n23474 & n23476;
  assign n23478 = pi0629 & ~n23271;
  assign n23479 = ~n23477 & n23478;
  assign n23480 = ~n23473 & ~n23479;
  assign n23481 = pi0792 & ~n23480;
  assign n23482 = ~pi0792 & n23464;
  assign n23483 = ~n23481 & ~n23482;
  assign n23484 = ~pi0647 & ~n23483;
  assign n23485 = ~n17779 & ~n23468;
  assign n23486 = n17779 & n23227;
  assign n23487 = ~n23485 & ~n23486;
  assign n23488 = pi0647 & n23487;
  assign n23489 = ~pi1157 & ~n23488;
  assign n23490 = ~n23484 & n23489;
  assign n23491 = ~pi0630 & ~n23279;
  assign n23492 = ~n23490 & n23491;
  assign n23493 = pi0647 & ~n23483;
  assign n23494 = ~pi0647 & n23487;
  assign n23495 = pi1157 & ~n23494;
  assign n23496 = ~n23493 & n23495;
  assign n23497 = pi0630 & ~n23283;
  assign n23498 = ~n23496 & n23497;
  assign n23499 = ~n23492 & ~n23498;
  assign n23500 = pi0787 & ~n23499;
  assign n23501 = ~pi0787 & ~n23483;
  assign n23502 = ~n23500 & ~n23501;
  assign n23503 = pi0644 & ~n23502;
  assign n23504 = pi0715 & ~n23287;
  assign n23505 = ~n23503 & n23504;
  assign n23506 = n17804 & ~n23227;
  assign n23507 = ~n17804 & n23487;
  assign n23508 = ~n23506 & ~n23507;
  assign n23509 = pi0644 & ~n23508;
  assign n23510 = ~pi0644 & ~n23227;
  assign n23511 = ~pi0715 & ~n23510;
  assign n23512 = ~n23509 & n23511;
  assign n23513 = pi1160 & ~n23512;
  assign n23514 = ~n23505 & n23513;
  assign n23515 = ~pi0644 & ~n23502;
  assign n23516 = pi0644 & n23286;
  assign n23517 = ~pi0715 & ~n23516;
  assign n23518 = ~n23515 & n23517;
  assign n23519 = ~pi0644 & ~n23508;
  assign n23520 = pi0644 & ~n23227;
  assign n23521 = pi0715 & ~n23520;
  assign n23522 = ~n23519 & n23521;
  assign n23523 = ~pi1160 & ~n23522;
  assign n23524 = ~n23518 & n23523;
  assign n23525 = pi0790 & ~n23514;
  assign n23526 = ~n23524 & n23525;
  assign n23527 = ~pi0790 & n23502;
  assign n23528 = n6305 & ~n23527;
  assign n23529 = ~n23526 & n23528;
  assign n23530 = ~pi0174 & ~n6305;
  assign n23531 = ~pi0057 & ~n23530;
  assign n23532 = ~n23529 & n23531;
  assign n23533 = pi0057 & pi0174;
  assign n23534 = ~pi0832 & ~n23533;
  assign n23535 = ~n23532 & n23534;
  assign n23536 = pi0174 & ~n2926;
  assign n23537 = pi0759 & n17244;
  assign n23538 = n17291 & n23537;
  assign n23539 = pi1155 & ~n23536;
  assign n23540 = ~n23538 & n23539;
  assign n23541 = pi0696 & n16645;
  assign n23542 = ~n23536 & ~n23541;
  assign n23543 = ~pi0778 & n23542;
  assign n23544 = pi0625 & n23541;
  assign n23545 = ~n23542 & ~n23544;
  assign n23546 = ~pi1153 & ~n23545;
  assign n23547 = pi1153 & ~n23536;
  assign n23548 = ~n23544 & n23547;
  assign n23549 = ~n23546 & ~n23548;
  assign n23550 = pi0778 & ~n23549;
  assign n23551 = ~n23543 & ~n23550;
  assign n23552 = pi0609 & n23551;
  assign n23553 = ~n23536 & ~n23537;
  assign n23554 = pi0696 & n17469;
  assign n23555 = n23553 & ~n23554;
  assign n23556 = pi0625 & n23554;
  assign n23557 = ~n23555 & ~n23556;
  assign n23558 = ~pi1153 & ~n23557;
  assign n23559 = ~pi0608 & ~n23548;
  assign n23560 = ~n23558 & n23559;
  assign n23561 = pi1153 & n23553;
  assign n23562 = ~n23556 & n23561;
  assign n23563 = pi0608 & ~n23546;
  assign n23564 = ~n23562 & n23563;
  assign n23565 = ~n23560 & ~n23564;
  assign n23566 = pi0778 & ~n23565;
  assign n23567 = ~pi0778 & ~n23555;
  assign n23568 = ~n23566 & ~n23567;
  assign n23569 = ~pi0609 & ~n23568;
  assign n23570 = ~pi1155 & ~n23552;
  assign n23571 = ~n23569 & n23570;
  assign n23572 = ~pi0660 & ~n23540;
  assign n23573 = ~n23571 & n23572;
  assign n23574 = n17296 & n23537;
  assign n23575 = ~pi1155 & ~n23536;
  assign n23576 = ~n23574 & n23575;
  assign n23577 = ~pi0609 & n23551;
  assign n23578 = pi0609 & ~n23568;
  assign n23579 = pi1155 & ~n23577;
  assign n23580 = ~n23578 & n23579;
  assign n23581 = pi0660 & ~n23576;
  assign n23582 = ~n23580 & n23581;
  assign n23583 = ~n23573 & ~n23582;
  assign n23584 = pi0785 & ~n23583;
  assign n23585 = ~pi0785 & ~n23568;
  assign n23586 = ~n23584 & ~n23585;
  assign n23587 = ~pi0781 & ~n23586;
  assign n23588 = ~n20225 & n23537;
  assign n23589 = n20270 & n23588;
  assign n23590 = pi1154 & ~n23536;
  assign n23591 = ~n23589 & n23590;
  assign n23592 = ~n17075 & n23551;
  assign n23593 = ~n23536 & ~n23592;
  assign n23594 = pi0618 & ~n23593;
  assign n23595 = ~pi0618 & ~n23586;
  assign n23596 = ~pi1154 & ~n23594;
  assign n23597 = ~n23595 & n23596;
  assign n23598 = ~pi0627 & ~n23591;
  assign n23599 = ~n23597 & n23598;
  assign n23600 = n20319 & n23588;
  assign n23601 = ~pi1154 & ~n23536;
  assign n23602 = ~n23600 & n23601;
  assign n23603 = ~pi0618 & ~n23593;
  assign n23604 = pi0618 & ~n23586;
  assign n23605 = pi1154 & ~n23603;
  assign n23606 = ~n23604 & n23605;
  assign n23607 = pi0627 & ~n23602;
  assign n23608 = ~n23606 & n23607;
  assign n23609 = ~n23599 & ~n23608;
  assign n23610 = pi0781 & ~n23609;
  assign n23611 = pi0648 & n20228;
  assign n23612 = ~pi0648 & n20229;
  assign n23613 = ~n23611 & ~n23612;
  assign n23614 = n16634 & n23613;
  assign n23615 = pi0789 & ~n23614;
  assign n23616 = ~n23587 & ~n23615;
  assign n23617 = ~n23610 & n23616;
  assign n23618 = ~n20235 & n23588;
  assign n23619 = n20345 & n23618;
  assign n23620 = n16633 & ~n23619;
  assign n23621 = n19150 & n23551;
  assign n23622 = ~n23613 & ~n23621;
  assign n23623 = n20335 & n23618;
  assign n23624 = n16632 & ~n23623;
  assign n23625 = ~n23620 & ~n23624;
  assign n23626 = ~n23622 & n23625;
  assign n23627 = pi0789 & ~n23536;
  assign n23628 = ~n23626 & n23627;
  assign n23629 = n17970 & ~n23628;
  assign n23630 = ~n23617 & n23629;
  assign n23631 = n20237 & n23588;
  assign n23632 = ~pi0626 & n23631;
  assign n23633 = ~n23536 & ~n23632;
  assign n23634 = ~pi1158 & ~n23633;
  assign n23635 = ~n16635 & n23621;
  assign n23636 = ~n23536 & ~n23635;
  assign n23637 = n17865 & ~n23636;
  assign n23638 = pi0641 & ~n23634;
  assign n23639 = ~n23637 & n23638;
  assign n23640 = n17866 & ~n23636;
  assign n23641 = pi0626 & n23631;
  assign n23642 = ~n23536 & ~n23641;
  assign n23643 = pi1158 & ~n23642;
  assign n23644 = ~pi0641 & ~n23643;
  assign n23645 = ~n23640 & n23644;
  assign n23646 = pi0788 & ~n23639;
  assign n23647 = ~n23645 & n23646;
  assign n23648 = ~n20364 & ~n23647;
  assign n23649 = ~n23630 & n23648;
  assign n23650 = ~n17969 & n23631;
  assign n23651 = ~pi0629 & n23650;
  assign n23652 = pi0628 & ~n23651;
  assign n23653 = n19151 & n23551;
  assign n23654 = pi0629 & ~n23653;
  assign n23655 = ~n23652 & ~n23654;
  assign n23656 = ~pi1156 & ~n23655;
  assign n23657 = ~pi0628 & ~n23650;
  assign n23658 = pi0629 & ~n23657;
  assign n23659 = pi0628 & n23653;
  assign n23660 = pi1156 & ~n23658;
  assign n23661 = ~n23659 & n23660;
  assign n23662 = ~n23656 & ~n23661;
  assign n23663 = pi0792 & ~n23536;
  assign n23664 = ~n23662 & n23663;
  assign n23665 = ~n23649 & ~n23664;
  assign n23666 = ~n20206 & ~n23665;
  assign n23667 = ~n17779 & n23650;
  assign n23668 = ~pi0630 & n23667;
  assign n23669 = pi0647 & ~n23668;
  assign n23670 = ~n19142 & n23653;
  assign n23671 = pi0630 & ~n23670;
  assign n23672 = ~n23669 & ~n23671;
  assign n23673 = ~pi1157 & ~n23672;
  assign n23674 = pi0630 & n23667;
  assign n23675 = ~pi0630 & ~n23670;
  assign n23676 = pi0647 & ~n23675;
  assign n23677 = pi1157 & ~n23674;
  assign n23678 = ~n23676 & n23677;
  assign n23679 = ~n23673 & ~n23678;
  assign n23680 = pi0787 & ~n23536;
  assign n23681 = ~n23679 & n23680;
  assign n23682 = ~n23666 & ~n23681;
  assign n23683 = ~pi0790 & n23682;
  assign n23684 = ~n17779 & ~n17804;
  assign n23685 = n23650 & n23684;
  assign n23686 = pi0644 & n23685;
  assign n23687 = ~pi0715 & ~n23536;
  assign n23688 = ~n23686 & n23687;
  assign n23689 = ~n19342 & n23670;
  assign n23690 = ~n23536 & ~n23689;
  assign n23691 = ~pi0644 & ~n23690;
  assign n23692 = pi0644 & n23682;
  assign n23693 = pi0715 & ~n23691;
  assign n23694 = ~n23692 & n23693;
  assign n23695 = pi1160 & ~n23688;
  assign n23696 = ~n23694 & n23695;
  assign n23697 = ~pi0644 & n23685;
  assign n23698 = pi0715 & ~n23536;
  assign n23699 = ~n23697 & n23698;
  assign n23700 = ~pi0644 & n23682;
  assign n23701 = pi0644 & ~n23690;
  assign n23702 = ~pi0715 & ~n23701;
  assign n23703 = ~n23700 & n23702;
  assign n23704 = ~pi1160 & ~n23699;
  assign n23705 = ~n23703 & n23704;
  assign n23706 = ~n23696 & ~n23705;
  assign n23707 = pi0790 & ~n23706;
  assign n23708 = pi0832 & ~n23683;
  assign n23709 = ~n23707 & n23708;
  assign po0331 = ~n23535 & ~n23709;
  assign n23711 = ~pi0175 & ~n2926;
  assign n23712 = pi0700 & n16645;
  assign n23713 = ~n23711 & ~n23712;
  assign n23714 = ~pi0778 & ~n23713;
  assign n23715 = ~pi0625 & n23712;
  assign n23716 = ~n23713 & ~n23715;
  assign n23717 = pi1153 & ~n23716;
  assign n23718 = ~pi1153 & ~n23711;
  assign n23719 = ~n23715 & n23718;
  assign n23720 = pi0778 & ~n23719;
  assign n23721 = ~n23717 & n23720;
  assign n23722 = ~n23714 & ~n23721;
  assign n23723 = ~n17845 & ~n23722;
  assign n23724 = ~n17847 & n23723;
  assign n23725 = ~n17849 & n23724;
  assign n23726 = ~n17851 & n23725;
  assign n23727 = ~n17857 & n23726;
  assign n23728 = ~pi0647 & n23727;
  assign n23729 = pi0647 & n23711;
  assign n23730 = ~pi1157 & ~n23729;
  assign n23731 = ~n23728 & n23730;
  assign n23732 = pi0630 & n23731;
  assign n23733 = pi0766 & n17244;
  assign n23734 = ~n23711 & ~n23733;
  assign n23735 = ~n17874 & ~n23734;
  assign n23736 = ~pi0785 & ~n23735;
  assign n23737 = n17296 & n23733;
  assign n23738 = n23735 & ~n23737;
  assign n23739 = pi1155 & ~n23738;
  assign n23740 = ~pi1155 & ~n23711;
  assign n23741 = ~n23737 & n23740;
  assign n23742 = ~n23739 & ~n23741;
  assign n23743 = pi0785 & ~n23742;
  assign n23744 = ~n23736 & ~n23743;
  assign n23745 = ~pi0781 & ~n23744;
  assign n23746 = ~n17889 & n23744;
  assign n23747 = pi1154 & ~n23746;
  assign n23748 = ~n17892 & n23744;
  assign n23749 = ~pi1154 & ~n23748;
  assign n23750 = ~n23747 & ~n23749;
  assign n23751 = pi0781 & ~n23750;
  assign n23752 = ~n23745 & ~n23751;
  assign n23753 = ~pi0789 & ~n23752;
  assign n23754 = ~n23078 & n23752;
  assign n23755 = pi1159 & ~n23754;
  assign n23756 = ~n23081 & n23752;
  assign n23757 = ~pi1159 & ~n23756;
  assign n23758 = ~n23755 & ~n23757;
  assign n23759 = pi0789 & ~n23758;
  assign n23760 = ~n23753 & ~n23759;
  assign n23761 = ~n17969 & n23760;
  assign n23762 = n17969 & n23711;
  assign n23763 = ~n23761 & ~n23762;
  assign n23764 = ~n17779 & ~n23763;
  assign n23765 = n17779 & n23711;
  assign n23766 = ~n23764 & ~n23765;
  assign n23767 = ~n20559 & n23766;
  assign n23768 = pi0647 & ~n23727;
  assign n23769 = ~pi0647 & ~n23711;
  assign n23770 = ~n23768 & ~n23769;
  assign n23771 = n17801 & ~n23770;
  assign n23772 = ~n23732 & ~n23771;
  assign n23773 = ~n23767 & n23772;
  assign n23774 = pi0787 & ~n23773;
  assign n23775 = n17871 & n23725;
  assign n23776 = ~pi0626 & ~n23760;
  assign n23777 = pi0626 & ~n23711;
  assign n23778 = n16629 & ~n23777;
  assign n23779 = ~n23776 & n23778;
  assign n23780 = pi0626 & ~n23760;
  assign n23781 = ~pi0626 & ~n23711;
  assign n23782 = n16628 & ~n23781;
  assign n23783 = ~n23780 & n23782;
  assign n23784 = ~n23775 & ~n23779;
  assign n23785 = ~n23783 & n23784;
  assign n23786 = pi0788 & ~n23785;
  assign n23787 = pi0618 & n23723;
  assign n23788 = ~n17168 & ~n23713;
  assign n23789 = pi0625 & n23788;
  assign n23790 = n23734 & ~n23788;
  assign n23791 = ~n23789 & ~n23790;
  assign n23792 = n23718 & ~n23791;
  assign n23793 = ~pi0608 & ~n23717;
  assign n23794 = ~n23792 & n23793;
  assign n23795 = pi1153 & n23734;
  assign n23796 = ~n23789 & n23795;
  assign n23797 = pi0608 & ~n23719;
  assign n23798 = ~n23796 & n23797;
  assign n23799 = ~n23794 & ~n23798;
  assign n23800 = pi0778 & ~n23799;
  assign n23801 = ~pi0778 & ~n23790;
  assign n23802 = ~n23800 & ~n23801;
  assign n23803 = ~pi0609 & ~n23802;
  assign n23804 = pi0609 & ~n23722;
  assign n23805 = ~pi1155 & ~n23804;
  assign n23806 = ~n23803 & n23805;
  assign n23807 = ~pi0660 & ~n23739;
  assign n23808 = ~n23806 & n23807;
  assign n23809 = pi0609 & ~n23802;
  assign n23810 = ~pi0609 & ~n23722;
  assign n23811 = pi1155 & ~n23810;
  assign n23812 = ~n23809 & n23811;
  assign n23813 = pi0660 & ~n23741;
  assign n23814 = ~n23812 & n23813;
  assign n23815 = ~n23808 & ~n23814;
  assign n23816 = pi0785 & ~n23815;
  assign n23817 = ~pi0785 & ~n23802;
  assign n23818 = ~n23816 & ~n23817;
  assign n23819 = ~pi0618 & ~n23818;
  assign n23820 = ~pi1154 & ~n23787;
  assign n23821 = ~n23819 & n23820;
  assign n23822 = ~pi0627 & ~n23747;
  assign n23823 = ~n23821 & n23822;
  assign n23824 = ~pi0618 & n23723;
  assign n23825 = pi0618 & ~n23818;
  assign n23826 = pi1154 & ~n23824;
  assign n23827 = ~n23825 & n23826;
  assign n23828 = pi0627 & ~n23749;
  assign n23829 = ~n23827 & n23828;
  assign n23830 = ~n23823 & ~n23829;
  assign n23831 = pi0781 & ~n23830;
  assign n23832 = ~pi0781 & ~n23818;
  assign n23833 = ~n23831 & ~n23832;
  assign n23834 = ~pi0789 & n23833;
  assign n23835 = ~pi0619 & ~n23833;
  assign n23836 = pi0619 & n23724;
  assign n23837 = ~pi1159 & ~n23836;
  assign n23838 = ~n23835 & n23837;
  assign n23839 = ~pi0648 & ~n23755;
  assign n23840 = ~n23838 & n23839;
  assign n23841 = pi0619 & ~n23833;
  assign n23842 = ~pi0619 & n23724;
  assign n23843 = pi1159 & ~n23842;
  assign n23844 = ~n23841 & n23843;
  assign n23845 = pi0648 & ~n23757;
  assign n23846 = ~n23844 & n23845;
  assign n23847 = pi0789 & ~n23840;
  assign n23848 = ~n23846 & n23847;
  assign n23849 = n17970 & ~n23834;
  assign n23850 = ~n23848 & n23849;
  assign n23851 = ~n23786 & ~n23850;
  assign n23852 = ~n20364 & ~n23851;
  assign n23853 = n17854 & ~n23763;
  assign n23854 = n20851 & n23726;
  assign n23855 = ~n23853 & ~n23854;
  assign n23856 = ~pi0629 & ~n23855;
  assign n23857 = n20855 & n23726;
  assign n23858 = n17853 & ~n23763;
  assign n23859 = ~n23857 & ~n23858;
  assign n23860 = pi0629 & ~n23859;
  assign n23861 = ~n23856 & ~n23860;
  assign n23862 = pi0792 & ~n23861;
  assign n23863 = ~n20206 & ~n23862;
  assign n23864 = ~n23852 & n23863;
  assign n23865 = ~n23774 & ~n23864;
  assign n23866 = ~pi0790 & n23865;
  assign n23867 = ~pi0787 & ~n23727;
  assign n23868 = pi1157 & ~n23770;
  assign n23869 = ~n23731 & ~n23868;
  assign n23870 = pi0787 & ~n23869;
  assign n23871 = ~n23867 & ~n23870;
  assign n23872 = ~pi0644 & n23871;
  assign n23873 = pi0644 & n23865;
  assign n23874 = pi0715 & ~n23872;
  assign n23875 = ~n23873 & n23874;
  assign n23876 = ~n17804 & ~n23766;
  assign n23877 = n17804 & n23711;
  assign n23878 = ~n23876 & ~n23877;
  assign n23879 = pi0644 & ~n23878;
  assign n23880 = ~pi0644 & n23711;
  assign n23881 = ~pi0715 & ~n23880;
  assign n23882 = ~n23879 & n23881;
  assign n23883 = pi1160 & ~n23882;
  assign n23884 = ~n23875 & n23883;
  assign n23885 = ~pi0644 & ~n23878;
  assign n23886 = pi0644 & n23711;
  assign n23887 = pi0715 & ~n23886;
  assign n23888 = ~n23885 & n23887;
  assign n23889 = pi0644 & n23871;
  assign n23890 = ~pi0644 & n23865;
  assign n23891 = ~pi0715 & ~n23889;
  assign n23892 = ~n23890 & n23891;
  assign n23893 = ~pi1160 & ~n23888;
  assign n23894 = ~n23892 & n23893;
  assign n23895 = ~n23884 & ~n23894;
  assign n23896 = pi0790 & ~n23895;
  assign n23897 = pi0832 & ~n23866;
  assign n23898 = ~n23896 & n23897;
  assign n23899 = ~pi0175 & po1038;
  assign n23900 = ~pi0175 & ~n17059;
  assign n23901 = n16635 & ~n23900;
  assign n23902 = pi0175 & ~n2571;
  assign n23903 = ~pi0175 & ~n16641;
  assign n23904 = n16647 & ~n23903;
  assign n23905 = ~pi0175 & n18072;
  assign n23906 = pi0175 & ~n18076;
  assign n23907 = ~pi0038 & ~n23906;
  assign n23908 = ~n23905 & n23907;
  assign n23909 = pi0700 & ~n23904;
  assign n23910 = ~n23908 & n23909;
  assign n23911 = ~pi0175 & ~pi0700;
  assign n23912 = ~n17052 & n23911;
  assign n23913 = n2571 & ~n23912;
  assign n23914 = ~n23910 & n23913;
  assign n23915 = ~n23902 & ~n23914;
  assign n23916 = ~pi0778 & ~n23915;
  assign n23917 = ~pi0625 & n23900;
  assign n23918 = pi0625 & n23915;
  assign n23919 = pi1153 & ~n23917;
  assign n23920 = ~n23918 & n23919;
  assign n23921 = ~pi0625 & n23915;
  assign n23922 = pi0625 & n23900;
  assign n23923 = ~pi1153 & ~n23922;
  assign n23924 = ~n23921 & n23923;
  assign n23925 = ~n23920 & ~n23924;
  assign n23926 = pi0778 & ~n23925;
  assign n23927 = ~n23916 & ~n23926;
  assign n23928 = ~n17075 & ~n23927;
  assign n23929 = n17075 & ~n23900;
  assign n23930 = ~n23928 & ~n23929;
  assign n23931 = ~n16639 & n23930;
  assign n23932 = n16639 & n23900;
  assign n23933 = ~n23931 & ~n23932;
  assign n23934 = ~n16635 & n23933;
  assign n23935 = ~n23901 & ~n23934;
  assign n23936 = ~n16631 & n23935;
  assign n23937 = n16631 & n23900;
  assign n23938 = ~n23936 & ~n23937;
  assign n23939 = ~pi0628 & ~n23938;
  assign n23940 = pi0628 & n23900;
  assign n23941 = ~n23939 & ~n23940;
  assign n23942 = ~pi1156 & ~n23941;
  assign n23943 = pi0628 & ~n23938;
  assign n23944 = ~pi0628 & n23900;
  assign n23945 = ~n23943 & ~n23944;
  assign n23946 = pi1156 & ~n23945;
  assign n23947 = ~n23942 & ~n23946;
  assign n23948 = pi0792 & ~n23947;
  assign n23949 = ~pi0792 & ~n23938;
  assign n23950 = ~n23948 & ~n23949;
  assign n23951 = ~pi0647 & ~n23950;
  assign n23952 = pi0647 & n23900;
  assign n23953 = ~n23951 & ~n23952;
  assign n23954 = ~pi1157 & ~n23953;
  assign n23955 = pi0647 & ~n23950;
  assign n23956 = ~pi0647 & n23900;
  assign n23957 = ~n23955 & ~n23956;
  assign n23958 = pi1157 & ~n23957;
  assign n23959 = ~n23954 & ~n23958;
  assign n23960 = pi0787 & ~n23959;
  assign n23961 = ~pi0787 & ~n23950;
  assign n23962 = ~n23960 & ~n23961;
  assign n23963 = ~pi0644 & ~n23962;
  assign n23964 = pi0715 & ~n23963;
  assign n23965 = ~pi0766 & n17046;
  assign n23966 = pi0175 & n17273;
  assign n23967 = ~n23965 & ~n23966;
  assign n23968 = pi0039 & ~n23967;
  assign n23969 = pi0766 & ~n17234;
  assign n23970 = pi0175 & ~n23969;
  assign n23971 = ~pi0175 & pi0766;
  assign n23972 = n17221 & n23971;
  assign n23973 = ~n21499 & ~n23970;
  assign n23974 = ~n23972 & n23973;
  assign n23975 = ~n23968 & n23974;
  assign n23976 = ~pi0038 & ~n23975;
  assign n23977 = pi0766 & n17280;
  assign n23978 = pi0038 & ~n23903;
  assign n23979 = ~n23977 & n23978;
  assign n23980 = ~n23976 & ~n23979;
  assign n23981 = n2571 & ~n23980;
  assign n23982 = ~n23902 & ~n23981;
  assign n23983 = ~n17117 & ~n23982;
  assign n23984 = n17117 & ~n23900;
  assign n23985 = ~n23983 & ~n23984;
  assign n23986 = ~pi0785 & ~n23985;
  assign n23987 = ~n17291 & ~n23900;
  assign n23988 = pi0609 & n23983;
  assign n23989 = ~n23987 & ~n23988;
  assign n23990 = pi1155 & ~n23989;
  assign n23991 = ~n17296 & ~n23900;
  assign n23992 = ~pi0609 & n23983;
  assign n23993 = ~n23991 & ~n23992;
  assign n23994 = ~pi1155 & ~n23993;
  assign n23995 = ~n23990 & ~n23994;
  assign n23996 = pi0785 & ~n23995;
  assign n23997 = ~n23986 & ~n23996;
  assign n23998 = ~pi0781 & ~n23997;
  assign n23999 = ~pi0618 & n23900;
  assign n24000 = pi0618 & n23997;
  assign n24001 = pi1154 & ~n23999;
  assign n24002 = ~n24000 & n24001;
  assign n24003 = ~pi0618 & n23997;
  assign n24004 = pi0618 & n23900;
  assign n24005 = ~pi1154 & ~n24004;
  assign n24006 = ~n24003 & n24005;
  assign n24007 = ~n24002 & ~n24006;
  assign n24008 = pi0781 & ~n24007;
  assign n24009 = ~n23998 & ~n24008;
  assign n24010 = ~pi0789 & ~n24009;
  assign n24011 = ~pi0619 & n23900;
  assign n24012 = pi0619 & n24009;
  assign n24013 = pi1159 & ~n24011;
  assign n24014 = ~n24012 & n24013;
  assign n24015 = ~pi0619 & n24009;
  assign n24016 = pi0619 & n23900;
  assign n24017 = ~pi1159 & ~n24016;
  assign n24018 = ~n24015 & n24017;
  assign n24019 = ~n24014 & ~n24018;
  assign n24020 = pi0789 & ~n24019;
  assign n24021 = ~n24010 & ~n24020;
  assign n24022 = ~n17969 & n24021;
  assign n24023 = n17969 & n23900;
  assign n24024 = ~n24022 & ~n24023;
  assign n24025 = ~n17779 & ~n24024;
  assign n24026 = n17779 & n23900;
  assign n24027 = ~n24025 & ~n24026;
  assign n24028 = ~n17804 & ~n24027;
  assign n24029 = n17804 & n23900;
  assign n24030 = ~n24028 & ~n24029;
  assign n24031 = pi0644 & ~n24030;
  assign n24032 = ~pi0644 & n23900;
  assign n24033 = ~pi0715 & ~n24032;
  assign n24034 = ~n24031 & n24033;
  assign n24035 = pi1160 & ~n24034;
  assign n24036 = ~n23964 & n24035;
  assign n24037 = pi0644 & ~n23962;
  assign n24038 = ~pi0715 & ~n24037;
  assign n24039 = ~pi0644 & ~n24030;
  assign n24040 = pi0644 & n23900;
  assign n24041 = pi0715 & ~n24040;
  assign n24042 = ~n24039 & n24041;
  assign n24043 = ~pi1160 & ~n24042;
  assign n24044 = ~n24038 & n24043;
  assign n24045 = ~n24036 & ~n24044;
  assign n24046 = pi0790 & ~n24045;
  assign n24047 = n17777 & n23941;
  assign n24048 = ~n20570 & n24024;
  assign n24049 = n17776 & n23945;
  assign n24050 = ~n24047 & ~n24049;
  assign n24051 = ~n24048 & n24050;
  assign n24052 = pi0792 & ~n24051;
  assign n24053 = pi0609 & n23927;
  assign n24054 = ~pi0700 & n23980;
  assign n24055 = n16667 & ~n17336;
  assign n24056 = ~pi0766 & n24055;
  assign n24057 = ~n17490 & ~n24056;
  assign n24058 = ~pi0039 & ~n24057;
  assign n24059 = ~pi0175 & ~n24058;
  assign n24060 = ~n17469 & ~n23733;
  assign n24061 = pi0175 & ~n24060;
  assign n24062 = n6284 & n24061;
  assign n24063 = pi0038 & ~n24062;
  assign n24064 = ~n24059 & n24063;
  assign n24065 = ~pi0175 & ~n17629;
  assign n24066 = pi0175 & ~n17631;
  assign n24067 = pi0766 & ~n24066;
  assign n24068 = ~n24065 & n24067;
  assign n24069 = ~pi0175 & n17612;
  assign n24070 = pi0175 & n17625;
  assign n24071 = ~pi0766 & ~n24069;
  assign n24072 = ~n24070 & n24071;
  assign n24073 = ~pi0039 & ~n24068;
  assign n24074 = ~n24072 & n24073;
  assign n24075 = pi0175 & n17605;
  assign n24076 = ~pi0175 & ~n17546;
  assign n24077 = pi0766 & ~n24076;
  assign n24078 = ~n24075 & n24077;
  assign n24079 = ~pi0175 & n17404;
  assign n24080 = pi0175 & n17485;
  assign n24081 = ~pi0766 & ~n24080;
  assign n24082 = ~n24079 & n24081;
  assign n24083 = pi0039 & ~n24078;
  assign n24084 = ~n24082 & n24083;
  assign n24085 = ~pi0038 & ~n24074;
  assign n24086 = ~n24084 & n24085;
  assign n24087 = pi0700 & ~n24064;
  assign n24088 = ~n24086 & n24087;
  assign n24089 = n2571 & ~n24088;
  assign n24090 = ~n24054 & n24089;
  assign n24091 = ~n23902 & ~n24090;
  assign n24092 = ~pi0625 & n24091;
  assign n24093 = pi0625 & n23982;
  assign n24094 = ~pi1153 & ~n24093;
  assign n24095 = ~n24092 & n24094;
  assign n24096 = ~pi0608 & ~n23920;
  assign n24097 = ~n24095 & n24096;
  assign n24098 = ~pi0625 & n23982;
  assign n24099 = pi0625 & n24091;
  assign n24100 = pi1153 & ~n24098;
  assign n24101 = ~n24099 & n24100;
  assign n24102 = pi0608 & ~n23924;
  assign n24103 = ~n24101 & n24102;
  assign n24104 = ~n24097 & ~n24103;
  assign n24105 = pi0778 & ~n24104;
  assign n24106 = ~pi0778 & n24091;
  assign n24107 = ~n24105 & ~n24106;
  assign n24108 = ~pi0609 & ~n24107;
  assign n24109 = ~pi1155 & ~n24053;
  assign n24110 = ~n24108 & n24109;
  assign n24111 = ~pi0660 & ~n23990;
  assign n24112 = ~n24110 & n24111;
  assign n24113 = ~pi0609 & n23927;
  assign n24114 = pi0609 & ~n24107;
  assign n24115 = pi1155 & ~n24113;
  assign n24116 = ~n24114 & n24115;
  assign n24117 = pi0660 & ~n23994;
  assign n24118 = ~n24116 & n24117;
  assign n24119 = ~n24112 & ~n24118;
  assign n24120 = pi0785 & ~n24119;
  assign n24121 = ~pi0785 & ~n24107;
  assign n24122 = ~n24120 & ~n24121;
  assign n24123 = ~pi0618 & ~n24122;
  assign n24124 = pi0618 & n23930;
  assign n24125 = ~pi1154 & ~n24124;
  assign n24126 = ~n24123 & n24125;
  assign n24127 = ~pi0627 & ~n24002;
  assign n24128 = ~n24126 & n24127;
  assign n24129 = ~pi0618 & n23930;
  assign n24130 = pi0618 & ~n24122;
  assign n24131 = pi1154 & ~n24129;
  assign n24132 = ~n24130 & n24131;
  assign n24133 = pi0627 & ~n24006;
  assign n24134 = ~n24132 & n24133;
  assign n24135 = ~n24128 & ~n24134;
  assign n24136 = pi0781 & ~n24135;
  assign n24137 = ~pi0781 & ~n24122;
  assign n24138 = ~n24136 & ~n24137;
  assign n24139 = ~pi0789 & n24138;
  assign n24140 = pi0619 & ~n23933;
  assign n24141 = ~pi0619 & ~n24138;
  assign n24142 = ~pi1159 & ~n24140;
  assign n24143 = ~n24141 & n24142;
  assign n24144 = ~pi0648 & ~n24014;
  assign n24145 = ~n24143 & n24144;
  assign n24146 = ~pi0619 & ~n23933;
  assign n24147 = pi0619 & ~n24138;
  assign n24148 = pi1159 & ~n24146;
  assign n24149 = ~n24147 & n24148;
  assign n24150 = pi0648 & ~n24018;
  assign n24151 = ~n24149 & n24150;
  assign n24152 = pi0789 & ~n24145;
  assign n24153 = ~n24151 & n24152;
  assign n24154 = n17970 & ~n24139;
  assign n24155 = ~n24153 & n24154;
  assign n24156 = n17871 & n23935;
  assign n24157 = ~pi0626 & ~n24021;
  assign n24158 = pi0626 & ~n23900;
  assign n24159 = n16629 & ~n24158;
  assign n24160 = ~n24157 & n24159;
  assign n24161 = pi0626 & ~n24021;
  assign n24162 = ~pi0626 & ~n23900;
  assign n24163 = n16628 & ~n24162;
  assign n24164 = ~n24161 & n24163;
  assign n24165 = ~n24156 & ~n24160;
  assign n24166 = ~n24164 & n24165;
  assign n24167 = pi0788 & ~n24166;
  assign n24168 = ~n20364 & ~n24167;
  assign n24169 = ~n24155 & n24168;
  assign n24170 = ~n24052 & ~n24169;
  assign n24171 = ~n20206 & ~n24170;
  assign n24172 = n17802 & n23953;
  assign n24173 = ~n20559 & n24027;
  assign n24174 = n17801 & n23957;
  assign n24175 = ~n24172 & ~n24173;
  assign n24176 = ~n24174 & n24175;
  assign n24177 = pi0787 & ~n24176;
  assign n24178 = ~pi0644 & n24043;
  assign n24179 = pi0644 & n24035;
  assign n24180 = pi0790 & ~n24178;
  assign n24181 = ~n24179 & n24180;
  assign n24182 = ~n24171 & ~n24177;
  assign n24183 = ~n24181 & n24182;
  assign n24184 = ~n24046 & ~n24183;
  assign n24185 = ~po1038 & ~n24184;
  assign n24186 = ~pi0832 & ~n23899;
  assign n24187 = ~n24185 & n24186;
  assign po0332 = ~n23898 & ~n24187;
  assign n24189 = ~pi0176 & ~n2926;
  assign n24190 = ~pi0704 & n16645;
  assign n24191 = ~n24189 & ~n24190;
  assign n24192 = ~pi0778 & n24191;
  assign n24193 = ~pi0625 & n24190;
  assign n24194 = ~n24191 & ~n24193;
  assign n24195 = pi1153 & ~n24194;
  assign n24196 = ~pi1153 & ~n24189;
  assign n24197 = ~n24193 & n24196;
  assign n24198 = ~n24195 & ~n24197;
  assign n24199 = pi0778 & ~n24198;
  assign n24200 = ~n24192 & ~n24199;
  assign n24201 = ~n17845 & n24200;
  assign n24202 = ~n17847 & n24201;
  assign n24203 = ~n17849 & n24202;
  assign n24204 = ~n17851 & n24203;
  assign n24205 = ~n17857 & n24204;
  assign n24206 = ~pi0647 & n24205;
  assign n24207 = pi0647 & n24189;
  assign n24208 = ~pi1157 & ~n24207;
  assign n24209 = ~n24206 & n24208;
  assign n24210 = pi0630 & n24209;
  assign n24211 = ~pi0742 & n17244;
  assign n24212 = ~n24189 & ~n24211;
  assign n24213 = ~n17874 & ~n24212;
  assign n24214 = ~pi0785 & ~n24213;
  assign n24215 = ~n17879 & ~n24212;
  assign n24216 = pi1155 & ~n24215;
  assign n24217 = ~n17882 & n24213;
  assign n24218 = ~pi1155 & ~n24217;
  assign n24219 = ~n24216 & ~n24218;
  assign n24220 = pi0785 & ~n24219;
  assign n24221 = ~n24214 & ~n24220;
  assign n24222 = ~pi0781 & ~n24221;
  assign n24223 = ~n17889 & n24221;
  assign n24224 = pi1154 & ~n24223;
  assign n24225 = ~n17892 & n24221;
  assign n24226 = ~pi1154 & ~n24225;
  assign n24227 = ~n24224 & ~n24226;
  assign n24228 = pi0781 & ~n24227;
  assign n24229 = ~n24222 & ~n24228;
  assign n24230 = ~pi0789 & ~n24229;
  assign n24231 = ~pi0619 & n24189;
  assign n24232 = pi0619 & n24229;
  assign n24233 = pi1159 & ~n24231;
  assign n24234 = ~n24232 & n24233;
  assign n24235 = ~pi0619 & n24229;
  assign n24236 = pi0619 & n24189;
  assign n24237 = ~pi1159 & ~n24236;
  assign n24238 = ~n24235 & n24237;
  assign n24239 = ~n24234 & ~n24238;
  assign n24240 = pi0789 & ~n24239;
  assign n24241 = ~n24230 & ~n24240;
  assign n24242 = ~n17969 & n24241;
  assign n24243 = n17969 & n24189;
  assign n24244 = ~n24242 & ~n24243;
  assign n24245 = ~n17779 & ~n24244;
  assign n24246 = n17779 & n24189;
  assign n24247 = ~n24245 & ~n24246;
  assign n24248 = ~n20559 & n24247;
  assign n24249 = pi0647 & ~n24205;
  assign n24250 = ~pi0647 & ~n24189;
  assign n24251 = ~n24249 & ~n24250;
  assign n24252 = n17801 & ~n24251;
  assign n24253 = ~n24210 & ~n24252;
  assign n24254 = ~n24248 & n24253;
  assign n24255 = pi0787 & ~n24254;
  assign n24256 = n17871 & n24203;
  assign n24257 = ~pi0626 & ~n24241;
  assign n24258 = pi0626 & ~n24189;
  assign n24259 = n16629 & ~n24258;
  assign n24260 = ~n24257 & n24259;
  assign n24261 = pi0626 & ~n24241;
  assign n24262 = ~pi0626 & ~n24189;
  assign n24263 = n16628 & ~n24262;
  assign n24264 = ~n24261 & n24263;
  assign n24265 = ~n24256 & ~n24260;
  assign n24266 = ~n24264 & n24265;
  assign n24267 = pi0788 & ~n24266;
  assign n24268 = pi0618 & n24201;
  assign n24269 = pi0609 & n24200;
  assign n24270 = ~n17168 & ~n24191;
  assign n24271 = pi0625 & n24270;
  assign n24272 = n24212 & ~n24270;
  assign n24273 = ~n24271 & ~n24272;
  assign n24274 = n24196 & ~n24273;
  assign n24275 = ~pi0608 & ~n24195;
  assign n24276 = ~n24274 & n24275;
  assign n24277 = pi1153 & n24212;
  assign n24278 = ~n24271 & n24277;
  assign n24279 = pi0608 & ~n24197;
  assign n24280 = ~n24278 & n24279;
  assign n24281 = ~n24276 & ~n24280;
  assign n24282 = pi0778 & ~n24281;
  assign n24283 = ~pi0778 & ~n24272;
  assign n24284 = ~n24282 & ~n24283;
  assign n24285 = ~pi0609 & ~n24284;
  assign n24286 = ~pi1155 & ~n24269;
  assign n24287 = ~n24285 & n24286;
  assign n24288 = ~pi0660 & ~n24216;
  assign n24289 = ~n24287 & n24288;
  assign n24290 = ~pi0609 & n24200;
  assign n24291 = pi0609 & ~n24284;
  assign n24292 = pi1155 & ~n24290;
  assign n24293 = ~n24291 & n24292;
  assign n24294 = pi0660 & ~n24218;
  assign n24295 = ~n24293 & n24294;
  assign n24296 = ~n24289 & ~n24295;
  assign n24297 = pi0785 & ~n24296;
  assign n24298 = ~pi0785 & ~n24284;
  assign n24299 = ~n24297 & ~n24298;
  assign n24300 = ~pi0618 & ~n24299;
  assign n24301 = ~pi1154 & ~n24268;
  assign n24302 = ~n24300 & n24301;
  assign n24303 = ~pi0627 & ~n24224;
  assign n24304 = ~n24302 & n24303;
  assign n24305 = ~pi0618 & n24201;
  assign n24306 = pi0618 & ~n24299;
  assign n24307 = pi1154 & ~n24305;
  assign n24308 = ~n24306 & n24307;
  assign n24309 = pi0627 & ~n24226;
  assign n24310 = ~n24308 & n24309;
  assign n24311 = ~n24304 & ~n24310;
  assign n24312 = pi0781 & ~n24311;
  assign n24313 = ~pi0781 & ~n24299;
  assign n24314 = ~n24312 & ~n24313;
  assign n24315 = ~pi0789 & n24314;
  assign n24316 = ~pi0619 & ~n24314;
  assign n24317 = pi0619 & n24202;
  assign n24318 = ~pi1159 & ~n24317;
  assign n24319 = ~n24316 & n24318;
  assign n24320 = ~pi0648 & ~n24234;
  assign n24321 = ~n24319 & n24320;
  assign n24322 = pi0619 & ~n24314;
  assign n24323 = ~pi0619 & n24202;
  assign n24324 = pi1159 & ~n24323;
  assign n24325 = ~n24322 & n24324;
  assign n24326 = pi0648 & ~n24238;
  assign n24327 = ~n24325 & n24326;
  assign n24328 = pi0789 & ~n24321;
  assign n24329 = ~n24327 & n24328;
  assign n24330 = n17970 & ~n24315;
  assign n24331 = ~n24329 & n24330;
  assign n24332 = ~n24267 & ~n24331;
  assign n24333 = ~n20364 & ~n24332;
  assign n24334 = n17854 & ~n24244;
  assign n24335 = n20851 & n24204;
  assign n24336 = ~n24334 & ~n24335;
  assign n24337 = ~pi0629 & ~n24336;
  assign n24338 = n20855 & n24204;
  assign n24339 = n17853 & ~n24244;
  assign n24340 = ~n24338 & ~n24339;
  assign n24341 = pi0629 & ~n24340;
  assign n24342 = ~n24337 & ~n24341;
  assign n24343 = pi0792 & ~n24342;
  assign n24344 = ~n20206 & ~n24343;
  assign n24345 = ~n24333 & n24344;
  assign n24346 = ~n24255 & ~n24345;
  assign n24347 = ~pi0790 & n24346;
  assign n24348 = ~pi0787 & ~n24205;
  assign n24349 = pi1157 & ~n24251;
  assign n24350 = ~n24209 & ~n24349;
  assign n24351 = pi0787 & ~n24350;
  assign n24352 = ~n24348 & ~n24351;
  assign n24353 = ~pi0644 & n24352;
  assign n24354 = pi0644 & n24346;
  assign n24355 = pi0715 & ~n24353;
  assign n24356 = ~n24354 & n24355;
  assign n24357 = ~n17804 & ~n24247;
  assign n24358 = n17804 & n24189;
  assign n24359 = ~n24357 & ~n24358;
  assign n24360 = pi0644 & ~n24359;
  assign n24361 = ~pi0644 & n24189;
  assign n24362 = ~pi0715 & ~n24361;
  assign n24363 = ~n24360 & n24362;
  assign n24364 = pi1160 & ~n24363;
  assign n24365 = ~n24356 & n24364;
  assign n24366 = ~pi0644 & ~n24359;
  assign n24367 = pi0644 & n24189;
  assign n24368 = pi0715 & ~n24367;
  assign n24369 = ~n24366 & n24368;
  assign n24370 = pi0644 & n24352;
  assign n24371 = ~pi0644 & n24346;
  assign n24372 = ~pi0715 & ~n24370;
  assign n24373 = ~n24371 & n24372;
  assign n24374 = ~pi1160 & ~n24369;
  assign n24375 = ~n24373 & n24374;
  assign n24376 = ~n24365 & ~n24375;
  assign n24377 = pi0790 & ~n24376;
  assign n24378 = pi0832 & ~n24347;
  assign n24379 = ~n24377 & n24378;
  assign n24380 = ~pi0176 & po1038;
  assign n24381 = ~pi0176 & ~n17059;
  assign n24382 = n16635 & ~n24381;
  assign n24383 = ~pi0038 & n18076;
  assign n24384 = n2571 & ~n16647;
  assign n24385 = ~n24383 & n24384;
  assign n24386 = pi0176 & ~n24385;
  assign n24387 = ~pi0038 & n18072;
  assign n24388 = ~n19899 & ~n24387;
  assign n24389 = ~pi0176 & n24388;
  assign n24390 = ~pi0704 & ~n24389;
  assign n24391 = ~pi0176 & ~n17052;
  assign n24392 = pi0704 & n24391;
  assign n24393 = n2571 & ~n24392;
  assign n24394 = ~n24390 & n24393;
  assign n24395 = ~n24386 & ~n24394;
  assign n24396 = ~pi0778 & ~n24395;
  assign n24397 = ~pi0625 & n24381;
  assign n24398 = pi0625 & n24395;
  assign n24399 = pi1153 & ~n24397;
  assign n24400 = ~n24398 & n24399;
  assign n24401 = ~pi0625 & n24395;
  assign n24402 = pi0625 & n24381;
  assign n24403 = ~pi1153 & ~n24402;
  assign n24404 = ~n24401 & n24403;
  assign n24405 = ~n24400 & ~n24404;
  assign n24406 = pi0778 & ~n24405;
  assign n24407 = ~n24396 & ~n24406;
  assign n24408 = ~n17075 & ~n24407;
  assign n24409 = n17075 & ~n24381;
  assign n24410 = ~n24408 & ~n24409;
  assign n24411 = ~n16639 & n24410;
  assign n24412 = n16639 & n24381;
  assign n24413 = ~n24411 & ~n24412;
  assign n24414 = ~n16635 & n24413;
  assign n24415 = ~n24382 & ~n24414;
  assign n24416 = ~n16631 & n24415;
  assign n24417 = n16631 & n24381;
  assign n24418 = ~n24416 & ~n24417;
  assign n24419 = ~pi0628 & ~n24418;
  assign n24420 = pi0628 & n24381;
  assign n24421 = ~n24419 & ~n24420;
  assign n24422 = ~pi1156 & ~n24421;
  assign n24423 = pi0628 & ~n24418;
  assign n24424 = ~pi0628 & n24381;
  assign n24425 = ~n24423 & ~n24424;
  assign n24426 = pi1156 & ~n24425;
  assign n24427 = ~n24422 & ~n24426;
  assign n24428 = pi0792 & ~n24427;
  assign n24429 = ~pi0792 & ~n24418;
  assign n24430 = ~n24428 & ~n24429;
  assign n24431 = ~pi0647 & ~n24430;
  assign n24432 = pi0647 & n24381;
  assign n24433 = ~n24431 & ~n24432;
  assign n24434 = ~pi1157 & ~n24433;
  assign n24435 = pi0647 & ~n24430;
  assign n24436 = ~pi0647 & n24381;
  assign n24437 = ~n24435 & ~n24436;
  assign n24438 = pi1157 & ~n24437;
  assign n24439 = ~n24434 & ~n24438;
  assign n24440 = pi0787 & ~n24439;
  assign n24441 = ~pi0787 & ~n24430;
  assign n24442 = ~n24440 & ~n24441;
  assign n24443 = ~pi0644 & ~n24442;
  assign n24444 = pi0715 & ~n24443;
  assign n24445 = pi0176 & ~n2571;
  assign n24446 = ~pi0176 & n19439;
  assign n24447 = ~n19433 & ~n19434;
  assign n24448 = pi0176 & n24447;
  assign n24449 = ~n24446 & ~n24448;
  assign n24450 = ~pi0742 & ~n24449;
  assign n24451 = pi0742 & ~n24391;
  assign n24452 = ~n24450 & ~n24451;
  assign n24453 = n2571 & ~n24452;
  assign n24454 = ~n24445 & ~n24453;
  assign n24455 = ~n17117 & ~n24454;
  assign n24456 = n17117 & ~n24381;
  assign n24457 = ~n24455 & ~n24456;
  assign n24458 = ~pi0785 & ~n24457;
  assign n24459 = ~n17291 & ~n24381;
  assign n24460 = pi0609 & n24455;
  assign n24461 = ~n24459 & ~n24460;
  assign n24462 = pi1155 & ~n24461;
  assign n24463 = ~n17296 & ~n24381;
  assign n24464 = ~pi0609 & n24455;
  assign n24465 = ~n24463 & ~n24464;
  assign n24466 = ~pi1155 & ~n24465;
  assign n24467 = ~n24462 & ~n24466;
  assign n24468 = pi0785 & ~n24467;
  assign n24469 = ~n24458 & ~n24468;
  assign n24470 = ~pi0781 & ~n24469;
  assign n24471 = ~pi0618 & n24381;
  assign n24472 = pi0618 & n24469;
  assign n24473 = pi1154 & ~n24471;
  assign n24474 = ~n24472 & n24473;
  assign n24475 = ~pi0618 & n24469;
  assign n24476 = pi0618 & n24381;
  assign n24477 = ~pi1154 & ~n24476;
  assign n24478 = ~n24475 & n24477;
  assign n24479 = ~n24474 & ~n24478;
  assign n24480 = pi0781 & ~n24479;
  assign n24481 = ~n24470 & ~n24480;
  assign n24482 = ~pi0789 & ~n24481;
  assign n24483 = ~pi0619 & n24381;
  assign n24484 = pi0619 & n24481;
  assign n24485 = pi1159 & ~n24483;
  assign n24486 = ~n24484 & n24485;
  assign n24487 = ~pi0619 & n24481;
  assign n24488 = pi0619 & n24381;
  assign n24489 = ~pi1159 & ~n24488;
  assign n24490 = ~n24487 & n24489;
  assign n24491 = ~n24486 & ~n24490;
  assign n24492 = pi0789 & ~n24491;
  assign n24493 = ~n24482 & ~n24492;
  assign n24494 = ~n17969 & n24493;
  assign n24495 = n17969 & n24381;
  assign n24496 = ~n24494 & ~n24495;
  assign n24497 = ~n17779 & ~n24496;
  assign n24498 = n17779 & n24381;
  assign n24499 = ~n24497 & ~n24498;
  assign n24500 = ~n17804 & ~n24499;
  assign n24501 = n17804 & n24381;
  assign n24502 = ~n24500 & ~n24501;
  assign n24503 = pi0644 & ~n24502;
  assign n24504 = ~pi0644 & n24381;
  assign n24505 = ~pi0715 & ~n24504;
  assign n24506 = ~n24503 & n24505;
  assign n24507 = pi1160 & ~n24506;
  assign n24508 = ~n24444 & n24507;
  assign n24509 = pi0644 & ~n24442;
  assign n24510 = ~pi0715 & ~n24509;
  assign n24511 = ~pi0644 & ~n24502;
  assign n24512 = pi0644 & n24381;
  assign n24513 = pi0715 & ~n24512;
  assign n24514 = ~n24511 & n24513;
  assign n24515 = ~pi1160 & ~n24514;
  assign n24516 = ~n24510 & n24515;
  assign n24517 = ~n24508 & ~n24516;
  assign n24518 = pi0790 & ~n24517;
  assign n24519 = n17802 & n24433;
  assign n24520 = ~n20559 & n24499;
  assign n24521 = n17801 & n24437;
  assign n24522 = ~n24519 & ~n24520;
  assign n24523 = ~n24521 & n24522;
  assign n24524 = pi0787 & ~n24523;
  assign n24525 = n17777 & n24421;
  assign n24526 = ~n20570 & n24496;
  assign n24527 = n17776 & n24425;
  assign n24528 = ~n24525 & ~n24527;
  assign n24529 = ~n24526 & n24528;
  assign n24530 = pi0792 & ~n24529;
  assign n24531 = n17871 & n24415;
  assign n24532 = ~pi0626 & ~n24493;
  assign n24533 = pi0626 & ~n24381;
  assign n24534 = n16629 & ~n24533;
  assign n24535 = ~n24532 & n24534;
  assign n24536 = pi0626 & ~n24493;
  assign n24537 = ~pi0626 & ~n24381;
  assign n24538 = n16628 & ~n24537;
  assign n24539 = ~n24536 & n24538;
  assign n24540 = ~n24531 & ~n24535;
  assign n24541 = ~n24539 & n24540;
  assign n24542 = pi0788 & ~n24541;
  assign n24543 = pi0609 & n24407;
  assign n24544 = ~pi0176 & ~n19488;
  assign n24545 = pi0176 & n19496;
  assign n24546 = ~pi0742 & ~n24544;
  assign n24547 = ~n24545 & n24546;
  assign n24548 = ~pi0176 & n19477;
  assign n24549 = ~n19468 & ~n19470;
  assign n24550 = pi0176 & ~n24549;
  assign n24551 = pi0742 & ~n24550;
  assign n24552 = ~n24548 & n24551;
  assign n24553 = ~pi0704 & ~n24547;
  assign n24554 = ~n24552 & n24553;
  assign n24555 = pi0704 & n24452;
  assign n24556 = n2571 & ~n24554;
  assign n24557 = ~n24555 & n24556;
  assign n24558 = ~n24445 & ~n24557;
  assign n24559 = ~pi0625 & n24558;
  assign n24560 = pi0625 & n24454;
  assign n24561 = ~pi1153 & ~n24560;
  assign n24562 = ~n24559 & n24561;
  assign n24563 = ~pi0608 & ~n24400;
  assign n24564 = ~n24562 & n24563;
  assign n24565 = ~pi0625 & n24454;
  assign n24566 = pi0625 & n24558;
  assign n24567 = pi1153 & ~n24565;
  assign n24568 = ~n24566 & n24567;
  assign n24569 = pi0608 & ~n24404;
  assign n24570 = ~n24568 & n24569;
  assign n24571 = ~n24564 & ~n24570;
  assign n24572 = pi0778 & ~n24571;
  assign n24573 = ~pi0778 & n24558;
  assign n24574 = ~n24572 & ~n24573;
  assign n24575 = ~pi0609 & ~n24574;
  assign n24576 = ~pi1155 & ~n24543;
  assign n24577 = ~n24575 & n24576;
  assign n24578 = ~pi0660 & ~n24462;
  assign n24579 = ~n24577 & n24578;
  assign n24580 = ~pi0609 & n24407;
  assign n24581 = pi0609 & ~n24574;
  assign n24582 = pi1155 & ~n24580;
  assign n24583 = ~n24581 & n24582;
  assign n24584 = pi0660 & ~n24466;
  assign n24585 = ~n24583 & n24584;
  assign n24586 = ~n24579 & ~n24585;
  assign n24587 = pi0785 & ~n24586;
  assign n24588 = ~pi0785 & ~n24574;
  assign n24589 = ~n24587 & ~n24588;
  assign n24590 = ~pi0618 & ~n24589;
  assign n24591 = pi0618 & n24410;
  assign n24592 = ~pi1154 & ~n24591;
  assign n24593 = ~n24590 & n24592;
  assign n24594 = ~pi0627 & ~n24474;
  assign n24595 = ~n24593 & n24594;
  assign n24596 = ~pi0618 & n24410;
  assign n24597 = pi0618 & ~n24589;
  assign n24598 = pi1154 & ~n24596;
  assign n24599 = ~n24597 & n24598;
  assign n24600 = pi0627 & ~n24478;
  assign n24601 = ~n24599 & n24600;
  assign n24602 = ~n24595 & ~n24601;
  assign n24603 = pi0781 & ~n24602;
  assign n24604 = ~pi0781 & ~n24589;
  assign n24605 = ~n24603 & ~n24604;
  assign n24606 = ~pi0789 & n24605;
  assign n24607 = pi0619 & ~n24413;
  assign n24608 = ~pi0619 & ~n24605;
  assign n24609 = ~pi1159 & ~n24607;
  assign n24610 = ~n24608 & n24609;
  assign n24611 = ~pi0648 & ~n24486;
  assign n24612 = ~n24610 & n24611;
  assign n24613 = pi0619 & ~n24605;
  assign n24614 = ~pi0619 & ~n24413;
  assign n24615 = pi1159 & ~n24614;
  assign n24616 = ~n24613 & n24615;
  assign n24617 = pi0648 & ~n24490;
  assign n24618 = ~n24616 & n24617;
  assign n24619 = pi0789 & ~n24612;
  assign n24620 = ~n24618 & n24619;
  assign n24621 = n17970 & ~n24606;
  assign n24622 = ~n24620 & n24621;
  assign n24623 = ~n24542 & ~n24622;
  assign n24624 = ~n24530 & ~n24623;
  assign n24625 = n20364 & n24529;
  assign n24626 = ~n20206 & ~n24625;
  assign n24627 = ~n24624 & n24626;
  assign n24628 = ~pi0644 & n24515;
  assign n24629 = pi0644 & n24507;
  assign n24630 = pi0790 & ~n24628;
  assign n24631 = ~n24629 & n24630;
  assign n24632 = ~n24524 & ~n24627;
  assign n24633 = ~n24631 & n24632;
  assign n24634 = ~n24518 & ~n24633;
  assign n24635 = ~po1038 & ~n24634;
  assign n24636 = ~pi0832 & ~n24380;
  assign n24637 = ~n24635 & n24636;
  assign po0333 = ~n24379 & ~n24637;
  assign n24639 = ~pi0177 & ~n17059;
  assign n24640 = n16635 & ~n24639;
  assign n24641 = pi0177 & ~n2571;
  assign n24642 = ~pi0177 & n18072;
  assign n24643 = pi0177 & ~n18076;
  assign n24644 = ~pi0038 & ~n24643;
  assign n24645 = ~n24642 & n24644;
  assign n24646 = ~pi0177 & ~n16641;
  assign n24647 = n16647 & ~n24646;
  assign n24648 = ~pi0686 & ~n24647;
  assign n24649 = ~n24645 & n24648;
  assign n24650 = ~pi0177 & pi0686;
  assign n24651 = ~n17052 & n24650;
  assign n24652 = n2571 & ~n24651;
  assign n24653 = ~n24649 & n24652;
  assign n24654 = ~n24641 & ~n24653;
  assign n24655 = ~pi0778 & ~n24654;
  assign n24656 = ~pi0625 & n24639;
  assign n24657 = pi0625 & n24654;
  assign n24658 = pi1153 & ~n24656;
  assign n24659 = ~n24657 & n24658;
  assign n24660 = ~pi0625 & n24654;
  assign n24661 = pi0625 & n24639;
  assign n24662 = ~pi1153 & ~n24661;
  assign n24663 = ~n24660 & n24662;
  assign n24664 = ~n24659 & ~n24663;
  assign n24665 = pi0778 & ~n24664;
  assign n24666 = ~n24655 & ~n24665;
  assign n24667 = ~n17075 & ~n24666;
  assign n24668 = n17075 & ~n24639;
  assign n24669 = ~n24667 & ~n24668;
  assign n24670 = ~n16639 & n24669;
  assign n24671 = n16639 & n24639;
  assign n24672 = ~n24670 & ~n24671;
  assign n24673 = ~n16635 & n24672;
  assign n24674 = ~n24640 & ~n24673;
  assign n24675 = ~n16631 & n24674;
  assign n24676 = n16631 & n24639;
  assign n24677 = ~n24675 & ~n24676;
  assign n24678 = ~pi0792 & n24677;
  assign n24679 = ~pi0628 & n24639;
  assign n24680 = pi0628 & ~n24677;
  assign n24681 = pi1156 & ~n24679;
  assign n24682 = ~n24680 & n24681;
  assign n24683 = pi0628 & n24639;
  assign n24684 = ~pi0628 & ~n24677;
  assign n24685 = ~pi1156 & ~n24683;
  assign n24686 = ~n24684 & n24685;
  assign n24687 = ~n24682 & ~n24686;
  assign n24688 = pi0792 & ~n24687;
  assign n24689 = ~n24678 & ~n24688;
  assign n24690 = ~pi0787 & ~n24689;
  assign n24691 = ~pi0647 & n24639;
  assign n24692 = pi0647 & n24689;
  assign n24693 = pi1157 & ~n24691;
  assign n24694 = ~n24692 & n24693;
  assign n24695 = ~pi0647 & n24689;
  assign n24696 = pi0647 & n24639;
  assign n24697 = ~pi1157 & ~n24696;
  assign n24698 = ~n24695 & n24697;
  assign n24699 = ~n24694 & ~n24698;
  assign n24700 = pi0787 & ~n24699;
  assign n24701 = ~n24690 & ~n24700;
  assign n24702 = ~pi0644 & n24701;
  assign n24703 = ~pi0619 & n24639;
  assign n24704 = ~pi0757 & ~n19439;
  assign n24705 = ~n21646 & ~n24704;
  assign n24706 = ~pi0177 & ~n24705;
  assign n24707 = ~pi0177 & ~n19433;
  assign n24708 = ~pi0757 & ~n24707;
  assign n24709 = ~n24447 & n24708;
  assign n24710 = ~n24706 & ~n24709;
  assign n24711 = n2571 & n24710;
  assign n24712 = ~n24641 & ~n24711;
  assign n24713 = ~n17117 & ~n24712;
  assign n24714 = n17117 & ~n24639;
  assign n24715 = ~n24713 & ~n24714;
  assign n24716 = ~pi0785 & ~n24715;
  assign n24717 = ~n17291 & ~n24639;
  assign n24718 = pi0609 & n24713;
  assign n24719 = ~n24717 & ~n24718;
  assign n24720 = pi1155 & ~n24719;
  assign n24721 = ~n17296 & ~n24639;
  assign n24722 = ~pi0609 & n24713;
  assign n24723 = ~n24721 & ~n24722;
  assign n24724 = ~pi1155 & ~n24723;
  assign n24725 = ~n24720 & ~n24724;
  assign n24726 = pi0785 & ~n24725;
  assign n24727 = ~n24716 & ~n24726;
  assign n24728 = ~pi0781 & ~n24727;
  assign n24729 = ~pi0618 & n24639;
  assign n24730 = pi0618 & n24727;
  assign n24731 = pi1154 & ~n24729;
  assign n24732 = ~n24730 & n24731;
  assign n24733 = ~pi0618 & n24727;
  assign n24734 = pi0618 & n24639;
  assign n24735 = ~pi1154 & ~n24734;
  assign n24736 = ~n24733 & n24735;
  assign n24737 = ~n24732 & ~n24736;
  assign n24738 = pi0781 & ~n24737;
  assign n24739 = ~n24728 & ~n24738;
  assign n24740 = pi0619 & n24739;
  assign n24741 = pi1159 & ~n24703;
  assign n24742 = ~n24740 & n24741;
  assign n24743 = n18176 & ~n24646;
  assign n24744 = ~pi0177 & n19475;
  assign n24745 = pi0177 & n19467;
  assign n24746 = ~pi0038 & ~n24745;
  assign n24747 = ~n24744 & n24746;
  assign n24748 = pi0757 & ~n24743;
  assign n24749 = ~n24747 & n24748;
  assign n24750 = ~pi0177 & ~n19485;
  assign n24751 = pi0177 & n19490;
  assign n24752 = pi0038 & ~n24751;
  assign n24753 = ~n24750 & n24752;
  assign n24754 = ~n19482 & ~n19484;
  assign n24755 = ~pi0177 & ~n24754;
  assign n24756 = pi0177 & n19494;
  assign n24757 = ~pi0038 & ~n24755;
  assign n24758 = ~n24756 & n24757;
  assign n24759 = ~pi0757 & ~n24753;
  assign n24760 = ~n24758 & n24759;
  assign n24761 = ~n24749 & ~n24760;
  assign n24762 = ~pi0686 & ~n24761;
  assign n24763 = pi0686 & ~n24710;
  assign n24764 = n2571 & ~n24762;
  assign n24765 = ~n24763 & n24764;
  assign n24766 = ~n24641 & ~n24765;
  assign n24767 = ~pi0625 & n24766;
  assign n24768 = pi0625 & n24712;
  assign n24769 = ~pi1153 & ~n24768;
  assign n24770 = ~n24767 & n24769;
  assign n24771 = ~pi0608 & ~n24659;
  assign n24772 = ~n24770 & n24771;
  assign n24773 = ~pi0625 & n24712;
  assign n24774 = pi0625 & n24766;
  assign n24775 = pi1153 & ~n24773;
  assign n24776 = ~n24774 & n24775;
  assign n24777 = pi0608 & ~n24663;
  assign n24778 = ~n24776 & n24777;
  assign n24779 = ~n24772 & ~n24778;
  assign n24780 = pi0778 & ~n24779;
  assign n24781 = ~pi0778 & n24766;
  assign n24782 = ~n24780 & ~n24781;
  assign n24783 = ~pi0609 & ~n24782;
  assign n24784 = pi0609 & n24666;
  assign n24785 = ~pi1155 & ~n24784;
  assign n24786 = ~n24783 & n24785;
  assign n24787 = ~pi0660 & ~n24720;
  assign n24788 = ~n24786 & n24787;
  assign n24789 = ~pi0609 & n24666;
  assign n24790 = pi0609 & ~n24782;
  assign n24791 = pi1155 & ~n24789;
  assign n24792 = ~n24790 & n24791;
  assign n24793 = pi0660 & ~n24724;
  assign n24794 = ~n24792 & n24793;
  assign n24795 = ~n24788 & ~n24794;
  assign n24796 = pi0785 & ~n24795;
  assign n24797 = ~pi0785 & ~n24782;
  assign n24798 = ~n24796 & ~n24797;
  assign n24799 = ~pi0618 & ~n24798;
  assign n24800 = pi0618 & n24669;
  assign n24801 = ~pi1154 & ~n24800;
  assign n24802 = ~n24799 & n24801;
  assign n24803 = ~pi0627 & ~n24732;
  assign n24804 = ~n24802 & n24803;
  assign n24805 = ~pi0618 & n24669;
  assign n24806 = pi0618 & ~n24798;
  assign n24807 = pi1154 & ~n24805;
  assign n24808 = ~n24806 & n24807;
  assign n24809 = pi0627 & ~n24736;
  assign n24810 = ~n24808 & n24809;
  assign n24811 = ~n24804 & ~n24810;
  assign n24812 = pi0781 & ~n24811;
  assign n24813 = ~pi0781 & ~n24798;
  assign n24814 = ~n24812 & ~n24813;
  assign n24815 = ~pi0619 & ~n24814;
  assign n24816 = pi0619 & ~n24672;
  assign n24817 = ~pi1159 & ~n24816;
  assign n24818 = ~n24815 & n24817;
  assign n24819 = ~pi0648 & ~n24742;
  assign n24820 = ~n24818 & n24819;
  assign n24821 = ~pi0619 & n24739;
  assign n24822 = pi0619 & n24639;
  assign n24823 = ~pi1159 & ~n24822;
  assign n24824 = ~n24821 & n24823;
  assign n24825 = pi0619 & ~n24814;
  assign n24826 = ~pi0619 & ~n24672;
  assign n24827 = pi1159 & ~n24826;
  assign n24828 = ~n24825 & n24827;
  assign n24829 = pi0648 & ~n24824;
  assign n24830 = ~n24828 & n24829;
  assign n24831 = ~n24820 & ~n24830;
  assign n24832 = pi0789 & ~n24831;
  assign n24833 = ~pi0789 & ~n24814;
  assign n24834 = ~n24832 & ~n24833;
  assign n24835 = ~pi0788 & n24834;
  assign n24836 = ~pi0626 & n24834;
  assign n24837 = pi0626 & ~n24674;
  assign n24838 = ~pi0641 & ~n24837;
  assign n24839 = ~n24836 & n24838;
  assign n24840 = ~pi0789 & ~n24739;
  assign n24841 = ~n24742 & ~n24824;
  assign n24842 = pi0789 & ~n24841;
  assign n24843 = ~n24840 & ~n24842;
  assign n24844 = ~pi0626 & ~n24843;
  assign n24845 = pi0626 & ~n24639;
  assign n24846 = pi0641 & ~n24845;
  assign n24847 = ~n24844 & n24846;
  assign n24848 = ~pi1158 & ~n24847;
  assign n24849 = ~n24839 & n24848;
  assign n24850 = pi0626 & n24834;
  assign n24851 = ~pi0626 & ~n24674;
  assign n24852 = pi0641 & ~n24851;
  assign n24853 = ~n24850 & n24852;
  assign n24854 = pi0626 & ~n24843;
  assign n24855 = ~pi0626 & ~n24639;
  assign n24856 = ~pi0641 & ~n24855;
  assign n24857 = ~n24854 & n24856;
  assign n24858 = pi1158 & ~n24857;
  assign n24859 = ~n24853 & n24858;
  assign n24860 = ~n24849 & ~n24859;
  assign n24861 = pi0788 & ~n24860;
  assign n24862 = ~n24835 & ~n24861;
  assign n24863 = ~pi0628 & n24862;
  assign n24864 = ~n17969 & n24843;
  assign n24865 = n17969 & n24639;
  assign n24866 = ~n24864 & ~n24865;
  assign n24867 = pi0628 & ~n24866;
  assign n24868 = ~pi1156 & ~n24867;
  assign n24869 = ~n24863 & n24868;
  assign n24870 = ~pi0629 & ~n24682;
  assign n24871 = ~n24869 & n24870;
  assign n24872 = pi0628 & n24862;
  assign n24873 = ~pi0628 & ~n24866;
  assign n24874 = pi1156 & ~n24873;
  assign n24875 = ~n24872 & n24874;
  assign n24876 = pi0629 & ~n24686;
  assign n24877 = ~n24875 & n24876;
  assign n24878 = ~n24871 & ~n24877;
  assign n24879 = pi0792 & ~n24878;
  assign n24880 = ~pi0792 & n24862;
  assign n24881 = ~n24879 & ~n24880;
  assign n24882 = ~pi0647 & ~n24881;
  assign n24883 = ~n17779 & ~n24866;
  assign n24884 = n17779 & n24639;
  assign n24885 = ~n24883 & ~n24884;
  assign n24886 = pi0647 & ~n24885;
  assign n24887 = ~pi1157 & ~n24886;
  assign n24888 = ~n24882 & n24887;
  assign n24889 = ~pi0630 & ~n24694;
  assign n24890 = ~n24888 & n24889;
  assign n24891 = pi0647 & ~n24881;
  assign n24892 = ~pi0647 & ~n24885;
  assign n24893 = pi1157 & ~n24892;
  assign n24894 = ~n24891 & n24893;
  assign n24895 = pi0630 & ~n24698;
  assign n24896 = ~n24894 & n24895;
  assign n24897 = ~n24890 & ~n24896;
  assign n24898 = pi0787 & ~n24897;
  assign n24899 = ~pi0787 & ~n24881;
  assign n24900 = ~n24898 & ~n24899;
  assign n24901 = pi0644 & ~n24900;
  assign n24902 = pi0715 & ~n24702;
  assign n24903 = ~n24901 & n24902;
  assign n24904 = n17804 & ~n24639;
  assign n24905 = ~n17804 & n24885;
  assign n24906 = ~n24904 & ~n24905;
  assign n24907 = pi0644 & n24906;
  assign n24908 = ~pi0644 & n24639;
  assign n24909 = ~pi0715 & ~n24908;
  assign n24910 = ~n24907 & n24909;
  assign n24911 = pi1160 & ~n24910;
  assign n24912 = ~n24903 & n24911;
  assign n24913 = ~pi0644 & ~n24900;
  assign n24914 = pi0644 & n24701;
  assign n24915 = ~pi0715 & ~n24914;
  assign n24916 = ~n24913 & n24915;
  assign n24917 = ~pi0644 & n24906;
  assign n24918 = pi0644 & n24639;
  assign n24919 = pi0715 & ~n24918;
  assign n24920 = ~n24917 & n24919;
  assign n24921 = ~pi1160 & ~n24920;
  assign n24922 = ~n24916 & n24921;
  assign n24923 = pi0790 & ~n24912;
  assign n24924 = ~n24922 & n24923;
  assign n24925 = ~pi0790 & n24900;
  assign n24926 = ~po1038 & ~n24925;
  assign n24927 = ~n24924 & n24926;
  assign n24928 = ~pi0177 & po1038;
  assign n24929 = ~pi0832 & ~n24928;
  assign n24930 = ~n24927 & n24929;
  assign n24931 = ~pi0177 & ~n2926;
  assign n24932 = ~pi0686 & n16645;
  assign n24933 = ~n24931 & ~n24932;
  assign n24934 = ~pi0778 & n24933;
  assign n24935 = ~pi0625 & n24932;
  assign n24936 = ~n24933 & ~n24935;
  assign n24937 = pi1153 & ~n24936;
  assign n24938 = ~pi1153 & ~n24931;
  assign n24939 = ~n24935 & n24938;
  assign n24940 = ~n24937 & ~n24939;
  assign n24941 = pi0778 & ~n24940;
  assign n24942 = ~n24934 & ~n24941;
  assign n24943 = ~n17845 & n24942;
  assign n24944 = ~n17847 & n24943;
  assign n24945 = ~n17849 & n24944;
  assign n24946 = ~n17851 & n24945;
  assign n24947 = ~n17857 & n24946;
  assign n24948 = ~pi0647 & n24947;
  assign n24949 = pi0647 & n24931;
  assign n24950 = ~pi1157 & ~n24949;
  assign n24951 = ~n24948 & n24950;
  assign n24952 = pi0630 & n24951;
  assign n24953 = ~pi0757 & n17244;
  assign n24954 = ~n24931 & ~n24953;
  assign n24955 = ~n17874 & ~n24954;
  assign n24956 = ~pi0785 & ~n24955;
  assign n24957 = ~n17879 & ~n24954;
  assign n24958 = pi1155 & ~n24957;
  assign n24959 = ~n17882 & n24955;
  assign n24960 = ~pi1155 & ~n24959;
  assign n24961 = ~n24958 & ~n24960;
  assign n24962 = pi0785 & ~n24961;
  assign n24963 = ~n24956 & ~n24962;
  assign n24964 = ~pi0781 & ~n24963;
  assign n24965 = ~n17889 & n24963;
  assign n24966 = pi1154 & ~n24965;
  assign n24967 = ~n17892 & n24963;
  assign n24968 = ~pi1154 & ~n24967;
  assign n24969 = ~n24966 & ~n24968;
  assign n24970 = pi0781 & ~n24969;
  assign n24971 = ~n24964 & ~n24970;
  assign n24972 = ~pi0789 & ~n24971;
  assign n24973 = ~pi0619 & n24931;
  assign n24974 = pi0619 & n24971;
  assign n24975 = pi1159 & ~n24973;
  assign n24976 = ~n24974 & n24975;
  assign n24977 = ~pi0619 & n24971;
  assign n24978 = pi0619 & n24931;
  assign n24979 = ~pi1159 & ~n24978;
  assign n24980 = ~n24977 & n24979;
  assign n24981 = ~n24976 & ~n24980;
  assign n24982 = pi0789 & ~n24981;
  assign n24983 = ~n24972 & ~n24982;
  assign n24984 = ~n17969 & n24983;
  assign n24985 = n17969 & n24931;
  assign n24986 = ~n24984 & ~n24985;
  assign n24987 = ~n17779 & ~n24986;
  assign n24988 = n17779 & n24931;
  assign n24989 = ~n24987 & ~n24988;
  assign n24990 = ~n20559 & n24989;
  assign n24991 = pi0647 & ~n24947;
  assign n24992 = ~pi0647 & ~n24931;
  assign n24993 = ~n24991 & ~n24992;
  assign n24994 = n17801 & ~n24993;
  assign n24995 = ~n24952 & ~n24994;
  assign n24996 = ~n24990 & n24995;
  assign n24997 = pi0787 & ~n24996;
  assign n24998 = n17871 & n24945;
  assign n24999 = ~pi0626 & ~n24983;
  assign n25000 = pi0626 & ~n24931;
  assign n25001 = n16629 & ~n25000;
  assign n25002 = ~n24999 & n25001;
  assign n25003 = pi0626 & ~n24983;
  assign n25004 = ~pi0626 & ~n24931;
  assign n25005 = n16628 & ~n25004;
  assign n25006 = ~n25003 & n25005;
  assign n25007 = ~n24998 & ~n25002;
  assign n25008 = ~n25006 & n25007;
  assign n25009 = pi0788 & ~n25008;
  assign n25010 = pi0618 & n24943;
  assign n25011 = pi0609 & n24942;
  assign n25012 = ~n17168 & ~n24933;
  assign n25013 = pi0625 & n25012;
  assign n25014 = n24954 & ~n25012;
  assign n25015 = ~n25013 & ~n25014;
  assign n25016 = n24938 & ~n25015;
  assign n25017 = ~pi0608 & ~n24937;
  assign n25018 = ~n25016 & n25017;
  assign n25019 = pi1153 & n24954;
  assign n25020 = ~n25013 & n25019;
  assign n25021 = pi0608 & ~n24939;
  assign n25022 = ~n25020 & n25021;
  assign n25023 = ~n25018 & ~n25022;
  assign n25024 = pi0778 & ~n25023;
  assign n25025 = ~pi0778 & ~n25014;
  assign n25026 = ~n25024 & ~n25025;
  assign n25027 = ~pi0609 & ~n25026;
  assign n25028 = ~pi1155 & ~n25011;
  assign n25029 = ~n25027 & n25028;
  assign n25030 = ~pi0660 & ~n24958;
  assign n25031 = ~n25029 & n25030;
  assign n25032 = ~pi0609 & n24942;
  assign n25033 = pi0609 & ~n25026;
  assign n25034 = pi1155 & ~n25032;
  assign n25035 = ~n25033 & n25034;
  assign n25036 = pi0660 & ~n24960;
  assign n25037 = ~n25035 & n25036;
  assign n25038 = ~n25031 & ~n25037;
  assign n25039 = pi0785 & ~n25038;
  assign n25040 = ~pi0785 & ~n25026;
  assign n25041 = ~n25039 & ~n25040;
  assign n25042 = ~pi0618 & ~n25041;
  assign n25043 = ~pi1154 & ~n25010;
  assign n25044 = ~n25042 & n25043;
  assign n25045 = ~pi0627 & ~n24966;
  assign n25046 = ~n25044 & n25045;
  assign n25047 = ~pi0618 & n24943;
  assign n25048 = pi0618 & ~n25041;
  assign n25049 = pi1154 & ~n25047;
  assign n25050 = ~n25048 & n25049;
  assign n25051 = pi0627 & ~n24968;
  assign n25052 = ~n25050 & n25051;
  assign n25053 = ~n25046 & ~n25052;
  assign n25054 = pi0781 & ~n25053;
  assign n25055 = ~pi0781 & ~n25041;
  assign n25056 = ~n25054 & ~n25055;
  assign n25057 = ~pi0789 & n25056;
  assign n25058 = ~pi0619 & ~n25056;
  assign n25059 = pi0619 & n24944;
  assign n25060 = ~pi1159 & ~n25059;
  assign n25061 = ~n25058 & n25060;
  assign n25062 = ~pi0648 & ~n24976;
  assign n25063 = ~n25061 & n25062;
  assign n25064 = pi0619 & ~n25056;
  assign n25065 = ~pi0619 & n24944;
  assign n25066 = pi1159 & ~n25065;
  assign n25067 = ~n25064 & n25066;
  assign n25068 = pi0648 & ~n24980;
  assign n25069 = ~n25067 & n25068;
  assign n25070 = pi0789 & ~n25063;
  assign n25071 = ~n25069 & n25070;
  assign n25072 = n17970 & ~n25057;
  assign n25073 = ~n25071 & n25072;
  assign n25074 = ~n25009 & ~n25073;
  assign n25075 = ~n20364 & ~n25074;
  assign n25076 = n17854 & ~n24986;
  assign n25077 = n20851 & n24946;
  assign n25078 = ~n25076 & ~n25077;
  assign n25079 = ~pi0629 & ~n25078;
  assign n25080 = n20855 & n24946;
  assign n25081 = n17853 & ~n24986;
  assign n25082 = ~n25080 & ~n25081;
  assign n25083 = pi0629 & ~n25082;
  assign n25084 = ~n25079 & ~n25083;
  assign n25085 = pi0792 & ~n25084;
  assign n25086 = ~n20206 & ~n25085;
  assign n25087 = ~n25075 & n25086;
  assign n25088 = ~n24997 & ~n25087;
  assign n25089 = ~pi0790 & n25088;
  assign n25090 = ~pi0787 & ~n24947;
  assign n25091 = pi1157 & ~n24993;
  assign n25092 = ~n24951 & ~n25091;
  assign n25093 = pi0787 & ~n25092;
  assign n25094 = ~n25090 & ~n25093;
  assign n25095 = ~pi0644 & n25094;
  assign n25096 = pi0644 & n25088;
  assign n25097 = pi0715 & ~n25095;
  assign n25098 = ~n25096 & n25097;
  assign n25099 = ~n17804 & ~n24989;
  assign n25100 = n17804 & n24931;
  assign n25101 = ~n25099 & ~n25100;
  assign n25102 = pi0644 & ~n25101;
  assign n25103 = ~pi0644 & n24931;
  assign n25104 = ~pi0715 & ~n25103;
  assign n25105 = ~n25102 & n25104;
  assign n25106 = pi1160 & ~n25105;
  assign n25107 = ~n25098 & n25106;
  assign n25108 = ~pi0644 & ~n25101;
  assign n25109 = pi0644 & n24931;
  assign n25110 = pi0715 & ~n25109;
  assign n25111 = ~n25108 & n25110;
  assign n25112 = pi0644 & n25094;
  assign n25113 = ~pi0644 & n25088;
  assign n25114 = ~pi0715 & ~n25112;
  assign n25115 = ~n25113 & n25114;
  assign n25116 = ~pi1160 & ~n25111;
  assign n25117 = ~n25115 & n25116;
  assign n25118 = ~n25107 & ~n25117;
  assign n25119 = pi0790 & ~n25118;
  assign n25120 = pi0832 & ~n25089;
  assign n25121 = ~n25119 & n25120;
  assign po0334 = ~n24930 & ~n25121;
  assign n25123 = ~pi0178 & ~n2926;
  assign n25124 = ~pi0688 & n16645;
  assign n25125 = ~n25123 & ~n25124;
  assign n25126 = ~pi0778 & ~n25125;
  assign n25127 = ~pi0625 & n25124;
  assign n25128 = ~n25125 & ~n25127;
  assign n25129 = pi1153 & ~n25128;
  assign n25130 = ~pi1153 & ~n25123;
  assign n25131 = ~n25127 & n25130;
  assign n25132 = pi0778 & ~n25131;
  assign n25133 = ~n25129 & n25132;
  assign n25134 = ~n25126 & ~n25133;
  assign n25135 = ~n17845 & ~n25134;
  assign n25136 = ~n17847 & n25135;
  assign n25137 = ~n17849 & n25136;
  assign n25138 = ~n17851 & n25137;
  assign n25139 = ~n17857 & n25138;
  assign n25140 = ~pi0647 & n25139;
  assign n25141 = pi0647 & n25123;
  assign n25142 = ~pi1157 & ~n25141;
  assign n25143 = ~n25140 & n25142;
  assign n25144 = pi0630 & n25143;
  assign n25145 = ~pi0760 & n17244;
  assign n25146 = ~n25123 & ~n25145;
  assign n25147 = ~n17874 & ~n25146;
  assign n25148 = ~pi0785 & ~n25147;
  assign n25149 = n17296 & n25145;
  assign n25150 = n25147 & ~n25149;
  assign n25151 = pi1155 & ~n25150;
  assign n25152 = ~pi1155 & ~n25123;
  assign n25153 = ~n25149 & n25152;
  assign n25154 = ~n25151 & ~n25153;
  assign n25155 = pi0785 & ~n25154;
  assign n25156 = ~n25148 & ~n25155;
  assign n25157 = ~pi0781 & ~n25156;
  assign n25158 = ~n17889 & n25156;
  assign n25159 = pi1154 & ~n25158;
  assign n25160 = ~n17892 & n25156;
  assign n25161 = ~pi1154 & ~n25160;
  assign n25162 = ~n25159 & ~n25161;
  assign n25163 = pi0781 & ~n25162;
  assign n25164 = ~n25157 & ~n25163;
  assign n25165 = ~pi0789 & ~n25164;
  assign n25166 = ~n23078 & n25164;
  assign n25167 = pi1159 & ~n25166;
  assign n25168 = ~n23081 & n25164;
  assign n25169 = ~pi1159 & ~n25168;
  assign n25170 = ~n25167 & ~n25169;
  assign n25171 = pi0789 & ~n25170;
  assign n25172 = ~n25165 & ~n25171;
  assign n25173 = ~n17969 & n25172;
  assign n25174 = n17969 & n25123;
  assign n25175 = ~n25173 & ~n25174;
  assign n25176 = ~n17779 & ~n25175;
  assign n25177 = n17779 & n25123;
  assign n25178 = ~n25176 & ~n25177;
  assign n25179 = ~n20559 & n25178;
  assign n25180 = pi0647 & ~n25139;
  assign n25181 = ~pi0647 & ~n25123;
  assign n25182 = ~n25180 & ~n25181;
  assign n25183 = n17801 & ~n25182;
  assign n25184 = ~n25144 & ~n25183;
  assign n25185 = ~n25179 & n25184;
  assign n25186 = pi0787 & ~n25185;
  assign n25187 = n17871 & n25137;
  assign n25188 = ~pi0626 & ~n25172;
  assign n25189 = pi0626 & ~n25123;
  assign n25190 = n16629 & ~n25189;
  assign n25191 = ~n25188 & n25190;
  assign n25192 = pi0626 & ~n25172;
  assign n25193 = ~pi0626 & ~n25123;
  assign n25194 = n16628 & ~n25193;
  assign n25195 = ~n25192 & n25194;
  assign n25196 = ~n25187 & ~n25191;
  assign n25197 = ~n25195 & n25196;
  assign n25198 = pi0788 & ~n25197;
  assign n25199 = pi0618 & n25135;
  assign n25200 = ~n17168 & ~n25125;
  assign n25201 = pi0625 & n25200;
  assign n25202 = n25146 & ~n25200;
  assign n25203 = ~n25201 & ~n25202;
  assign n25204 = n25130 & ~n25203;
  assign n25205 = ~pi0608 & ~n25129;
  assign n25206 = ~n25204 & n25205;
  assign n25207 = pi1153 & n25146;
  assign n25208 = ~n25201 & n25207;
  assign n25209 = pi0608 & ~n25131;
  assign n25210 = ~n25208 & n25209;
  assign n25211 = ~n25206 & ~n25210;
  assign n25212 = pi0778 & ~n25211;
  assign n25213 = ~pi0778 & ~n25202;
  assign n25214 = ~n25212 & ~n25213;
  assign n25215 = ~pi0609 & ~n25214;
  assign n25216 = pi0609 & ~n25134;
  assign n25217 = ~pi1155 & ~n25216;
  assign n25218 = ~n25215 & n25217;
  assign n25219 = ~pi0660 & ~n25151;
  assign n25220 = ~n25218 & n25219;
  assign n25221 = pi0609 & ~n25214;
  assign n25222 = ~pi0609 & ~n25134;
  assign n25223 = pi1155 & ~n25222;
  assign n25224 = ~n25221 & n25223;
  assign n25225 = pi0660 & ~n25153;
  assign n25226 = ~n25224 & n25225;
  assign n25227 = ~n25220 & ~n25226;
  assign n25228 = pi0785 & ~n25227;
  assign n25229 = ~pi0785 & ~n25214;
  assign n25230 = ~n25228 & ~n25229;
  assign n25231 = ~pi0618 & ~n25230;
  assign n25232 = ~pi1154 & ~n25199;
  assign n25233 = ~n25231 & n25232;
  assign n25234 = ~pi0627 & ~n25159;
  assign n25235 = ~n25233 & n25234;
  assign n25236 = ~pi0618 & n25135;
  assign n25237 = pi0618 & ~n25230;
  assign n25238 = pi1154 & ~n25236;
  assign n25239 = ~n25237 & n25238;
  assign n25240 = pi0627 & ~n25161;
  assign n25241 = ~n25239 & n25240;
  assign n25242 = ~n25235 & ~n25241;
  assign n25243 = pi0781 & ~n25242;
  assign n25244 = ~pi0781 & ~n25230;
  assign n25245 = ~n25243 & ~n25244;
  assign n25246 = ~pi0789 & n25245;
  assign n25247 = ~pi0619 & ~n25245;
  assign n25248 = pi0619 & n25136;
  assign n25249 = ~pi1159 & ~n25248;
  assign n25250 = ~n25247 & n25249;
  assign n25251 = ~pi0648 & ~n25167;
  assign n25252 = ~n25250 & n25251;
  assign n25253 = pi0619 & ~n25245;
  assign n25254 = ~pi0619 & n25136;
  assign n25255 = pi1159 & ~n25254;
  assign n25256 = ~n25253 & n25255;
  assign n25257 = pi0648 & ~n25169;
  assign n25258 = ~n25256 & n25257;
  assign n25259 = pi0789 & ~n25252;
  assign n25260 = ~n25258 & n25259;
  assign n25261 = n17970 & ~n25246;
  assign n25262 = ~n25260 & n25261;
  assign n25263 = ~n25198 & ~n25262;
  assign n25264 = ~n20364 & ~n25263;
  assign n25265 = n17854 & ~n25175;
  assign n25266 = n20851 & n25138;
  assign n25267 = ~n25265 & ~n25266;
  assign n25268 = ~pi0629 & ~n25267;
  assign n25269 = n20855 & n25138;
  assign n25270 = n17853 & ~n25175;
  assign n25271 = ~n25269 & ~n25270;
  assign n25272 = pi0629 & ~n25271;
  assign n25273 = ~n25268 & ~n25272;
  assign n25274 = pi0792 & ~n25273;
  assign n25275 = ~n20206 & ~n25274;
  assign n25276 = ~n25264 & n25275;
  assign n25277 = ~n25186 & ~n25276;
  assign n25278 = ~pi0790 & n25277;
  assign n25279 = ~pi0787 & ~n25139;
  assign n25280 = pi1157 & ~n25182;
  assign n25281 = ~n25143 & ~n25280;
  assign n25282 = pi0787 & ~n25281;
  assign n25283 = ~n25279 & ~n25282;
  assign n25284 = ~pi0644 & n25283;
  assign n25285 = pi0644 & n25277;
  assign n25286 = pi0715 & ~n25284;
  assign n25287 = ~n25285 & n25286;
  assign n25288 = ~n17804 & ~n25178;
  assign n25289 = n17804 & n25123;
  assign n25290 = ~n25288 & ~n25289;
  assign n25291 = pi0644 & ~n25290;
  assign n25292 = ~pi0644 & n25123;
  assign n25293 = ~pi0715 & ~n25292;
  assign n25294 = ~n25291 & n25293;
  assign n25295 = pi1160 & ~n25294;
  assign n25296 = ~n25287 & n25295;
  assign n25297 = ~pi0644 & ~n25290;
  assign n25298 = pi0644 & n25123;
  assign n25299 = pi0715 & ~n25298;
  assign n25300 = ~n25297 & n25299;
  assign n25301 = pi0644 & n25283;
  assign n25302 = ~pi0644 & n25277;
  assign n25303 = ~pi0715 & ~n25301;
  assign n25304 = ~n25302 & n25303;
  assign n25305 = ~pi1160 & ~n25300;
  assign n25306 = ~n25304 & n25305;
  assign n25307 = ~n25296 & ~n25306;
  assign n25308 = pi0790 & ~n25307;
  assign n25309 = pi0832 & ~n25278;
  assign n25310 = ~n25308 & n25309;
  assign n25311 = ~pi0178 & po1038;
  assign n25312 = ~pi0178 & ~n17059;
  assign n25313 = n16635 & ~n25312;
  assign n25314 = ~pi0688 & n2571;
  assign n25315 = n25312 & ~n25314;
  assign n25316 = ~pi0178 & ~n16641;
  assign n25317 = n16647 & ~n25316;
  assign n25318 = pi0178 & ~n18076;
  assign n25319 = ~pi0038 & ~n25318;
  assign n25320 = n2571 & ~n25319;
  assign n25321 = ~pi0178 & n18072;
  assign n25322 = ~n25320 & ~n25321;
  assign n25323 = ~pi0688 & ~n25317;
  assign n25324 = ~n25322 & n25323;
  assign n25325 = ~n25315 & ~n25324;
  assign n25326 = ~pi0778 & n25325;
  assign n25327 = ~pi0625 & n25312;
  assign n25328 = pi0625 & ~n25325;
  assign n25329 = pi1153 & ~n25327;
  assign n25330 = ~n25328 & n25329;
  assign n25331 = pi0625 & n25312;
  assign n25332 = ~pi0625 & ~n25325;
  assign n25333 = ~pi1153 & ~n25331;
  assign n25334 = ~n25332 & n25333;
  assign n25335 = ~n25330 & ~n25334;
  assign n25336 = pi0778 & ~n25335;
  assign n25337 = ~n25326 & ~n25336;
  assign n25338 = ~n17075 & ~n25337;
  assign n25339 = n17075 & ~n25312;
  assign n25340 = ~n25338 & ~n25339;
  assign n25341 = ~n16639 & n25340;
  assign n25342 = n16639 & n25312;
  assign n25343 = ~n25341 & ~n25342;
  assign n25344 = ~n16635 & n25343;
  assign n25345 = ~n25313 & ~n25344;
  assign n25346 = ~n16631 & n25345;
  assign n25347 = n16631 & n25312;
  assign n25348 = ~n25346 & ~n25347;
  assign n25349 = ~pi0792 & n25348;
  assign n25350 = pi0628 & ~n25348;
  assign n25351 = ~pi0628 & n25312;
  assign n25352 = pi1156 & ~n25351;
  assign n25353 = ~n25350 & n25352;
  assign n25354 = pi0628 & n25312;
  assign n25355 = ~pi0628 & ~n25348;
  assign n25356 = ~pi1156 & ~n25354;
  assign n25357 = ~n25355 & n25356;
  assign n25358 = ~n25353 & ~n25357;
  assign n25359 = pi0792 & ~n25358;
  assign n25360 = ~n25349 & ~n25359;
  assign n25361 = ~pi0647 & ~n25360;
  assign n25362 = pi0647 & ~n25312;
  assign n25363 = ~n25361 & ~n25362;
  assign n25364 = ~pi1157 & n25363;
  assign n25365 = pi0647 & ~n25360;
  assign n25366 = ~pi0647 & ~n25312;
  assign n25367 = ~n25365 & ~n25366;
  assign n25368 = pi1157 & n25367;
  assign n25369 = ~n25364 & ~n25368;
  assign n25370 = pi0787 & ~n25369;
  assign n25371 = ~pi0787 & n25360;
  assign n25372 = ~n25370 & ~n25371;
  assign n25373 = ~pi0644 & ~n25372;
  assign n25374 = pi0715 & ~n25373;
  assign n25375 = pi0178 & ~n2571;
  assign n25376 = ~pi0760 & n17280;
  assign n25377 = ~n25316 & ~n25376;
  assign n25378 = pi0038 & ~n25377;
  assign n25379 = ~pi0178 & n17221;
  assign n25380 = pi0178 & ~n17275;
  assign n25381 = ~pi0760 & ~n25380;
  assign n25382 = ~n25379 & n25381;
  assign n25383 = ~pi0178 & pi0760;
  assign n25384 = ~n17048 & n25383;
  assign n25385 = ~n25382 & ~n25384;
  assign n25386 = ~pi0038 & ~n25385;
  assign n25387 = ~n25378 & ~n25386;
  assign n25388 = n2571 & n25387;
  assign n25389 = ~n25375 & ~n25388;
  assign n25390 = ~n17117 & ~n25389;
  assign n25391 = n17117 & ~n25312;
  assign n25392 = ~n25390 & ~n25391;
  assign n25393 = ~pi0785 & ~n25392;
  assign n25394 = ~n17291 & ~n25312;
  assign n25395 = pi0609 & n25390;
  assign n25396 = ~n25394 & ~n25395;
  assign n25397 = pi1155 & ~n25396;
  assign n25398 = ~n17296 & ~n25312;
  assign n25399 = ~pi0609 & n25390;
  assign n25400 = ~n25398 & ~n25399;
  assign n25401 = ~pi1155 & ~n25400;
  assign n25402 = ~n25397 & ~n25401;
  assign n25403 = pi0785 & ~n25402;
  assign n25404 = ~n25393 & ~n25403;
  assign n25405 = ~pi0781 & ~n25404;
  assign n25406 = ~pi0618 & n25312;
  assign n25407 = pi0618 & n25404;
  assign n25408 = pi1154 & ~n25406;
  assign n25409 = ~n25407 & n25408;
  assign n25410 = ~pi0618 & n25404;
  assign n25411 = pi0618 & n25312;
  assign n25412 = ~pi1154 & ~n25411;
  assign n25413 = ~n25410 & n25412;
  assign n25414 = ~n25409 & ~n25413;
  assign n25415 = pi0781 & ~n25414;
  assign n25416 = ~n25405 & ~n25415;
  assign n25417 = ~pi0789 & ~n25416;
  assign n25418 = ~pi0619 & n25312;
  assign n25419 = pi0619 & n25416;
  assign n25420 = pi1159 & ~n25418;
  assign n25421 = ~n25419 & n25420;
  assign n25422 = ~pi0619 & n25416;
  assign n25423 = pi0619 & n25312;
  assign n25424 = ~pi1159 & ~n25423;
  assign n25425 = ~n25422 & n25424;
  assign n25426 = ~n25421 & ~n25425;
  assign n25427 = pi0789 & ~n25426;
  assign n25428 = ~n25417 & ~n25427;
  assign n25429 = ~n17969 & n25428;
  assign n25430 = n17969 & n25312;
  assign n25431 = ~n25429 & ~n25430;
  assign n25432 = ~n17779 & ~n25431;
  assign n25433 = n17779 & n25312;
  assign n25434 = ~n25432 & ~n25433;
  assign n25435 = ~n17804 & ~n25434;
  assign n25436 = n17804 & n25312;
  assign n25437 = ~n25435 & ~n25436;
  assign n25438 = pi0644 & ~n25437;
  assign n25439 = ~pi0644 & n25312;
  assign n25440 = ~pi0715 & ~n25439;
  assign n25441 = ~n25438 & n25440;
  assign n25442 = pi1160 & ~n25441;
  assign n25443 = ~n25374 & n25442;
  assign n25444 = pi0644 & ~n25372;
  assign n25445 = ~pi0715 & ~n25444;
  assign n25446 = ~pi0644 & ~n25437;
  assign n25447 = pi0644 & n25312;
  assign n25448 = pi0715 & ~n25447;
  assign n25449 = ~n25446 & n25448;
  assign n25450 = ~pi1160 & ~n25449;
  assign n25451 = ~n25445 & n25450;
  assign n25452 = ~n25443 & ~n25451;
  assign n25453 = pi0790 & ~n25452;
  assign n25454 = ~pi0629 & n25353;
  assign n25455 = ~n20570 & n25431;
  assign n25456 = pi0629 & n25357;
  assign n25457 = ~n25454 & ~n25456;
  assign n25458 = ~n25455 & n25457;
  assign n25459 = pi0792 & ~n25458;
  assign n25460 = pi0609 & n25337;
  assign n25461 = pi0178 & ~n17625;
  assign n25462 = ~pi0178 & ~n17612;
  assign n25463 = pi0760 & ~n25461;
  assign n25464 = ~n25462 & n25463;
  assign n25465 = ~pi0178 & n17629;
  assign n25466 = pi0178 & n17631;
  assign n25467 = ~pi0760 & ~n25466;
  assign n25468 = ~n25465 & n25467;
  assign n25469 = ~n25464 & ~n25468;
  assign n25470 = ~pi0039 & ~n25469;
  assign n25471 = pi0178 & n17605;
  assign n25472 = ~pi0178 & ~n17546;
  assign n25473 = ~pi0760 & ~n25472;
  assign n25474 = ~n25471 & n25473;
  assign n25475 = ~pi0178 & n17404;
  assign n25476 = pi0178 & n17485;
  assign n25477 = pi0760 & ~n25476;
  assign n25478 = ~n25475 & n25477;
  assign n25479 = pi0039 & ~n25474;
  assign n25480 = ~n25478 & n25479;
  assign n25481 = ~pi0038 & ~n25470;
  assign n25482 = ~n25480 & n25481;
  assign n25483 = ~pi0760 & ~n17490;
  assign n25484 = n19471 & ~n25483;
  assign n25485 = ~pi0178 & ~n25484;
  assign n25486 = ~n17469 & ~n25145;
  assign n25487 = pi0178 & ~n25486;
  assign n25488 = n6284 & n25487;
  assign n25489 = pi0038 & ~n25488;
  assign n25490 = ~n25485 & n25489;
  assign n25491 = ~pi0688 & ~n25490;
  assign n25492 = ~n25482 & n25491;
  assign n25493 = pi0688 & ~n25387;
  assign n25494 = n2571 & ~n25492;
  assign n25495 = ~n25493 & n25494;
  assign n25496 = ~n25375 & ~n25495;
  assign n25497 = ~pi0625 & n25496;
  assign n25498 = pi0625 & n25389;
  assign n25499 = ~pi1153 & ~n25498;
  assign n25500 = ~n25497 & n25499;
  assign n25501 = ~pi0608 & ~n25330;
  assign n25502 = ~n25500 & n25501;
  assign n25503 = ~pi0625 & n25389;
  assign n25504 = pi0625 & n25496;
  assign n25505 = pi1153 & ~n25503;
  assign n25506 = ~n25504 & n25505;
  assign n25507 = pi0608 & ~n25334;
  assign n25508 = ~n25506 & n25507;
  assign n25509 = ~n25502 & ~n25508;
  assign n25510 = pi0778 & ~n25509;
  assign n25511 = ~pi0778 & n25496;
  assign n25512 = ~n25510 & ~n25511;
  assign n25513 = ~pi0609 & ~n25512;
  assign n25514 = ~pi1155 & ~n25460;
  assign n25515 = ~n25513 & n25514;
  assign n25516 = ~pi0660 & ~n25397;
  assign n25517 = ~n25515 & n25516;
  assign n25518 = ~pi0609 & n25337;
  assign n25519 = pi0609 & ~n25512;
  assign n25520 = pi1155 & ~n25518;
  assign n25521 = ~n25519 & n25520;
  assign n25522 = pi0660 & ~n25401;
  assign n25523 = ~n25521 & n25522;
  assign n25524 = ~n25517 & ~n25523;
  assign n25525 = pi0785 & ~n25524;
  assign n25526 = ~pi0785 & ~n25512;
  assign n25527 = ~n25525 & ~n25526;
  assign n25528 = ~pi0618 & ~n25527;
  assign n25529 = pi0618 & n25340;
  assign n25530 = ~pi1154 & ~n25529;
  assign n25531 = ~n25528 & n25530;
  assign n25532 = ~pi0627 & ~n25409;
  assign n25533 = ~n25531 & n25532;
  assign n25534 = ~pi0618 & n25340;
  assign n25535 = pi0618 & ~n25527;
  assign n25536 = pi1154 & ~n25534;
  assign n25537 = ~n25535 & n25536;
  assign n25538 = pi0627 & ~n25413;
  assign n25539 = ~n25537 & n25538;
  assign n25540 = ~n25533 & ~n25539;
  assign n25541 = pi0781 & ~n25540;
  assign n25542 = ~pi0781 & ~n25527;
  assign n25543 = ~n25541 & ~n25542;
  assign n25544 = ~pi0789 & n25543;
  assign n25545 = pi0619 & ~n25343;
  assign n25546 = ~pi0619 & ~n25543;
  assign n25547 = ~pi1159 & ~n25545;
  assign n25548 = ~n25546 & n25547;
  assign n25549 = ~pi0648 & ~n25421;
  assign n25550 = ~n25548 & n25549;
  assign n25551 = ~pi0619 & ~n25343;
  assign n25552 = pi0619 & ~n25543;
  assign n25553 = pi1159 & ~n25551;
  assign n25554 = ~n25552 & n25553;
  assign n25555 = pi0648 & ~n25425;
  assign n25556 = ~n25554 & n25555;
  assign n25557 = pi0789 & ~n25550;
  assign n25558 = ~n25556 & n25557;
  assign n25559 = n17970 & ~n25544;
  assign n25560 = ~n25558 & n25559;
  assign n25561 = n17871 & n25345;
  assign n25562 = ~pi0626 & ~n25428;
  assign n25563 = pi0626 & ~n25312;
  assign n25564 = n16629 & ~n25563;
  assign n25565 = ~n25562 & n25564;
  assign n25566 = pi0626 & ~n25428;
  assign n25567 = ~pi0626 & ~n25312;
  assign n25568 = n16628 & ~n25567;
  assign n25569 = ~n25566 & n25568;
  assign n25570 = ~n25561 & ~n25565;
  assign n25571 = ~n25569 & n25570;
  assign n25572 = pi0788 & ~n25571;
  assign n25573 = ~n20364 & ~n25572;
  assign n25574 = ~n25560 & n25573;
  assign n25575 = ~n25459 & ~n25574;
  assign n25576 = ~n20206 & ~n25575;
  assign n25577 = n17802 & ~n25363;
  assign n25578 = ~n20559 & n25434;
  assign n25579 = n17801 & ~n25367;
  assign n25580 = ~n25577 & ~n25579;
  assign n25581 = ~n25578 & n25580;
  assign n25582 = pi0787 & ~n25581;
  assign n25583 = ~pi0644 & n25450;
  assign n25584 = pi0644 & n25442;
  assign n25585 = pi0790 & ~n25583;
  assign n25586 = ~n25584 & n25585;
  assign n25587 = ~n25576 & ~n25582;
  assign n25588 = ~n25586 & n25587;
  assign n25589 = ~n25453 & ~n25588;
  assign n25590 = ~po1038 & ~n25589;
  assign n25591 = ~pi0832 & ~n25311;
  assign n25592 = ~n25590 & n25591;
  assign po0335 = ~n25310 & ~n25592;
  assign n25594 = ~pi0179 & ~n17059;
  assign n25595 = n16635 & ~n25594;
  assign n25596 = ~pi0724 & n2571;
  assign n25597 = n25594 & ~n25596;
  assign n25598 = ~pi0179 & ~n16641;
  assign n25599 = n16647 & ~n25598;
  assign n25600 = ~pi0179 & n18072;
  assign n25601 = pi0179 & ~n18076;
  assign n25602 = ~pi0038 & ~n25601;
  assign n25603 = n2571 & ~n25602;
  assign n25604 = ~n25600 & ~n25603;
  assign n25605 = ~pi0724 & ~n25599;
  assign n25606 = ~n25604 & n25605;
  assign n25607 = ~n25597 & ~n25606;
  assign n25608 = ~pi0778 & n25607;
  assign n25609 = ~pi0625 & n25594;
  assign n25610 = pi0625 & ~n25607;
  assign n25611 = pi1153 & ~n25609;
  assign n25612 = ~n25610 & n25611;
  assign n25613 = pi0625 & n25594;
  assign n25614 = ~pi0625 & ~n25607;
  assign n25615 = ~pi1153 & ~n25613;
  assign n25616 = ~n25614 & n25615;
  assign n25617 = ~n25612 & ~n25616;
  assign n25618 = pi0778 & ~n25617;
  assign n25619 = ~n25608 & ~n25618;
  assign n25620 = ~n17075 & ~n25619;
  assign n25621 = n17075 & ~n25594;
  assign n25622 = ~n25620 & ~n25621;
  assign n25623 = ~n16639 & n25622;
  assign n25624 = n16639 & n25594;
  assign n25625 = ~n25623 & ~n25624;
  assign n25626 = ~n16635 & n25625;
  assign n25627 = ~n25595 & ~n25626;
  assign n25628 = ~n16631 & n25627;
  assign n25629 = n16631 & n25594;
  assign n25630 = ~n25628 & ~n25629;
  assign n25631 = ~pi0792 & n25630;
  assign n25632 = ~pi0628 & n25594;
  assign n25633 = pi0628 & ~n25630;
  assign n25634 = pi1156 & ~n25632;
  assign n25635 = ~n25633 & n25634;
  assign n25636 = pi0628 & n25594;
  assign n25637 = ~pi0628 & ~n25630;
  assign n25638 = ~pi1156 & ~n25636;
  assign n25639 = ~n25637 & n25638;
  assign n25640 = ~n25635 & ~n25639;
  assign n25641 = pi0792 & ~n25640;
  assign n25642 = ~n25631 & ~n25641;
  assign n25643 = ~pi0787 & ~n25642;
  assign n25644 = ~pi0647 & n25594;
  assign n25645 = pi0647 & n25642;
  assign n25646 = pi1157 & ~n25644;
  assign n25647 = ~n25645 & n25646;
  assign n25648 = ~pi0647 & n25642;
  assign n25649 = pi0647 & n25594;
  assign n25650 = ~pi1157 & ~n25649;
  assign n25651 = ~n25648 & n25650;
  assign n25652 = ~n25647 & ~n25651;
  assign n25653 = pi0787 & ~n25652;
  assign n25654 = ~n25643 & ~n25653;
  assign n25655 = ~pi0644 & n25654;
  assign n25656 = ~pi0618 & n25594;
  assign n25657 = pi0179 & ~n2571;
  assign n25658 = ~pi0741 & ~n24447;
  assign n25659 = pi0179 & ~n25658;
  assign n25660 = ~pi0179 & ~pi0741;
  assign n25661 = ~n19433 & n25660;
  assign n25662 = n19439 & n25661;
  assign n25663 = ~n25659 & ~n25662;
  assign n25664 = ~n21674 & n25663;
  assign n25665 = n2571 & ~n25664;
  assign n25666 = ~n25657 & ~n25665;
  assign n25667 = ~n17117 & ~n25666;
  assign n25668 = n17117 & ~n25594;
  assign n25669 = ~n25667 & ~n25668;
  assign n25670 = ~pi0785 & ~n25669;
  assign n25671 = ~n17291 & ~n25594;
  assign n25672 = pi0609 & n25667;
  assign n25673 = ~n25671 & ~n25672;
  assign n25674 = pi1155 & ~n25673;
  assign n25675 = ~n17296 & ~n25594;
  assign n25676 = ~pi0609 & n25667;
  assign n25677 = ~n25675 & ~n25676;
  assign n25678 = ~pi1155 & ~n25677;
  assign n25679 = ~n25674 & ~n25678;
  assign n25680 = pi0785 & ~n25679;
  assign n25681 = ~n25670 & ~n25680;
  assign n25682 = pi0618 & n25681;
  assign n25683 = pi1154 & ~n25656;
  assign n25684 = ~n25682 & n25683;
  assign n25685 = n18176 & ~n25598;
  assign n25686 = ~pi0179 & n17404;
  assign n25687 = pi0179 & n17485;
  assign n25688 = pi0039 & ~n25687;
  assign n25689 = ~n25686 & n25688;
  assign n25690 = ~pi0179 & n17612;
  assign n25691 = pi0179 & n17625;
  assign n25692 = ~pi0039 & ~n25690;
  assign n25693 = ~n25691 & n25692;
  assign n25694 = ~n25689 & ~n25693;
  assign n25695 = ~pi0038 & ~n25694;
  assign n25696 = ~n25685 & ~n25695;
  assign n25697 = pi0741 & ~n25696;
  assign n25698 = ~pi0179 & ~n19488;
  assign n25699 = pi0179 & n19496;
  assign n25700 = ~pi0741 & ~n25698;
  assign n25701 = ~n25699 & n25700;
  assign n25702 = ~pi0724 & ~n25701;
  assign n25703 = ~n25697 & n25702;
  assign n25704 = pi0724 & n25664;
  assign n25705 = n2571 & ~n25704;
  assign n25706 = ~n25703 & n25705;
  assign n25707 = ~n25657 & ~n25706;
  assign n25708 = ~pi0625 & n25707;
  assign n25709 = pi0625 & n25666;
  assign n25710 = ~pi1153 & ~n25709;
  assign n25711 = ~n25708 & n25710;
  assign n25712 = ~pi0608 & ~n25612;
  assign n25713 = ~n25711 & n25712;
  assign n25714 = ~pi0625 & n25666;
  assign n25715 = pi0625 & n25707;
  assign n25716 = pi1153 & ~n25714;
  assign n25717 = ~n25715 & n25716;
  assign n25718 = pi0608 & ~n25616;
  assign n25719 = ~n25717 & n25718;
  assign n25720 = ~n25713 & ~n25719;
  assign n25721 = pi0778 & ~n25720;
  assign n25722 = ~pi0778 & n25707;
  assign n25723 = ~n25721 & ~n25722;
  assign n25724 = ~pi0609 & ~n25723;
  assign n25725 = pi0609 & n25619;
  assign n25726 = ~pi1155 & ~n25725;
  assign n25727 = ~n25724 & n25726;
  assign n25728 = ~pi0660 & ~n25674;
  assign n25729 = ~n25727 & n25728;
  assign n25730 = ~pi0609 & n25619;
  assign n25731 = pi0609 & ~n25723;
  assign n25732 = pi1155 & ~n25730;
  assign n25733 = ~n25731 & n25732;
  assign n25734 = pi0660 & ~n25678;
  assign n25735 = ~n25733 & n25734;
  assign n25736 = ~n25729 & ~n25735;
  assign n25737 = pi0785 & ~n25736;
  assign n25738 = ~pi0785 & ~n25723;
  assign n25739 = ~n25737 & ~n25738;
  assign n25740 = ~pi0618 & ~n25739;
  assign n25741 = pi0618 & n25622;
  assign n25742 = ~pi1154 & ~n25741;
  assign n25743 = ~n25740 & n25742;
  assign n25744 = ~pi0627 & ~n25684;
  assign n25745 = ~n25743 & n25744;
  assign n25746 = ~pi0618 & n25681;
  assign n25747 = pi0618 & n25594;
  assign n25748 = ~pi1154 & ~n25747;
  assign n25749 = ~n25746 & n25748;
  assign n25750 = ~pi0618 & n25622;
  assign n25751 = pi0618 & ~n25739;
  assign n25752 = pi1154 & ~n25750;
  assign n25753 = ~n25751 & n25752;
  assign n25754 = pi0627 & ~n25749;
  assign n25755 = ~n25753 & n25754;
  assign n25756 = ~n25745 & ~n25755;
  assign n25757 = pi0781 & ~n25756;
  assign n25758 = ~pi0781 & ~n25739;
  assign n25759 = ~n25757 & ~n25758;
  assign n25760 = ~pi0619 & ~n25759;
  assign n25761 = pi0619 & ~n25625;
  assign n25762 = ~pi1159 & ~n25761;
  assign n25763 = ~n25760 & n25762;
  assign n25764 = ~pi0619 & n25594;
  assign n25765 = ~pi0781 & ~n25681;
  assign n25766 = ~n25684 & ~n25749;
  assign n25767 = pi0781 & ~n25766;
  assign n25768 = ~n25765 & ~n25767;
  assign n25769 = pi0619 & n25768;
  assign n25770 = pi1159 & ~n25764;
  assign n25771 = ~n25769 & n25770;
  assign n25772 = ~pi0648 & ~n25771;
  assign n25773 = ~n25763 & n25772;
  assign n25774 = pi0619 & ~n25759;
  assign n25775 = ~pi0619 & ~n25625;
  assign n25776 = pi1159 & ~n25775;
  assign n25777 = ~n25774 & n25776;
  assign n25778 = ~pi0619 & n25768;
  assign n25779 = pi0619 & n25594;
  assign n25780 = ~pi1159 & ~n25779;
  assign n25781 = ~n25778 & n25780;
  assign n25782 = pi0648 & ~n25781;
  assign n25783 = ~n25777 & n25782;
  assign n25784 = ~n25773 & ~n25783;
  assign n25785 = pi0789 & ~n25784;
  assign n25786 = ~pi0789 & ~n25759;
  assign n25787 = ~n25785 & ~n25786;
  assign n25788 = ~pi0788 & n25787;
  assign n25789 = ~pi0626 & n25787;
  assign n25790 = pi0626 & ~n25627;
  assign n25791 = ~pi0641 & ~n25790;
  assign n25792 = ~n25789 & n25791;
  assign n25793 = ~pi0789 & ~n25768;
  assign n25794 = ~n25771 & ~n25781;
  assign n25795 = pi0789 & ~n25794;
  assign n25796 = ~n25793 & ~n25795;
  assign n25797 = ~pi0626 & ~n25796;
  assign n25798 = pi0626 & ~n25594;
  assign n25799 = pi0641 & ~n25798;
  assign n25800 = ~n25797 & n25799;
  assign n25801 = ~pi1158 & ~n25800;
  assign n25802 = ~n25792 & n25801;
  assign n25803 = pi0626 & n25787;
  assign n25804 = ~pi0626 & ~n25627;
  assign n25805 = pi0641 & ~n25804;
  assign n25806 = ~n25803 & n25805;
  assign n25807 = pi0626 & ~n25796;
  assign n25808 = ~pi0626 & ~n25594;
  assign n25809 = ~pi0641 & ~n25808;
  assign n25810 = ~n25807 & n25809;
  assign n25811 = pi1158 & ~n25810;
  assign n25812 = ~n25806 & n25811;
  assign n25813 = ~n25802 & ~n25812;
  assign n25814 = pi0788 & ~n25813;
  assign n25815 = ~n25788 & ~n25814;
  assign n25816 = ~pi0628 & n25815;
  assign n25817 = ~n17969 & n25796;
  assign n25818 = n17969 & n25594;
  assign n25819 = ~n25817 & ~n25818;
  assign n25820 = pi0628 & ~n25819;
  assign n25821 = ~pi1156 & ~n25820;
  assign n25822 = ~n25816 & n25821;
  assign n25823 = ~pi0629 & ~n25635;
  assign n25824 = ~n25822 & n25823;
  assign n25825 = pi0628 & n25815;
  assign n25826 = ~pi0628 & ~n25819;
  assign n25827 = pi1156 & ~n25826;
  assign n25828 = ~n25825 & n25827;
  assign n25829 = pi0629 & ~n25639;
  assign n25830 = ~n25828 & n25829;
  assign n25831 = ~n25824 & ~n25830;
  assign n25832 = pi0792 & ~n25831;
  assign n25833 = ~pi0792 & n25815;
  assign n25834 = ~n25832 & ~n25833;
  assign n25835 = ~pi0647 & ~n25834;
  assign n25836 = ~n17779 & ~n25819;
  assign n25837 = n17779 & n25594;
  assign n25838 = ~n25836 & ~n25837;
  assign n25839 = pi0647 & ~n25838;
  assign n25840 = ~pi1157 & ~n25839;
  assign n25841 = ~n25835 & n25840;
  assign n25842 = ~pi0630 & ~n25647;
  assign n25843 = ~n25841 & n25842;
  assign n25844 = pi0647 & ~n25834;
  assign n25845 = ~pi0647 & ~n25838;
  assign n25846 = pi1157 & ~n25845;
  assign n25847 = ~n25844 & n25846;
  assign n25848 = pi0630 & ~n25651;
  assign n25849 = ~n25847 & n25848;
  assign n25850 = ~n25843 & ~n25849;
  assign n25851 = pi0787 & ~n25850;
  assign n25852 = ~pi0787 & ~n25834;
  assign n25853 = ~n25851 & ~n25852;
  assign n25854 = pi0644 & ~n25853;
  assign n25855 = pi0715 & ~n25655;
  assign n25856 = ~n25854 & n25855;
  assign n25857 = n17804 & ~n25594;
  assign n25858 = ~n17804 & n25838;
  assign n25859 = ~n25857 & ~n25858;
  assign n25860 = pi0644 & n25859;
  assign n25861 = ~pi0644 & n25594;
  assign n25862 = ~pi0715 & ~n25861;
  assign n25863 = ~n25860 & n25862;
  assign n25864 = pi1160 & ~n25863;
  assign n25865 = ~n25856 & n25864;
  assign n25866 = ~pi0644 & ~n25853;
  assign n25867 = pi0644 & n25654;
  assign n25868 = ~pi0715 & ~n25867;
  assign n25869 = ~n25866 & n25868;
  assign n25870 = ~pi0644 & n25859;
  assign n25871 = pi0644 & n25594;
  assign n25872 = pi0715 & ~n25871;
  assign n25873 = ~n25870 & n25872;
  assign n25874 = ~pi1160 & ~n25873;
  assign n25875 = ~n25869 & n25874;
  assign n25876 = pi0790 & ~n25865;
  assign n25877 = ~n25875 & n25876;
  assign n25878 = ~pi0790 & n25853;
  assign n25879 = ~po1038 & ~n25878;
  assign n25880 = ~n25877 & n25879;
  assign n25881 = ~pi0179 & po1038;
  assign n25882 = ~pi0832 & ~n25881;
  assign n25883 = ~n25880 & n25882;
  assign n25884 = ~pi0179 & ~n2926;
  assign n25885 = ~pi0724 & n16645;
  assign n25886 = ~n25884 & ~n25885;
  assign n25887 = ~pi0778 & n25886;
  assign n25888 = ~pi0625 & n25885;
  assign n25889 = ~n25886 & ~n25888;
  assign n25890 = pi1153 & ~n25889;
  assign n25891 = ~pi1153 & ~n25884;
  assign n25892 = ~n25888 & n25891;
  assign n25893 = ~n25890 & ~n25892;
  assign n25894 = pi0778 & ~n25893;
  assign n25895 = ~n25887 & ~n25894;
  assign n25896 = ~n17845 & n25895;
  assign n25897 = ~n17847 & n25896;
  assign n25898 = ~n17849 & n25897;
  assign n25899 = ~n17851 & n25898;
  assign n25900 = ~n17857 & n25899;
  assign n25901 = ~pi0647 & n25900;
  assign n25902 = pi0647 & n25884;
  assign n25903 = ~pi1157 & ~n25902;
  assign n25904 = ~n25901 & n25903;
  assign n25905 = pi0630 & n25904;
  assign n25906 = ~pi0741 & n17244;
  assign n25907 = ~n25884 & ~n25906;
  assign n25908 = ~n17874 & ~n25907;
  assign n25909 = ~pi0785 & ~n25908;
  assign n25910 = ~n17879 & ~n25907;
  assign n25911 = pi1155 & ~n25910;
  assign n25912 = ~n17882 & n25908;
  assign n25913 = ~pi1155 & ~n25912;
  assign n25914 = ~n25911 & ~n25913;
  assign n25915 = pi0785 & ~n25914;
  assign n25916 = ~n25909 & ~n25915;
  assign n25917 = ~pi0781 & ~n25916;
  assign n25918 = ~n17889 & n25916;
  assign n25919 = pi1154 & ~n25918;
  assign n25920 = ~n17892 & n25916;
  assign n25921 = ~pi1154 & ~n25920;
  assign n25922 = ~n25919 & ~n25921;
  assign n25923 = pi0781 & ~n25922;
  assign n25924 = ~n25917 & ~n25923;
  assign n25925 = ~pi0789 & ~n25924;
  assign n25926 = ~pi0619 & n25884;
  assign n25927 = pi0619 & n25924;
  assign n25928 = pi1159 & ~n25926;
  assign n25929 = ~n25927 & n25928;
  assign n25930 = ~pi0619 & n25924;
  assign n25931 = pi0619 & n25884;
  assign n25932 = ~pi1159 & ~n25931;
  assign n25933 = ~n25930 & n25932;
  assign n25934 = ~n25929 & ~n25933;
  assign n25935 = pi0789 & ~n25934;
  assign n25936 = ~n25925 & ~n25935;
  assign n25937 = ~n17969 & n25936;
  assign n25938 = n17969 & n25884;
  assign n25939 = ~n25937 & ~n25938;
  assign n25940 = ~n17779 & ~n25939;
  assign n25941 = n17779 & n25884;
  assign n25942 = ~n25940 & ~n25941;
  assign n25943 = ~n20559 & n25942;
  assign n25944 = pi0647 & ~n25900;
  assign n25945 = ~pi0647 & ~n25884;
  assign n25946 = ~n25944 & ~n25945;
  assign n25947 = n17801 & ~n25946;
  assign n25948 = ~n25905 & ~n25947;
  assign n25949 = ~n25943 & n25948;
  assign n25950 = pi0787 & ~n25949;
  assign n25951 = n17871 & n25898;
  assign n25952 = ~pi0626 & ~n25936;
  assign n25953 = pi0626 & ~n25884;
  assign n25954 = n16629 & ~n25953;
  assign n25955 = ~n25952 & n25954;
  assign n25956 = pi0626 & ~n25936;
  assign n25957 = ~pi0626 & ~n25884;
  assign n25958 = n16628 & ~n25957;
  assign n25959 = ~n25956 & n25958;
  assign n25960 = ~n25951 & ~n25955;
  assign n25961 = ~n25959 & n25960;
  assign n25962 = pi0788 & ~n25961;
  assign n25963 = pi0618 & n25896;
  assign n25964 = pi0609 & n25895;
  assign n25965 = ~n17168 & ~n25886;
  assign n25966 = pi0625 & n25965;
  assign n25967 = n25907 & ~n25965;
  assign n25968 = ~n25966 & ~n25967;
  assign n25969 = n25891 & ~n25968;
  assign n25970 = ~pi0608 & ~n25890;
  assign n25971 = ~n25969 & n25970;
  assign n25972 = pi1153 & n25907;
  assign n25973 = ~n25966 & n25972;
  assign n25974 = pi0608 & ~n25892;
  assign n25975 = ~n25973 & n25974;
  assign n25976 = ~n25971 & ~n25975;
  assign n25977 = pi0778 & ~n25976;
  assign n25978 = ~pi0778 & ~n25967;
  assign n25979 = ~n25977 & ~n25978;
  assign n25980 = ~pi0609 & ~n25979;
  assign n25981 = ~pi1155 & ~n25964;
  assign n25982 = ~n25980 & n25981;
  assign n25983 = ~pi0660 & ~n25911;
  assign n25984 = ~n25982 & n25983;
  assign n25985 = ~pi0609 & n25895;
  assign n25986 = pi0609 & ~n25979;
  assign n25987 = pi1155 & ~n25985;
  assign n25988 = ~n25986 & n25987;
  assign n25989 = pi0660 & ~n25913;
  assign n25990 = ~n25988 & n25989;
  assign n25991 = ~n25984 & ~n25990;
  assign n25992 = pi0785 & ~n25991;
  assign n25993 = ~pi0785 & ~n25979;
  assign n25994 = ~n25992 & ~n25993;
  assign n25995 = ~pi0618 & ~n25994;
  assign n25996 = ~pi1154 & ~n25963;
  assign n25997 = ~n25995 & n25996;
  assign n25998 = ~pi0627 & ~n25919;
  assign n25999 = ~n25997 & n25998;
  assign n26000 = ~pi0618 & n25896;
  assign n26001 = pi0618 & ~n25994;
  assign n26002 = pi1154 & ~n26000;
  assign n26003 = ~n26001 & n26002;
  assign n26004 = pi0627 & ~n25921;
  assign n26005 = ~n26003 & n26004;
  assign n26006 = ~n25999 & ~n26005;
  assign n26007 = pi0781 & ~n26006;
  assign n26008 = ~pi0781 & ~n25994;
  assign n26009 = ~n26007 & ~n26008;
  assign n26010 = ~pi0789 & n26009;
  assign n26011 = ~pi0619 & ~n26009;
  assign n26012 = pi0619 & n25897;
  assign n26013 = ~pi1159 & ~n26012;
  assign n26014 = ~n26011 & n26013;
  assign n26015 = ~pi0648 & ~n25929;
  assign n26016 = ~n26014 & n26015;
  assign n26017 = pi0619 & ~n26009;
  assign n26018 = ~pi0619 & n25897;
  assign n26019 = pi1159 & ~n26018;
  assign n26020 = ~n26017 & n26019;
  assign n26021 = pi0648 & ~n25933;
  assign n26022 = ~n26020 & n26021;
  assign n26023 = pi0789 & ~n26016;
  assign n26024 = ~n26022 & n26023;
  assign n26025 = n17970 & ~n26010;
  assign n26026 = ~n26024 & n26025;
  assign n26027 = ~n25962 & ~n26026;
  assign n26028 = ~n20364 & ~n26027;
  assign n26029 = n17854 & ~n25939;
  assign n26030 = n20851 & n25899;
  assign n26031 = ~n26029 & ~n26030;
  assign n26032 = ~pi0629 & ~n26031;
  assign n26033 = n20855 & n25899;
  assign n26034 = n17853 & ~n25939;
  assign n26035 = ~n26033 & ~n26034;
  assign n26036 = pi0629 & ~n26035;
  assign n26037 = ~n26032 & ~n26036;
  assign n26038 = pi0792 & ~n26037;
  assign n26039 = ~n20206 & ~n26038;
  assign n26040 = ~n26028 & n26039;
  assign n26041 = ~n25950 & ~n26040;
  assign n26042 = ~pi0790 & n26041;
  assign n26043 = ~pi0787 & ~n25900;
  assign n26044 = pi1157 & ~n25946;
  assign n26045 = ~n25904 & ~n26044;
  assign n26046 = pi0787 & ~n26045;
  assign n26047 = ~n26043 & ~n26046;
  assign n26048 = ~pi0644 & n26047;
  assign n26049 = pi0644 & n26041;
  assign n26050 = pi0715 & ~n26048;
  assign n26051 = ~n26049 & n26050;
  assign n26052 = ~n17804 & ~n25942;
  assign n26053 = n17804 & n25884;
  assign n26054 = ~n26052 & ~n26053;
  assign n26055 = pi0644 & ~n26054;
  assign n26056 = ~pi0644 & n25884;
  assign n26057 = ~pi0715 & ~n26056;
  assign n26058 = ~n26055 & n26057;
  assign n26059 = pi1160 & ~n26058;
  assign n26060 = ~n26051 & n26059;
  assign n26061 = ~pi0644 & ~n26054;
  assign n26062 = pi0644 & n25884;
  assign n26063 = pi0715 & ~n26062;
  assign n26064 = ~n26061 & n26063;
  assign n26065 = pi0644 & n26047;
  assign n26066 = ~pi0644 & n26041;
  assign n26067 = ~pi0715 & ~n26065;
  assign n26068 = ~n26066 & n26067;
  assign n26069 = ~pi1160 & ~n26064;
  assign n26070 = ~n26068 & n26069;
  assign n26071 = ~n26060 & ~n26070;
  assign n26072 = pi0790 & ~n26071;
  assign n26073 = pi0832 & ~n26042;
  assign n26074 = ~n26072 & n26073;
  assign po0336 = ~n25883 & ~n26074;
  assign n26076 = ~pi0180 & ~n2926;
  assign n26077 = ~pi0702 & n16645;
  assign n26078 = ~n26076 & ~n26077;
  assign n26079 = ~pi0778 & ~n26078;
  assign n26080 = ~pi0625 & n26077;
  assign n26081 = ~n26078 & ~n26080;
  assign n26082 = pi1153 & ~n26081;
  assign n26083 = ~pi1153 & ~n26076;
  assign n26084 = ~n26080 & n26083;
  assign n26085 = pi0778 & ~n26084;
  assign n26086 = ~n26082 & n26085;
  assign n26087 = ~n26079 & ~n26086;
  assign n26088 = ~n17845 & ~n26087;
  assign n26089 = ~n17847 & n26088;
  assign n26090 = ~n17849 & n26089;
  assign n26091 = ~n17851 & n26090;
  assign n26092 = ~n17857 & n26091;
  assign n26093 = ~pi0647 & n26092;
  assign n26094 = pi0647 & n26076;
  assign n26095 = ~pi1157 & ~n26094;
  assign n26096 = ~n26093 & n26095;
  assign n26097 = pi0630 & n26096;
  assign n26098 = ~pi0753 & n17244;
  assign n26099 = ~n26076 & ~n26098;
  assign n26100 = ~n17874 & ~n26099;
  assign n26101 = ~pi0785 & ~n26100;
  assign n26102 = n17296 & n26098;
  assign n26103 = n26100 & ~n26102;
  assign n26104 = pi1155 & ~n26103;
  assign n26105 = ~pi1155 & ~n26076;
  assign n26106 = ~n26102 & n26105;
  assign n26107 = ~n26104 & ~n26106;
  assign n26108 = pi0785 & ~n26107;
  assign n26109 = ~n26101 & ~n26108;
  assign n26110 = ~pi0781 & ~n26109;
  assign n26111 = ~n17889 & n26109;
  assign n26112 = pi1154 & ~n26111;
  assign n26113 = ~n17892 & n26109;
  assign n26114 = ~pi1154 & ~n26113;
  assign n26115 = ~n26112 & ~n26114;
  assign n26116 = pi0781 & ~n26115;
  assign n26117 = ~n26110 & ~n26116;
  assign n26118 = ~pi0789 & ~n26117;
  assign n26119 = ~n23078 & n26117;
  assign n26120 = pi1159 & ~n26119;
  assign n26121 = ~n23081 & n26117;
  assign n26122 = ~pi1159 & ~n26121;
  assign n26123 = ~n26120 & ~n26122;
  assign n26124 = pi0789 & ~n26123;
  assign n26125 = ~n26118 & ~n26124;
  assign n26126 = ~n17969 & n26125;
  assign n26127 = n17969 & n26076;
  assign n26128 = ~n26126 & ~n26127;
  assign n26129 = ~n17779 & ~n26128;
  assign n26130 = n17779 & n26076;
  assign n26131 = ~n26129 & ~n26130;
  assign n26132 = ~n20559 & n26131;
  assign n26133 = pi0647 & ~n26092;
  assign n26134 = ~pi0647 & ~n26076;
  assign n26135 = ~n26133 & ~n26134;
  assign n26136 = n17801 & ~n26135;
  assign n26137 = ~n26097 & ~n26136;
  assign n26138 = ~n26132 & n26137;
  assign n26139 = pi0787 & ~n26138;
  assign n26140 = n17871 & n26090;
  assign n26141 = ~pi0626 & ~n26125;
  assign n26142 = pi0626 & ~n26076;
  assign n26143 = n16629 & ~n26142;
  assign n26144 = ~n26141 & n26143;
  assign n26145 = pi0626 & ~n26125;
  assign n26146 = ~pi0626 & ~n26076;
  assign n26147 = n16628 & ~n26146;
  assign n26148 = ~n26145 & n26147;
  assign n26149 = ~n26140 & ~n26144;
  assign n26150 = ~n26148 & n26149;
  assign n26151 = pi0788 & ~n26150;
  assign n26152 = pi0618 & n26088;
  assign n26153 = ~n17168 & ~n26078;
  assign n26154 = pi0625 & n26153;
  assign n26155 = n26099 & ~n26153;
  assign n26156 = ~n26154 & ~n26155;
  assign n26157 = n26083 & ~n26156;
  assign n26158 = ~pi0608 & ~n26082;
  assign n26159 = ~n26157 & n26158;
  assign n26160 = pi1153 & n26099;
  assign n26161 = ~n26154 & n26160;
  assign n26162 = pi0608 & ~n26084;
  assign n26163 = ~n26161 & n26162;
  assign n26164 = ~n26159 & ~n26163;
  assign n26165 = pi0778 & ~n26164;
  assign n26166 = ~pi0778 & ~n26155;
  assign n26167 = ~n26165 & ~n26166;
  assign n26168 = ~pi0609 & ~n26167;
  assign n26169 = pi0609 & ~n26087;
  assign n26170 = ~pi1155 & ~n26169;
  assign n26171 = ~n26168 & n26170;
  assign n26172 = ~pi0660 & ~n26104;
  assign n26173 = ~n26171 & n26172;
  assign n26174 = pi0609 & ~n26167;
  assign n26175 = ~pi0609 & ~n26087;
  assign n26176 = pi1155 & ~n26175;
  assign n26177 = ~n26174 & n26176;
  assign n26178 = pi0660 & ~n26106;
  assign n26179 = ~n26177 & n26178;
  assign n26180 = ~n26173 & ~n26179;
  assign n26181 = pi0785 & ~n26180;
  assign n26182 = ~pi0785 & ~n26167;
  assign n26183 = ~n26181 & ~n26182;
  assign n26184 = ~pi0618 & ~n26183;
  assign n26185 = ~pi1154 & ~n26152;
  assign n26186 = ~n26184 & n26185;
  assign n26187 = ~pi0627 & ~n26112;
  assign n26188 = ~n26186 & n26187;
  assign n26189 = ~pi0618 & n26088;
  assign n26190 = pi0618 & ~n26183;
  assign n26191 = pi1154 & ~n26189;
  assign n26192 = ~n26190 & n26191;
  assign n26193 = pi0627 & ~n26114;
  assign n26194 = ~n26192 & n26193;
  assign n26195 = ~n26188 & ~n26194;
  assign n26196 = pi0781 & ~n26195;
  assign n26197 = ~pi0781 & ~n26183;
  assign n26198 = ~n26196 & ~n26197;
  assign n26199 = ~pi0789 & n26198;
  assign n26200 = ~pi0619 & ~n26198;
  assign n26201 = pi0619 & n26089;
  assign n26202 = ~pi1159 & ~n26201;
  assign n26203 = ~n26200 & n26202;
  assign n26204 = ~pi0648 & ~n26120;
  assign n26205 = ~n26203 & n26204;
  assign n26206 = pi0619 & ~n26198;
  assign n26207 = ~pi0619 & n26089;
  assign n26208 = pi1159 & ~n26207;
  assign n26209 = ~n26206 & n26208;
  assign n26210 = pi0648 & ~n26122;
  assign n26211 = ~n26209 & n26210;
  assign n26212 = pi0789 & ~n26205;
  assign n26213 = ~n26211 & n26212;
  assign n26214 = n17970 & ~n26199;
  assign n26215 = ~n26213 & n26214;
  assign n26216 = ~n26151 & ~n26215;
  assign n26217 = ~n20364 & ~n26216;
  assign n26218 = n17854 & ~n26128;
  assign n26219 = n20851 & n26091;
  assign n26220 = ~n26218 & ~n26219;
  assign n26221 = ~pi0629 & ~n26220;
  assign n26222 = n20855 & n26091;
  assign n26223 = n17853 & ~n26128;
  assign n26224 = ~n26222 & ~n26223;
  assign n26225 = pi0629 & ~n26224;
  assign n26226 = ~n26221 & ~n26225;
  assign n26227 = pi0792 & ~n26226;
  assign n26228 = ~n20206 & ~n26227;
  assign n26229 = ~n26217 & n26228;
  assign n26230 = ~n26139 & ~n26229;
  assign n26231 = ~pi0790 & n26230;
  assign n26232 = ~pi0787 & ~n26092;
  assign n26233 = pi1157 & ~n26135;
  assign n26234 = ~n26096 & ~n26233;
  assign n26235 = pi0787 & ~n26234;
  assign n26236 = ~n26232 & ~n26235;
  assign n26237 = ~pi0644 & n26236;
  assign n26238 = pi0644 & n26230;
  assign n26239 = pi0715 & ~n26237;
  assign n26240 = ~n26238 & n26239;
  assign n26241 = ~n17804 & ~n26131;
  assign n26242 = n17804 & n26076;
  assign n26243 = ~n26241 & ~n26242;
  assign n26244 = pi0644 & ~n26243;
  assign n26245 = ~pi0644 & n26076;
  assign n26246 = ~pi0715 & ~n26245;
  assign n26247 = ~n26244 & n26246;
  assign n26248 = pi1160 & ~n26247;
  assign n26249 = ~n26240 & n26248;
  assign n26250 = ~pi0644 & ~n26243;
  assign n26251 = pi0644 & n26076;
  assign n26252 = pi0715 & ~n26251;
  assign n26253 = ~n26250 & n26252;
  assign n26254 = pi0644 & n26236;
  assign n26255 = ~pi0644 & n26230;
  assign n26256 = ~pi0715 & ~n26254;
  assign n26257 = ~n26255 & n26256;
  assign n26258 = ~pi1160 & ~n26253;
  assign n26259 = ~n26257 & n26258;
  assign n26260 = ~n26249 & ~n26259;
  assign n26261 = pi0790 & ~n26260;
  assign n26262 = pi0832 & ~n26231;
  assign n26263 = ~n26261 & n26262;
  assign n26264 = ~pi0180 & po1038;
  assign n26265 = ~pi0180 & ~n17059;
  assign n26266 = n16635 & ~n26265;
  assign n26267 = ~pi0702 & n2571;
  assign n26268 = n26265 & ~n26267;
  assign n26269 = ~pi0180 & ~n16641;
  assign n26270 = n16647 & ~n26269;
  assign n26271 = pi0180 & ~n18076;
  assign n26272 = ~pi0038 & ~n26271;
  assign n26273 = n2571 & ~n26272;
  assign n26274 = ~pi0180 & n18072;
  assign n26275 = ~n26273 & ~n26274;
  assign n26276 = ~pi0702 & ~n26270;
  assign n26277 = ~n26275 & n26276;
  assign n26278 = ~n26268 & ~n26277;
  assign n26279 = ~pi0778 & n26278;
  assign n26280 = ~pi0625 & n26265;
  assign n26281 = pi0625 & ~n26278;
  assign n26282 = pi1153 & ~n26280;
  assign n26283 = ~n26281 & n26282;
  assign n26284 = pi0625 & n26265;
  assign n26285 = ~pi0625 & ~n26278;
  assign n26286 = ~pi1153 & ~n26284;
  assign n26287 = ~n26285 & n26286;
  assign n26288 = ~n26283 & ~n26287;
  assign n26289 = pi0778 & ~n26288;
  assign n26290 = ~n26279 & ~n26289;
  assign n26291 = ~n17075 & ~n26290;
  assign n26292 = n17075 & ~n26265;
  assign n26293 = ~n26291 & ~n26292;
  assign n26294 = ~n16639 & n26293;
  assign n26295 = n16639 & n26265;
  assign n26296 = ~n26294 & ~n26295;
  assign n26297 = ~n16635 & n26296;
  assign n26298 = ~n26266 & ~n26297;
  assign n26299 = ~n16631 & n26298;
  assign n26300 = n16631 & n26265;
  assign n26301 = ~n26299 & ~n26300;
  assign n26302 = ~pi0792 & n26301;
  assign n26303 = pi0628 & ~n26301;
  assign n26304 = ~pi0628 & n26265;
  assign n26305 = pi1156 & ~n26304;
  assign n26306 = ~n26303 & n26305;
  assign n26307 = pi0628 & n26265;
  assign n26308 = ~pi0628 & ~n26301;
  assign n26309 = ~pi1156 & ~n26307;
  assign n26310 = ~n26308 & n26309;
  assign n26311 = ~n26306 & ~n26310;
  assign n26312 = pi0792 & ~n26311;
  assign n26313 = ~n26302 & ~n26312;
  assign n26314 = ~pi0647 & ~n26313;
  assign n26315 = pi0647 & ~n26265;
  assign n26316 = ~n26314 & ~n26315;
  assign n26317 = ~pi1157 & n26316;
  assign n26318 = pi0647 & ~n26313;
  assign n26319 = ~pi0647 & ~n26265;
  assign n26320 = ~n26318 & ~n26319;
  assign n26321 = pi1157 & n26320;
  assign n26322 = ~n26317 & ~n26321;
  assign n26323 = pi0787 & ~n26322;
  assign n26324 = ~pi0787 & n26313;
  assign n26325 = ~n26323 & ~n26324;
  assign n26326 = ~pi0644 & ~n26325;
  assign n26327 = pi0715 & ~n26326;
  assign n26328 = pi0180 & ~n2571;
  assign n26329 = pi0180 & pi0753;
  assign n26330 = pi0753 & n17046;
  assign n26331 = pi0180 & n17273;
  assign n26332 = ~n26330 & ~n26331;
  assign n26333 = pi0039 & ~n26332;
  assign n26334 = pi0180 & ~n17233;
  assign n26335 = ~n21756 & ~n26334;
  assign n26336 = ~pi0039 & ~n26335;
  assign n26337 = ~pi0180 & ~pi0753;
  assign n26338 = n17221 & n26337;
  assign n26339 = ~n26329 & ~n26336;
  assign n26340 = ~n26338 & n26339;
  assign n26341 = ~n26333 & n26340;
  assign n26342 = ~pi0038 & ~n26341;
  assign n26343 = ~pi0753 & n17280;
  assign n26344 = pi0038 & ~n26269;
  assign n26345 = ~n26343 & n26344;
  assign n26346 = ~n26342 & ~n26345;
  assign n26347 = n2571 & ~n26346;
  assign n26348 = ~n26328 & ~n26347;
  assign n26349 = ~n17117 & ~n26348;
  assign n26350 = n17117 & ~n26265;
  assign n26351 = ~n26349 & ~n26350;
  assign n26352 = ~pi0785 & ~n26351;
  assign n26353 = ~n17291 & ~n26265;
  assign n26354 = pi0609 & n26349;
  assign n26355 = ~n26353 & ~n26354;
  assign n26356 = pi1155 & ~n26355;
  assign n26357 = ~n17296 & ~n26265;
  assign n26358 = ~pi0609 & n26349;
  assign n26359 = ~n26357 & ~n26358;
  assign n26360 = ~pi1155 & ~n26359;
  assign n26361 = ~n26356 & ~n26360;
  assign n26362 = pi0785 & ~n26361;
  assign n26363 = ~n26352 & ~n26362;
  assign n26364 = ~pi0781 & ~n26363;
  assign n26365 = ~pi0618 & n26265;
  assign n26366 = pi0618 & n26363;
  assign n26367 = pi1154 & ~n26365;
  assign n26368 = ~n26366 & n26367;
  assign n26369 = ~pi0618 & n26363;
  assign n26370 = pi0618 & n26265;
  assign n26371 = ~pi1154 & ~n26370;
  assign n26372 = ~n26369 & n26371;
  assign n26373 = ~n26368 & ~n26372;
  assign n26374 = pi0781 & ~n26373;
  assign n26375 = ~n26364 & ~n26374;
  assign n26376 = ~pi0789 & ~n26375;
  assign n26377 = ~pi0619 & n26265;
  assign n26378 = pi0619 & n26375;
  assign n26379 = pi1159 & ~n26377;
  assign n26380 = ~n26378 & n26379;
  assign n26381 = ~pi0619 & n26375;
  assign n26382 = pi0619 & n26265;
  assign n26383 = ~pi1159 & ~n26382;
  assign n26384 = ~n26381 & n26383;
  assign n26385 = ~n26380 & ~n26384;
  assign n26386 = pi0789 & ~n26385;
  assign n26387 = ~n26376 & ~n26386;
  assign n26388 = ~n17969 & n26387;
  assign n26389 = n17969 & n26265;
  assign n26390 = ~n26388 & ~n26389;
  assign n26391 = ~n17779 & ~n26390;
  assign n26392 = n17779 & n26265;
  assign n26393 = ~n26391 & ~n26392;
  assign n26394 = ~n17804 & ~n26393;
  assign n26395 = n17804 & n26265;
  assign n26396 = ~n26394 & ~n26395;
  assign n26397 = pi0644 & ~n26396;
  assign n26398 = ~pi0644 & n26265;
  assign n26399 = ~pi0715 & ~n26398;
  assign n26400 = ~n26397 & n26399;
  assign n26401 = pi1160 & ~n26400;
  assign n26402 = ~n26327 & n26401;
  assign n26403 = pi0644 & ~n26325;
  assign n26404 = ~pi0715 & ~n26403;
  assign n26405 = ~pi0644 & ~n26396;
  assign n26406 = pi0644 & n26265;
  assign n26407 = pi0715 & ~n26406;
  assign n26408 = ~n26405 & n26407;
  assign n26409 = ~pi1160 & ~n26408;
  assign n26410 = ~n26404 & n26409;
  assign n26411 = ~n26402 & ~n26410;
  assign n26412 = pi0790 & ~n26411;
  assign n26413 = ~pi0629 & n26306;
  assign n26414 = ~n20570 & n26390;
  assign n26415 = pi0629 & n26310;
  assign n26416 = ~n26413 & ~n26415;
  assign n26417 = ~n26414 & n26416;
  assign n26418 = pi0792 & ~n26417;
  assign n26419 = pi0609 & n26290;
  assign n26420 = pi0180 & ~n17625;
  assign n26421 = ~pi0180 & ~n17612;
  assign n26422 = pi0753 & ~n26420;
  assign n26423 = ~n26421 & n26422;
  assign n26424 = ~pi0180 & n17629;
  assign n26425 = pi0180 & n17631;
  assign n26426 = ~pi0753 & ~n26425;
  assign n26427 = ~n26424 & n26426;
  assign n26428 = ~n26423 & ~n26427;
  assign n26429 = ~pi0039 & ~n26428;
  assign n26430 = pi0180 & n17605;
  assign n26431 = ~pi0180 & ~n17546;
  assign n26432 = ~pi0753 & ~n26431;
  assign n26433 = ~n26430 & n26432;
  assign n26434 = ~pi0180 & n17404;
  assign n26435 = pi0180 & n17485;
  assign n26436 = pi0753 & ~n26435;
  assign n26437 = ~n26434 & n26436;
  assign n26438 = pi0039 & ~n26433;
  assign n26439 = ~n26437 & n26438;
  assign n26440 = ~pi0038 & ~n26429;
  assign n26441 = ~n26439 & n26440;
  assign n26442 = ~n17469 & ~n26098;
  assign n26443 = pi0180 & ~n26442;
  assign n26444 = n6284 & n26443;
  assign n26445 = ~pi0753 & ~n17490;
  assign n26446 = n19471 & ~n26445;
  assign n26447 = ~pi0180 & ~n26446;
  assign n26448 = pi0038 & ~n26444;
  assign n26449 = ~n26447 & n26448;
  assign n26450 = ~pi0702 & ~n26449;
  assign n26451 = ~n26441 & n26450;
  assign n26452 = pi0702 & n26346;
  assign n26453 = n2571 & ~n26451;
  assign n26454 = ~n26452 & n26453;
  assign n26455 = ~n26328 & ~n26454;
  assign n26456 = ~pi0625 & n26455;
  assign n26457 = pi0625 & n26348;
  assign n26458 = ~pi1153 & ~n26457;
  assign n26459 = ~n26456 & n26458;
  assign n26460 = ~pi0608 & ~n26283;
  assign n26461 = ~n26459 & n26460;
  assign n26462 = ~pi0625 & n26348;
  assign n26463 = pi0625 & n26455;
  assign n26464 = pi1153 & ~n26462;
  assign n26465 = ~n26463 & n26464;
  assign n26466 = pi0608 & ~n26287;
  assign n26467 = ~n26465 & n26466;
  assign n26468 = ~n26461 & ~n26467;
  assign n26469 = pi0778 & ~n26468;
  assign n26470 = ~pi0778 & n26455;
  assign n26471 = ~n26469 & ~n26470;
  assign n26472 = ~pi0609 & ~n26471;
  assign n26473 = ~pi1155 & ~n26419;
  assign n26474 = ~n26472 & n26473;
  assign n26475 = ~pi0660 & ~n26356;
  assign n26476 = ~n26474 & n26475;
  assign n26477 = ~pi0609 & n26290;
  assign n26478 = pi0609 & ~n26471;
  assign n26479 = pi1155 & ~n26477;
  assign n26480 = ~n26478 & n26479;
  assign n26481 = pi0660 & ~n26360;
  assign n26482 = ~n26480 & n26481;
  assign n26483 = ~n26476 & ~n26482;
  assign n26484 = pi0785 & ~n26483;
  assign n26485 = ~pi0785 & ~n26471;
  assign n26486 = ~n26484 & ~n26485;
  assign n26487 = ~pi0618 & ~n26486;
  assign n26488 = pi0618 & n26293;
  assign n26489 = ~pi1154 & ~n26488;
  assign n26490 = ~n26487 & n26489;
  assign n26491 = ~pi0627 & ~n26368;
  assign n26492 = ~n26490 & n26491;
  assign n26493 = ~pi0618 & n26293;
  assign n26494 = pi0618 & ~n26486;
  assign n26495 = pi1154 & ~n26493;
  assign n26496 = ~n26494 & n26495;
  assign n26497 = pi0627 & ~n26372;
  assign n26498 = ~n26496 & n26497;
  assign n26499 = ~n26492 & ~n26498;
  assign n26500 = pi0781 & ~n26499;
  assign n26501 = ~pi0781 & ~n26486;
  assign n26502 = ~n26500 & ~n26501;
  assign n26503 = ~pi0789 & n26502;
  assign n26504 = pi0619 & ~n26296;
  assign n26505 = ~pi0619 & ~n26502;
  assign n26506 = ~pi1159 & ~n26504;
  assign n26507 = ~n26505 & n26506;
  assign n26508 = ~pi0648 & ~n26380;
  assign n26509 = ~n26507 & n26508;
  assign n26510 = ~pi0619 & ~n26296;
  assign n26511 = pi0619 & ~n26502;
  assign n26512 = pi1159 & ~n26510;
  assign n26513 = ~n26511 & n26512;
  assign n26514 = pi0648 & ~n26384;
  assign n26515 = ~n26513 & n26514;
  assign n26516 = pi0789 & ~n26509;
  assign n26517 = ~n26515 & n26516;
  assign n26518 = n17970 & ~n26503;
  assign n26519 = ~n26517 & n26518;
  assign n26520 = n17871 & n26298;
  assign n26521 = ~pi0626 & ~n26387;
  assign n26522 = pi0626 & ~n26265;
  assign n26523 = n16629 & ~n26522;
  assign n26524 = ~n26521 & n26523;
  assign n26525 = pi0626 & ~n26387;
  assign n26526 = ~pi0626 & ~n26265;
  assign n26527 = n16628 & ~n26526;
  assign n26528 = ~n26525 & n26527;
  assign n26529 = ~n26520 & ~n26524;
  assign n26530 = ~n26528 & n26529;
  assign n26531 = pi0788 & ~n26530;
  assign n26532 = ~n20364 & ~n26531;
  assign n26533 = ~n26519 & n26532;
  assign n26534 = ~n26418 & ~n26533;
  assign n26535 = ~n20206 & ~n26534;
  assign n26536 = n17802 & ~n26316;
  assign n26537 = ~n20559 & n26393;
  assign n26538 = n17801 & ~n26320;
  assign n26539 = ~n26536 & ~n26538;
  assign n26540 = ~n26537 & n26539;
  assign n26541 = pi0787 & ~n26540;
  assign n26542 = ~pi0644 & n26409;
  assign n26543 = pi0644 & n26401;
  assign n26544 = pi0790 & ~n26542;
  assign n26545 = ~n26543 & n26544;
  assign n26546 = ~n26535 & ~n26541;
  assign n26547 = ~n26545 & n26546;
  assign n26548 = ~n26412 & ~n26547;
  assign n26549 = ~po1038 & ~n26548;
  assign n26550 = ~pi0832 & ~n26264;
  assign n26551 = ~n26549 & n26550;
  assign po0337 = ~n26263 & ~n26551;
  assign n26553 = ~pi0181 & ~n2926;
  assign n26554 = ~pi0709 & n16645;
  assign n26555 = ~n26553 & ~n26554;
  assign n26556 = ~pi0778 & ~n26555;
  assign n26557 = ~pi0625 & n26554;
  assign n26558 = ~n26555 & ~n26557;
  assign n26559 = pi1153 & ~n26558;
  assign n26560 = ~pi1153 & ~n26553;
  assign n26561 = ~n26557 & n26560;
  assign n26562 = pi0778 & ~n26561;
  assign n26563 = ~n26559 & n26562;
  assign n26564 = ~n26556 & ~n26563;
  assign n26565 = ~n17845 & ~n26564;
  assign n26566 = ~n17847 & n26565;
  assign n26567 = ~n17849 & n26566;
  assign n26568 = ~n17851 & n26567;
  assign n26569 = ~n17857 & n26568;
  assign n26570 = ~pi0647 & n26569;
  assign n26571 = pi0647 & n26553;
  assign n26572 = ~pi1157 & ~n26571;
  assign n26573 = ~n26570 & n26572;
  assign n26574 = pi0630 & n26573;
  assign n26575 = ~pi0754 & n17244;
  assign n26576 = ~n26553 & ~n26575;
  assign n26577 = ~n17874 & ~n26576;
  assign n26578 = ~pi0785 & ~n26577;
  assign n26579 = n17296 & n26575;
  assign n26580 = n26577 & ~n26579;
  assign n26581 = pi1155 & ~n26580;
  assign n26582 = ~pi1155 & ~n26553;
  assign n26583 = ~n26579 & n26582;
  assign n26584 = ~n26581 & ~n26583;
  assign n26585 = pi0785 & ~n26584;
  assign n26586 = ~n26578 & ~n26585;
  assign n26587 = ~pi0781 & ~n26586;
  assign n26588 = ~n17889 & n26586;
  assign n26589 = pi1154 & ~n26588;
  assign n26590 = ~n17892 & n26586;
  assign n26591 = ~pi1154 & ~n26590;
  assign n26592 = ~n26589 & ~n26591;
  assign n26593 = pi0781 & ~n26592;
  assign n26594 = ~n26587 & ~n26593;
  assign n26595 = ~pi0789 & ~n26594;
  assign n26596 = ~n23078 & n26594;
  assign n26597 = pi1159 & ~n26596;
  assign n26598 = ~n23081 & n26594;
  assign n26599 = ~pi1159 & ~n26598;
  assign n26600 = ~n26597 & ~n26599;
  assign n26601 = pi0789 & ~n26600;
  assign n26602 = ~n26595 & ~n26601;
  assign n26603 = ~n17969 & n26602;
  assign n26604 = n17969 & n26553;
  assign n26605 = ~n26603 & ~n26604;
  assign n26606 = ~n17779 & ~n26605;
  assign n26607 = n17779 & n26553;
  assign n26608 = ~n26606 & ~n26607;
  assign n26609 = ~n20559 & n26608;
  assign n26610 = pi0647 & ~n26569;
  assign n26611 = ~pi0647 & ~n26553;
  assign n26612 = ~n26610 & ~n26611;
  assign n26613 = n17801 & ~n26612;
  assign n26614 = ~n26574 & ~n26613;
  assign n26615 = ~n26609 & n26614;
  assign n26616 = pi0787 & ~n26615;
  assign n26617 = n17871 & n26567;
  assign n26618 = ~pi0626 & ~n26602;
  assign n26619 = pi0626 & ~n26553;
  assign n26620 = n16629 & ~n26619;
  assign n26621 = ~n26618 & n26620;
  assign n26622 = pi0626 & ~n26602;
  assign n26623 = ~pi0626 & ~n26553;
  assign n26624 = n16628 & ~n26623;
  assign n26625 = ~n26622 & n26624;
  assign n26626 = ~n26617 & ~n26621;
  assign n26627 = ~n26625 & n26626;
  assign n26628 = pi0788 & ~n26627;
  assign n26629 = pi0618 & n26565;
  assign n26630 = ~n17168 & ~n26555;
  assign n26631 = pi0625 & n26630;
  assign n26632 = n26576 & ~n26630;
  assign n26633 = ~n26631 & ~n26632;
  assign n26634 = n26560 & ~n26633;
  assign n26635 = ~pi0608 & ~n26559;
  assign n26636 = ~n26634 & n26635;
  assign n26637 = pi1153 & n26576;
  assign n26638 = ~n26631 & n26637;
  assign n26639 = pi0608 & ~n26561;
  assign n26640 = ~n26638 & n26639;
  assign n26641 = ~n26636 & ~n26640;
  assign n26642 = pi0778 & ~n26641;
  assign n26643 = ~pi0778 & ~n26632;
  assign n26644 = ~n26642 & ~n26643;
  assign n26645 = ~pi0609 & ~n26644;
  assign n26646 = pi0609 & ~n26564;
  assign n26647 = ~pi1155 & ~n26646;
  assign n26648 = ~n26645 & n26647;
  assign n26649 = ~pi0660 & ~n26581;
  assign n26650 = ~n26648 & n26649;
  assign n26651 = pi0609 & ~n26644;
  assign n26652 = ~pi0609 & ~n26564;
  assign n26653 = pi1155 & ~n26652;
  assign n26654 = ~n26651 & n26653;
  assign n26655 = pi0660 & ~n26583;
  assign n26656 = ~n26654 & n26655;
  assign n26657 = ~n26650 & ~n26656;
  assign n26658 = pi0785 & ~n26657;
  assign n26659 = ~pi0785 & ~n26644;
  assign n26660 = ~n26658 & ~n26659;
  assign n26661 = ~pi0618 & ~n26660;
  assign n26662 = ~pi1154 & ~n26629;
  assign n26663 = ~n26661 & n26662;
  assign n26664 = ~pi0627 & ~n26589;
  assign n26665 = ~n26663 & n26664;
  assign n26666 = ~pi0618 & n26565;
  assign n26667 = pi0618 & ~n26660;
  assign n26668 = pi1154 & ~n26666;
  assign n26669 = ~n26667 & n26668;
  assign n26670 = pi0627 & ~n26591;
  assign n26671 = ~n26669 & n26670;
  assign n26672 = ~n26665 & ~n26671;
  assign n26673 = pi0781 & ~n26672;
  assign n26674 = ~pi0781 & ~n26660;
  assign n26675 = ~n26673 & ~n26674;
  assign n26676 = ~pi0789 & n26675;
  assign n26677 = ~pi0619 & ~n26675;
  assign n26678 = pi0619 & n26566;
  assign n26679 = ~pi1159 & ~n26678;
  assign n26680 = ~n26677 & n26679;
  assign n26681 = ~pi0648 & ~n26597;
  assign n26682 = ~n26680 & n26681;
  assign n26683 = pi0619 & ~n26675;
  assign n26684 = ~pi0619 & n26566;
  assign n26685 = pi1159 & ~n26684;
  assign n26686 = ~n26683 & n26685;
  assign n26687 = pi0648 & ~n26599;
  assign n26688 = ~n26686 & n26687;
  assign n26689 = pi0789 & ~n26682;
  assign n26690 = ~n26688 & n26689;
  assign n26691 = n17970 & ~n26676;
  assign n26692 = ~n26690 & n26691;
  assign n26693 = ~n26628 & ~n26692;
  assign n26694 = ~n20364 & ~n26693;
  assign n26695 = n17854 & ~n26605;
  assign n26696 = n20851 & n26568;
  assign n26697 = ~n26695 & ~n26696;
  assign n26698 = ~pi0629 & ~n26697;
  assign n26699 = n20855 & n26568;
  assign n26700 = n17853 & ~n26605;
  assign n26701 = ~n26699 & ~n26700;
  assign n26702 = pi0629 & ~n26701;
  assign n26703 = ~n26698 & ~n26702;
  assign n26704 = pi0792 & ~n26703;
  assign n26705 = ~n20206 & ~n26704;
  assign n26706 = ~n26694 & n26705;
  assign n26707 = ~n26616 & ~n26706;
  assign n26708 = ~pi0790 & n26707;
  assign n26709 = ~pi0787 & ~n26569;
  assign n26710 = pi1157 & ~n26612;
  assign n26711 = ~n26573 & ~n26710;
  assign n26712 = pi0787 & ~n26711;
  assign n26713 = ~n26709 & ~n26712;
  assign n26714 = ~pi0644 & n26713;
  assign n26715 = pi0644 & n26707;
  assign n26716 = pi0715 & ~n26714;
  assign n26717 = ~n26715 & n26716;
  assign n26718 = ~n17804 & ~n26608;
  assign n26719 = n17804 & n26553;
  assign n26720 = ~n26718 & ~n26719;
  assign n26721 = pi0644 & ~n26720;
  assign n26722 = ~pi0644 & n26553;
  assign n26723 = ~pi0715 & ~n26722;
  assign n26724 = ~n26721 & n26723;
  assign n26725 = pi1160 & ~n26724;
  assign n26726 = ~n26717 & n26725;
  assign n26727 = ~pi0644 & ~n26720;
  assign n26728 = pi0644 & n26553;
  assign n26729 = pi0715 & ~n26728;
  assign n26730 = ~n26727 & n26729;
  assign n26731 = pi0644 & n26713;
  assign n26732 = ~pi0644 & n26707;
  assign n26733 = ~pi0715 & ~n26731;
  assign n26734 = ~n26732 & n26733;
  assign n26735 = ~pi1160 & ~n26730;
  assign n26736 = ~n26734 & n26735;
  assign n26737 = ~n26726 & ~n26736;
  assign n26738 = pi0790 & ~n26737;
  assign n26739 = pi0832 & ~n26708;
  assign n26740 = ~n26738 & n26739;
  assign n26741 = ~pi0181 & po1038;
  assign n26742 = ~pi0181 & ~n17059;
  assign n26743 = n16635 & ~n26742;
  assign n26744 = ~pi0709 & n2571;
  assign n26745 = n26742 & ~n26744;
  assign n26746 = ~pi0181 & ~n16641;
  assign n26747 = n16647 & ~n26746;
  assign n26748 = pi0181 & ~n18076;
  assign n26749 = ~pi0038 & ~n26748;
  assign n26750 = n2571 & ~n26749;
  assign n26751 = ~pi0181 & n18072;
  assign n26752 = ~n26750 & ~n26751;
  assign n26753 = ~pi0709 & ~n26747;
  assign n26754 = ~n26752 & n26753;
  assign n26755 = ~n26745 & ~n26754;
  assign n26756 = ~pi0778 & n26755;
  assign n26757 = ~pi0625 & n26742;
  assign n26758 = pi0625 & ~n26755;
  assign n26759 = pi1153 & ~n26757;
  assign n26760 = ~n26758 & n26759;
  assign n26761 = pi0625 & n26742;
  assign n26762 = ~pi0625 & ~n26755;
  assign n26763 = ~pi1153 & ~n26761;
  assign n26764 = ~n26762 & n26763;
  assign n26765 = ~n26760 & ~n26764;
  assign n26766 = pi0778 & ~n26765;
  assign n26767 = ~n26756 & ~n26766;
  assign n26768 = ~n17075 & ~n26767;
  assign n26769 = n17075 & ~n26742;
  assign n26770 = ~n26768 & ~n26769;
  assign n26771 = ~n16639 & n26770;
  assign n26772 = n16639 & n26742;
  assign n26773 = ~n26771 & ~n26772;
  assign n26774 = ~n16635 & n26773;
  assign n26775 = ~n26743 & ~n26774;
  assign n26776 = ~n16631 & n26775;
  assign n26777 = n16631 & n26742;
  assign n26778 = ~n26776 & ~n26777;
  assign n26779 = ~pi0792 & n26778;
  assign n26780 = pi0628 & ~n26778;
  assign n26781 = ~pi0628 & n26742;
  assign n26782 = pi1156 & ~n26781;
  assign n26783 = ~n26780 & n26782;
  assign n26784 = pi0628 & n26742;
  assign n26785 = ~pi0628 & ~n26778;
  assign n26786 = ~pi1156 & ~n26784;
  assign n26787 = ~n26785 & n26786;
  assign n26788 = ~n26783 & ~n26787;
  assign n26789 = pi0792 & ~n26788;
  assign n26790 = ~n26779 & ~n26789;
  assign n26791 = ~pi0647 & ~n26790;
  assign n26792 = pi0647 & ~n26742;
  assign n26793 = ~n26791 & ~n26792;
  assign n26794 = ~pi1157 & n26793;
  assign n26795 = pi0647 & ~n26790;
  assign n26796 = ~pi0647 & ~n26742;
  assign n26797 = ~n26795 & ~n26796;
  assign n26798 = pi1157 & n26797;
  assign n26799 = ~n26794 & ~n26798;
  assign n26800 = pi0787 & ~n26799;
  assign n26801 = ~pi0787 & n26790;
  assign n26802 = ~n26800 & ~n26801;
  assign n26803 = ~pi0644 & ~n26802;
  assign n26804 = pi0715 & ~n26803;
  assign n26805 = pi0181 & ~n2571;
  assign n26806 = pi0181 & pi0754;
  assign n26807 = pi0754 & n17046;
  assign n26808 = pi0181 & n17273;
  assign n26809 = ~n26807 & ~n26808;
  assign n26810 = pi0039 & ~n26809;
  assign n26811 = pi0181 & ~n17233;
  assign n26812 = ~n21812 & ~n26811;
  assign n26813 = ~pi0039 & ~n26812;
  assign n26814 = ~pi0181 & ~pi0754;
  assign n26815 = n17221 & n26814;
  assign n26816 = ~n26806 & ~n26813;
  assign n26817 = ~n26815 & n26816;
  assign n26818 = ~n26810 & n26817;
  assign n26819 = ~pi0038 & ~n26818;
  assign n26820 = ~pi0754 & n17280;
  assign n26821 = pi0038 & ~n26746;
  assign n26822 = ~n26820 & n26821;
  assign n26823 = ~n26819 & ~n26822;
  assign n26824 = n2571 & ~n26823;
  assign n26825 = ~n26805 & ~n26824;
  assign n26826 = ~n17117 & ~n26825;
  assign n26827 = n17117 & ~n26742;
  assign n26828 = ~n26826 & ~n26827;
  assign n26829 = ~pi0785 & ~n26828;
  assign n26830 = ~n17291 & ~n26742;
  assign n26831 = pi0609 & n26826;
  assign n26832 = ~n26830 & ~n26831;
  assign n26833 = pi1155 & ~n26832;
  assign n26834 = ~n17296 & ~n26742;
  assign n26835 = ~pi0609 & n26826;
  assign n26836 = ~n26834 & ~n26835;
  assign n26837 = ~pi1155 & ~n26836;
  assign n26838 = ~n26833 & ~n26837;
  assign n26839 = pi0785 & ~n26838;
  assign n26840 = ~n26829 & ~n26839;
  assign n26841 = ~pi0781 & ~n26840;
  assign n26842 = ~pi0618 & n26742;
  assign n26843 = pi0618 & n26840;
  assign n26844 = pi1154 & ~n26842;
  assign n26845 = ~n26843 & n26844;
  assign n26846 = ~pi0618 & n26840;
  assign n26847 = pi0618 & n26742;
  assign n26848 = ~pi1154 & ~n26847;
  assign n26849 = ~n26846 & n26848;
  assign n26850 = ~n26845 & ~n26849;
  assign n26851 = pi0781 & ~n26850;
  assign n26852 = ~n26841 & ~n26851;
  assign n26853 = ~pi0789 & ~n26852;
  assign n26854 = ~pi0619 & n26742;
  assign n26855 = pi0619 & n26852;
  assign n26856 = pi1159 & ~n26854;
  assign n26857 = ~n26855 & n26856;
  assign n26858 = ~pi0619 & n26852;
  assign n26859 = pi0619 & n26742;
  assign n26860 = ~pi1159 & ~n26859;
  assign n26861 = ~n26858 & n26860;
  assign n26862 = ~n26857 & ~n26861;
  assign n26863 = pi0789 & ~n26862;
  assign n26864 = ~n26853 & ~n26863;
  assign n26865 = ~n17969 & n26864;
  assign n26866 = n17969 & n26742;
  assign n26867 = ~n26865 & ~n26866;
  assign n26868 = ~n17779 & ~n26867;
  assign n26869 = n17779 & n26742;
  assign n26870 = ~n26868 & ~n26869;
  assign n26871 = ~n17804 & ~n26870;
  assign n26872 = n17804 & n26742;
  assign n26873 = ~n26871 & ~n26872;
  assign n26874 = pi0644 & ~n26873;
  assign n26875 = ~pi0644 & n26742;
  assign n26876 = ~pi0715 & ~n26875;
  assign n26877 = ~n26874 & n26876;
  assign n26878 = pi1160 & ~n26877;
  assign n26879 = ~n26804 & n26878;
  assign n26880 = pi0644 & ~n26802;
  assign n26881 = ~pi0715 & ~n26880;
  assign n26882 = ~pi0644 & ~n26873;
  assign n26883 = pi0644 & n26742;
  assign n26884 = pi0715 & ~n26883;
  assign n26885 = ~n26882 & n26884;
  assign n26886 = ~pi1160 & ~n26885;
  assign n26887 = ~n26881 & n26886;
  assign n26888 = ~n26879 & ~n26887;
  assign n26889 = pi0790 & ~n26888;
  assign n26890 = ~pi0629 & n26783;
  assign n26891 = ~n20570 & n26867;
  assign n26892 = pi0629 & n26787;
  assign n26893 = ~n26890 & ~n26892;
  assign n26894 = ~n26891 & n26893;
  assign n26895 = pi0792 & ~n26894;
  assign n26896 = pi0609 & n26767;
  assign n26897 = pi0181 & ~n17625;
  assign n26898 = ~pi0181 & ~n17612;
  assign n26899 = pi0754 & ~n26897;
  assign n26900 = ~n26898 & n26899;
  assign n26901 = ~pi0181 & n17629;
  assign n26902 = pi0181 & n17631;
  assign n26903 = ~pi0754 & ~n26902;
  assign n26904 = ~n26901 & n26903;
  assign n26905 = ~n26900 & ~n26904;
  assign n26906 = ~pi0039 & ~n26905;
  assign n26907 = pi0181 & n17605;
  assign n26908 = ~pi0181 & ~n17546;
  assign n26909 = ~pi0754 & ~n26908;
  assign n26910 = ~n26907 & n26909;
  assign n26911 = ~pi0181 & n17404;
  assign n26912 = pi0181 & n17485;
  assign n26913 = pi0754 & ~n26912;
  assign n26914 = ~n26911 & n26913;
  assign n26915 = pi0039 & ~n26910;
  assign n26916 = ~n26914 & n26915;
  assign n26917 = ~pi0038 & ~n26906;
  assign n26918 = ~n26916 & n26917;
  assign n26919 = ~n17469 & ~n26575;
  assign n26920 = pi0181 & ~n26919;
  assign n26921 = n6284 & n26920;
  assign n26922 = ~pi0754 & ~n17490;
  assign n26923 = n19471 & ~n26922;
  assign n26924 = ~pi0181 & ~n26923;
  assign n26925 = pi0038 & ~n26921;
  assign n26926 = ~n26924 & n26925;
  assign n26927 = ~pi0709 & ~n26926;
  assign n26928 = ~n26918 & n26927;
  assign n26929 = pi0709 & n26823;
  assign n26930 = n2571 & ~n26928;
  assign n26931 = ~n26929 & n26930;
  assign n26932 = ~n26805 & ~n26931;
  assign n26933 = ~pi0625 & n26932;
  assign n26934 = pi0625 & n26825;
  assign n26935 = ~pi1153 & ~n26934;
  assign n26936 = ~n26933 & n26935;
  assign n26937 = ~pi0608 & ~n26760;
  assign n26938 = ~n26936 & n26937;
  assign n26939 = ~pi0625 & n26825;
  assign n26940 = pi0625 & n26932;
  assign n26941 = pi1153 & ~n26939;
  assign n26942 = ~n26940 & n26941;
  assign n26943 = pi0608 & ~n26764;
  assign n26944 = ~n26942 & n26943;
  assign n26945 = ~n26938 & ~n26944;
  assign n26946 = pi0778 & ~n26945;
  assign n26947 = ~pi0778 & n26932;
  assign n26948 = ~n26946 & ~n26947;
  assign n26949 = ~pi0609 & ~n26948;
  assign n26950 = ~pi1155 & ~n26896;
  assign n26951 = ~n26949 & n26950;
  assign n26952 = ~pi0660 & ~n26833;
  assign n26953 = ~n26951 & n26952;
  assign n26954 = ~pi0609 & n26767;
  assign n26955 = pi0609 & ~n26948;
  assign n26956 = pi1155 & ~n26954;
  assign n26957 = ~n26955 & n26956;
  assign n26958 = pi0660 & ~n26837;
  assign n26959 = ~n26957 & n26958;
  assign n26960 = ~n26953 & ~n26959;
  assign n26961 = pi0785 & ~n26960;
  assign n26962 = ~pi0785 & ~n26948;
  assign n26963 = ~n26961 & ~n26962;
  assign n26964 = ~pi0618 & ~n26963;
  assign n26965 = pi0618 & n26770;
  assign n26966 = ~pi1154 & ~n26965;
  assign n26967 = ~n26964 & n26966;
  assign n26968 = ~pi0627 & ~n26845;
  assign n26969 = ~n26967 & n26968;
  assign n26970 = ~pi0618 & n26770;
  assign n26971 = pi0618 & ~n26963;
  assign n26972 = pi1154 & ~n26970;
  assign n26973 = ~n26971 & n26972;
  assign n26974 = pi0627 & ~n26849;
  assign n26975 = ~n26973 & n26974;
  assign n26976 = ~n26969 & ~n26975;
  assign n26977 = pi0781 & ~n26976;
  assign n26978 = ~pi0781 & ~n26963;
  assign n26979 = ~n26977 & ~n26978;
  assign n26980 = ~pi0789 & n26979;
  assign n26981 = pi0619 & ~n26773;
  assign n26982 = ~pi0619 & ~n26979;
  assign n26983 = ~pi1159 & ~n26981;
  assign n26984 = ~n26982 & n26983;
  assign n26985 = ~pi0648 & ~n26857;
  assign n26986 = ~n26984 & n26985;
  assign n26987 = ~pi0619 & ~n26773;
  assign n26988 = pi0619 & ~n26979;
  assign n26989 = pi1159 & ~n26987;
  assign n26990 = ~n26988 & n26989;
  assign n26991 = pi0648 & ~n26861;
  assign n26992 = ~n26990 & n26991;
  assign n26993 = pi0789 & ~n26986;
  assign n26994 = ~n26992 & n26993;
  assign n26995 = n17970 & ~n26980;
  assign n26996 = ~n26994 & n26995;
  assign n26997 = n17871 & n26775;
  assign n26998 = ~pi0626 & ~n26864;
  assign n26999 = pi0626 & ~n26742;
  assign n27000 = n16629 & ~n26999;
  assign n27001 = ~n26998 & n27000;
  assign n27002 = pi0626 & ~n26864;
  assign n27003 = ~pi0626 & ~n26742;
  assign n27004 = n16628 & ~n27003;
  assign n27005 = ~n27002 & n27004;
  assign n27006 = ~n26997 & ~n27001;
  assign n27007 = ~n27005 & n27006;
  assign n27008 = pi0788 & ~n27007;
  assign n27009 = ~n20364 & ~n27008;
  assign n27010 = ~n26996 & n27009;
  assign n27011 = ~n26895 & ~n27010;
  assign n27012 = ~n20206 & ~n27011;
  assign n27013 = n17802 & ~n26793;
  assign n27014 = ~n20559 & n26870;
  assign n27015 = n17801 & ~n26797;
  assign n27016 = ~n27013 & ~n27015;
  assign n27017 = ~n27014 & n27016;
  assign n27018 = pi0787 & ~n27017;
  assign n27019 = ~pi0644 & n26886;
  assign n27020 = pi0644 & n26878;
  assign n27021 = pi0790 & ~n27019;
  assign n27022 = ~n27020 & n27021;
  assign n27023 = ~n27012 & ~n27018;
  assign n27024 = ~n27022 & n27023;
  assign n27025 = ~n26889 & ~n27024;
  assign n27026 = ~po1038 & ~n27025;
  assign n27027 = ~pi0832 & ~n26741;
  assign n27028 = ~n27026 & n27027;
  assign po0338 = ~n26740 & ~n27028;
  assign n27030 = ~pi0182 & ~n2926;
  assign n27031 = ~pi0734 & n16645;
  assign n27032 = ~n27030 & ~n27031;
  assign n27033 = ~pi0778 & ~n27032;
  assign n27034 = ~pi0625 & n27031;
  assign n27035 = ~n27032 & ~n27034;
  assign n27036 = pi1153 & ~n27035;
  assign n27037 = ~pi1153 & ~n27030;
  assign n27038 = ~n27034 & n27037;
  assign n27039 = pi0778 & ~n27038;
  assign n27040 = ~n27036 & n27039;
  assign n27041 = ~n27033 & ~n27040;
  assign n27042 = ~n17845 & ~n27041;
  assign n27043 = ~n17847 & n27042;
  assign n27044 = ~n17849 & n27043;
  assign n27045 = ~n17851 & n27044;
  assign n27046 = ~n17857 & n27045;
  assign n27047 = ~pi0647 & n27046;
  assign n27048 = pi0647 & n27030;
  assign n27049 = ~pi1157 & ~n27048;
  assign n27050 = ~n27047 & n27049;
  assign n27051 = pi0630 & n27050;
  assign n27052 = ~pi0756 & n17244;
  assign n27053 = ~n27030 & ~n27052;
  assign n27054 = ~n17874 & ~n27053;
  assign n27055 = ~pi0785 & ~n27054;
  assign n27056 = n17296 & n27052;
  assign n27057 = n27054 & ~n27056;
  assign n27058 = pi1155 & ~n27057;
  assign n27059 = ~pi1155 & ~n27030;
  assign n27060 = ~n27056 & n27059;
  assign n27061 = ~n27058 & ~n27060;
  assign n27062 = pi0785 & ~n27061;
  assign n27063 = ~n27055 & ~n27062;
  assign n27064 = ~pi0781 & ~n27063;
  assign n27065 = ~n17889 & n27063;
  assign n27066 = pi1154 & ~n27065;
  assign n27067 = ~n17892 & n27063;
  assign n27068 = ~pi1154 & ~n27067;
  assign n27069 = ~n27066 & ~n27068;
  assign n27070 = pi0781 & ~n27069;
  assign n27071 = ~n27064 & ~n27070;
  assign n27072 = ~pi0789 & ~n27071;
  assign n27073 = ~n23078 & n27071;
  assign n27074 = pi1159 & ~n27073;
  assign n27075 = ~n23081 & n27071;
  assign n27076 = ~pi1159 & ~n27075;
  assign n27077 = ~n27074 & ~n27076;
  assign n27078 = pi0789 & ~n27077;
  assign n27079 = ~n27072 & ~n27078;
  assign n27080 = ~n17969 & n27079;
  assign n27081 = n17969 & n27030;
  assign n27082 = ~n27080 & ~n27081;
  assign n27083 = ~n17779 & ~n27082;
  assign n27084 = n17779 & n27030;
  assign n27085 = ~n27083 & ~n27084;
  assign n27086 = ~n20559 & n27085;
  assign n27087 = pi0647 & ~n27046;
  assign n27088 = ~pi0647 & ~n27030;
  assign n27089 = ~n27087 & ~n27088;
  assign n27090 = n17801 & ~n27089;
  assign n27091 = ~n27051 & ~n27090;
  assign n27092 = ~n27086 & n27091;
  assign n27093 = pi0787 & ~n27092;
  assign n27094 = n17871 & n27044;
  assign n27095 = ~pi0626 & ~n27079;
  assign n27096 = pi0626 & ~n27030;
  assign n27097 = n16629 & ~n27096;
  assign n27098 = ~n27095 & n27097;
  assign n27099 = pi0626 & ~n27079;
  assign n27100 = ~pi0626 & ~n27030;
  assign n27101 = n16628 & ~n27100;
  assign n27102 = ~n27099 & n27101;
  assign n27103 = ~n27094 & ~n27098;
  assign n27104 = ~n27102 & n27103;
  assign n27105 = pi0788 & ~n27104;
  assign n27106 = pi0618 & n27042;
  assign n27107 = ~n17168 & ~n27032;
  assign n27108 = pi0625 & n27107;
  assign n27109 = n27053 & ~n27107;
  assign n27110 = ~n27108 & ~n27109;
  assign n27111 = n27037 & ~n27110;
  assign n27112 = ~pi0608 & ~n27036;
  assign n27113 = ~n27111 & n27112;
  assign n27114 = pi1153 & n27053;
  assign n27115 = ~n27108 & n27114;
  assign n27116 = pi0608 & ~n27038;
  assign n27117 = ~n27115 & n27116;
  assign n27118 = ~n27113 & ~n27117;
  assign n27119 = pi0778 & ~n27118;
  assign n27120 = ~pi0778 & ~n27109;
  assign n27121 = ~n27119 & ~n27120;
  assign n27122 = ~pi0609 & ~n27121;
  assign n27123 = pi0609 & ~n27041;
  assign n27124 = ~pi1155 & ~n27123;
  assign n27125 = ~n27122 & n27124;
  assign n27126 = ~pi0660 & ~n27058;
  assign n27127 = ~n27125 & n27126;
  assign n27128 = pi0609 & ~n27121;
  assign n27129 = ~pi0609 & ~n27041;
  assign n27130 = pi1155 & ~n27129;
  assign n27131 = ~n27128 & n27130;
  assign n27132 = pi0660 & ~n27060;
  assign n27133 = ~n27131 & n27132;
  assign n27134 = ~n27127 & ~n27133;
  assign n27135 = pi0785 & ~n27134;
  assign n27136 = ~pi0785 & ~n27121;
  assign n27137 = ~n27135 & ~n27136;
  assign n27138 = ~pi0618 & ~n27137;
  assign n27139 = ~pi1154 & ~n27106;
  assign n27140 = ~n27138 & n27139;
  assign n27141 = ~pi0627 & ~n27066;
  assign n27142 = ~n27140 & n27141;
  assign n27143 = ~pi0618 & n27042;
  assign n27144 = pi0618 & ~n27137;
  assign n27145 = pi1154 & ~n27143;
  assign n27146 = ~n27144 & n27145;
  assign n27147 = pi0627 & ~n27068;
  assign n27148 = ~n27146 & n27147;
  assign n27149 = ~n27142 & ~n27148;
  assign n27150 = pi0781 & ~n27149;
  assign n27151 = ~pi0781 & ~n27137;
  assign n27152 = ~n27150 & ~n27151;
  assign n27153 = ~pi0789 & n27152;
  assign n27154 = ~pi0619 & ~n27152;
  assign n27155 = pi0619 & n27043;
  assign n27156 = ~pi1159 & ~n27155;
  assign n27157 = ~n27154 & n27156;
  assign n27158 = ~pi0648 & ~n27074;
  assign n27159 = ~n27157 & n27158;
  assign n27160 = pi0619 & ~n27152;
  assign n27161 = ~pi0619 & n27043;
  assign n27162 = pi1159 & ~n27161;
  assign n27163 = ~n27160 & n27162;
  assign n27164 = pi0648 & ~n27076;
  assign n27165 = ~n27163 & n27164;
  assign n27166 = pi0789 & ~n27159;
  assign n27167 = ~n27165 & n27166;
  assign n27168 = n17970 & ~n27153;
  assign n27169 = ~n27167 & n27168;
  assign n27170 = ~n27105 & ~n27169;
  assign n27171 = ~n20364 & ~n27170;
  assign n27172 = n17854 & ~n27082;
  assign n27173 = n20851 & n27045;
  assign n27174 = ~n27172 & ~n27173;
  assign n27175 = ~pi0629 & ~n27174;
  assign n27176 = n20855 & n27045;
  assign n27177 = n17853 & ~n27082;
  assign n27178 = ~n27176 & ~n27177;
  assign n27179 = pi0629 & ~n27178;
  assign n27180 = ~n27175 & ~n27179;
  assign n27181 = pi0792 & ~n27180;
  assign n27182 = ~n20206 & ~n27181;
  assign n27183 = ~n27171 & n27182;
  assign n27184 = ~n27093 & ~n27183;
  assign n27185 = ~pi0790 & n27184;
  assign n27186 = ~pi0787 & ~n27046;
  assign n27187 = pi1157 & ~n27089;
  assign n27188 = ~n27050 & ~n27187;
  assign n27189 = pi0787 & ~n27188;
  assign n27190 = ~n27186 & ~n27189;
  assign n27191 = ~pi0644 & n27190;
  assign n27192 = pi0644 & n27184;
  assign n27193 = pi0715 & ~n27191;
  assign n27194 = ~n27192 & n27193;
  assign n27195 = ~n17804 & ~n27085;
  assign n27196 = n17804 & n27030;
  assign n27197 = ~n27195 & ~n27196;
  assign n27198 = pi0644 & ~n27197;
  assign n27199 = ~pi0644 & n27030;
  assign n27200 = ~pi0715 & ~n27199;
  assign n27201 = ~n27198 & n27200;
  assign n27202 = pi1160 & ~n27201;
  assign n27203 = ~n27194 & n27202;
  assign n27204 = ~pi0644 & ~n27197;
  assign n27205 = pi0644 & n27030;
  assign n27206 = pi0715 & ~n27205;
  assign n27207 = ~n27204 & n27206;
  assign n27208 = pi0644 & n27190;
  assign n27209 = ~pi0644 & n27184;
  assign n27210 = ~pi0715 & ~n27208;
  assign n27211 = ~n27209 & n27210;
  assign n27212 = ~pi1160 & ~n27207;
  assign n27213 = ~n27211 & n27212;
  assign n27214 = ~n27203 & ~n27213;
  assign n27215 = pi0790 & ~n27214;
  assign n27216 = pi0832 & ~n27185;
  assign n27217 = ~n27215 & n27216;
  assign n27218 = ~pi0182 & po1038;
  assign n27219 = ~pi0182 & ~n17059;
  assign n27220 = n16635 & ~n27219;
  assign n27221 = ~pi0734 & n2571;
  assign n27222 = n27219 & ~n27221;
  assign n27223 = ~pi0182 & ~n16641;
  assign n27224 = n16647 & ~n27223;
  assign n27225 = pi0182 & ~n18076;
  assign n27226 = ~pi0038 & ~n27225;
  assign n27227 = n2571 & ~n27226;
  assign n27228 = ~pi0182 & n18072;
  assign n27229 = ~n27227 & ~n27228;
  assign n27230 = ~pi0734 & ~n27224;
  assign n27231 = ~n27229 & n27230;
  assign n27232 = ~n27222 & ~n27231;
  assign n27233 = ~pi0778 & n27232;
  assign n27234 = ~pi0625 & n27219;
  assign n27235 = pi0625 & ~n27232;
  assign n27236 = pi1153 & ~n27234;
  assign n27237 = ~n27235 & n27236;
  assign n27238 = pi0625 & n27219;
  assign n27239 = ~pi0625 & ~n27232;
  assign n27240 = ~pi1153 & ~n27238;
  assign n27241 = ~n27239 & n27240;
  assign n27242 = ~n27237 & ~n27241;
  assign n27243 = pi0778 & ~n27242;
  assign n27244 = ~n27233 & ~n27243;
  assign n27245 = ~n17075 & ~n27244;
  assign n27246 = n17075 & ~n27219;
  assign n27247 = ~n27245 & ~n27246;
  assign n27248 = ~n16639 & n27247;
  assign n27249 = n16639 & n27219;
  assign n27250 = ~n27248 & ~n27249;
  assign n27251 = ~n16635 & n27250;
  assign n27252 = ~n27220 & ~n27251;
  assign n27253 = ~n16631 & n27252;
  assign n27254 = n16631 & n27219;
  assign n27255 = ~n27253 & ~n27254;
  assign n27256 = ~pi0792 & n27255;
  assign n27257 = pi0628 & ~n27255;
  assign n27258 = ~pi0628 & n27219;
  assign n27259 = pi1156 & ~n27258;
  assign n27260 = ~n27257 & n27259;
  assign n27261 = pi0628 & n27219;
  assign n27262 = ~pi0628 & ~n27255;
  assign n27263 = ~pi1156 & ~n27261;
  assign n27264 = ~n27262 & n27263;
  assign n27265 = ~n27260 & ~n27264;
  assign n27266 = pi0792 & ~n27265;
  assign n27267 = ~n27256 & ~n27266;
  assign n27268 = ~pi0647 & ~n27267;
  assign n27269 = pi0647 & ~n27219;
  assign n27270 = ~n27268 & ~n27269;
  assign n27271 = ~pi1157 & n27270;
  assign n27272 = pi0647 & ~n27267;
  assign n27273 = ~pi0647 & ~n27219;
  assign n27274 = ~n27272 & ~n27273;
  assign n27275 = pi1157 & n27274;
  assign n27276 = ~n27271 & ~n27275;
  assign n27277 = pi0787 & ~n27276;
  assign n27278 = ~pi0787 & n27267;
  assign n27279 = ~n27277 & ~n27278;
  assign n27280 = ~pi0644 & ~n27279;
  assign n27281 = pi0715 & ~n27280;
  assign n27282 = pi0182 & ~n2571;
  assign n27283 = ~pi0756 & n17280;
  assign n27284 = ~n27223 & ~n27283;
  assign n27285 = pi0038 & ~n27284;
  assign n27286 = ~pi0182 & n17221;
  assign n27287 = pi0182 & ~n17275;
  assign n27288 = ~pi0756 & ~n27287;
  assign n27289 = ~n27286 & n27288;
  assign n27290 = ~pi0182 & pi0756;
  assign n27291 = ~n17048 & n27290;
  assign n27292 = ~n27289 & ~n27291;
  assign n27293 = ~pi0038 & ~n27292;
  assign n27294 = ~n27285 & ~n27293;
  assign n27295 = n2571 & n27294;
  assign n27296 = ~n27282 & ~n27295;
  assign n27297 = ~n17117 & ~n27296;
  assign n27298 = n17117 & ~n27219;
  assign n27299 = ~n27297 & ~n27298;
  assign n27300 = ~pi0785 & ~n27299;
  assign n27301 = ~n17291 & ~n27219;
  assign n27302 = pi0609 & n27297;
  assign n27303 = ~n27301 & ~n27302;
  assign n27304 = pi1155 & ~n27303;
  assign n27305 = ~n17296 & ~n27219;
  assign n27306 = ~pi0609 & n27297;
  assign n27307 = ~n27305 & ~n27306;
  assign n27308 = ~pi1155 & ~n27307;
  assign n27309 = ~n27304 & ~n27308;
  assign n27310 = pi0785 & ~n27309;
  assign n27311 = ~n27300 & ~n27310;
  assign n27312 = ~pi0781 & ~n27311;
  assign n27313 = ~pi0618 & n27219;
  assign n27314 = pi0618 & n27311;
  assign n27315 = pi1154 & ~n27313;
  assign n27316 = ~n27314 & n27315;
  assign n27317 = ~pi0618 & n27311;
  assign n27318 = pi0618 & n27219;
  assign n27319 = ~pi1154 & ~n27318;
  assign n27320 = ~n27317 & n27319;
  assign n27321 = ~n27316 & ~n27320;
  assign n27322 = pi0781 & ~n27321;
  assign n27323 = ~n27312 & ~n27322;
  assign n27324 = ~pi0789 & ~n27323;
  assign n27325 = ~pi0619 & n27219;
  assign n27326 = pi0619 & n27323;
  assign n27327 = pi1159 & ~n27325;
  assign n27328 = ~n27326 & n27327;
  assign n27329 = ~pi0619 & n27323;
  assign n27330 = pi0619 & n27219;
  assign n27331 = ~pi1159 & ~n27330;
  assign n27332 = ~n27329 & n27331;
  assign n27333 = ~n27328 & ~n27332;
  assign n27334 = pi0789 & ~n27333;
  assign n27335 = ~n27324 & ~n27334;
  assign n27336 = ~n17969 & n27335;
  assign n27337 = n17969 & n27219;
  assign n27338 = ~n27336 & ~n27337;
  assign n27339 = ~n17779 & ~n27338;
  assign n27340 = n17779 & n27219;
  assign n27341 = ~n27339 & ~n27340;
  assign n27342 = ~n17804 & ~n27341;
  assign n27343 = n17804 & n27219;
  assign n27344 = ~n27342 & ~n27343;
  assign n27345 = pi0644 & ~n27344;
  assign n27346 = ~pi0644 & n27219;
  assign n27347 = ~pi0715 & ~n27346;
  assign n27348 = ~n27345 & n27347;
  assign n27349 = pi1160 & ~n27348;
  assign n27350 = ~n27281 & n27349;
  assign n27351 = pi0644 & ~n27279;
  assign n27352 = ~pi0715 & ~n27351;
  assign n27353 = ~pi0644 & ~n27344;
  assign n27354 = pi0644 & n27219;
  assign n27355 = pi0715 & ~n27354;
  assign n27356 = ~n27353 & n27355;
  assign n27357 = ~pi1160 & ~n27356;
  assign n27358 = ~n27352 & n27357;
  assign n27359 = ~n27350 & ~n27358;
  assign n27360 = pi0790 & ~n27359;
  assign n27361 = ~pi0629 & n27260;
  assign n27362 = ~n20570 & n27338;
  assign n27363 = pi0629 & n27264;
  assign n27364 = ~n27361 & ~n27363;
  assign n27365 = ~n27362 & n27364;
  assign n27366 = pi0792 & ~n27365;
  assign n27367 = pi0609 & n27244;
  assign n27368 = pi0182 & ~n17625;
  assign n27369 = ~pi0182 & ~n17612;
  assign n27370 = pi0756 & ~n27368;
  assign n27371 = ~n27369 & n27370;
  assign n27372 = ~pi0182 & n17629;
  assign n27373 = pi0182 & n17631;
  assign n27374 = ~pi0756 & ~n27373;
  assign n27375 = ~n27372 & n27374;
  assign n27376 = ~n27371 & ~n27375;
  assign n27377 = ~pi0039 & ~n27376;
  assign n27378 = pi0182 & n17605;
  assign n27379 = ~pi0182 & ~n17546;
  assign n27380 = ~pi0756 & ~n27379;
  assign n27381 = ~n27378 & n27380;
  assign n27382 = ~pi0182 & n17404;
  assign n27383 = pi0182 & n17485;
  assign n27384 = pi0756 & ~n27383;
  assign n27385 = ~n27382 & n27384;
  assign n27386 = pi0039 & ~n27381;
  assign n27387 = ~n27385 & n27386;
  assign n27388 = ~pi0038 & ~n27377;
  assign n27389 = ~n27387 & n27388;
  assign n27390 = ~pi0756 & ~n17490;
  assign n27391 = n19471 & ~n27390;
  assign n27392 = ~pi0182 & ~n27391;
  assign n27393 = ~n17469 & ~n27052;
  assign n27394 = pi0182 & ~n27393;
  assign n27395 = n6284 & n27394;
  assign n27396 = pi0038 & ~n27395;
  assign n27397 = ~n27392 & n27396;
  assign n27398 = ~pi0734 & ~n27397;
  assign n27399 = ~n27389 & n27398;
  assign n27400 = pi0734 & ~n27294;
  assign n27401 = n2571 & ~n27399;
  assign n27402 = ~n27400 & n27401;
  assign n27403 = ~n27282 & ~n27402;
  assign n27404 = ~pi0625 & n27403;
  assign n27405 = pi0625 & n27296;
  assign n27406 = ~pi1153 & ~n27405;
  assign n27407 = ~n27404 & n27406;
  assign n27408 = ~pi0608 & ~n27237;
  assign n27409 = ~n27407 & n27408;
  assign n27410 = ~pi0625 & n27296;
  assign n27411 = pi0625 & n27403;
  assign n27412 = pi1153 & ~n27410;
  assign n27413 = ~n27411 & n27412;
  assign n27414 = pi0608 & ~n27241;
  assign n27415 = ~n27413 & n27414;
  assign n27416 = ~n27409 & ~n27415;
  assign n27417 = pi0778 & ~n27416;
  assign n27418 = ~pi0778 & n27403;
  assign n27419 = ~n27417 & ~n27418;
  assign n27420 = ~pi0609 & ~n27419;
  assign n27421 = ~pi1155 & ~n27367;
  assign n27422 = ~n27420 & n27421;
  assign n27423 = ~pi0660 & ~n27304;
  assign n27424 = ~n27422 & n27423;
  assign n27425 = ~pi0609 & n27244;
  assign n27426 = pi0609 & ~n27419;
  assign n27427 = pi1155 & ~n27425;
  assign n27428 = ~n27426 & n27427;
  assign n27429 = pi0660 & ~n27308;
  assign n27430 = ~n27428 & n27429;
  assign n27431 = ~n27424 & ~n27430;
  assign n27432 = pi0785 & ~n27431;
  assign n27433 = ~pi0785 & ~n27419;
  assign n27434 = ~n27432 & ~n27433;
  assign n27435 = ~pi0618 & ~n27434;
  assign n27436 = pi0618 & n27247;
  assign n27437 = ~pi1154 & ~n27436;
  assign n27438 = ~n27435 & n27437;
  assign n27439 = ~pi0627 & ~n27316;
  assign n27440 = ~n27438 & n27439;
  assign n27441 = ~pi0618 & n27247;
  assign n27442 = pi0618 & ~n27434;
  assign n27443 = pi1154 & ~n27441;
  assign n27444 = ~n27442 & n27443;
  assign n27445 = pi0627 & ~n27320;
  assign n27446 = ~n27444 & n27445;
  assign n27447 = ~n27440 & ~n27446;
  assign n27448 = pi0781 & ~n27447;
  assign n27449 = ~pi0781 & ~n27434;
  assign n27450 = ~n27448 & ~n27449;
  assign n27451 = ~pi0789 & n27450;
  assign n27452 = pi0619 & ~n27250;
  assign n27453 = ~pi0619 & ~n27450;
  assign n27454 = ~pi1159 & ~n27452;
  assign n27455 = ~n27453 & n27454;
  assign n27456 = ~pi0648 & ~n27328;
  assign n27457 = ~n27455 & n27456;
  assign n27458 = ~pi0619 & ~n27250;
  assign n27459 = pi0619 & ~n27450;
  assign n27460 = pi1159 & ~n27458;
  assign n27461 = ~n27459 & n27460;
  assign n27462 = pi0648 & ~n27332;
  assign n27463 = ~n27461 & n27462;
  assign n27464 = pi0789 & ~n27457;
  assign n27465 = ~n27463 & n27464;
  assign n27466 = n17970 & ~n27451;
  assign n27467 = ~n27465 & n27466;
  assign n27468 = n17871 & n27252;
  assign n27469 = ~pi0626 & ~n27335;
  assign n27470 = pi0626 & ~n27219;
  assign n27471 = n16629 & ~n27470;
  assign n27472 = ~n27469 & n27471;
  assign n27473 = pi0626 & ~n27335;
  assign n27474 = ~pi0626 & ~n27219;
  assign n27475 = n16628 & ~n27474;
  assign n27476 = ~n27473 & n27475;
  assign n27477 = ~n27468 & ~n27472;
  assign n27478 = ~n27476 & n27477;
  assign n27479 = pi0788 & ~n27478;
  assign n27480 = ~n20364 & ~n27479;
  assign n27481 = ~n27467 & n27480;
  assign n27482 = ~n27366 & ~n27481;
  assign n27483 = ~n20206 & ~n27482;
  assign n27484 = n17802 & ~n27270;
  assign n27485 = ~n20559 & n27341;
  assign n27486 = n17801 & ~n27274;
  assign n27487 = ~n27484 & ~n27486;
  assign n27488 = ~n27485 & n27487;
  assign n27489 = pi0787 & ~n27488;
  assign n27490 = ~pi0644 & n27357;
  assign n27491 = pi0644 & n27349;
  assign n27492 = pi0790 & ~n27490;
  assign n27493 = ~n27491 & n27492;
  assign n27494 = ~n27483 & ~n27489;
  assign n27495 = ~n27493 & n27494;
  assign n27496 = ~n27360 & ~n27495;
  assign n27497 = ~po1038 & ~n27496;
  assign n27498 = ~pi0832 & ~n27218;
  assign n27499 = ~n27497 & n27498;
  assign po0339 = ~n27217 & ~n27499;
  assign n27501 = ~pi0183 & ~n2926;
  assign n27502 = ~pi0725 & n16645;
  assign n27503 = ~n27501 & ~n27502;
  assign n27504 = ~pi0778 & ~n27503;
  assign n27505 = ~pi0625 & n27502;
  assign n27506 = ~n27503 & ~n27505;
  assign n27507 = pi1153 & ~n27506;
  assign n27508 = ~pi1153 & ~n27501;
  assign n27509 = ~n27505 & n27508;
  assign n27510 = pi0778 & ~n27509;
  assign n27511 = ~n27507 & n27510;
  assign n27512 = ~n27504 & ~n27511;
  assign n27513 = ~n17845 & ~n27512;
  assign n27514 = ~n17847 & n27513;
  assign n27515 = ~n17849 & n27514;
  assign n27516 = ~n17851 & n27515;
  assign n27517 = ~n17857 & n27516;
  assign n27518 = ~pi0647 & n27517;
  assign n27519 = pi0647 & n27501;
  assign n27520 = ~pi1157 & ~n27519;
  assign n27521 = ~n27518 & n27520;
  assign n27522 = pi0630 & n27521;
  assign n27523 = ~pi0755 & n17244;
  assign n27524 = ~n27501 & ~n27523;
  assign n27525 = ~n17874 & ~n27524;
  assign n27526 = ~pi0785 & ~n27525;
  assign n27527 = n17296 & n27523;
  assign n27528 = n27525 & ~n27527;
  assign n27529 = pi1155 & ~n27528;
  assign n27530 = ~pi1155 & ~n27501;
  assign n27531 = ~n27527 & n27530;
  assign n27532 = ~n27529 & ~n27531;
  assign n27533 = pi0785 & ~n27532;
  assign n27534 = ~n27526 & ~n27533;
  assign n27535 = ~pi0781 & ~n27534;
  assign n27536 = ~n17889 & n27534;
  assign n27537 = pi1154 & ~n27536;
  assign n27538 = ~n17892 & n27534;
  assign n27539 = ~pi1154 & ~n27538;
  assign n27540 = ~n27537 & ~n27539;
  assign n27541 = pi0781 & ~n27540;
  assign n27542 = ~n27535 & ~n27541;
  assign n27543 = ~pi0789 & ~n27542;
  assign n27544 = ~n23078 & n27542;
  assign n27545 = pi1159 & ~n27544;
  assign n27546 = ~n23081 & n27542;
  assign n27547 = ~pi1159 & ~n27546;
  assign n27548 = ~n27545 & ~n27547;
  assign n27549 = pi0789 & ~n27548;
  assign n27550 = ~n27543 & ~n27549;
  assign n27551 = ~n17969 & n27550;
  assign n27552 = n17969 & n27501;
  assign n27553 = ~n27551 & ~n27552;
  assign n27554 = ~n17779 & ~n27553;
  assign n27555 = n17779 & n27501;
  assign n27556 = ~n27554 & ~n27555;
  assign n27557 = ~n20559 & n27556;
  assign n27558 = pi0647 & ~n27517;
  assign n27559 = ~pi0647 & ~n27501;
  assign n27560 = ~n27558 & ~n27559;
  assign n27561 = n17801 & ~n27560;
  assign n27562 = ~n27522 & ~n27561;
  assign n27563 = ~n27557 & n27562;
  assign n27564 = pi0787 & ~n27563;
  assign n27565 = n17871 & n27515;
  assign n27566 = ~pi0626 & ~n27550;
  assign n27567 = pi0626 & ~n27501;
  assign n27568 = n16629 & ~n27567;
  assign n27569 = ~n27566 & n27568;
  assign n27570 = pi0626 & ~n27550;
  assign n27571 = ~pi0626 & ~n27501;
  assign n27572 = n16628 & ~n27571;
  assign n27573 = ~n27570 & n27572;
  assign n27574 = ~n27565 & ~n27569;
  assign n27575 = ~n27573 & n27574;
  assign n27576 = pi0788 & ~n27575;
  assign n27577 = pi0618 & n27513;
  assign n27578 = ~n17168 & ~n27503;
  assign n27579 = pi0625 & n27578;
  assign n27580 = n27524 & ~n27578;
  assign n27581 = ~n27579 & ~n27580;
  assign n27582 = n27508 & ~n27581;
  assign n27583 = ~pi0608 & ~n27507;
  assign n27584 = ~n27582 & n27583;
  assign n27585 = pi1153 & n27524;
  assign n27586 = ~n27579 & n27585;
  assign n27587 = pi0608 & ~n27509;
  assign n27588 = ~n27586 & n27587;
  assign n27589 = ~n27584 & ~n27588;
  assign n27590 = pi0778 & ~n27589;
  assign n27591 = ~pi0778 & ~n27580;
  assign n27592 = ~n27590 & ~n27591;
  assign n27593 = ~pi0609 & ~n27592;
  assign n27594 = pi0609 & ~n27512;
  assign n27595 = ~pi1155 & ~n27594;
  assign n27596 = ~n27593 & n27595;
  assign n27597 = ~pi0660 & ~n27529;
  assign n27598 = ~n27596 & n27597;
  assign n27599 = pi0609 & ~n27592;
  assign n27600 = ~pi0609 & ~n27512;
  assign n27601 = pi1155 & ~n27600;
  assign n27602 = ~n27599 & n27601;
  assign n27603 = pi0660 & ~n27531;
  assign n27604 = ~n27602 & n27603;
  assign n27605 = ~n27598 & ~n27604;
  assign n27606 = pi0785 & ~n27605;
  assign n27607 = ~pi0785 & ~n27592;
  assign n27608 = ~n27606 & ~n27607;
  assign n27609 = ~pi0618 & ~n27608;
  assign n27610 = ~pi1154 & ~n27577;
  assign n27611 = ~n27609 & n27610;
  assign n27612 = ~pi0627 & ~n27537;
  assign n27613 = ~n27611 & n27612;
  assign n27614 = ~pi0618 & n27513;
  assign n27615 = pi0618 & ~n27608;
  assign n27616 = pi1154 & ~n27614;
  assign n27617 = ~n27615 & n27616;
  assign n27618 = pi0627 & ~n27539;
  assign n27619 = ~n27617 & n27618;
  assign n27620 = ~n27613 & ~n27619;
  assign n27621 = pi0781 & ~n27620;
  assign n27622 = ~pi0781 & ~n27608;
  assign n27623 = ~n27621 & ~n27622;
  assign n27624 = ~pi0789 & n27623;
  assign n27625 = ~pi0619 & ~n27623;
  assign n27626 = pi0619 & n27514;
  assign n27627 = ~pi1159 & ~n27626;
  assign n27628 = ~n27625 & n27627;
  assign n27629 = ~pi0648 & ~n27545;
  assign n27630 = ~n27628 & n27629;
  assign n27631 = pi0619 & ~n27623;
  assign n27632 = ~pi0619 & n27514;
  assign n27633 = pi1159 & ~n27632;
  assign n27634 = ~n27631 & n27633;
  assign n27635 = pi0648 & ~n27547;
  assign n27636 = ~n27634 & n27635;
  assign n27637 = pi0789 & ~n27630;
  assign n27638 = ~n27636 & n27637;
  assign n27639 = n17970 & ~n27624;
  assign n27640 = ~n27638 & n27639;
  assign n27641 = ~n27576 & ~n27640;
  assign n27642 = ~n20364 & ~n27641;
  assign n27643 = n17854 & ~n27553;
  assign n27644 = n20851 & n27516;
  assign n27645 = ~n27643 & ~n27644;
  assign n27646 = ~pi0629 & ~n27645;
  assign n27647 = n20855 & n27516;
  assign n27648 = n17853 & ~n27553;
  assign n27649 = ~n27647 & ~n27648;
  assign n27650 = pi0629 & ~n27649;
  assign n27651 = ~n27646 & ~n27650;
  assign n27652 = pi0792 & ~n27651;
  assign n27653 = ~n20206 & ~n27652;
  assign n27654 = ~n27642 & n27653;
  assign n27655 = ~n27564 & ~n27654;
  assign n27656 = ~pi0790 & n27655;
  assign n27657 = ~pi0787 & ~n27517;
  assign n27658 = pi1157 & ~n27560;
  assign n27659 = ~n27521 & ~n27658;
  assign n27660 = pi0787 & ~n27659;
  assign n27661 = ~n27657 & ~n27660;
  assign n27662 = ~pi0644 & n27661;
  assign n27663 = pi0644 & n27655;
  assign n27664 = pi0715 & ~n27662;
  assign n27665 = ~n27663 & n27664;
  assign n27666 = ~n17804 & ~n27556;
  assign n27667 = n17804 & n27501;
  assign n27668 = ~n27666 & ~n27667;
  assign n27669 = pi0644 & ~n27668;
  assign n27670 = ~pi0644 & n27501;
  assign n27671 = ~pi0715 & ~n27670;
  assign n27672 = ~n27669 & n27671;
  assign n27673 = pi1160 & ~n27672;
  assign n27674 = ~n27665 & n27673;
  assign n27675 = ~pi0644 & ~n27668;
  assign n27676 = pi0644 & n27501;
  assign n27677 = pi0715 & ~n27676;
  assign n27678 = ~n27675 & n27677;
  assign n27679 = pi0644 & n27661;
  assign n27680 = ~pi0644 & n27655;
  assign n27681 = ~pi0715 & ~n27679;
  assign n27682 = ~n27680 & n27681;
  assign n27683 = ~pi1160 & ~n27678;
  assign n27684 = ~n27682 & n27683;
  assign n27685 = ~n27674 & ~n27684;
  assign n27686 = pi0790 & ~n27685;
  assign n27687 = pi0832 & ~n27656;
  assign n27688 = ~n27686 & n27687;
  assign n27689 = ~pi0183 & po1038;
  assign n27690 = ~pi0183 & ~n17059;
  assign n27691 = n16635 & ~n27690;
  assign n27692 = ~pi0725 & n2571;
  assign n27693 = n27690 & ~n27692;
  assign n27694 = ~pi0183 & ~n16641;
  assign n27695 = n16647 & ~n27694;
  assign n27696 = pi0183 & ~n18076;
  assign n27697 = ~pi0038 & ~n27696;
  assign n27698 = n2571 & ~n27697;
  assign n27699 = ~pi0183 & n18072;
  assign n27700 = ~n27698 & ~n27699;
  assign n27701 = ~pi0725 & ~n27695;
  assign n27702 = ~n27700 & n27701;
  assign n27703 = ~n27693 & ~n27702;
  assign n27704 = ~pi0778 & n27703;
  assign n27705 = ~pi0625 & n27690;
  assign n27706 = pi0625 & ~n27703;
  assign n27707 = pi1153 & ~n27705;
  assign n27708 = ~n27706 & n27707;
  assign n27709 = pi0625 & n27690;
  assign n27710 = ~pi0625 & ~n27703;
  assign n27711 = ~pi1153 & ~n27709;
  assign n27712 = ~n27710 & n27711;
  assign n27713 = ~n27708 & ~n27712;
  assign n27714 = pi0778 & ~n27713;
  assign n27715 = ~n27704 & ~n27714;
  assign n27716 = ~n17075 & ~n27715;
  assign n27717 = n17075 & ~n27690;
  assign n27718 = ~n27716 & ~n27717;
  assign n27719 = ~n16639 & n27718;
  assign n27720 = n16639 & n27690;
  assign n27721 = ~n27719 & ~n27720;
  assign n27722 = ~n16635 & n27721;
  assign n27723 = ~n27691 & ~n27722;
  assign n27724 = ~n16631 & n27723;
  assign n27725 = n16631 & n27690;
  assign n27726 = ~n27724 & ~n27725;
  assign n27727 = ~pi0792 & n27726;
  assign n27728 = pi0628 & ~n27726;
  assign n27729 = ~pi0628 & n27690;
  assign n27730 = pi1156 & ~n27729;
  assign n27731 = ~n27728 & n27730;
  assign n27732 = pi0628 & n27690;
  assign n27733 = ~pi0628 & ~n27726;
  assign n27734 = ~pi1156 & ~n27732;
  assign n27735 = ~n27733 & n27734;
  assign n27736 = ~n27731 & ~n27735;
  assign n27737 = pi0792 & ~n27736;
  assign n27738 = ~n27727 & ~n27737;
  assign n27739 = ~pi0647 & ~n27738;
  assign n27740 = pi0647 & ~n27690;
  assign n27741 = ~n27739 & ~n27740;
  assign n27742 = ~pi1157 & n27741;
  assign n27743 = pi0647 & ~n27738;
  assign n27744 = ~pi0647 & ~n27690;
  assign n27745 = ~n27743 & ~n27744;
  assign n27746 = pi1157 & n27745;
  assign n27747 = ~n27742 & ~n27746;
  assign n27748 = pi0787 & ~n27747;
  assign n27749 = ~pi0787 & n27738;
  assign n27750 = ~n27748 & ~n27749;
  assign n27751 = ~pi0644 & ~n27750;
  assign n27752 = pi0715 & ~n27751;
  assign n27753 = pi0183 & ~n2571;
  assign n27754 = ~pi0755 & n17280;
  assign n27755 = ~n27694 & ~n27754;
  assign n27756 = pi0038 & ~n27755;
  assign n27757 = ~pi0183 & n17221;
  assign n27758 = pi0183 & ~n17275;
  assign n27759 = ~pi0755 & ~n27758;
  assign n27760 = ~n27757 & n27759;
  assign n27761 = ~pi0183 & pi0755;
  assign n27762 = ~n17048 & n27761;
  assign n27763 = ~n27760 & ~n27762;
  assign n27764 = ~pi0038 & ~n27763;
  assign n27765 = ~n27756 & ~n27764;
  assign n27766 = n2571 & n27765;
  assign n27767 = ~n27753 & ~n27766;
  assign n27768 = ~n17117 & ~n27767;
  assign n27769 = n17117 & ~n27690;
  assign n27770 = ~n27768 & ~n27769;
  assign n27771 = ~pi0785 & ~n27770;
  assign n27772 = ~n17291 & ~n27690;
  assign n27773 = pi0609 & n27768;
  assign n27774 = ~n27772 & ~n27773;
  assign n27775 = pi1155 & ~n27774;
  assign n27776 = ~n17296 & ~n27690;
  assign n27777 = ~pi0609 & n27768;
  assign n27778 = ~n27776 & ~n27777;
  assign n27779 = ~pi1155 & ~n27778;
  assign n27780 = ~n27775 & ~n27779;
  assign n27781 = pi0785 & ~n27780;
  assign n27782 = ~n27771 & ~n27781;
  assign n27783 = ~pi0781 & ~n27782;
  assign n27784 = ~pi0618 & n27690;
  assign n27785 = pi0618 & n27782;
  assign n27786 = pi1154 & ~n27784;
  assign n27787 = ~n27785 & n27786;
  assign n27788 = ~pi0618 & n27782;
  assign n27789 = pi0618 & n27690;
  assign n27790 = ~pi1154 & ~n27789;
  assign n27791 = ~n27788 & n27790;
  assign n27792 = ~n27787 & ~n27791;
  assign n27793 = pi0781 & ~n27792;
  assign n27794 = ~n27783 & ~n27793;
  assign n27795 = ~pi0789 & ~n27794;
  assign n27796 = ~pi0619 & n27690;
  assign n27797 = pi0619 & n27794;
  assign n27798 = pi1159 & ~n27796;
  assign n27799 = ~n27797 & n27798;
  assign n27800 = ~pi0619 & n27794;
  assign n27801 = pi0619 & n27690;
  assign n27802 = ~pi1159 & ~n27801;
  assign n27803 = ~n27800 & n27802;
  assign n27804 = ~n27799 & ~n27803;
  assign n27805 = pi0789 & ~n27804;
  assign n27806 = ~n27795 & ~n27805;
  assign n27807 = ~n17969 & n27806;
  assign n27808 = n17969 & n27690;
  assign n27809 = ~n27807 & ~n27808;
  assign n27810 = ~n17779 & ~n27809;
  assign n27811 = n17779 & n27690;
  assign n27812 = ~n27810 & ~n27811;
  assign n27813 = ~n17804 & ~n27812;
  assign n27814 = n17804 & n27690;
  assign n27815 = ~n27813 & ~n27814;
  assign n27816 = pi0644 & ~n27815;
  assign n27817 = ~pi0644 & n27690;
  assign n27818 = ~pi0715 & ~n27817;
  assign n27819 = ~n27816 & n27818;
  assign n27820 = pi1160 & ~n27819;
  assign n27821 = ~n27752 & n27820;
  assign n27822 = pi0644 & ~n27750;
  assign n27823 = ~pi0715 & ~n27822;
  assign n27824 = ~pi0644 & ~n27815;
  assign n27825 = pi0644 & n27690;
  assign n27826 = pi0715 & ~n27825;
  assign n27827 = ~n27824 & n27826;
  assign n27828 = ~pi1160 & ~n27827;
  assign n27829 = ~n27823 & n27828;
  assign n27830 = ~n27821 & ~n27829;
  assign n27831 = pi0790 & ~n27830;
  assign n27832 = ~pi0629 & n27731;
  assign n27833 = ~n20570 & n27809;
  assign n27834 = pi0629 & n27735;
  assign n27835 = ~n27832 & ~n27834;
  assign n27836 = ~n27833 & n27835;
  assign n27837 = pi0792 & ~n27836;
  assign n27838 = pi0609 & n27715;
  assign n27839 = pi0183 & ~n17625;
  assign n27840 = ~pi0183 & ~n17612;
  assign n27841 = pi0755 & ~n27839;
  assign n27842 = ~n27840 & n27841;
  assign n27843 = ~pi0183 & n17629;
  assign n27844 = pi0183 & n17631;
  assign n27845 = ~pi0755 & ~n27844;
  assign n27846 = ~n27843 & n27845;
  assign n27847 = ~n27842 & ~n27846;
  assign n27848 = ~pi0039 & ~n27847;
  assign n27849 = pi0183 & n17605;
  assign n27850 = ~pi0183 & ~n17546;
  assign n27851 = ~pi0755 & ~n27850;
  assign n27852 = ~n27849 & n27851;
  assign n27853 = ~pi0183 & n17404;
  assign n27854 = pi0183 & n17485;
  assign n27855 = pi0755 & ~n27854;
  assign n27856 = ~n27853 & n27855;
  assign n27857 = pi0039 & ~n27852;
  assign n27858 = ~n27856 & n27857;
  assign n27859 = ~pi0038 & ~n27848;
  assign n27860 = ~n27858 & n27859;
  assign n27861 = ~pi0755 & ~n17490;
  assign n27862 = n19471 & ~n27861;
  assign n27863 = ~pi0183 & ~n27862;
  assign n27864 = ~n17469 & ~n27523;
  assign n27865 = pi0183 & ~n27864;
  assign n27866 = n6284 & n27865;
  assign n27867 = pi0038 & ~n27866;
  assign n27868 = ~n27863 & n27867;
  assign n27869 = ~pi0725 & ~n27868;
  assign n27870 = ~n27860 & n27869;
  assign n27871 = pi0725 & ~n27765;
  assign n27872 = n2571 & ~n27870;
  assign n27873 = ~n27871 & n27872;
  assign n27874 = ~n27753 & ~n27873;
  assign n27875 = ~pi0625 & n27874;
  assign n27876 = pi0625 & n27767;
  assign n27877 = ~pi1153 & ~n27876;
  assign n27878 = ~n27875 & n27877;
  assign n27879 = ~pi0608 & ~n27708;
  assign n27880 = ~n27878 & n27879;
  assign n27881 = ~pi0625 & n27767;
  assign n27882 = pi0625 & n27874;
  assign n27883 = pi1153 & ~n27881;
  assign n27884 = ~n27882 & n27883;
  assign n27885 = pi0608 & ~n27712;
  assign n27886 = ~n27884 & n27885;
  assign n27887 = ~n27880 & ~n27886;
  assign n27888 = pi0778 & ~n27887;
  assign n27889 = ~pi0778 & n27874;
  assign n27890 = ~n27888 & ~n27889;
  assign n27891 = ~pi0609 & ~n27890;
  assign n27892 = ~pi1155 & ~n27838;
  assign n27893 = ~n27891 & n27892;
  assign n27894 = ~pi0660 & ~n27775;
  assign n27895 = ~n27893 & n27894;
  assign n27896 = ~pi0609 & n27715;
  assign n27897 = pi0609 & ~n27890;
  assign n27898 = pi1155 & ~n27896;
  assign n27899 = ~n27897 & n27898;
  assign n27900 = pi0660 & ~n27779;
  assign n27901 = ~n27899 & n27900;
  assign n27902 = ~n27895 & ~n27901;
  assign n27903 = pi0785 & ~n27902;
  assign n27904 = ~pi0785 & ~n27890;
  assign n27905 = ~n27903 & ~n27904;
  assign n27906 = ~pi0618 & ~n27905;
  assign n27907 = pi0618 & n27718;
  assign n27908 = ~pi1154 & ~n27907;
  assign n27909 = ~n27906 & n27908;
  assign n27910 = ~pi0627 & ~n27787;
  assign n27911 = ~n27909 & n27910;
  assign n27912 = ~pi0618 & n27718;
  assign n27913 = pi0618 & ~n27905;
  assign n27914 = pi1154 & ~n27912;
  assign n27915 = ~n27913 & n27914;
  assign n27916 = pi0627 & ~n27791;
  assign n27917 = ~n27915 & n27916;
  assign n27918 = ~n27911 & ~n27917;
  assign n27919 = pi0781 & ~n27918;
  assign n27920 = ~pi0781 & ~n27905;
  assign n27921 = ~n27919 & ~n27920;
  assign n27922 = ~pi0789 & n27921;
  assign n27923 = pi0619 & ~n27721;
  assign n27924 = ~pi0619 & ~n27921;
  assign n27925 = ~pi1159 & ~n27923;
  assign n27926 = ~n27924 & n27925;
  assign n27927 = ~pi0648 & ~n27799;
  assign n27928 = ~n27926 & n27927;
  assign n27929 = ~pi0619 & ~n27721;
  assign n27930 = pi0619 & ~n27921;
  assign n27931 = pi1159 & ~n27929;
  assign n27932 = ~n27930 & n27931;
  assign n27933 = pi0648 & ~n27803;
  assign n27934 = ~n27932 & n27933;
  assign n27935 = pi0789 & ~n27928;
  assign n27936 = ~n27934 & n27935;
  assign n27937 = n17970 & ~n27922;
  assign n27938 = ~n27936 & n27937;
  assign n27939 = n17871 & n27723;
  assign n27940 = ~pi0626 & ~n27806;
  assign n27941 = pi0626 & ~n27690;
  assign n27942 = n16629 & ~n27941;
  assign n27943 = ~n27940 & n27942;
  assign n27944 = pi0626 & ~n27806;
  assign n27945 = ~pi0626 & ~n27690;
  assign n27946 = n16628 & ~n27945;
  assign n27947 = ~n27944 & n27946;
  assign n27948 = ~n27939 & ~n27943;
  assign n27949 = ~n27947 & n27948;
  assign n27950 = pi0788 & ~n27949;
  assign n27951 = ~n20364 & ~n27950;
  assign n27952 = ~n27938 & n27951;
  assign n27953 = ~n27837 & ~n27952;
  assign n27954 = ~n20206 & ~n27953;
  assign n27955 = n17802 & ~n27741;
  assign n27956 = ~n20559 & n27812;
  assign n27957 = n17801 & ~n27745;
  assign n27958 = ~n27955 & ~n27957;
  assign n27959 = ~n27956 & n27958;
  assign n27960 = pi0787 & ~n27959;
  assign n27961 = ~pi0644 & n27828;
  assign n27962 = pi0644 & n27820;
  assign n27963 = pi0790 & ~n27961;
  assign n27964 = ~n27962 & n27963;
  assign n27965 = ~n27954 & ~n27960;
  assign n27966 = ~n27964 & n27965;
  assign n27967 = ~n27831 & ~n27966;
  assign n27968 = ~po1038 & ~n27967;
  assign n27969 = ~pi0832 & ~n27689;
  assign n27970 = ~n27968 & n27969;
  assign po0340 = ~n27688 & ~n27970;
  assign n27972 = ~pi0184 & ~n2926;
  assign n27973 = ~pi0737 & n16645;
  assign n27974 = ~n27972 & ~n27973;
  assign n27975 = ~pi0778 & ~n27974;
  assign n27976 = ~pi0625 & n27973;
  assign n27977 = ~n27974 & ~n27976;
  assign n27978 = pi1153 & ~n27977;
  assign n27979 = ~pi1153 & ~n27972;
  assign n27980 = ~n27976 & n27979;
  assign n27981 = pi0778 & ~n27980;
  assign n27982 = ~n27978 & n27981;
  assign n27983 = ~n27975 & ~n27982;
  assign n27984 = ~n17845 & ~n27983;
  assign n27985 = ~n17847 & n27984;
  assign n27986 = ~n17849 & n27985;
  assign n27987 = ~n17851 & n27986;
  assign n27988 = ~n17857 & n27987;
  assign n27989 = ~pi0647 & n27988;
  assign n27990 = pi0647 & n27972;
  assign n27991 = ~pi1157 & ~n27990;
  assign n27992 = ~n27989 & n27991;
  assign n27993 = pi0630 & n27992;
  assign n27994 = ~pi0777 & n17244;
  assign n27995 = ~n27972 & ~n27994;
  assign n27996 = ~n17874 & ~n27995;
  assign n27997 = ~pi0785 & ~n27996;
  assign n27998 = n17296 & n27994;
  assign n27999 = n27996 & ~n27998;
  assign n28000 = pi1155 & ~n27999;
  assign n28001 = ~pi1155 & ~n27972;
  assign n28002 = ~n27998 & n28001;
  assign n28003 = ~n28000 & ~n28002;
  assign n28004 = pi0785 & ~n28003;
  assign n28005 = ~n27997 & ~n28004;
  assign n28006 = ~pi0781 & ~n28005;
  assign n28007 = ~n17889 & n28005;
  assign n28008 = pi1154 & ~n28007;
  assign n28009 = ~n17892 & n28005;
  assign n28010 = ~pi1154 & ~n28009;
  assign n28011 = ~n28008 & ~n28010;
  assign n28012 = pi0781 & ~n28011;
  assign n28013 = ~n28006 & ~n28012;
  assign n28014 = ~pi0789 & ~n28013;
  assign n28015 = ~n23078 & n28013;
  assign n28016 = pi1159 & ~n28015;
  assign n28017 = ~n23081 & n28013;
  assign n28018 = ~pi1159 & ~n28017;
  assign n28019 = ~n28016 & ~n28018;
  assign n28020 = pi0789 & ~n28019;
  assign n28021 = ~n28014 & ~n28020;
  assign n28022 = ~n17969 & n28021;
  assign n28023 = n17969 & n27972;
  assign n28024 = ~n28022 & ~n28023;
  assign n28025 = ~n17779 & ~n28024;
  assign n28026 = n17779 & n27972;
  assign n28027 = ~n28025 & ~n28026;
  assign n28028 = ~n20559 & n28027;
  assign n28029 = pi0647 & ~n27988;
  assign n28030 = ~pi0647 & ~n27972;
  assign n28031 = ~n28029 & ~n28030;
  assign n28032 = n17801 & ~n28031;
  assign n28033 = ~n27993 & ~n28032;
  assign n28034 = ~n28028 & n28033;
  assign n28035 = pi0787 & ~n28034;
  assign n28036 = n17871 & n27986;
  assign n28037 = ~pi0626 & ~n28021;
  assign n28038 = pi0626 & ~n27972;
  assign n28039 = n16629 & ~n28038;
  assign n28040 = ~n28037 & n28039;
  assign n28041 = pi0626 & ~n28021;
  assign n28042 = ~pi0626 & ~n27972;
  assign n28043 = n16628 & ~n28042;
  assign n28044 = ~n28041 & n28043;
  assign n28045 = ~n28036 & ~n28040;
  assign n28046 = ~n28044 & n28045;
  assign n28047 = pi0788 & ~n28046;
  assign n28048 = pi0618 & n27984;
  assign n28049 = ~n17168 & ~n27974;
  assign n28050 = pi0625 & n28049;
  assign n28051 = n27995 & ~n28049;
  assign n28052 = ~n28050 & ~n28051;
  assign n28053 = n27979 & ~n28052;
  assign n28054 = ~pi0608 & ~n27978;
  assign n28055 = ~n28053 & n28054;
  assign n28056 = pi1153 & n27995;
  assign n28057 = ~n28050 & n28056;
  assign n28058 = pi0608 & ~n27980;
  assign n28059 = ~n28057 & n28058;
  assign n28060 = ~n28055 & ~n28059;
  assign n28061 = pi0778 & ~n28060;
  assign n28062 = ~pi0778 & ~n28051;
  assign n28063 = ~n28061 & ~n28062;
  assign n28064 = ~pi0609 & ~n28063;
  assign n28065 = pi0609 & ~n27983;
  assign n28066 = ~pi1155 & ~n28065;
  assign n28067 = ~n28064 & n28066;
  assign n28068 = ~pi0660 & ~n28000;
  assign n28069 = ~n28067 & n28068;
  assign n28070 = pi0609 & ~n28063;
  assign n28071 = ~pi0609 & ~n27983;
  assign n28072 = pi1155 & ~n28071;
  assign n28073 = ~n28070 & n28072;
  assign n28074 = pi0660 & ~n28002;
  assign n28075 = ~n28073 & n28074;
  assign n28076 = ~n28069 & ~n28075;
  assign n28077 = pi0785 & ~n28076;
  assign n28078 = ~pi0785 & ~n28063;
  assign n28079 = ~n28077 & ~n28078;
  assign n28080 = ~pi0618 & ~n28079;
  assign n28081 = ~pi1154 & ~n28048;
  assign n28082 = ~n28080 & n28081;
  assign n28083 = ~pi0627 & ~n28008;
  assign n28084 = ~n28082 & n28083;
  assign n28085 = ~pi0618 & n27984;
  assign n28086 = pi0618 & ~n28079;
  assign n28087 = pi1154 & ~n28085;
  assign n28088 = ~n28086 & n28087;
  assign n28089 = pi0627 & ~n28010;
  assign n28090 = ~n28088 & n28089;
  assign n28091 = ~n28084 & ~n28090;
  assign n28092 = pi0781 & ~n28091;
  assign n28093 = ~pi0781 & ~n28079;
  assign n28094 = ~n28092 & ~n28093;
  assign n28095 = ~pi0789 & n28094;
  assign n28096 = ~pi0619 & ~n28094;
  assign n28097 = pi0619 & n27985;
  assign n28098 = ~pi1159 & ~n28097;
  assign n28099 = ~n28096 & n28098;
  assign n28100 = ~pi0648 & ~n28016;
  assign n28101 = ~n28099 & n28100;
  assign n28102 = pi0619 & ~n28094;
  assign n28103 = ~pi0619 & n27985;
  assign n28104 = pi1159 & ~n28103;
  assign n28105 = ~n28102 & n28104;
  assign n28106 = pi0648 & ~n28018;
  assign n28107 = ~n28105 & n28106;
  assign n28108 = pi0789 & ~n28101;
  assign n28109 = ~n28107 & n28108;
  assign n28110 = n17970 & ~n28095;
  assign n28111 = ~n28109 & n28110;
  assign n28112 = ~n28047 & ~n28111;
  assign n28113 = ~n20364 & ~n28112;
  assign n28114 = n17854 & ~n28024;
  assign n28115 = n20851 & n27987;
  assign n28116 = ~n28114 & ~n28115;
  assign n28117 = ~pi0629 & ~n28116;
  assign n28118 = n20855 & n27987;
  assign n28119 = n17853 & ~n28024;
  assign n28120 = ~n28118 & ~n28119;
  assign n28121 = pi0629 & ~n28120;
  assign n28122 = ~n28117 & ~n28121;
  assign n28123 = pi0792 & ~n28122;
  assign n28124 = ~n20206 & ~n28123;
  assign n28125 = ~n28113 & n28124;
  assign n28126 = ~n28035 & ~n28125;
  assign n28127 = ~pi0790 & n28126;
  assign n28128 = ~pi0787 & ~n27988;
  assign n28129 = pi1157 & ~n28031;
  assign n28130 = ~n27992 & ~n28129;
  assign n28131 = pi0787 & ~n28130;
  assign n28132 = ~n28128 & ~n28131;
  assign n28133 = ~pi0644 & n28132;
  assign n28134 = pi0644 & n28126;
  assign n28135 = pi0715 & ~n28133;
  assign n28136 = ~n28134 & n28135;
  assign n28137 = ~n17804 & ~n28027;
  assign n28138 = n17804 & n27972;
  assign n28139 = ~n28137 & ~n28138;
  assign n28140 = pi0644 & ~n28139;
  assign n28141 = ~pi0644 & n27972;
  assign n28142 = ~pi0715 & ~n28141;
  assign n28143 = ~n28140 & n28142;
  assign n28144 = pi1160 & ~n28143;
  assign n28145 = ~n28136 & n28144;
  assign n28146 = ~pi0644 & ~n28139;
  assign n28147 = pi0644 & n27972;
  assign n28148 = pi0715 & ~n28147;
  assign n28149 = ~n28146 & n28148;
  assign n28150 = pi0644 & n28132;
  assign n28151 = ~pi0644 & n28126;
  assign n28152 = ~pi0715 & ~n28150;
  assign n28153 = ~n28151 & n28152;
  assign n28154 = ~pi1160 & ~n28149;
  assign n28155 = ~n28153 & n28154;
  assign n28156 = ~n28145 & ~n28155;
  assign n28157 = pi0790 & ~n28156;
  assign n28158 = pi0832 & ~n28127;
  assign n28159 = ~n28157 & n28158;
  assign n28160 = ~pi0184 & po1038;
  assign n28161 = ~pi0184 & ~n17059;
  assign n28162 = n16635 & ~n28161;
  assign n28163 = ~pi0737 & n2571;
  assign n28164 = n28161 & ~n28163;
  assign n28165 = ~pi0184 & ~n16641;
  assign n28166 = n16647 & ~n28165;
  assign n28167 = pi0184 & ~n18076;
  assign n28168 = ~pi0038 & ~n28167;
  assign n28169 = n2571 & ~n28168;
  assign n28170 = ~pi0184 & n18072;
  assign n28171 = ~n28169 & ~n28170;
  assign n28172 = ~pi0737 & ~n28166;
  assign n28173 = ~n28171 & n28172;
  assign n28174 = ~n28164 & ~n28173;
  assign n28175 = ~pi0778 & n28174;
  assign n28176 = ~pi0625 & n28161;
  assign n28177 = pi0625 & ~n28174;
  assign n28178 = pi1153 & ~n28176;
  assign n28179 = ~n28177 & n28178;
  assign n28180 = pi0625 & n28161;
  assign n28181 = ~pi0625 & ~n28174;
  assign n28182 = ~pi1153 & ~n28180;
  assign n28183 = ~n28181 & n28182;
  assign n28184 = ~n28179 & ~n28183;
  assign n28185 = pi0778 & ~n28184;
  assign n28186 = ~n28175 & ~n28185;
  assign n28187 = ~n17075 & ~n28186;
  assign n28188 = n17075 & ~n28161;
  assign n28189 = ~n28187 & ~n28188;
  assign n28190 = ~n16639 & n28189;
  assign n28191 = n16639 & n28161;
  assign n28192 = ~n28190 & ~n28191;
  assign n28193 = ~n16635 & n28192;
  assign n28194 = ~n28162 & ~n28193;
  assign n28195 = ~n16631 & n28194;
  assign n28196 = n16631 & n28161;
  assign n28197 = ~n28195 & ~n28196;
  assign n28198 = ~pi0792 & n28197;
  assign n28199 = pi0628 & ~n28197;
  assign n28200 = ~pi0628 & n28161;
  assign n28201 = pi1156 & ~n28200;
  assign n28202 = ~n28199 & n28201;
  assign n28203 = pi0628 & n28161;
  assign n28204 = ~pi0628 & ~n28197;
  assign n28205 = ~pi1156 & ~n28203;
  assign n28206 = ~n28204 & n28205;
  assign n28207 = ~n28202 & ~n28206;
  assign n28208 = pi0792 & ~n28207;
  assign n28209 = ~n28198 & ~n28208;
  assign n28210 = ~pi0647 & ~n28209;
  assign n28211 = pi0647 & ~n28161;
  assign n28212 = ~n28210 & ~n28211;
  assign n28213 = ~pi1157 & n28212;
  assign n28214 = pi0647 & ~n28209;
  assign n28215 = ~pi0647 & ~n28161;
  assign n28216 = ~n28214 & ~n28215;
  assign n28217 = pi1157 & n28216;
  assign n28218 = ~n28213 & ~n28217;
  assign n28219 = pi0787 & ~n28218;
  assign n28220 = ~pi0787 & n28209;
  assign n28221 = ~n28219 & ~n28220;
  assign n28222 = ~pi0644 & ~n28221;
  assign n28223 = pi0715 & ~n28222;
  assign n28224 = pi0184 & ~n2571;
  assign n28225 = ~pi0777 & n17280;
  assign n28226 = ~n28165 & ~n28225;
  assign n28227 = pi0038 & ~n28226;
  assign n28228 = ~pi0184 & n17221;
  assign n28229 = pi0184 & ~n17275;
  assign n28230 = ~pi0777 & ~n28229;
  assign n28231 = ~n28228 & n28230;
  assign n28232 = ~pi0184 & pi0777;
  assign n28233 = ~n17048 & n28232;
  assign n28234 = ~n28231 & ~n28233;
  assign n28235 = ~pi0038 & ~n28234;
  assign n28236 = ~n28227 & ~n28235;
  assign n28237 = n2571 & n28236;
  assign n28238 = ~n28224 & ~n28237;
  assign n28239 = ~n17117 & ~n28238;
  assign n28240 = n17117 & ~n28161;
  assign n28241 = ~n28239 & ~n28240;
  assign n28242 = ~pi0785 & ~n28241;
  assign n28243 = ~n17291 & ~n28161;
  assign n28244 = pi0609 & n28239;
  assign n28245 = ~n28243 & ~n28244;
  assign n28246 = pi1155 & ~n28245;
  assign n28247 = ~n17296 & ~n28161;
  assign n28248 = ~pi0609 & n28239;
  assign n28249 = ~n28247 & ~n28248;
  assign n28250 = ~pi1155 & ~n28249;
  assign n28251 = ~n28246 & ~n28250;
  assign n28252 = pi0785 & ~n28251;
  assign n28253 = ~n28242 & ~n28252;
  assign n28254 = ~pi0781 & ~n28253;
  assign n28255 = ~pi0618 & n28161;
  assign n28256 = pi0618 & n28253;
  assign n28257 = pi1154 & ~n28255;
  assign n28258 = ~n28256 & n28257;
  assign n28259 = ~pi0618 & n28253;
  assign n28260 = pi0618 & n28161;
  assign n28261 = ~pi1154 & ~n28260;
  assign n28262 = ~n28259 & n28261;
  assign n28263 = ~n28258 & ~n28262;
  assign n28264 = pi0781 & ~n28263;
  assign n28265 = ~n28254 & ~n28264;
  assign n28266 = ~pi0789 & ~n28265;
  assign n28267 = ~pi0619 & n28161;
  assign n28268 = pi0619 & n28265;
  assign n28269 = pi1159 & ~n28267;
  assign n28270 = ~n28268 & n28269;
  assign n28271 = ~pi0619 & n28265;
  assign n28272 = pi0619 & n28161;
  assign n28273 = ~pi1159 & ~n28272;
  assign n28274 = ~n28271 & n28273;
  assign n28275 = ~n28270 & ~n28274;
  assign n28276 = pi0789 & ~n28275;
  assign n28277 = ~n28266 & ~n28276;
  assign n28278 = ~n17969 & n28277;
  assign n28279 = n17969 & n28161;
  assign n28280 = ~n28278 & ~n28279;
  assign n28281 = ~n17779 & ~n28280;
  assign n28282 = n17779 & n28161;
  assign n28283 = ~n28281 & ~n28282;
  assign n28284 = ~n17804 & ~n28283;
  assign n28285 = n17804 & n28161;
  assign n28286 = ~n28284 & ~n28285;
  assign n28287 = pi0644 & ~n28286;
  assign n28288 = ~pi0644 & n28161;
  assign n28289 = ~pi0715 & ~n28288;
  assign n28290 = ~n28287 & n28289;
  assign n28291 = pi1160 & ~n28290;
  assign n28292 = ~n28223 & n28291;
  assign n28293 = pi0644 & ~n28221;
  assign n28294 = ~pi0715 & ~n28293;
  assign n28295 = ~pi0644 & ~n28286;
  assign n28296 = pi0644 & n28161;
  assign n28297 = pi0715 & ~n28296;
  assign n28298 = ~n28295 & n28297;
  assign n28299 = ~pi1160 & ~n28298;
  assign n28300 = ~n28294 & n28299;
  assign n28301 = ~n28292 & ~n28300;
  assign n28302 = pi0790 & ~n28301;
  assign n28303 = ~pi0629 & n28202;
  assign n28304 = ~n20570 & n28280;
  assign n28305 = pi0629 & n28206;
  assign n28306 = ~n28303 & ~n28305;
  assign n28307 = ~n28304 & n28306;
  assign n28308 = pi0792 & ~n28307;
  assign n28309 = pi0609 & n28186;
  assign n28310 = pi0184 & ~n17625;
  assign n28311 = ~pi0184 & ~n17612;
  assign n28312 = pi0777 & ~n28310;
  assign n28313 = ~n28311 & n28312;
  assign n28314 = ~pi0184 & n17629;
  assign n28315 = pi0184 & n17631;
  assign n28316 = ~pi0777 & ~n28315;
  assign n28317 = ~n28314 & n28316;
  assign n28318 = ~n28313 & ~n28317;
  assign n28319 = ~pi0039 & ~n28318;
  assign n28320 = pi0184 & n17605;
  assign n28321 = ~pi0184 & ~n17546;
  assign n28322 = ~pi0777 & ~n28321;
  assign n28323 = ~n28320 & n28322;
  assign n28324 = ~pi0184 & n17404;
  assign n28325 = pi0184 & n17485;
  assign n28326 = pi0777 & ~n28325;
  assign n28327 = ~n28324 & n28326;
  assign n28328 = pi0039 & ~n28323;
  assign n28329 = ~n28327 & n28328;
  assign n28330 = ~pi0038 & ~n28319;
  assign n28331 = ~n28329 & n28330;
  assign n28332 = ~pi0777 & ~n17490;
  assign n28333 = n19471 & ~n28332;
  assign n28334 = ~pi0184 & ~n28333;
  assign n28335 = ~n17469 & ~n27994;
  assign n28336 = pi0184 & ~n28335;
  assign n28337 = n6284 & n28336;
  assign n28338 = pi0038 & ~n28337;
  assign n28339 = ~n28334 & n28338;
  assign n28340 = ~pi0737 & ~n28339;
  assign n28341 = ~n28331 & n28340;
  assign n28342 = pi0737 & ~n28236;
  assign n28343 = n2571 & ~n28341;
  assign n28344 = ~n28342 & n28343;
  assign n28345 = ~n28224 & ~n28344;
  assign n28346 = ~pi0625 & n28345;
  assign n28347 = pi0625 & n28238;
  assign n28348 = ~pi1153 & ~n28347;
  assign n28349 = ~n28346 & n28348;
  assign n28350 = ~pi0608 & ~n28179;
  assign n28351 = ~n28349 & n28350;
  assign n28352 = ~pi0625 & n28238;
  assign n28353 = pi0625 & n28345;
  assign n28354 = pi1153 & ~n28352;
  assign n28355 = ~n28353 & n28354;
  assign n28356 = pi0608 & ~n28183;
  assign n28357 = ~n28355 & n28356;
  assign n28358 = ~n28351 & ~n28357;
  assign n28359 = pi0778 & ~n28358;
  assign n28360 = ~pi0778 & n28345;
  assign n28361 = ~n28359 & ~n28360;
  assign n28362 = ~pi0609 & ~n28361;
  assign n28363 = ~pi1155 & ~n28309;
  assign n28364 = ~n28362 & n28363;
  assign n28365 = ~pi0660 & ~n28246;
  assign n28366 = ~n28364 & n28365;
  assign n28367 = ~pi0609 & n28186;
  assign n28368 = pi0609 & ~n28361;
  assign n28369 = pi1155 & ~n28367;
  assign n28370 = ~n28368 & n28369;
  assign n28371 = pi0660 & ~n28250;
  assign n28372 = ~n28370 & n28371;
  assign n28373 = ~n28366 & ~n28372;
  assign n28374 = pi0785 & ~n28373;
  assign n28375 = ~pi0785 & ~n28361;
  assign n28376 = ~n28374 & ~n28375;
  assign n28377 = ~pi0618 & ~n28376;
  assign n28378 = pi0618 & n28189;
  assign n28379 = ~pi1154 & ~n28378;
  assign n28380 = ~n28377 & n28379;
  assign n28381 = ~pi0627 & ~n28258;
  assign n28382 = ~n28380 & n28381;
  assign n28383 = ~pi0618 & n28189;
  assign n28384 = pi0618 & ~n28376;
  assign n28385 = pi1154 & ~n28383;
  assign n28386 = ~n28384 & n28385;
  assign n28387 = pi0627 & ~n28262;
  assign n28388 = ~n28386 & n28387;
  assign n28389 = ~n28382 & ~n28388;
  assign n28390 = pi0781 & ~n28389;
  assign n28391 = ~pi0781 & ~n28376;
  assign n28392 = ~n28390 & ~n28391;
  assign n28393 = ~pi0789 & n28392;
  assign n28394 = pi0619 & ~n28192;
  assign n28395 = ~pi0619 & ~n28392;
  assign n28396 = ~pi1159 & ~n28394;
  assign n28397 = ~n28395 & n28396;
  assign n28398 = ~pi0648 & ~n28270;
  assign n28399 = ~n28397 & n28398;
  assign n28400 = ~pi0619 & ~n28192;
  assign n28401 = pi0619 & ~n28392;
  assign n28402 = pi1159 & ~n28400;
  assign n28403 = ~n28401 & n28402;
  assign n28404 = pi0648 & ~n28274;
  assign n28405 = ~n28403 & n28404;
  assign n28406 = pi0789 & ~n28399;
  assign n28407 = ~n28405 & n28406;
  assign n28408 = n17970 & ~n28393;
  assign n28409 = ~n28407 & n28408;
  assign n28410 = n17871 & n28194;
  assign n28411 = ~pi0626 & ~n28277;
  assign n28412 = pi0626 & ~n28161;
  assign n28413 = n16629 & ~n28412;
  assign n28414 = ~n28411 & n28413;
  assign n28415 = pi0626 & ~n28277;
  assign n28416 = ~pi0626 & ~n28161;
  assign n28417 = n16628 & ~n28416;
  assign n28418 = ~n28415 & n28417;
  assign n28419 = ~n28410 & ~n28414;
  assign n28420 = ~n28418 & n28419;
  assign n28421 = pi0788 & ~n28420;
  assign n28422 = ~n20364 & ~n28421;
  assign n28423 = ~n28409 & n28422;
  assign n28424 = ~n28308 & ~n28423;
  assign n28425 = ~n20206 & ~n28424;
  assign n28426 = n17802 & ~n28212;
  assign n28427 = ~n20559 & n28283;
  assign n28428 = n17801 & ~n28216;
  assign n28429 = ~n28426 & ~n28428;
  assign n28430 = ~n28427 & n28429;
  assign n28431 = pi0787 & ~n28430;
  assign n28432 = ~pi0644 & n28299;
  assign n28433 = pi0644 & n28291;
  assign n28434 = pi0790 & ~n28432;
  assign n28435 = ~n28433 & n28434;
  assign n28436 = ~n28425 & ~n28431;
  assign n28437 = ~n28435 & n28436;
  assign n28438 = ~n28302 & ~n28437;
  assign n28439 = ~po1038 & ~n28438;
  assign n28440 = ~pi0832 & ~n28160;
  assign n28441 = ~n28439 & n28440;
  assign po0341 = ~n28159 & ~n28441;
  assign n28443 = ~pi0185 & ~n2926;
  assign n28444 = ~pi0701 & n16645;
  assign n28445 = ~n28443 & ~n28444;
  assign n28446 = ~pi0778 & ~n28445;
  assign n28447 = ~pi0625 & n28444;
  assign n28448 = ~n28445 & ~n28447;
  assign n28449 = pi1153 & ~n28448;
  assign n28450 = ~pi1153 & ~n28443;
  assign n28451 = ~n28447 & n28450;
  assign n28452 = pi0778 & ~n28451;
  assign n28453 = ~n28449 & n28452;
  assign n28454 = ~n28446 & ~n28453;
  assign n28455 = ~n17845 & ~n28454;
  assign n28456 = ~n17847 & n28455;
  assign n28457 = ~n17849 & n28456;
  assign n28458 = ~n17851 & n28457;
  assign n28459 = ~n17857 & n28458;
  assign n28460 = ~pi0647 & n28459;
  assign n28461 = pi0647 & n28443;
  assign n28462 = ~pi1157 & ~n28461;
  assign n28463 = ~n28460 & n28462;
  assign n28464 = pi0630 & n28463;
  assign n28465 = ~pi0751 & n17244;
  assign n28466 = ~n28443 & ~n28465;
  assign n28467 = ~n17874 & ~n28466;
  assign n28468 = ~pi0785 & ~n28467;
  assign n28469 = n17296 & n28465;
  assign n28470 = n28467 & ~n28469;
  assign n28471 = pi1155 & ~n28470;
  assign n28472 = ~pi1155 & ~n28443;
  assign n28473 = ~n28469 & n28472;
  assign n28474 = ~n28471 & ~n28473;
  assign n28475 = pi0785 & ~n28474;
  assign n28476 = ~n28468 & ~n28475;
  assign n28477 = ~pi0781 & ~n28476;
  assign n28478 = ~n17889 & n28476;
  assign n28479 = pi1154 & ~n28478;
  assign n28480 = ~n17892 & n28476;
  assign n28481 = ~pi1154 & ~n28480;
  assign n28482 = ~n28479 & ~n28481;
  assign n28483 = pi0781 & ~n28482;
  assign n28484 = ~n28477 & ~n28483;
  assign n28485 = ~pi0789 & ~n28484;
  assign n28486 = ~n23078 & n28484;
  assign n28487 = pi1159 & ~n28486;
  assign n28488 = ~n23081 & n28484;
  assign n28489 = ~pi1159 & ~n28488;
  assign n28490 = ~n28487 & ~n28489;
  assign n28491 = pi0789 & ~n28490;
  assign n28492 = ~n28485 & ~n28491;
  assign n28493 = ~n17969 & n28492;
  assign n28494 = n17969 & n28443;
  assign n28495 = ~n28493 & ~n28494;
  assign n28496 = ~n17779 & ~n28495;
  assign n28497 = n17779 & n28443;
  assign n28498 = ~n28496 & ~n28497;
  assign n28499 = ~n20559 & n28498;
  assign n28500 = pi0647 & ~n28459;
  assign n28501 = ~pi0647 & ~n28443;
  assign n28502 = ~n28500 & ~n28501;
  assign n28503 = n17801 & ~n28502;
  assign n28504 = ~n28464 & ~n28503;
  assign n28505 = ~n28499 & n28504;
  assign n28506 = pi0787 & ~n28505;
  assign n28507 = n17871 & n28457;
  assign n28508 = ~pi0626 & ~n28492;
  assign n28509 = pi0626 & ~n28443;
  assign n28510 = n16629 & ~n28509;
  assign n28511 = ~n28508 & n28510;
  assign n28512 = pi0626 & ~n28492;
  assign n28513 = ~pi0626 & ~n28443;
  assign n28514 = n16628 & ~n28513;
  assign n28515 = ~n28512 & n28514;
  assign n28516 = ~n28507 & ~n28511;
  assign n28517 = ~n28515 & n28516;
  assign n28518 = pi0788 & ~n28517;
  assign n28519 = pi0618 & n28455;
  assign n28520 = ~n17168 & ~n28445;
  assign n28521 = pi0625 & n28520;
  assign n28522 = n28466 & ~n28520;
  assign n28523 = ~n28521 & ~n28522;
  assign n28524 = n28450 & ~n28523;
  assign n28525 = ~pi0608 & ~n28449;
  assign n28526 = ~n28524 & n28525;
  assign n28527 = pi1153 & n28466;
  assign n28528 = ~n28521 & n28527;
  assign n28529 = pi0608 & ~n28451;
  assign n28530 = ~n28528 & n28529;
  assign n28531 = ~n28526 & ~n28530;
  assign n28532 = pi0778 & ~n28531;
  assign n28533 = ~pi0778 & ~n28522;
  assign n28534 = ~n28532 & ~n28533;
  assign n28535 = ~pi0609 & ~n28534;
  assign n28536 = pi0609 & ~n28454;
  assign n28537 = ~pi1155 & ~n28536;
  assign n28538 = ~n28535 & n28537;
  assign n28539 = ~pi0660 & ~n28471;
  assign n28540 = ~n28538 & n28539;
  assign n28541 = pi0609 & ~n28534;
  assign n28542 = ~pi0609 & ~n28454;
  assign n28543 = pi1155 & ~n28542;
  assign n28544 = ~n28541 & n28543;
  assign n28545 = pi0660 & ~n28473;
  assign n28546 = ~n28544 & n28545;
  assign n28547 = ~n28540 & ~n28546;
  assign n28548 = pi0785 & ~n28547;
  assign n28549 = ~pi0785 & ~n28534;
  assign n28550 = ~n28548 & ~n28549;
  assign n28551 = ~pi0618 & ~n28550;
  assign n28552 = ~pi1154 & ~n28519;
  assign n28553 = ~n28551 & n28552;
  assign n28554 = ~pi0627 & ~n28479;
  assign n28555 = ~n28553 & n28554;
  assign n28556 = ~pi0618 & n28455;
  assign n28557 = pi0618 & ~n28550;
  assign n28558 = pi1154 & ~n28556;
  assign n28559 = ~n28557 & n28558;
  assign n28560 = pi0627 & ~n28481;
  assign n28561 = ~n28559 & n28560;
  assign n28562 = ~n28555 & ~n28561;
  assign n28563 = pi0781 & ~n28562;
  assign n28564 = ~pi0781 & ~n28550;
  assign n28565 = ~n28563 & ~n28564;
  assign n28566 = ~pi0789 & n28565;
  assign n28567 = ~pi0619 & ~n28565;
  assign n28568 = pi0619 & n28456;
  assign n28569 = ~pi1159 & ~n28568;
  assign n28570 = ~n28567 & n28569;
  assign n28571 = ~pi0648 & ~n28487;
  assign n28572 = ~n28570 & n28571;
  assign n28573 = pi0619 & ~n28565;
  assign n28574 = ~pi0619 & n28456;
  assign n28575 = pi1159 & ~n28574;
  assign n28576 = ~n28573 & n28575;
  assign n28577 = pi0648 & ~n28489;
  assign n28578 = ~n28576 & n28577;
  assign n28579 = pi0789 & ~n28572;
  assign n28580 = ~n28578 & n28579;
  assign n28581 = n17970 & ~n28566;
  assign n28582 = ~n28580 & n28581;
  assign n28583 = ~n28518 & ~n28582;
  assign n28584 = ~n20364 & ~n28583;
  assign n28585 = n17854 & ~n28495;
  assign n28586 = n20851 & n28458;
  assign n28587 = ~n28585 & ~n28586;
  assign n28588 = ~pi0629 & ~n28587;
  assign n28589 = n20855 & n28458;
  assign n28590 = n17853 & ~n28495;
  assign n28591 = ~n28589 & ~n28590;
  assign n28592 = pi0629 & ~n28591;
  assign n28593 = ~n28588 & ~n28592;
  assign n28594 = pi0792 & ~n28593;
  assign n28595 = ~n20206 & ~n28594;
  assign n28596 = ~n28584 & n28595;
  assign n28597 = ~n28506 & ~n28596;
  assign n28598 = ~pi0790 & n28597;
  assign n28599 = ~pi0787 & ~n28459;
  assign n28600 = pi1157 & ~n28502;
  assign n28601 = ~n28463 & ~n28600;
  assign n28602 = pi0787 & ~n28601;
  assign n28603 = ~n28599 & ~n28602;
  assign n28604 = ~pi0644 & n28603;
  assign n28605 = pi0644 & n28597;
  assign n28606 = pi0715 & ~n28604;
  assign n28607 = ~n28605 & n28606;
  assign n28608 = ~n17804 & ~n28498;
  assign n28609 = n17804 & n28443;
  assign n28610 = ~n28608 & ~n28609;
  assign n28611 = pi0644 & ~n28610;
  assign n28612 = ~pi0644 & n28443;
  assign n28613 = ~pi0715 & ~n28612;
  assign n28614 = ~n28611 & n28613;
  assign n28615 = pi1160 & ~n28614;
  assign n28616 = ~n28607 & n28615;
  assign n28617 = ~pi0644 & ~n28610;
  assign n28618 = pi0644 & n28443;
  assign n28619 = pi0715 & ~n28618;
  assign n28620 = ~n28617 & n28619;
  assign n28621 = pi0644 & n28603;
  assign n28622 = ~pi0644 & n28597;
  assign n28623 = ~pi0715 & ~n28621;
  assign n28624 = ~n28622 & n28623;
  assign n28625 = ~pi1160 & ~n28620;
  assign n28626 = ~n28624 & n28625;
  assign n28627 = ~n28616 & ~n28626;
  assign n28628 = pi0790 & ~n28627;
  assign n28629 = pi0832 & ~n28598;
  assign n28630 = ~n28628 & n28629;
  assign n28631 = ~pi0185 & po1038;
  assign n28632 = ~pi0185 & ~n17059;
  assign n28633 = n16635 & ~n28632;
  assign n28634 = ~pi0701 & n2571;
  assign n28635 = n28632 & ~n28634;
  assign n28636 = ~pi0185 & ~n16641;
  assign n28637 = n16647 & ~n28636;
  assign n28638 = pi0185 & ~n18076;
  assign n28639 = ~pi0038 & ~n28638;
  assign n28640 = n2571 & ~n28639;
  assign n28641 = ~pi0185 & n18072;
  assign n28642 = ~n28640 & ~n28641;
  assign n28643 = ~pi0701 & ~n28637;
  assign n28644 = ~n28642 & n28643;
  assign n28645 = ~n28635 & ~n28644;
  assign n28646 = ~pi0778 & n28645;
  assign n28647 = ~pi0625 & n28632;
  assign n28648 = pi0625 & ~n28645;
  assign n28649 = pi1153 & ~n28647;
  assign n28650 = ~n28648 & n28649;
  assign n28651 = pi0625 & n28632;
  assign n28652 = ~pi0625 & ~n28645;
  assign n28653 = ~pi1153 & ~n28651;
  assign n28654 = ~n28652 & n28653;
  assign n28655 = ~n28650 & ~n28654;
  assign n28656 = pi0778 & ~n28655;
  assign n28657 = ~n28646 & ~n28656;
  assign n28658 = ~n17075 & ~n28657;
  assign n28659 = n17075 & ~n28632;
  assign n28660 = ~n28658 & ~n28659;
  assign n28661 = ~n16639 & n28660;
  assign n28662 = n16639 & n28632;
  assign n28663 = ~n28661 & ~n28662;
  assign n28664 = ~n16635 & n28663;
  assign n28665 = ~n28633 & ~n28664;
  assign n28666 = ~n16631 & n28665;
  assign n28667 = n16631 & n28632;
  assign n28668 = ~n28666 & ~n28667;
  assign n28669 = ~pi0792 & n28668;
  assign n28670 = pi0628 & ~n28668;
  assign n28671 = ~pi0628 & n28632;
  assign n28672 = pi1156 & ~n28671;
  assign n28673 = ~n28670 & n28672;
  assign n28674 = pi0628 & n28632;
  assign n28675 = ~pi0628 & ~n28668;
  assign n28676 = ~pi1156 & ~n28674;
  assign n28677 = ~n28675 & n28676;
  assign n28678 = ~n28673 & ~n28677;
  assign n28679 = pi0792 & ~n28678;
  assign n28680 = ~n28669 & ~n28679;
  assign n28681 = ~pi0647 & ~n28680;
  assign n28682 = pi0647 & ~n28632;
  assign n28683 = ~n28681 & ~n28682;
  assign n28684 = ~pi1157 & n28683;
  assign n28685 = pi0647 & ~n28680;
  assign n28686 = ~pi0647 & ~n28632;
  assign n28687 = ~n28685 & ~n28686;
  assign n28688 = pi1157 & n28687;
  assign n28689 = ~n28684 & ~n28688;
  assign n28690 = pi0787 & ~n28689;
  assign n28691 = ~pi0787 & n28680;
  assign n28692 = ~n28690 & ~n28691;
  assign n28693 = ~pi0644 & ~n28692;
  assign n28694 = pi0715 & ~n28693;
  assign n28695 = pi0185 & ~n2571;
  assign n28696 = pi0185 & pi0751;
  assign n28697 = pi0751 & n17046;
  assign n28698 = pi0185 & n17273;
  assign n28699 = ~n28697 & ~n28698;
  assign n28700 = pi0039 & ~n28699;
  assign n28701 = pi0185 & ~n17233;
  assign n28702 = ~n21259 & ~n28701;
  assign n28703 = ~pi0039 & ~n28702;
  assign n28704 = ~pi0185 & ~pi0751;
  assign n28705 = n17221 & n28704;
  assign n28706 = ~n28696 & ~n28703;
  assign n28707 = ~n28705 & n28706;
  assign n28708 = ~n28700 & n28707;
  assign n28709 = ~pi0038 & ~n28708;
  assign n28710 = ~pi0751 & n17280;
  assign n28711 = pi0038 & ~n28636;
  assign n28712 = ~n28710 & n28711;
  assign n28713 = ~n28709 & ~n28712;
  assign n28714 = n2571 & ~n28713;
  assign n28715 = ~n28695 & ~n28714;
  assign n28716 = ~n17117 & ~n28715;
  assign n28717 = n17117 & ~n28632;
  assign n28718 = ~n28716 & ~n28717;
  assign n28719 = ~pi0785 & ~n28718;
  assign n28720 = ~n17291 & ~n28632;
  assign n28721 = pi0609 & n28716;
  assign n28722 = ~n28720 & ~n28721;
  assign n28723 = pi1155 & ~n28722;
  assign n28724 = ~n17296 & ~n28632;
  assign n28725 = ~pi0609 & n28716;
  assign n28726 = ~n28724 & ~n28725;
  assign n28727 = ~pi1155 & ~n28726;
  assign n28728 = ~n28723 & ~n28727;
  assign n28729 = pi0785 & ~n28728;
  assign n28730 = ~n28719 & ~n28729;
  assign n28731 = ~pi0781 & ~n28730;
  assign n28732 = ~pi0618 & n28632;
  assign n28733 = pi0618 & n28730;
  assign n28734 = pi1154 & ~n28732;
  assign n28735 = ~n28733 & n28734;
  assign n28736 = ~pi0618 & n28730;
  assign n28737 = pi0618 & n28632;
  assign n28738 = ~pi1154 & ~n28737;
  assign n28739 = ~n28736 & n28738;
  assign n28740 = ~n28735 & ~n28739;
  assign n28741 = pi0781 & ~n28740;
  assign n28742 = ~n28731 & ~n28741;
  assign n28743 = ~pi0789 & ~n28742;
  assign n28744 = ~pi0619 & n28632;
  assign n28745 = pi0619 & n28742;
  assign n28746 = pi1159 & ~n28744;
  assign n28747 = ~n28745 & n28746;
  assign n28748 = ~pi0619 & n28742;
  assign n28749 = pi0619 & n28632;
  assign n28750 = ~pi1159 & ~n28749;
  assign n28751 = ~n28748 & n28750;
  assign n28752 = ~n28747 & ~n28751;
  assign n28753 = pi0789 & ~n28752;
  assign n28754 = ~n28743 & ~n28753;
  assign n28755 = ~n17969 & n28754;
  assign n28756 = n17969 & n28632;
  assign n28757 = ~n28755 & ~n28756;
  assign n28758 = ~n17779 & ~n28757;
  assign n28759 = n17779 & n28632;
  assign n28760 = ~n28758 & ~n28759;
  assign n28761 = ~n17804 & ~n28760;
  assign n28762 = n17804 & n28632;
  assign n28763 = ~n28761 & ~n28762;
  assign n28764 = pi0644 & ~n28763;
  assign n28765 = ~pi0644 & n28632;
  assign n28766 = ~pi0715 & ~n28765;
  assign n28767 = ~n28764 & n28766;
  assign n28768 = pi1160 & ~n28767;
  assign n28769 = ~n28694 & n28768;
  assign n28770 = pi0644 & ~n28692;
  assign n28771 = ~pi0715 & ~n28770;
  assign n28772 = ~pi0644 & ~n28763;
  assign n28773 = pi0644 & n28632;
  assign n28774 = pi0715 & ~n28773;
  assign n28775 = ~n28772 & n28774;
  assign n28776 = ~pi1160 & ~n28775;
  assign n28777 = ~n28771 & n28776;
  assign n28778 = ~n28769 & ~n28777;
  assign n28779 = pi0790 & ~n28778;
  assign n28780 = ~pi0629 & n28673;
  assign n28781 = ~n20570 & n28757;
  assign n28782 = pi0629 & n28677;
  assign n28783 = ~n28780 & ~n28782;
  assign n28784 = ~n28781 & n28783;
  assign n28785 = pi0792 & ~n28784;
  assign n28786 = pi0609 & n28657;
  assign n28787 = pi0185 & ~n17625;
  assign n28788 = ~pi0185 & ~n17612;
  assign n28789 = pi0751 & ~n28787;
  assign n28790 = ~n28788 & n28789;
  assign n28791 = ~pi0185 & n17629;
  assign n28792 = pi0185 & n17631;
  assign n28793 = ~pi0751 & ~n28792;
  assign n28794 = ~n28791 & n28793;
  assign n28795 = ~n28790 & ~n28794;
  assign n28796 = ~pi0039 & ~n28795;
  assign n28797 = pi0185 & n17605;
  assign n28798 = ~pi0185 & ~n17546;
  assign n28799 = ~pi0751 & ~n28798;
  assign n28800 = ~n28797 & n28799;
  assign n28801 = ~pi0185 & n17404;
  assign n28802 = pi0185 & n17485;
  assign n28803 = pi0751 & ~n28802;
  assign n28804 = ~n28801 & n28803;
  assign n28805 = pi0039 & ~n28800;
  assign n28806 = ~n28804 & n28805;
  assign n28807 = ~pi0038 & ~n28796;
  assign n28808 = ~n28806 & n28807;
  assign n28809 = ~n17469 & ~n28465;
  assign n28810 = pi0185 & ~n28809;
  assign n28811 = n6284 & n28810;
  assign n28812 = ~pi0751 & ~n17490;
  assign n28813 = n19471 & ~n28812;
  assign n28814 = ~pi0185 & ~n28813;
  assign n28815 = pi0038 & ~n28811;
  assign n28816 = ~n28814 & n28815;
  assign n28817 = ~pi0701 & ~n28816;
  assign n28818 = ~n28808 & n28817;
  assign n28819 = pi0701 & n28713;
  assign n28820 = n2571 & ~n28818;
  assign n28821 = ~n28819 & n28820;
  assign n28822 = ~n28695 & ~n28821;
  assign n28823 = ~pi0625 & n28822;
  assign n28824 = pi0625 & n28715;
  assign n28825 = ~pi1153 & ~n28824;
  assign n28826 = ~n28823 & n28825;
  assign n28827 = ~pi0608 & ~n28650;
  assign n28828 = ~n28826 & n28827;
  assign n28829 = ~pi0625 & n28715;
  assign n28830 = pi0625 & n28822;
  assign n28831 = pi1153 & ~n28829;
  assign n28832 = ~n28830 & n28831;
  assign n28833 = pi0608 & ~n28654;
  assign n28834 = ~n28832 & n28833;
  assign n28835 = ~n28828 & ~n28834;
  assign n28836 = pi0778 & ~n28835;
  assign n28837 = ~pi0778 & n28822;
  assign n28838 = ~n28836 & ~n28837;
  assign n28839 = ~pi0609 & ~n28838;
  assign n28840 = ~pi1155 & ~n28786;
  assign n28841 = ~n28839 & n28840;
  assign n28842 = ~pi0660 & ~n28723;
  assign n28843 = ~n28841 & n28842;
  assign n28844 = ~pi0609 & n28657;
  assign n28845 = pi0609 & ~n28838;
  assign n28846 = pi1155 & ~n28844;
  assign n28847 = ~n28845 & n28846;
  assign n28848 = pi0660 & ~n28727;
  assign n28849 = ~n28847 & n28848;
  assign n28850 = ~n28843 & ~n28849;
  assign n28851 = pi0785 & ~n28850;
  assign n28852 = ~pi0785 & ~n28838;
  assign n28853 = ~n28851 & ~n28852;
  assign n28854 = ~pi0618 & ~n28853;
  assign n28855 = pi0618 & n28660;
  assign n28856 = ~pi1154 & ~n28855;
  assign n28857 = ~n28854 & n28856;
  assign n28858 = ~pi0627 & ~n28735;
  assign n28859 = ~n28857 & n28858;
  assign n28860 = ~pi0618 & n28660;
  assign n28861 = pi0618 & ~n28853;
  assign n28862 = pi1154 & ~n28860;
  assign n28863 = ~n28861 & n28862;
  assign n28864 = pi0627 & ~n28739;
  assign n28865 = ~n28863 & n28864;
  assign n28866 = ~n28859 & ~n28865;
  assign n28867 = pi0781 & ~n28866;
  assign n28868 = ~pi0781 & ~n28853;
  assign n28869 = ~n28867 & ~n28868;
  assign n28870 = ~pi0789 & n28869;
  assign n28871 = pi0619 & ~n28663;
  assign n28872 = ~pi0619 & ~n28869;
  assign n28873 = ~pi1159 & ~n28871;
  assign n28874 = ~n28872 & n28873;
  assign n28875 = ~pi0648 & ~n28747;
  assign n28876 = ~n28874 & n28875;
  assign n28877 = ~pi0619 & ~n28663;
  assign n28878 = pi0619 & ~n28869;
  assign n28879 = pi1159 & ~n28877;
  assign n28880 = ~n28878 & n28879;
  assign n28881 = pi0648 & ~n28751;
  assign n28882 = ~n28880 & n28881;
  assign n28883 = pi0789 & ~n28876;
  assign n28884 = ~n28882 & n28883;
  assign n28885 = n17970 & ~n28870;
  assign n28886 = ~n28884 & n28885;
  assign n28887 = n17871 & n28665;
  assign n28888 = ~pi0626 & ~n28754;
  assign n28889 = pi0626 & ~n28632;
  assign n28890 = n16629 & ~n28889;
  assign n28891 = ~n28888 & n28890;
  assign n28892 = pi0626 & ~n28754;
  assign n28893 = ~pi0626 & ~n28632;
  assign n28894 = n16628 & ~n28893;
  assign n28895 = ~n28892 & n28894;
  assign n28896 = ~n28887 & ~n28891;
  assign n28897 = ~n28895 & n28896;
  assign n28898 = pi0788 & ~n28897;
  assign n28899 = ~n20364 & ~n28898;
  assign n28900 = ~n28886 & n28899;
  assign n28901 = ~n28785 & ~n28900;
  assign n28902 = ~n20206 & ~n28901;
  assign n28903 = n17802 & ~n28683;
  assign n28904 = ~n20559 & n28760;
  assign n28905 = n17801 & ~n28687;
  assign n28906 = ~n28903 & ~n28905;
  assign n28907 = ~n28904 & n28906;
  assign n28908 = pi0787 & ~n28907;
  assign n28909 = ~pi0644 & n28776;
  assign n28910 = pi0644 & n28768;
  assign n28911 = pi0790 & ~n28909;
  assign n28912 = ~n28910 & n28911;
  assign n28913 = ~n28902 & ~n28908;
  assign n28914 = ~n28912 & n28913;
  assign n28915 = ~n28779 & ~n28914;
  assign n28916 = ~po1038 & ~n28915;
  assign n28917 = ~pi0832 & ~n28631;
  assign n28918 = ~n28916 & n28917;
  assign po0342 = ~n28630 & ~n28918;
  assign n28920 = ~pi0186 & ~n17059;
  assign n28921 = n16635 & ~n28920;
  assign n28922 = pi0186 & ~n2571;
  assign n28923 = ~pi0186 & ~n17052;
  assign n28924 = ~pi0703 & n28923;
  assign n28925 = ~pi0186 & ~n16641;
  assign n28926 = n16647 & ~n28925;
  assign n28927 = ~pi0186 & n18072;
  assign n28928 = pi0186 & ~n18076;
  assign n28929 = ~pi0038 & ~n28928;
  assign n28930 = ~n28927 & n28929;
  assign n28931 = pi0703 & ~n28926;
  assign n28932 = ~n28930 & n28931;
  assign n28933 = n2571 & ~n28924;
  assign n28934 = ~n28932 & n28933;
  assign n28935 = ~n28922 & ~n28934;
  assign n28936 = ~pi0778 & ~n28935;
  assign n28937 = ~pi0625 & n28920;
  assign n28938 = pi0625 & n28935;
  assign n28939 = pi1153 & ~n28937;
  assign n28940 = ~n28938 & n28939;
  assign n28941 = ~pi0625 & n28935;
  assign n28942 = pi0625 & n28920;
  assign n28943 = ~pi1153 & ~n28942;
  assign n28944 = ~n28941 & n28943;
  assign n28945 = ~n28940 & ~n28944;
  assign n28946 = pi0778 & ~n28945;
  assign n28947 = ~n28936 & ~n28946;
  assign n28948 = ~n17075 & ~n28947;
  assign n28949 = n17075 & ~n28920;
  assign n28950 = ~n28948 & ~n28949;
  assign n28951 = ~n16639 & n28950;
  assign n28952 = n16639 & n28920;
  assign n28953 = ~n28951 & ~n28952;
  assign n28954 = ~n16635 & n28953;
  assign n28955 = ~n28921 & ~n28954;
  assign n28956 = ~n16631 & n28955;
  assign n28957 = n16631 & n28920;
  assign n28958 = ~n28956 & ~n28957;
  assign n28959 = ~pi0792 & n28958;
  assign n28960 = ~pi0628 & n28920;
  assign n28961 = pi0628 & ~n28958;
  assign n28962 = pi1156 & ~n28960;
  assign n28963 = ~n28961 & n28962;
  assign n28964 = pi0628 & n28920;
  assign n28965 = ~pi0628 & ~n28958;
  assign n28966 = ~pi1156 & ~n28964;
  assign n28967 = ~n28965 & n28966;
  assign n28968 = ~n28963 & ~n28967;
  assign n28969 = pi0792 & ~n28968;
  assign n28970 = ~n28959 & ~n28969;
  assign n28971 = ~pi0787 & ~n28970;
  assign n28972 = ~pi0647 & n28920;
  assign n28973 = pi0647 & n28970;
  assign n28974 = pi1157 & ~n28972;
  assign n28975 = ~n28973 & n28974;
  assign n28976 = ~pi0647 & n28970;
  assign n28977 = pi0647 & n28920;
  assign n28978 = ~pi1157 & ~n28977;
  assign n28979 = ~n28976 & n28978;
  assign n28980 = ~n28975 & ~n28979;
  assign n28981 = pi0787 & ~n28980;
  assign n28982 = ~n28971 & ~n28981;
  assign n28983 = ~pi0644 & n28982;
  assign n28984 = ~pi0618 & n28920;
  assign n28985 = pi0752 & ~n28923;
  assign n28986 = pi0186 & ~n19434;
  assign n28987 = ~pi0186 & ~pi0752;
  assign n28988 = n19439 & n28987;
  assign n28989 = ~n28986 & ~n28988;
  assign n28990 = ~n19433 & ~n28989;
  assign n28991 = ~n28985 & ~n28990;
  assign n28992 = n2571 & ~n28991;
  assign n28993 = ~n28922 & ~n28992;
  assign n28994 = ~n17117 & ~n28993;
  assign n28995 = n17117 & ~n28920;
  assign n28996 = ~n28994 & ~n28995;
  assign n28997 = ~pi0785 & ~n28996;
  assign n28998 = ~n17291 & ~n28920;
  assign n28999 = pi0609 & n28994;
  assign n29000 = ~n28998 & ~n28999;
  assign n29001 = pi1155 & ~n29000;
  assign n29002 = ~n17296 & ~n28920;
  assign n29003 = ~pi0609 & n28994;
  assign n29004 = ~n29002 & ~n29003;
  assign n29005 = ~pi1155 & ~n29004;
  assign n29006 = ~n29001 & ~n29005;
  assign n29007 = pi0785 & ~n29006;
  assign n29008 = ~n28997 & ~n29007;
  assign n29009 = pi0618 & n29008;
  assign n29010 = pi1154 & ~n28984;
  assign n29011 = ~n29009 & n29010;
  assign n29012 = pi0186 & n19468;
  assign n29013 = ~pi0186 & n19477;
  assign n29014 = pi0752 & ~n19470;
  assign n29015 = ~n29012 & n29014;
  assign n29016 = ~n29013 & n29015;
  assign n29017 = ~pi0186 & ~n19488;
  assign n29018 = pi0186 & n19496;
  assign n29019 = ~pi0752 & ~n29017;
  assign n29020 = ~n29018 & n29019;
  assign n29021 = pi0703 & ~n29020;
  assign n29022 = ~n29016 & n29021;
  assign n29023 = ~pi0703 & n28991;
  assign n29024 = n2571 & ~n29022;
  assign n29025 = ~n29023 & n29024;
  assign n29026 = ~n28922 & ~n29025;
  assign n29027 = ~pi0625 & n29026;
  assign n29028 = pi0625 & n28993;
  assign n29029 = ~pi1153 & ~n29028;
  assign n29030 = ~n29027 & n29029;
  assign n29031 = ~pi0608 & ~n28940;
  assign n29032 = ~n29030 & n29031;
  assign n29033 = ~pi0625 & n28993;
  assign n29034 = pi0625 & n29026;
  assign n29035 = pi1153 & ~n29033;
  assign n29036 = ~n29034 & n29035;
  assign n29037 = pi0608 & ~n28944;
  assign n29038 = ~n29036 & n29037;
  assign n29039 = ~n29032 & ~n29038;
  assign n29040 = pi0778 & ~n29039;
  assign n29041 = ~pi0778 & n29026;
  assign n29042 = ~n29040 & ~n29041;
  assign n29043 = ~pi0609 & ~n29042;
  assign n29044 = pi0609 & n28947;
  assign n29045 = ~pi1155 & ~n29044;
  assign n29046 = ~n29043 & n29045;
  assign n29047 = ~pi0660 & ~n29001;
  assign n29048 = ~n29046 & n29047;
  assign n29049 = ~pi0609 & n28947;
  assign n29050 = pi0609 & ~n29042;
  assign n29051 = pi1155 & ~n29049;
  assign n29052 = ~n29050 & n29051;
  assign n29053 = pi0660 & ~n29005;
  assign n29054 = ~n29052 & n29053;
  assign n29055 = ~n29048 & ~n29054;
  assign n29056 = pi0785 & ~n29055;
  assign n29057 = ~pi0785 & ~n29042;
  assign n29058 = ~n29056 & ~n29057;
  assign n29059 = ~pi0618 & ~n29058;
  assign n29060 = pi0618 & n28950;
  assign n29061 = ~pi1154 & ~n29060;
  assign n29062 = ~n29059 & n29061;
  assign n29063 = ~pi0627 & ~n29011;
  assign n29064 = ~n29062 & n29063;
  assign n29065 = ~pi0618 & n29008;
  assign n29066 = pi0618 & n28920;
  assign n29067 = ~pi1154 & ~n29066;
  assign n29068 = ~n29065 & n29067;
  assign n29069 = ~pi0618 & n28950;
  assign n29070 = pi0618 & ~n29058;
  assign n29071 = pi1154 & ~n29069;
  assign n29072 = ~n29070 & n29071;
  assign n29073 = pi0627 & ~n29068;
  assign n29074 = ~n29072 & n29073;
  assign n29075 = ~n29064 & ~n29074;
  assign n29076 = pi0781 & ~n29075;
  assign n29077 = ~pi0781 & ~n29058;
  assign n29078 = ~n29076 & ~n29077;
  assign n29079 = ~pi0619 & ~n29078;
  assign n29080 = pi0619 & ~n28953;
  assign n29081 = ~pi1159 & ~n29080;
  assign n29082 = ~n29079 & n29081;
  assign n29083 = ~pi0619 & n28920;
  assign n29084 = ~pi0781 & ~n29008;
  assign n29085 = ~n29011 & ~n29068;
  assign n29086 = pi0781 & ~n29085;
  assign n29087 = ~n29084 & ~n29086;
  assign n29088 = pi0619 & n29087;
  assign n29089 = pi1159 & ~n29083;
  assign n29090 = ~n29088 & n29089;
  assign n29091 = ~pi0648 & ~n29090;
  assign n29092 = ~n29082 & n29091;
  assign n29093 = pi0619 & ~n29078;
  assign n29094 = ~pi0619 & ~n28953;
  assign n29095 = pi1159 & ~n29094;
  assign n29096 = ~n29093 & n29095;
  assign n29097 = ~pi0619 & n29087;
  assign n29098 = pi0619 & n28920;
  assign n29099 = ~pi1159 & ~n29098;
  assign n29100 = ~n29097 & n29099;
  assign n29101 = pi0648 & ~n29100;
  assign n29102 = ~n29096 & n29101;
  assign n29103 = ~n29092 & ~n29102;
  assign n29104 = pi0789 & ~n29103;
  assign n29105 = ~pi0789 & ~n29078;
  assign n29106 = ~n29104 & ~n29105;
  assign n29107 = ~pi0788 & n29106;
  assign n29108 = ~pi0626 & n29106;
  assign n29109 = pi0626 & ~n28955;
  assign n29110 = ~pi0641 & ~n29109;
  assign n29111 = ~n29108 & n29110;
  assign n29112 = ~pi0789 & ~n29087;
  assign n29113 = ~n29090 & ~n29100;
  assign n29114 = pi0789 & ~n29113;
  assign n29115 = ~n29112 & ~n29114;
  assign n29116 = ~pi0626 & ~n29115;
  assign n29117 = pi0626 & ~n28920;
  assign n29118 = pi0641 & ~n29117;
  assign n29119 = ~n29116 & n29118;
  assign n29120 = ~pi1158 & ~n29119;
  assign n29121 = ~n29111 & n29120;
  assign n29122 = pi0626 & n29106;
  assign n29123 = ~pi0626 & ~n28955;
  assign n29124 = pi0641 & ~n29123;
  assign n29125 = ~n29122 & n29124;
  assign n29126 = pi0626 & ~n29115;
  assign n29127 = ~pi0626 & ~n28920;
  assign n29128 = ~pi0641 & ~n29127;
  assign n29129 = ~n29126 & n29128;
  assign n29130 = pi1158 & ~n29129;
  assign n29131 = ~n29125 & n29130;
  assign n29132 = ~n29121 & ~n29131;
  assign n29133 = pi0788 & ~n29132;
  assign n29134 = ~n29107 & ~n29133;
  assign n29135 = ~pi0628 & n29134;
  assign n29136 = ~n17969 & n29115;
  assign n29137 = n17969 & n28920;
  assign n29138 = ~n29136 & ~n29137;
  assign n29139 = pi0628 & ~n29138;
  assign n29140 = ~pi1156 & ~n29139;
  assign n29141 = ~n29135 & n29140;
  assign n29142 = ~pi0629 & ~n28963;
  assign n29143 = ~n29141 & n29142;
  assign n29144 = pi0628 & n29134;
  assign n29145 = ~pi0628 & ~n29138;
  assign n29146 = pi1156 & ~n29145;
  assign n29147 = ~n29144 & n29146;
  assign n29148 = pi0629 & ~n28967;
  assign n29149 = ~n29147 & n29148;
  assign n29150 = ~n29143 & ~n29149;
  assign n29151 = pi0792 & ~n29150;
  assign n29152 = ~pi0792 & n29134;
  assign n29153 = ~n29151 & ~n29152;
  assign n29154 = ~pi0647 & ~n29153;
  assign n29155 = ~n17779 & ~n29138;
  assign n29156 = n17779 & n28920;
  assign n29157 = ~n29155 & ~n29156;
  assign n29158 = pi0647 & ~n29157;
  assign n29159 = ~pi1157 & ~n29158;
  assign n29160 = ~n29154 & n29159;
  assign n29161 = ~pi0630 & ~n28975;
  assign n29162 = ~n29160 & n29161;
  assign n29163 = pi0647 & ~n29153;
  assign n29164 = ~pi0647 & ~n29157;
  assign n29165 = pi1157 & ~n29164;
  assign n29166 = ~n29163 & n29165;
  assign n29167 = pi0630 & ~n28979;
  assign n29168 = ~n29166 & n29167;
  assign n29169 = ~n29162 & ~n29168;
  assign n29170 = pi0787 & ~n29169;
  assign n29171 = ~pi0787 & ~n29153;
  assign n29172 = ~n29170 & ~n29171;
  assign n29173 = pi0644 & ~n29172;
  assign n29174 = pi0715 & ~n28983;
  assign n29175 = ~n29173 & n29174;
  assign n29176 = n17804 & ~n28920;
  assign n29177 = ~n17804 & n29157;
  assign n29178 = ~n29176 & ~n29177;
  assign n29179 = pi0644 & n29178;
  assign n29180 = ~pi0644 & n28920;
  assign n29181 = ~pi0715 & ~n29180;
  assign n29182 = ~n29179 & n29181;
  assign n29183 = pi1160 & ~n29182;
  assign n29184 = ~n29175 & n29183;
  assign n29185 = ~pi0644 & ~n29172;
  assign n29186 = pi0644 & n28982;
  assign n29187 = ~pi0715 & ~n29186;
  assign n29188 = ~n29185 & n29187;
  assign n29189 = ~pi0644 & n29178;
  assign n29190 = pi0644 & n28920;
  assign n29191 = pi0715 & ~n29190;
  assign n29192 = ~n29189 & n29191;
  assign n29193 = ~pi1160 & ~n29192;
  assign n29194 = ~n29188 & n29193;
  assign n29195 = pi0790 & ~n29184;
  assign n29196 = ~n29194 & n29195;
  assign n29197 = ~pi0790 & n29172;
  assign n29198 = ~po1038 & ~n29197;
  assign n29199 = ~n29196 & n29198;
  assign n29200 = ~pi0186 & po1038;
  assign n29201 = ~pi0832 & ~n29200;
  assign n29202 = ~n29199 & n29201;
  assign n29203 = ~pi0186 & ~n2926;
  assign n29204 = pi0703 & n16645;
  assign n29205 = ~n29203 & ~n29204;
  assign n29206 = ~pi0778 & n29205;
  assign n29207 = ~pi0625 & n29204;
  assign n29208 = ~n29205 & ~n29207;
  assign n29209 = pi1153 & ~n29208;
  assign n29210 = ~pi1153 & ~n29203;
  assign n29211 = ~n29207 & n29210;
  assign n29212 = ~n29209 & ~n29211;
  assign n29213 = pi0778 & ~n29212;
  assign n29214 = ~n29206 & ~n29213;
  assign n29215 = ~n17845 & n29214;
  assign n29216 = ~n17847 & n29215;
  assign n29217 = ~n17849 & n29216;
  assign n29218 = ~n17851 & n29217;
  assign n29219 = ~n17857 & n29218;
  assign n29220 = ~pi0647 & n29219;
  assign n29221 = pi0647 & n29203;
  assign n29222 = ~pi1157 & ~n29221;
  assign n29223 = ~n29220 & n29222;
  assign n29224 = pi0630 & n29223;
  assign n29225 = ~pi0752 & n17244;
  assign n29226 = ~n29203 & ~n29225;
  assign n29227 = ~n17874 & ~n29226;
  assign n29228 = ~pi0785 & ~n29227;
  assign n29229 = ~n17879 & ~n29226;
  assign n29230 = pi1155 & ~n29229;
  assign n29231 = ~n17882 & n29227;
  assign n29232 = ~pi1155 & ~n29231;
  assign n29233 = ~n29230 & ~n29232;
  assign n29234 = pi0785 & ~n29233;
  assign n29235 = ~n29228 & ~n29234;
  assign n29236 = ~pi0781 & ~n29235;
  assign n29237 = ~n17889 & n29235;
  assign n29238 = pi1154 & ~n29237;
  assign n29239 = ~n17892 & n29235;
  assign n29240 = ~pi1154 & ~n29239;
  assign n29241 = ~n29238 & ~n29240;
  assign n29242 = pi0781 & ~n29241;
  assign n29243 = ~n29236 & ~n29242;
  assign n29244 = ~pi0789 & ~n29243;
  assign n29245 = ~pi0619 & n29203;
  assign n29246 = pi0619 & n29243;
  assign n29247 = pi1159 & ~n29245;
  assign n29248 = ~n29246 & n29247;
  assign n29249 = ~pi0619 & n29243;
  assign n29250 = pi0619 & n29203;
  assign n29251 = ~pi1159 & ~n29250;
  assign n29252 = ~n29249 & n29251;
  assign n29253 = ~n29248 & ~n29252;
  assign n29254 = pi0789 & ~n29253;
  assign n29255 = ~n29244 & ~n29254;
  assign n29256 = ~n17969 & n29255;
  assign n29257 = n17969 & n29203;
  assign n29258 = ~n29256 & ~n29257;
  assign n29259 = ~n17779 & ~n29258;
  assign n29260 = n17779 & n29203;
  assign n29261 = ~n29259 & ~n29260;
  assign n29262 = ~n20559 & n29261;
  assign n29263 = pi0647 & ~n29219;
  assign n29264 = ~pi0647 & ~n29203;
  assign n29265 = ~n29263 & ~n29264;
  assign n29266 = n17801 & ~n29265;
  assign n29267 = ~n29224 & ~n29266;
  assign n29268 = ~n29262 & n29267;
  assign n29269 = pi0787 & ~n29268;
  assign n29270 = n17871 & n29217;
  assign n29271 = ~pi0626 & ~n29255;
  assign n29272 = pi0626 & ~n29203;
  assign n29273 = n16629 & ~n29272;
  assign n29274 = ~n29271 & n29273;
  assign n29275 = pi0626 & ~n29255;
  assign n29276 = ~pi0626 & ~n29203;
  assign n29277 = n16628 & ~n29276;
  assign n29278 = ~n29275 & n29277;
  assign n29279 = ~n29270 & ~n29274;
  assign n29280 = ~n29278 & n29279;
  assign n29281 = pi0788 & ~n29280;
  assign n29282 = pi0618 & n29215;
  assign n29283 = pi0609 & n29214;
  assign n29284 = ~n17168 & ~n29205;
  assign n29285 = pi0625 & n29284;
  assign n29286 = n29226 & ~n29284;
  assign n29287 = ~n29285 & ~n29286;
  assign n29288 = n29210 & ~n29287;
  assign n29289 = ~pi0608 & ~n29209;
  assign n29290 = ~n29288 & n29289;
  assign n29291 = pi1153 & n29226;
  assign n29292 = ~n29285 & n29291;
  assign n29293 = pi0608 & ~n29211;
  assign n29294 = ~n29292 & n29293;
  assign n29295 = ~n29290 & ~n29294;
  assign n29296 = pi0778 & ~n29295;
  assign n29297 = ~pi0778 & ~n29286;
  assign n29298 = ~n29296 & ~n29297;
  assign n29299 = ~pi0609 & ~n29298;
  assign n29300 = ~pi1155 & ~n29283;
  assign n29301 = ~n29299 & n29300;
  assign n29302 = ~pi0660 & ~n29230;
  assign n29303 = ~n29301 & n29302;
  assign n29304 = ~pi0609 & n29214;
  assign n29305 = pi0609 & ~n29298;
  assign n29306 = pi1155 & ~n29304;
  assign n29307 = ~n29305 & n29306;
  assign n29308 = pi0660 & ~n29232;
  assign n29309 = ~n29307 & n29308;
  assign n29310 = ~n29303 & ~n29309;
  assign n29311 = pi0785 & ~n29310;
  assign n29312 = ~pi0785 & ~n29298;
  assign n29313 = ~n29311 & ~n29312;
  assign n29314 = ~pi0618 & ~n29313;
  assign n29315 = ~pi1154 & ~n29282;
  assign n29316 = ~n29314 & n29315;
  assign n29317 = ~pi0627 & ~n29238;
  assign n29318 = ~n29316 & n29317;
  assign n29319 = ~pi0618 & n29215;
  assign n29320 = pi0618 & ~n29313;
  assign n29321 = pi1154 & ~n29319;
  assign n29322 = ~n29320 & n29321;
  assign n29323 = pi0627 & ~n29240;
  assign n29324 = ~n29322 & n29323;
  assign n29325 = ~n29318 & ~n29324;
  assign n29326 = pi0781 & ~n29325;
  assign n29327 = ~pi0781 & ~n29313;
  assign n29328 = ~n29326 & ~n29327;
  assign n29329 = ~pi0789 & n29328;
  assign n29330 = ~pi0619 & ~n29328;
  assign n29331 = pi0619 & n29216;
  assign n29332 = ~pi1159 & ~n29331;
  assign n29333 = ~n29330 & n29332;
  assign n29334 = ~pi0648 & ~n29248;
  assign n29335 = ~n29333 & n29334;
  assign n29336 = pi0619 & ~n29328;
  assign n29337 = ~pi0619 & n29216;
  assign n29338 = pi1159 & ~n29337;
  assign n29339 = ~n29336 & n29338;
  assign n29340 = pi0648 & ~n29252;
  assign n29341 = ~n29339 & n29340;
  assign n29342 = pi0789 & ~n29335;
  assign n29343 = ~n29341 & n29342;
  assign n29344 = n17970 & ~n29329;
  assign n29345 = ~n29343 & n29344;
  assign n29346 = ~n29281 & ~n29345;
  assign n29347 = ~n20364 & ~n29346;
  assign n29348 = n17854 & ~n29258;
  assign n29349 = n20851 & n29218;
  assign n29350 = ~n29348 & ~n29349;
  assign n29351 = ~pi0629 & ~n29350;
  assign n29352 = n20855 & n29218;
  assign n29353 = n17853 & ~n29258;
  assign n29354 = ~n29352 & ~n29353;
  assign n29355 = pi0629 & ~n29354;
  assign n29356 = ~n29351 & ~n29355;
  assign n29357 = pi0792 & ~n29356;
  assign n29358 = ~n20206 & ~n29357;
  assign n29359 = ~n29347 & n29358;
  assign n29360 = ~n29269 & ~n29359;
  assign n29361 = ~pi0790 & n29360;
  assign n29362 = ~pi0787 & ~n29219;
  assign n29363 = pi1157 & ~n29265;
  assign n29364 = ~n29223 & ~n29363;
  assign n29365 = pi0787 & ~n29364;
  assign n29366 = ~n29362 & ~n29365;
  assign n29367 = ~pi0644 & n29366;
  assign n29368 = pi0644 & n29360;
  assign n29369 = pi0715 & ~n29367;
  assign n29370 = ~n29368 & n29369;
  assign n29371 = ~n17804 & ~n29261;
  assign n29372 = n17804 & n29203;
  assign n29373 = ~n29371 & ~n29372;
  assign n29374 = pi0644 & ~n29373;
  assign n29375 = ~pi0644 & n29203;
  assign n29376 = ~pi0715 & ~n29375;
  assign n29377 = ~n29374 & n29376;
  assign n29378 = pi1160 & ~n29377;
  assign n29379 = ~n29370 & n29378;
  assign n29380 = ~pi0644 & ~n29373;
  assign n29381 = pi0644 & n29203;
  assign n29382 = pi0715 & ~n29381;
  assign n29383 = ~n29380 & n29382;
  assign n29384 = pi0644 & n29366;
  assign n29385 = ~pi0644 & n29360;
  assign n29386 = ~pi0715 & ~n29384;
  assign n29387 = ~n29385 & n29386;
  assign n29388 = ~pi1160 & ~n29383;
  assign n29389 = ~n29387 & n29388;
  assign n29390 = ~n29379 & ~n29389;
  assign n29391 = pi0790 & ~n29390;
  assign n29392 = pi0832 & ~n29361;
  assign n29393 = ~n29391 & n29392;
  assign po0343 = ~n29202 & ~n29393;
  assign n29395 = ~pi0187 & ~n17059;
  assign n29396 = n16635 & ~n29395;
  assign n29397 = pi0187 & ~n2571;
  assign n29398 = ~pi0187 & ~pi0726;
  assign n29399 = ~n17052 & n29398;
  assign n29400 = ~pi0187 & ~n16641;
  assign n29401 = n16647 & ~n29400;
  assign n29402 = ~pi0187 & n18072;
  assign n29403 = pi0187 & ~n18076;
  assign n29404 = ~pi0038 & ~n29403;
  assign n29405 = ~n29402 & n29404;
  assign n29406 = pi0726 & ~n29401;
  assign n29407 = ~n29405 & n29406;
  assign n29408 = n2571 & ~n29399;
  assign n29409 = ~n29407 & n29408;
  assign n29410 = ~n29397 & ~n29409;
  assign n29411 = ~pi0778 & ~n29410;
  assign n29412 = ~pi0625 & n29395;
  assign n29413 = pi0625 & n29410;
  assign n29414 = pi1153 & ~n29412;
  assign n29415 = ~n29413 & n29414;
  assign n29416 = ~pi0625 & n29410;
  assign n29417 = pi0625 & n29395;
  assign n29418 = ~pi1153 & ~n29417;
  assign n29419 = ~n29416 & n29418;
  assign n29420 = ~n29415 & ~n29419;
  assign n29421 = pi0778 & ~n29420;
  assign n29422 = ~n29411 & ~n29421;
  assign n29423 = ~n17075 & ~n29422;
  assign n29424 = n17075 & ~n29395;
  assign n29425 = ~n29423 & ~n29424;
  assign n29426 = ~n16639 & n29425;
  assign n29427 = n16639 & n29395;
  assign n29428 = ~n29426 & ~n29427;
  assign n29429 = ~n16635 & n29428;
  assign n29430 = ~n29396 & ~n29429;
  assign n29431 = ~n16631 & n29430;
  assign n29432 = n16631 & n29395;
  assign n29433 = ~n29431 & ~n29432;
  assign n29434 = ~pi0792 & n29433;
  assign n29435 = ~pi0628 & n29395;
  assign n29436 = pi0628 & ~n29433;
  assign n29437 = pi1156 & ~n29435;
  assign n29438 = ~n29436 & n29437;
  assign n29439 = pi0628 & n29395;
  assign n29440 = ~pi0628 & ~n29433;
  assign n29441 = ~pi1156 & ~n29439;
  assign n29442 = ~n29440 & n29441;
  assign n29443 = ~n29438 & ~n29442;
  assign n29444 = pi0792 & ~n29443;
  assign n29445 = ~n29434 & ~n29444;
  assign n29446 = ~pi0787 & ~n29445;
  assign n29447 = ~pi0647 & n29395;
  assign n29448 = pi0647 & n29445;
  assign n29449 = pi1157 & ~n29447;
  assign n29450 = ~n29448 & n29449;
  assign n29451 = ~pi0647 & n29445;
  assign n29452 = pi0647 & n29395;
  assign n29453 = ~pi1157 & ~n29452;
  assign n29454 = ~n29451 & n29453;
  assign n29455 = ~n29450 & ~n29454;
  assign n29456 = pi0787 & ~n29455;
  assign n29457 = ~n29446 & ~n29456;
  assign n29458 = ~pi0644 & n29457;
  assign n29459 = ~pi0618 & n29395;
  assign n29460 = ~pi0770 & ~n19439;
  assign n29461 = ~n21012 & ~n29460;
  assign n29462 = ~pi0187 & ~n29461;
  assign n29463 = ~pi0187 & ~n19433;
  assign n29464 = ~pi0770 & ~n29463;
  assign n29465 = ~n24447 & n29464;
  assign n29466 = ~n29462 & ~n29465;
  assign n29467 = n2571 & n29466;
  assign n29468 = ~n29397 & ~n29467;
  assign n29469 = ~n17117 & ~n29468;
  assign n29470 = n17117 & ~n29395;
  assign n29471 = ~n29469 & ~n29470;
  assign n29472 = ~pi0785 & ~n29471;
  assign n29473 = ~n17291 & ~n29395;
  assign n29474 = pi0609 & n29469;
  assign n29475 = ~n29473 & ~n29474;
  assign n29476 = pi1155 & ~n29475;
  assign n29477 = ~n17296 & ~n29395;
  assign n29478 = ~pi0609 & n29469;
  assign n29479 = ~n29477 & ~n29478;
  assign n29480 = ~pi1155 & ~n29479;
  assign n29481 = ~n29476 & ~n29480;
  assign n29482 = pi0785 & ~n29481;
  assign n29483 = ~n29472 & ~n29482;
  assign n29484 = pi0618 & n29483;
  assign n29485 = pi1154 & ~n29459;
  assign n29486 = ~n29484 & n29485;
  assign n29487 = pi0187 & n19468;
  assign n29488 = ~pi0187 & n19477;
  assign n29489 = pi0770 & ~n19470;
  assign n29490 = ~n29487 & n29489;
  assign n29491 = ~n29488 & n29490;
  assign n29492 = ~pi0187 & ~n19488;
  assign n29493 = pi0187 & n19496;
  assign n29494 = ~pi0770 & ~n29492;
  assign n29495 = ~n29493 & n29494;
  assign n29496 = pi0726 & ~n29495;
  assign n29497 = ~n29491 & n29496;
  assign n29498 = ~pi0726 & ~n29466;
  assign n29499 = n2571 & ~n29497;
  assign n29500 = ~n29498 & n29499;
  assign n29501 = ~n29397 & ~n29500;
  assign n29502 = ~pi0625 & n29501;
  assign n29503 = pi0625 & n29468;
  assign n29504 = ~pi1153 & ~n29503;
  assign n29505 = ~n29502 & n29504;
  assign n29506 = ~pi0608 & ~n29415;
  assign n29507 = ~n29505 & n29506;
  assign n29508 = ~pi0625 & n29468;
  assign n29509 = pi0625 & n29501;
  assign n29510 = pi1153 & ~n29508;
  assign n29511 = ~n29509 & n29510;
  assign n29512 = pi0608 & ~n29419;
  assign n29513 = ~n29511 & n29512;
  assign n29514 = ~n29507 & ~n29513;
  assign n29515 = pi0778 & ~n29514;
  assign n29516 = ~pi0778 & n29501;
  assign n29517 = ~n29515 & ~n29516;
  assign n29518 = ~pi0609 & ~n29517;
  assign n29519 = pi0609 & n29422;
  assign n29520 = ~pi1155 & ~n29519;
  assign n29521 = ~n29518 & n29520;
  assign n29522 = ~pi0660 & ~n29476;
  assign n29523 = ~n29521 & n29522;
  assign n29524 = ~pi0609 & n29422;
  assign n29525 = pi0609 & ~n29517;
  assign n29526 = pi1155 & ~n29524;
  assign n29527 = ~n29525 & n29526;
  assign n29528 = pi0660 & ~n29480;
  assign n29529 = ~n29527 & n29528;
  assign n29530 = ~n29523 & ~n29529;
  assign n29531 = pi0785 & ~n29530;
  assign n29532 = ~pi0785 & ~n29517;
  assign n29533 = ~n29531 & ~n29532;
  assign n29534 = ~pi0618 & ~n29533;
  assign n29535 = pi0618 & n29425;
  assign n29536 = ~pi1154 & ~n29535;
  assign n29537 = ~n29534 & n29536;
  assign n29538 = ~pi0627 & ~n29486;
  assign n29539 = ~n29537 & n29538;
  assign n29540 = ~pi0618 & n29483;
  assign n29541 = pi0618 & n29395;
  assign n29542 = ~pi1154 & ~n29541;
  assign n29543 = ~n29540 & n29542;
  assign n29544 = ~pi0618 & n29425;
  assign n29545 = pi0618 & ~n29533;
  assign n29546 = pi1154 & ~n29544;
  assign n29547 = ~n29545 & n29546;
  assign n29548 = pi0627 & ~n29543;
  assign n29549 = ~n29547 & n29548;
  assign n29550 = ~n29539 & ~n29549;
  assign n29551 = pi0781 & ~n29550;
  assign n29552 = ~pi0781 & ~n29533;
  assign n29553 = ~n29551 & ~n29552;
  assign n29554 = ~pi0619 & ~n29553;
  assign n29555 = pi0619 & ~n29428;
  assign n29556 = ~pi1159 & ~n29555;
  assign n29557 = ~n29554 & n29556;
  assign n29558 = ~pi0619 & n29395;
  assign n29559 = ~pi0781 & ~n29483;
  assign n29560 = ~n29486 & ~n29543;
  assign n29561 = pi0781 & ~n29560;
  assign n29562 = ~n29559 & ~n29561;
  assign n29563 = pi0619 & n29562;
  assign n29564 = pi1159 & ~n29558;
  assign n29565 = ~n29563 & n29564;
  assign n29566 = ~pi0648 & ~n29565;
  assign n29567 = ~n29557 & n29566;
  assign n29568 = pi0619 & ~n29553;
  assign n29569 = ~pi0619 & ~n29428;
  assign n29570 = pi1159 & ~n29569;
  assign n29571 = ~n29568 & n29570;
  assign n29572 = ~pi0619 & n29562;
  assign n29573 = pi0619 & n29395;
  assign n29574 = ~pi1159 & ~n29573;
  assign n29575 = ~n29572 & n29574;
  assign n29576 = pi0648 & ~n29575;
  assign n29577 = ~n29571 & n29576;
  assign n29578 = ~n29567 & ~n29577;
  assign n29579 = pi0789 & ~n29578;
  assign n29580 = ~pi0789 & ~n29553;
  assign n29581 = ~n29579 & ~n29580;
  assign n29582 = ~pi0788 & n29581;
  assign n29583 = ~pi0626 & n29581;
  assign n29584 = pi0626 & ~n29430;
  assign n29585 = ~pi0641 & ~n29584;
  assign n29586 = ~n29583 & n29585;
  assign n29587 = ~pi0789 & ~n29562;
  assign n29588 = ~n29565 & ~n29575;
  assign n29589 = pi0789 & ~n29588;
  assign n29590 = ~n29587 & ~n29589;
  assign n29591 = ~pi0626 & ~n29590;
  assign n29592 = pi0626 & ~n29395;
  assign n29593 = pi0641 & ~n29592;
  assign n29594 = ~n29591 & n29593;
  assign n29595 = ~pi1158 & ~n29594;
  assign n29596 = ~n29586 & n29595;
  assign n29597 = pi0626 & n29581;
  assign n29598 = ~pi0626 & ~n29430;
  assign n29599 = pi0641 & ~n29598;
  assign n29600 = ~n29597 & n29599;
  assign n29601 = pi0626 & ~n29590;
  assign n29602 = ~pi0626 & ~n29395;
  assign n29603 = ~pi0641 & ~n29602;
  assign n29604 = ~n29601 & n29603;
  assign n29605 = pi1158 & ~n29604;
  assign n29606 = ~n29600 & n29605;
  assign n29607 = ~n29596 & ~n29606;
  assign n29608 = pi0788 & ~n29607;
  assign n29609 = ~n29582 & ~n29608;
  assign n29610 = ~pi0628 & n29609;
  assign n29611 = ~n17969 & n29590;
  assign n29612 = n17969 & n29395;
  assign n29613 = ~n29611 & ~n29612;
  assign n29614 = pi0628 & ~n29613;
  assign n29615 = ~pi1156 & ~n29614;
  assign n29616 = ~n29610 & n29615;
  assign n29617 = ~pi0629 & ~n29438;
  assign n29618 = ~n29616 & n29617;
  assign n29619 = pi0628 & n29609;
  assign n29620 = ~pi0628 & ~n29613;
  assign n29621 = pi1156 & ~n29620;
  assign n29622 = ~n29619 & n29621;
  assign n29623 = pi0629 & ~n29442;
  assign n29624 = ~n29622 & n29623;
  assign n29625 = ~n29618 & ~n29624;
  assign n29626 = pi0792 & ~n29625;
  assign n29627 = ~pi0792 & n29609;
  assign n29628 = ~n29626 & ~n29627;
  assign n29629 = ~pi0647 & ~n29628;
  assign n29630 = ~n17779 & ~n29613;
  assign n29631 = n17779 & n29395;
  assign n29632 = ~n29630 & ~n29631;
  assign n29633 = pi0647 & ~n29632;
  assign n29634 = ~pi1157 & ~n29633;
  assign n29635 = ~n29629 & n29634;
  assign n29636 = ~pi0630 & ~n29450;
  assign n29637 = ~n29635 & n29636;
  assign n29638 = pi0647 & ~n29628;
  assign n29639 = ~pi0647 & ~n29632;
  assign n29640 = pi1157 & ~n29639;
  assign n29641 = ~n29638 & n29640;
  assign n29642 = pi0630 & ~n29454;
  assign n29643 = ~n29641 & n29642;
  assign n29644 = ~n29637 & ~n29643;
  assign n29645 = pi0787 & ~n29644;
  assign n29646 = ~pi0787 & ~n29628;
  assign n29647 = ~n29645 & ~n29646;
  assign n29648 = pi0644 & ~n29647;
  assign n29649 = pi0715 & ~n29458;
  assign n29650 = ~n29648 & n29649;
  assign n29651 = n17804 & ~n29395;
  assign n29652 = ~n17804 & n29632;
  assign n29653 = ~n29651 & ~n29652;
  assign n29654 = pi0644 & n29653;
  assign n29655 = ~pi0644 & n29395;
  assign n29656 = ~pi0715 & ~n29655;
  assign n29657 = ~n29654 & n29656;
  assign n29658 = pi1160 & ~n29657;
  assign n29659 = ~n29650 & n29658;
  assign n29660 = ~pi0644 & ~n29647;
  assign n29661 = pi0644 & n29457;
  assign n29662 = ~pi0715 & ~n29661;
  assign n29663 = ~n29660 & n29662;
  assign n29664 = ~pi0644 & n29653;
  assign n29665 = pi0644 & n29395;
  assign n29666 = pi0715 & ~n29665;
  assign n29667 = ~n29664 & n29666;
  assign n29668 = ~pi1160 & ~n29667;
  assign n29669 = ~n29663 & n29668;
  assign n29670 = pi0790 & ~n29659;
  assign n29671 = ~n29669 & n29670;
  assign n29672 = ~pi0790 & n29647;
  assign n29673 = ~po1038 & ~n29672;
  assign n29674 = ~n29671 & n29673;
  assign n29675 = ~pi0187 & po1038;
  assign n29676 = ~pi0832 & ~n29675;
  assign n29677 = ~n29674 & n29676;
  assign n29678 = ~pi0187 & ~n2926;
  assign n29679 = pi0726 & n16645;
  assign n29680 = ~n29678 & ~n29679;
  assign n29681 = ~pi0778 & n29680;
  assign n29682 = ~pi0625 & n29679;
  assign n29683 = ~n29680 & ~n29682;
  assign n29684 = pi1153 & ~n29683;
  assign n29685 = ~pi1153 & ~n29678;
  assign n29686 = ~n29682 & n29685;
  assign n29687 = ~n29684 & ~n29686;
  assign n29688 = pi0778 & ~n29687;
  assign n29689 = ~n29681 & ~n29688;
  assign n29690 = ~n17845 & n29689;
  assign n29691 = ~n17847 & n29690;
  assign n29692 = ~n17849 & n29691;
  assign n29693 = ~n17851 & n29692;
  assign n29694 = ~n17857 & n29693;
  assign n29695 = ~pi0647 & n29694;
  assign n29696 = pi0647 & n29678;
  assign n29697 = ~pi1157 & ~n29696;
  assign n29698 = ~n29695 & n29697;
  assign n29699 = pi0630 & n29698;
  assign n29700 = ~pi0770 & n17244;
  assign n29701 = ~n29678 & ~n29700;
  assign n29702 = ~n17874 & ~n29701;
  assign n29703 = ~pi0785 & ~n29702;
  assign n29704 = ~n17879 & ~n29701;
  assign n29705 = pi1155 & ~n29704;
  assign n29706 = ~n17882 & n29702;
  assign n29707 = ~pi1155 & ~n29706;
  assign n29708 = ~n29705 & ~n29707;
  assign n29709 = pi0785 & ~n29708;
  assign n29710 = ~n29703 & ~n29709;
  assign n29711 = ~pi0781 & ~n29710;
  assign n29712 = ~n17889 & n29710;
  assign n29713 = pi1154 & ~n29712;
  assign n29714 = ~n17892 & n29710;
  assign n29715 = ~pi1154 & ~n29714;
  assign n29716 = ~n29713 & ~n29715;
  assign n29717 = pi0781 & ~n29716;
  assign n29718 = ~n29711 & ~n29717;
  assign n29719 = ~pi0789 & ~n29718;
  assign n29720 = ~pi0619 & n29678;
  assign n29721 = pi0619 & n29718;
  assign n29722 = pi1159 & ~n29720;
  assign n29723 = ~n29721 & n29722;
  assign n29724 = ~pi0619 & n29718;
  assign n29725 = pi0619 & n29678;
  assign n29726 = ~pi1159 & ~n29725;
  assign n29727 = ~n29724 & n29726;
  assign n29728 = ~n29723 & ~n29727;
  assign n29729 = pi0789 & ~n29728;
  assign n29730 = ~n29719 & ~n29729;
  assign n29731 = ~n17969 & n29730;
  assign n29732 = n17969 & n29678;
  assign n29733 = ~n29731 & ~n29732;
  assign n29734 = ~n17779 & ~n29733;
  assign n29735 = n17779 & n29678;
  assign n29736 = ~n29734 & ~n29735;
  assign n29737 = ~n20559 & n29736;
  assign n29738 = pi0647 & ~n29694;
  assign n29739 = ~pi0647 & ~n29678;
  assign n29740 = ~n29738 & ~n29739;
  assign n29741 = n17801 & ~n29740;
  assign n29742 = ~n29699 & ~n29741;
  assign n29743 = ~n29737 & n29742;
  assign n29744 = pi0787 & ~n29743;
  assign n29745 = n17871 & n29692;
  assign n29746 = ~pi0626 & ~n29730;
  assign n29747 = pi0626 & ~n29678;
  assign n29748 = n16629 & ~n29747;
  assign n29749 = ~n29746 & n29748;
  assign n29750 = pi0626 & ~n29730;
  assign n29751 = ~pi0626 & ~n29678;
  assign n29752 = n16628 & ~n29751;
  assign n29753 = ~n29750 & n29752;
  assign n29754 = ~n29745 & ~n29749;
  assign n29755 = ~n29753 & n29754;
  assign n29756 = pi0788 & ~n29755;
  assign n29757 = pi0618 & n29690;
  assign n29758 = pi0609 & n29689;
  assign n29759 = ~n17168 & ~n29680;
  assign n29760 = pi0625 & n29759;
  assign n29761 = n29701 & ~n29759;
  assign n29762 = ~n29760 & ~n29761;
  assign n29763 = n29685 & ~n29762;
  assign n29764 = ~pi0608 & ~n29684;
  assign n29765 = ~n29763 & n29764;
  assign n29766 = pi1153 & n29701;
  assign n29767 = ~n29760 & n29766;
  assign n29768 = pi0608 & ~n29686;
  assign n29769 = ~n29767 & n29768;
  assign n29770 = ~n29765 & ~n29769;
  assign n29771 = pi0778 & ~n29770;
  assign n29772 = ~pi0778 & ~n29761;
  assign n29773 = ~n29771 & ~n29772;
  assign n29774 = ~pi0609 & ~n29773;
  assign n29775 = ~pi1155 & ~n29758;
  assign n29776 = ~n29774 & n29775;
  assign n29777 = ~pi0660 & ~n29705;
  assign n29778 = ~n29776 & n29777;
  assign n29779 = ~pi0609 & n29689;
  assign n29780 = pi0609 & ~n29773;
  assign n29781 = pi1155 & ~n29779;
  assign n29782 = ~n29780 & n29781;
  assign n29783 = pi0660 & ~n29707;
  assign n29784 = ~n29782 & n29783;
  assign n29785 = ~n29778 & ~n29784;
  assign n29786 = pi0785 & ~n29785;
  assign n29787 = ~pi0785 & ~n29773;
  assign n29788 = ~n29786 & ~n29787;
  assign n29789 = ~pi0618 & ~n29788;
  assign n29790 = ~pi1154 & ~n29757;
  assign n29791 = ~n29789 & n29790;
  assign n29792 = ~pi0627 & ~n29713;
  assign n29793 = ~n29791 & n29792;
  assign n29794 = ~pi0618 & n29690;
  assign n29795 = pi0618 & ~n29788;
  assign n29796 = pi1154 & ~n29794;
  assign n29797 = ~n29795 & n29796;
  assign n29798 = pi0627 & ~n29715;
  assign n29799 = ~n29797 & n29798;
  assign n29800 = ~n29793 & ~n29799;
  assign n29801 = pi0781 & ~n29800;
  assign n29802 = ~pi0781 & ~n29788;
  assign n29803 = ~n29801 & ~n29802;
  assign n29804 = ~pi0789 & n29803;
  assign n29805 = ~pi0619 & ~n29803;
  assign n29806 = pi0619 & n29691;
  assign n29807 = ~pi1159 & ~n29806;
  assign n29808 = ~n29805 & n29807;
  assign n29809 = ~pi0648 & ~n29723;
  assign n29810 = ~n29808 & n29809;
  assign n29811 = pi0619 & ~n29803;
  assign n29812 = ~pi0619 & n29691;
  assign n29813 = pi1159 & ~n29812;
  assign n29814 = ~n29811 & n29813;
  assign n29815 = pi0648 & ~n29727;
  assign n29816 = ~n29814 & n29815;
  assign n29817 = pi0789 & ~n29810;
  assign n29818 = ~n29816 & n29817;
  assign n29819 = n17970 & ~n29804;
  assign n29820 = ~n29818 & n29819;
  assign n29821 = ~n29756 & ~n29820;
  assign n29822 = ~n20364 & ~n29821;
  assign n29823 = n17854 & ~n29733;
  assign n29824 = n20851 & n29693;
  assign n29825 = ~n29823 & ~n29824;
  assign n29826 = ~pi0629 & ~n29825;
  assign n29827 = n20855 & n29693;
  assign n29828 = n17853 & ~n29733;
  assign n29829 = ~n29827 & ~n29828;
  assign n29830 = pi0629 & ~n29829;
  assign n29831 = ~n29826 & ~n29830;
  assign n29832 = pi0792 & ~n29831;
  assign n29833 = ~n20206 & ~n29832;
  assign n29834 = ~n29822 & n29833;
  assign n29835 = ~n29744 & ~n29834;
  assign n29836 = ~pi0790 & n29835;
  assign n29837 = ~pi0787 & ~n29694;
  assign n29838 = pi1157 & ~n29740;
  assign n29839 = ~n29698 & ~n29838;
  assign n29840 = pi0787 & ~n29839;
  assign n29841 = ~n29837 & ~n29840;
  assign n29842 = ~pi0644 & n29841;
  assign n29843 = pi0644 & n29835;
  assign n29844 = pi0715 & ~n29842;
  assign n29845 = ~n29843 & n29844;
  assign n29846 = ~n17804 & ~n29736;
  assign n29847 = n17804 & n29678;
  assign n29848 = ~n29846 & ~n29847;
  assign n29849 = pi0644 & ~n29848;
  assign n29850 = ~pi0644 & n29678;
  assign n29851 = ~pi0715 & ~n29850;
  assign n29852 = ~n29849 & n29851;
  assign n29853 = pi1160 & ~n29852;
  assign n29854 = ~n29845 & n29853;
  assign n29855 = ~pi0644 & ~n29848;
  assign n29856 = pi0644 & n29678;
  assign n29857 = pi0715 & ~n29856;
  assign n29858 = ~n29855 & n29857;
  assign n29859 = pi0644 & n29841;
  assign n29860 = ~pi0644 & n29835;
  assign n29861 = ~pi0715 & ~n29859;
  assign n29862 = ~n29860 & n29861;
  assign n29863 = ~pi1160 & ~n29858;
  assign n29864 = ~n29862 & n29863;
  assign n29865 = ~n29854 & ~n29864;
  assign n29866 = pi0790 & ~n29865;
  assign n29867 = pi0832 & ~n29836;
  assign n29868 = ~n29866 & n29867;
  assign po0344 = ~n29677 & ~n29868;
  assign n29870 = ~pi0188 & ~n17059;
  assign n29871 = n16635 & ~n29870;
  assign n29872 = pi0188 & ~n2571;
  assign n29873 = ~pi0188 & ~pi0705;
  assign n29874 = ~n17052 & n29873;
  assign n29875 = ~pi0188 & ~n16641;
  assign n29876 = n16647 & ~n29875;
  assign n29877 = ~pi0188 & n18072;
  assign n29878 = pi0188 & ~n18076;
  assign n29879 = ~pi0038 & ~n29878;
  assign n29880 = ~n29877 & n29879;
  assign n29881 = pi0705 & ~n29876;
  assign n29882 = ~n29880 & n29881;
  assign n29883 = n2571 & ~n29874;
  assign n29884 = ~n29882 & n29883;
  assign n29885 = ~n29872 & ~n29884;
  assign n29886 = ~pi0778 & ~n29885;
  assign n29887 = ~pi0625 & n29870;
  assign n29888 = pi0625 & n29885;
  assign n29889 = pi1153 & ~n29887;
  assign n29890 = ~n29888 & n29889;
  assign n29891 = ~pi0625 & n29885;
  assign n29892 = pi0625 & n29870;
  assign n29893 = ~pi1153 & ~n29892;
  assign n29894 = ~n29891 & n29893;
  assign n29895 = ~n29890 & ~n29894;
  assign n29896 = pi0778 & ~n29895;
  assign n29897 = ~n29886 & ~n29896;
  assign n29898 = ~n17075 & ~n29897;
  assign n29899 = n17075 & ~n29870;
  assign n29900 = ~n29898 & ~n29899;
  assign n29901 = ~n16639 & n29900;
  assign n29902 = n16639 & n29870;
  assign n29903 = ~n29901 & ~n29902;
  assign n29904 = ~n16635 & n29903;
  assign n29905 = ~n29871 & ~n29904;
  assign n29906 = ~n16631 & n29905;
  assign n29907 = n16631 & n29870;
  assign n29908 = ~n29906 & ~n29907;
  assign n29909 = ~pi0792 & n29908;
  assign n29910 = ~pi0628 & n29870;
  assign n29911 = pi0628 & ~n29908;
  assign n29912 = pi1156 & ~n29910;
  assign n29913 = ~n29911 & n29912;
  assign n29914 = pi0628 & n29870;
  assign n29915 = ~pi0628 & ~n29908;
  assign n29916 = ~pi1156 & ~n29914;
  assign n29917 = ~n29915 & n29916;
  assign n29918 = ~n29913 & ~n29917;
  assign n29919 = pi0792 & ~n29918;
  assign n29920 = ~n29909 & ~n29919;
  assign n29921 = ~pi0787 & ~n29920;
  assign n29922 = ~pi0647 & n29870;
  assign n29923 = pi0647 & n29920;
  assign n29924 = pi1157 & ~n29922;
  assign n29925 = ~n29923 & n29924;
  assign n29926 = ~pi0647 & n29920;
  assign n29927 = pi0647 & n29870;
  assign n29928 = ~pi1157 & ~n29927;
  assign n29929 = ~n29926 & n29928;
  assign n29930 = ~n29925 & ~n29929;
  assign n29931 = pi0787 & ~n29930;
  assign n29932 = ~n29921 & ~n29931;
  assign n29933 = ~pi0644 & n29932;
  assign n29934 = ~pi0618 & n29870;
  assign n29935 = ~pi0768 & ~n19439;
  assign n29936 = ~n22313 & ~n29935;
  assign n29937 = ~pi0188 & ~n29936;
  assign n29938 = ~pi0188 & ~n19433;
  assign n29939 = ~pi0768 & ~n29938;
  assign n29940 = ~n24447 & n29939;
  assign n29941 = ~n29937 & ~n29940;
  assign n29942 = n2571 & n29941;
  assign n29943 = ~n29872 & ~n29942;
  assign n29944 = ~n17117 & ~n29943;
  assign n29945 = n17117 & ~n29870;
  assign n29946 = ~n29944 & ~n29945;
  assign n29947 = ~pi0785 & ~n29946;
  assign n29948 = ~n17291 & ~n29870;
  assign n29949 = pi0609 & n29944;
  assign n29950 = ~n29948 & ~n29949;
  assign n29951 = pi1155 & ~n29950;
  assign n29952 = ~n17296 & ~n29870;
  assign n29953 = ~pi0609 & n29944;
  assign n29954 = ~n29952 & ~n29953;
  assign n29955 = ~pi1155 & ~n29954;
  assign n29956 = ~n29951 & ~n29955;
  assign n29957 = pi0785 & ~n29956;
  assign n29958 = ~n29947 & ~n29957;
  assign n29959 = pi0618 & n29958;
  assign n29960 = pi1154 & ~n29934;
  assign n29961 = ~n29959 & n29960;
  assign n29962 = pi0188 & n19468;
  assign n29963 = ~pi0188 & n19477;
  assign n29964 = pi0768 & ~n19470;
  assign n29965 = ~n29962 & n29964;
  assign n29966 = ~n29963 & n29965;
  assign n29967 = ~pi0188 & ~n19488;
  assign n29968 = pi0188 & n19496;
  assign n29969 = ~pi0768 & ~n29967;
  assign n29970 = ~n29968 & n29969;
  assign n29971 = pi0705 & ~n29970;
  assign n29972 = ~n29966 & n29971;
  assign n29973 = ~pi0705 & ~n29941;
  assign n29974 = n2571 & ~n29972;
  assign n29975 = ~n29973 & n29974;
  assign n29976 = ~n29872 & ~n29975;
  assign n29977 = ~pi0625 & n29976;
  assign n29978 = pi0625 & n29943;
  assign n29979 = ~pi1153 & ~n29978;
  assign n29980 = ~n29977 & n29979;
  assign n29981 = ~pi0608 & ~n29890;
  assign n29982 = ~n29980 & n29981;
  assign n29983 = ~pi0625 & n29943;
  assign n29984 = pi0625 & n29976;
  assign n29985 = pi1153 & ~n29983;
  assign n29986 = ~n29984 & n29985;
  assign n29987 = pi0608 & ~n29894;
  assign n29988 = ~n29986 & n29987;
  assign n29989 = ~n29982 & ~n29988;
  assign n29990 = pi0778 & ~n29989;
  assign n29991 = ~pi0778 & n29976;
  assign n29992 = ~n29990 & ~n29991;
  assign n29993 = ~pi0609 & ~n29992;
  assign n29994 = pi0609 & n29897;
  assign n29995 = ~pi1155 & ~n29994;
  assign n29996 = ~n29993 & n29995;
  assign n29997 = ~pi0660 & ~n29951;
  assign n29998 = ~n29996 & n29997;
  assign n29999 = ~pi0609 & n29897;
  assign n30000 = pi0609 & ~n29992;
  assign n30001 = pi1155 & ~n29999;
  assign n30002 = ~n30000 & n30001;
  assign n30003 = pi0660 & ~n29955;
  assign n30004 = ~n30002 & n30003;
  assign n30005 = ~n29998 & ~n30004;
  assign n30006 = pi0785 & ~n30005;
  assign n30007 = ~pi0785 & ~n29992;
  assign n30008 = ~n30006 & ~n30007;
  assign n30009 = ~pi0618 & ~n30008;
  assign n30010 = pi0618 & n29900;
  assign n30011 = ~pi1154 & ~n30010;
  assign n30012 = ~n30009 & n30011;
  assign n30013 = ~pi0627 & ~n29961;
  assign n30014 = ~n30012 & n30013;
  assign n30015 = ~pi0618 & n29958;
  assign n30016 = pi0618 & n29870;
  assign n30017 = ~pi1154 & ~n30016;
  assign n30018 = ~n30015 & n30017;
  assign n30019 = ~pi0618 & n29900;
  assign n30020 = pi0618 & ~n30008;
  assign n30021 = pi1154 & ~n30019;
  assign n30022 = ~n30020 & n30021;
  assign n30023 = pi0627 & ~n30018;
  assign n30024 = ~n30022 & n30023;
  assign n30025 = ~n30014 & ~n30024;
  assign n30026 = pi0781 & ~n30025;
  assign n30027 = ~pi0781 & ~n30008;
  assign n30028 = ~n30026 & ~n30027;
  assign n30029 = ~pi0619 & ~n30028;
  assign n30030 = pi0619 & ~n29903;
  assign n30031 = ~pi1159 & ~n30030;
  assign n30032 = ~n30029 & n30031;
  assign n30033 = ~pi0619 & n29870;
  assign n30034 = ~pi0781 & ~n29958;
  assign n30035 = ~n29961 & ~n30018;
  assign n30036 = pi0781 & ~n30035;
  assign n30037 = ~n30034 & ~n30036;
  assign n30038 = pi0619 & n30037;
  assign n30039 = pi1159 & ~n30033;
  assign n30040 = ~n30038 & n30039;
  assign n30041 = ~pi0648 & ~n30040;
  assign n30042 = ~n30032 & n30041;
  assign n30043 = pi0619 & ~n30028;
  assign n30044 = ~pi0619 & ~n29903;
  assign n30045 = pi1159 & ~n30044;
  assign n30046 = ~n30043 & n30045;
  assign n30047 = ~pi0619 & n30037;
  assign n30048 = pi0619 & n29870;
  assign n30049 = ~pi1159 & ~n30048;
  assign n30050 = ~n30047 & n30049;
  assign n30051 = pi0648 & ~n30050;
  assign n30052 = ~n30046 & n30051;
  assign n30053 = ~n30042 & ~n30052;
  assign n30054 = pi0789 & ~n30053;
  assign n30055 = ~pi0789 & ~n30028;
  assign n30056 = ~n30054 & ~n30055;
  assign n30057 = ~pi0788 & n30056;
  assign n30058 = ~pi0626 & n30056;
  assign n30059 = pi0626 & ~n29905;
  assign n30060 = ~pi0641 & ~n30059;
  assign n30061 = ~n30058 & n30060;
  assign n30062 = ~pi0789 & ~n30037;
  assign n30063 = ~n30040 & ~n30050;
  assign n30064 = pi0789 & ~n30063;
  assign n30065 = ~n30062 & ~n30064;
  assign n30066 = ~pi0626 & ~n30065;
  assign n30067 = pi0626 & ~n29870;
  assign n30068 = pi0641 & ~n30067;
  assign n30069 = ~n30066 & n30068;
  assign n30070 = ~pi1158 & ~n30069;
  assign n30071 = ~n30061 & n30070;
  assign n30072 = pi0626 & n30056;
  assign n30073 = ~pi0626 & ~n29905;
  assign n30074 = pi0641 & ~n30073;
  assign n30075 = ~n30072 & n30074;
  assign n30076 = pi0626 & ~n30065;
  assign n30077 = ~pi0626 & ~n29870;
  assign n30078 = ~pi0641 & ~n30077;
  assign n30079 = ~n30076 & n30078;
  assign n30080 = pi1158 & ~n30079;
  assign n30081 = ~n30075 & n30080;
  assign n30082 = ~n30071 & ~n30081;
  assign n30083 = pi0788 & ~n30082;
  assign n30084 = ~n30057 & ~n30083;
  assign n30085 = ~pi0628 & n30084;
  assign n30086 = ~n17969 & n30065;
  assign n30087 = n17969 & n29870;
  assign n30088 = ~n30086 & ~n30087;
  assign n30089 = pi0628 & ~n30088;
  assign n30090 = ~pi1156 & ~n30089;
  assign n30091 = ~n30085 & n30090;
  assign n30092 = ~pi0629 & ~n29913;
  assign n30093 = ~n30091 & n30092;
  assign n30094 = pi0628 & n30084;
  assign n30095 = ~pi0628 & ~n30088;
  assign n30096 = pi1156 & ~n30095;
  assign n30097 = ~n30094 & n30096;
  assign n30098 = pi0629 & ~n29917;
  assign n30099 = ~n30097 & n30098;
  assign n30100 = ~n30093 & ~n30099;
  assign n30101 = pi0792 & ~n30100;
  assign n30102 = ~pi0792 & n30084;
  assign n30103 = ~n30101 & ~n30102;
  assign n30104 = ~pi0647 & ~n30103;
  assign n30105 = ~n17779 & ~n30088;
  assign n30106 = n17779 & n29870;
  assign n30107 = ~n30105 & ~n30106;
  assign n30108 = pi0647 & ~n30107;
  assign n30109 = ~pi1157 & ~n30108;
  assign n30110 = ~n30104 & n30109;
  assign n30111 = ~pi0630 & ~n29925;
  assign n30112 = ~n30110 & n30111;
  assign n30113 = pi0647 & ~n30103;
  assign n30114 = ~pi0647 & ~n30107;
  assign n30115 = pi1157 & ~n30114;
  assign n30116 = ~n30113 & n30115;
  assign n30117 = pi0630 & ~n29929;
  assign n30118 = ~n30116 & n30117;
  assign n30119 = ~n30112 & ~n30118;
  assign n30120 = pi0787 & ~n30119;
  assign n30121 = ~pi0787 & ~n30103;
  assign n30122 = ~n30120 & ~n30121;
  assign n30123 = pi0644 & ~n30122;
  assign n30124 = pi0715 & ~n29933;
  assign n30125 = ~n30123 & n30124;
  assign n30126 = n17804 & ~n29870;
  assign n30127 = ~n17804 & n30107;
  assign n30128 = ~n30126 & ~n30127;
  assign n30129 = pi0644 & n30128;
  assign n30130 = ~pi0644 & n29870;
  assign n30131 = ~pi0715 & ~n30130;
  assign n30132 = ~n30129 & n30131;
  assign n30133 = pi1160 & ~n30132;
  assign n30134 = ~n30125 & n30133;
  assign n30135 = ~pi0644 & ~n30122;
  assign n30136 = pi0644 & n29932;
  assign n30137 = ~pi0715 & ~n30136;
  assign n30138 = ~n30135 & n30137;
  assign n30139 = ~pi0644 & n30128;
  assign n30140 = pi0644 & n29870;
  assign n30141 = pi0715 & ~n30140;
  assign n30142 = ~n30139 & n30141;
  assign n30143 = ~pi1160 & ~n30142;
  assign n30144 = ~n30138 & n30143;
  assign n30145 = pi0790 & ~n30134;
  assign n30146 = ~n30144 & n30145;
  assign n30147 = ~pi0790 & n30122;
  assign n30148 = ~po1038 & ~n30147;
  assign n30149 = ~n30146 & n30148;
  assign n30150 = ~pi0188 & po1038;
  assign n30151 = ~pi0832 & ~n30150;
  assign n30152 = ~n30149 & n30151;
  assign n30153 = ~pi0188 & ~n2926;
  assign n30154 = pi0705 & n16645;
  assign n30155 = ~n30153 & ~n30154;
  assign n30156 = ~pi0778 & n30155;
  assign n30157 = ~pi0625 & n30154;
  assign n30158 = ~n30155 & ~n30157;
  assign n30159 = pi1153 & ~n30158;
  assign n30160 = ~pi1153 & ~n30153;
  assign n30161 = ~n30157 & n30160;
  assign n30162 = ~n30159 & ~n30161;
  assign n30163 = pi0778 & ~n30162;
  assign n30164 = ~n30156 & ~n30163;
  assign n30165 = ~n17845 & n30164;
  assign n30166 = ~n17847 & n30165;
  assign n30167 = ~n17849 & n30166;
  assign n30168 = ~n17851 & n30167;
  assign n30169 = ~n17857 & n30168;
  assign n30170 = ~pi0647 & n30169;
  assign n30171 = pi0647 & n30153;
  assign n30172 = ~pi1157 & ~n30171;
  assign n30173 = ~n30170 & n30172;
  assign n30174 = pi0630 & n30173;
  assign n30175 = ~pi0768 & n17244;
  assign n30176 = ~n30153 & ~n30175;
  assign n30177 = ~n17874 & ~n30176;
  assign n30178 = ~pi0785 & ~n30177;
  assign n30179 = ~n17879 & ~n30176;
  assign n30180 = pi1155 & ~n30179;
  assign n30181 = ~n17882 & n30177;
  assign n30182 = ~pi1155 & ~n30181;
  assign n30183 = ~n30180 & ~n30182;
  assign n30184 = pi0785 & ~n30183;
  assign n30185 = ~n30178 & ~n30184;
  assign n30186 = ~pi0781 & ~n30185;
  assign n30187 = ~n17889 & n30185;
  assign n30188 = pi1154 & ~n30187;
  assign n30189 = ~n17892 & n30185;
  assign n30190 = ~pi1154 & ~n30189;
  assign n30191 = ~n30188 & ~n30190;
  assign n30192 = pi0781 & ~n30191;
  assign n30193 = ~n30186 & ~n30192;
  assign n30194 = ~pi0789 & ~n30193;
  assign n30195 = ~pi0619 & n30153;
  assign n30196 = pi0619 & n30193;
  assign n30197 = pi1159 & ~n30195;
  assign n30198 = ~n30196 & n30197;
  assign n30199 = ~pi0619 & n30193;
  assign n30200 = pi0619 & n30153;
  assign n30201 = ~pi1159 & ~n30200;
  assign n30202 = ~n30199 & n30201;
  assign n30203 = ~n30198 & ~n30202;
  assign n30204 = pi0789 & ~n30203;
  assign n30205 = ~n30194 & ~n30204;
  assign n30206 = ~n17969 & n30205;
  assign n30207 = n17969 & n30153;
  assign n30208 = ~n30206 & ~n30207;
  assign n30209 = ~n17779 & ~n30208;
  assign n30210 = n17779 & n30153;
  assign n30211 = ~n30209 & ~n30210;
  assign n30212 = ~n20559 & n30211;
  assign n30213 = pi0647 & ~n30169;
  assign n30214 = ~pi0647 & ~n30153;
  assign n30215 = ~n30213 & ~n30214;
  assign n30216 = n17801 & ~n30215;
  assign n30217 = ~n30174 & ~n30216;
  assign n30218 = ~n30212 & n30217;
  assign n30219 = pi0787 & ~n30218;
  assign n30220 = n17871 & n30167;
  assign n30221 = ~pi0626 & ~n30205;
  assign n30222 = pi0626 & ~n30153;
  assign n30223 = n16629 & ~n30222;
  assign n30224 = ~n30221 & n30223;
  assign n30225 = pi0626 & ~n30205;
  assign n30226 = ~pi0626 & ~n30153;
  assign n30227 = n16628 & ~n30226;
  assign n30228 = ~n30225 & n30227;
  assign n30229 = ~n30220 & ~n30224;
  assign n30230 = ~n30228 & n30229;
  assign n30231 = pi0788 & ~n30230;
  assign n30232 = pi0618 & n30165;
  assign n30233 = pi0609 & n30164;
  assign n30234 = ~n17168 & ~n30155;
  assign n30235 = pi0625 & n30234;
  assign n30236 = n30176 & ~n30234;
  assign n30237 = ~n30235 & ~n30236;
  assign n30238 = n30160 & ~n30237;
  assign n30239 = ~pi0608 & ~n30159;
  assign n30240 = ~n30238 & n30239;
  assign n30241 = pi1153 & n30176;
  assign n30242 = ~n30235 & n30241;
  assign n30243 = pi0608 & ~n30161;
  assign n30244 = ~n30242 & n30243;
  assign n30245 = ~n30240 & ~n30244;
  assign n30246 = pi0778 & ~n30245;
  assign n30247 = ~pi0778 & ~n30236;
  assign n30248 = ~n30246 & ~n30247;
  assign n30249 = ~pi0609 & ~n30248;
  assign n30250 = ~pi1155 & ~n30233;
  assign n30251 = ~n30249 & n30250;
  assign n30252 = ~pi0660 & ~n30180;
  assign n30253 = ~n30251 & n30252;
  assign n30254 = ~pi0609 & n30164;
  assign n30255 = pi0609 & ~n30248;
  assign n30256 = pi1155 & ~n30254;
  assign n30257 = ~n30255 & n30256;
  assign n30258 = pi0660 & ~n30182;
  assign n30259 = ~n30257 & n30258;
  assign n30260 = ~n30253 & ~n30259;
  assign n30261 = pi0785 & ~n30260;
  assign n30262 = ~pi0785 & ~n30248;
  assign n30263 = ~n30261 & ~n30262;
  assign n30264 = ~pi0618 & ~n30263;
  assign n30265 = ~pi1154 & ~n30232;
  assign n30266 = ~n30264 & n30265;
  assign n30267 = ~pi0627 & ~n30188;
  assign n30268 = ~n30266 & n30267;
  assign n30269 = ~pi0618 & n30165;
  assign n30270 = pi0618 & ~n30263;
  assign n30271 = pi1154 & ~n30269;
  assign n30272 = ~n30270 & n30271;
  assign n30273 = pi0627 & ~n30190;
  assign n30274 = ~n30272 & n30273;
  assign n30275 = ~n30268 & ~n30274;
  assign n30276 = pi0781 & ~n30275;
  assign n30277 = ~pi0781 & ~n30263;
  assign n30278 = ~n30276 & ~n30277;
  assign n30279 = ~pi0789 & n30278;
  assign n30280 = ~pi0619 & ~n30278;
  assign n30281 = pi0619 & n30166;
  assign n30282 = ~pi1159 & ~n30281;
  assign n30283 = ~n30280 & n30282;
  assign n30284 = ~pi0648 & ~n30198;
  assign n30285 = ~n30283 & n30284;
  assign n30286 = pi0619 & ~n30278;
  assign n30287 = ~pi0619 & n30166;
  assign n30288 = pi1159 & ~n30287;
  assign n30289 = ~n30286 & n30288;
  assign n30290 = pi0648 & ~n30202;
  assign n30291 = ~n30289 & n30290;
  assign n30292 = pi0789 & ~n30285;
  assign n30293 = ~n30291 & n30292;
  assign n30294 = n17970 & ~n30279;
  assign n30295 = ~n30293 & n30294;
  assign n30296 = ~n30231 & ~n30295;
  assign n30297 = ~n20364 & ~n30296;
  assign n30298 = n17854 & ~n30208;
  assign n30299 = n20851 & n30168;
  assign n30300 = ~n30298 & ~n30299;
  assign n30301 = ~pi0629 & ~n30300;
  assign n30302 = n20855 & n30168;
  assign n30303 = n17853 & ~n30208;
  assign n30304 = ~n30302 & ~n30303;
  assign n30305 = pi0629 & ~n30304;
  assign n30306 = ~n30301 & ~n30305;
  assign n30307 = pi0792 & ~n30306;
  assign n30308 = ~n20206 & ~n30307;
  assign n30309 = ~n30297 & n30308;
  assign n30310 = ~n30219 & ~n30309;
  assign n30311 = ~pi0790 & n30310;
  assign n30312 = ~pi0787 & ~n30169;
  assign n30313 = pi1157 & ~n30215;
  assign n30314 = ~n30173 & ~n30313;
  assign n30315 = pi0787 & ~n30314;
  assign n30316 = ~n30312 & ~n30315;
  assign n30317 = ~pi0644 & n30316;
  assign n30318 = pi0644 & n30310;
  assign n30319 = pi0715 & ~n30317;
  assign n30320 = ~n30318 & n30319;
  assign n30321 = ~n17804 & ~n30211;
  assign n30322 = n17804 & n30153;
  assign n30323 = ~n30321 & ~n30322;
  assign n30324 = pi0644 & ~n30323;
  assign n30325 = ~pi0644 & n30153;
  assign n30326 = ~pi0715 & ~n30325;
  assign n30327 = ~n30324 & n30326;
  assign n30328 = pi1160 & ~n30327;
  assign n30329 = ~n30320 & n30328;
  assign n30330 = ~pi0644 & ~n30323;
  assign n30331 = pi0644 & n30153;
  assign n30332 = pi0715 & ~n30331;
  assign n30333 = ~n30330 & n30332;
  assign n30334 = pi0644 & n30316;
  assign n30335 = ~pi0644 & n30310;
  assign n30336 = ~pi0715 & ~n30334;
  assign n30337 = ~n30335 & n30336;
  assign n30338 = ~pi1160 & ~n30333;
  assign n30339 = ~n30337 & n30338;
  assign n30340 = ~n30329 & ~n30339;
  assign n30341 = pi0790 & ~n30340;
  assign n30342 = pi0832 & ~n30311;
  assign n30343 = ~n30341 & n30342;
  assign po0345 = ~n30152 & ~n30343;
  assign n30345 = pi0189 & ~n17059;
  assign n30346 = n16635 & ~n30345;
  assign n30347 = n17075 & ~n30345;
  assign n30348 = pi0727 & n2571;
  assign n30349 = ~n30345 & ~n30348;
  assign n30350 = ~pi0189 & ~n16641;
  assign n30351 = n19899 & ~n30350;
  assign n30352 = ~pi0189 & n18076;
  assign n30353 = pi0189 & ~n18072;
  assign n30354 = ~pi0038 & ~n30352;
  assign n30355 = ~n30353 & n30354;
  assign n30356 = n30348 & ~n30351;
  assign n30357 = ~n30355 & n30356;
  assign n30358 = ~n30349 & ~n30357;
  assign n30359 = ~pi0778 & n30358;
  assign n30360 = ~pi0625 & ~n30345;
  assign n30361 = pi0625 & ~n30358;
  assign n30362 = pi1153 & ~n30360;
  assign n30363 = ~n30361 & n30362;
  assign n30364 = ~pi0625 & ~n30358;
  assign n30365 = pi0625 & ~n30345;
  assign n30366 = ~pi1153 & ~n30365;
  assign n30367 = ~n30364 & n30366;
  assign n30368 = ~n30363 & ~n30367;
  assign n30369 = pi0778 & ~n30368;
  assign n30370 = ~n30359 & ~n30369;
  assign n30371 = ~n17075 & n30370;
  assign n30372 = ~n30347 & ~n30371;
  assign n30373 = ~n16639 & n30372;
  assign n30374 = n16639 & n30345;
  assign n30375 = ~n30373 & ~n30374;
  assign n30376 = ~n16635 & n30375;
  assign n30377 = ~n30346 & ~n30376;
  assign n30378 = ~n16631 & n30377;
  assign n30379 = n16631 & n30345;
  assign n30380 = ~n30378 & ~n30379;
  assign n30381 = ~pi0792 & ~n30380;
  assign n30382 = ~pi0628 & ~n30345;
  assign n30383 = pi0628 & n30380;
  assign n30384 = pi1156 & ~n30382;
  assign n30385 = ~n30383 & n30384;
  assign n30386 = pi0628 & ~n30345;
  assign n30387 = ~pi0628 & n30380;
  assign n30388 = ~pi1156 & ~n30386;
  assign n30389 = ~n30387 & n30388;
  assign n30390 = ~n30385 & ~n30389;
  assign n30391 = pi0792 & ~n30390;
  assign n30392 = ~n30381 & ~n30391;
  assign n30393 = ~pi0787 & ~n30392;
  assign n30394 = ~pi0647 & ~n30345;
  assign n30395 = pi0647 & n30392;
  assign n30396 = pi1157 & ~n30394;
  assign n30397 = ~n30395 & n30396;
  assign n30398 = pi0647 & ~n30345;
  assign n30399 = ~pi0647 & n30392;
  assign n30400 = ~pi1157 & ~n30398;
  assign n30401 = ~n30399 & n30400;
  assign n30402 = ~n30397 & ~n30401;
  assign n30403 = pi0787 & ~n30402;
  assign n30404 = ~n30393 & ~n30403;
  assign n30405 = ~pi0644 & n30404;
  assign n30406 = ~pi0619 & ~n30345;
  assign n30407 = n17117 & ~n30345;
  assign n30408 = pi0189 & ~n2571;
  assign n30409 = pi0772 & n17219;
  assign n30410 = ~n22241 & ~n30409;
  assign n30411 = pi0039 & ~n30410;
  assign n30412 = ~pi0772 & n16958;
  assign n30413 = pi0772 & n17139;
  assign n30414 = ~pi0039 & ~n30412;
  assign n30415 = ~n30413 & n30414;
  assign n30416 = ~n30411 & ~n30415;
  assign n30417 = pi0189 & ~n30416;
  assign n30418 = ~pi0189 & pi0772;
  assign n30419 = n17275 & n30418;
  assign n30420 = ~n30417 & ~n30419;
  assign n30421 = ~pi0038 & ~n30420;
  assign n30422 = pi0772 & n17168;
  assign n30423 = n16641 & ~n30422;
  assign n30424 = pi0038 & ~n30350;
  assign n30425 = ~n30423 & n30424;
  assign n30426 = ~n30421 & ~n30425;
  assign n30427 = n2571 & ~n30426;
  assign n30428 = ~n30408 & ~n30427;
  assign n30429 = ~n17117 & n30428;
  assign n30430 = ~n30407 & ~n30429;
  assign n30431 = ~pi0785 & n30430;
  assign n30432 = ~pi0609 & ~n30345;
  assign n30433 = pi0609 & ~n30430;
  assign n30434 = pi1155 & ~n30432;
  assign n30435 = ~n30433 & n30434;
  assign n30436 = ~pi0609 & ~n30430;
  assign n30437 = pi0609 & ~n30345;
  assign n30438 = ~pi1155 & ~n30437;
  assign n30439 = ~n30436 & n30438;
  assign n30440 = ~n30435 & ~n30439;
  assign n30441 = pi0785 & ~n30440;
  assign n30442 = ~n30431 & ~n30441;
  assign n30443 = ~pi0781 & ~n30442;
  assign n30444 = ~pi0618 & ~n30345;
  assign n30445 = pi0618 & n30442;
  assign n30446 = pi1154 & ~n30444;
  assign n30447 = ~n30445 & n30446;
  assign n30448 = pi0618 & ~n30345;
  assign n30449 = ~pi0618 & n30442;
  assign n30450 = ~pi1154 & ~n30448;
  assign n30451 = ~n30449 & n30450;
  assign n30452 = ~n30447 & ~n30451;
  assign n30453 = pi0781 & ~n30452;
  assign n30454 = ~n30443 & ~n30453;
  assign n30455 = pi0619 & n30454;
  assign n30456 = pi1159 & ~n30406;
  assign n30457 = ~n30455 & n30456;
  assign n30458 = ~pi0727 & n30426;
  assign n30459 = ~pi0189 & ~n17605;
  assign n30460 = pi0189 & n17546;
  assign n30461 = pi0772 & ~n30460;
  assign n30462 = ~n30459 & n30461;
  assign n30463 = pi0189 & ~n17404;
  assign n30464 = ~pi0189 & ~n17485;
  assign n30465 = ~pi0772 & ~n30464;
  assign n30466 = ~n30463 & n30465;
  assign n30467 = pi0039 & ~n30462;
  assign n30468 = ~n30466 & n30467;
  assign n30469 = ~pi0189 & n17631;
  assign n30470 = pi0189 & n17629;
  assign n30471 = pi0772 & ~n30469;
  assign n30472 = ~n30470 & n30471;
  assign n30473 = ~pi0189 & ~n17625;
  assign n30474 = pi0189 & ~n17612;
  assign n30475 = ~pi0772 & ~n30473;
  assign n30476 = ~n30474 & n30475;
  assign n30477 = ~pi0039 & ~n30472;
  assign n30478 = ~n30476 & n30477;
  assign n30479 = ~pi0038 & ~n30478;
  assign n30480 = ~n30468 & n30479;
  assign n30481 = pi0727 & ~n19470;
  assign n30482 = ~n30425 & n30481;
  assign n30483 = ~n30480 & n30482;
  assign n30484 = n2571 & ~n30483;
  assign n30485 = ~n30458 & n30484;
  assign n30486 = ~n30408 & ~n30485;
  assign n30487 = ~pi0625 & n30486;
  assign n30488 = pi0625 & n30428;
  assign n30489 = ~pi1153 & ~n30488;
  assign n30490 = ~n30487 & n30489;
  assign n30491 = ~pi0608 & ~n30363;
  assign n30492 = ~n30490 & n30491;
  assign n30493 = ~pi0625 & n30428;
  assign n30494 = pi0625 & n30486;
  assign n30495 = pi1153 & ~n30493;
  assign n30496 = ~n30494 & n30495;
  assign n30497 = pi0608 & ~n30367;
  assign n30498 = ~n30496 & n30497;
  assign n30499 = ~n30492 & ~n30498;
  assign n30500 = pi0778 & ~n30499;
  assign n30501 = ~pi0778 & n30486;
  assign n30502 = ~n30500 & ~n30501;
  assign n30503 = ~pi0609 & ~n30502;
  assign n30504 = pi0609 & n30370;
  assign n30505 = ~pi1155 & ~n30504;
  assign n30506 = ~n30503 & n30505;
  assign n30507 = ~pi0660 & ~n30435;
  assign n30508 = ~n30506 & n30507;
  assign n30509 = ~pi0609 & n30370;
  assign n30510 = pi0609 & ~n30502;
  assign n30511 = pi1155 & ~n30509;
  assign n30512 = ~n30510 & n30511;
  assign n30513 = pi0660 & ~n30439;
  assign n30514 = ~n30512 & n30513;
  assign n30515 = ~n30508 & ~n30514;
  assign n30516 = pi0785 & ~n30515;
  assign n30517 = ~pi0785 & ~n30502;
  assign n30518 = ~n30516 & ~n30517;
  assign n30519 = ~pi0618 & ~n30518;
  assign n30520 = pi0618 & ~n30372;
  assign n30521 = ~pi1154 & ~n30520;
  assign n30522 = ~n30519 & n30521;
  assign n30523 = ~pi0627 & ~n30447;
  assign n30524 = ~n30522 & n30523;
  assign n30525 = pi0618 & ~n30518;
  assign n30526 = ~pi0618 & ~n30372;
  assign n30527 = pi1154 & ~n30526;
  assign n30528 = ~n30525 & n30527;
  assign n30529 = pi0627 & ~n30451;
  assign n30530 = ~n30528 & n30529;
  assign n30531 = ~n30524 & ~n30530;
  assign n30532 = pi0781 & ~n30531;
  assign n30533 = ~pi0781 & ~n30518;
  assign n30534 = ~n30532 & ~n30533;
  assign n30535 = ~pi0619 & ~n30534;
  assign n30536 = pi0619 & n30375;
  assign n30537 = ~pi1159 & ~n30536;
  assign n30538 = ~n30535 & n30537;
  assign n30539 = ~pi0648 & ~n30457;
  assign n30540 = ~n30538 & n30539;
  assign n30541 = pi0619 & ~n30345;
  assign n30542 = ~pi0619 & n30454;
  assign n30543 = ~pi1159 & ~n30541;
  assign n30544 = ~n30542 & n30543;
  assign n30545 = ~pi0619 & n30375;
  assign n30546 = pi0619 & ~n30534;
  assign n30547 = pi1159 & ~n30545;
  assign n30548 = ~n30546 & n30547;
  assign n30549 = pi0648 & ~n30544;
  assign n30550 = ~n30548 & n30549;
  assign n30551 = ~n30540 & ~n30550;
  assign n30552 = pi0789 & ~n30551;
  assign n30553 = ~pi0789 & ~n30534;
  assign n30554 = ~n30552 & ~n30553;
  assign n30555 = ~pi0788 & n30554;
  assign n30556 = ~pi0626 & n30554;
  assign n30557 = pi0626 & n30377;
  assign n30558 = ~pi0641 & ~n30557;
  assign n30559 = ~n30556 & n30558;
  assign n30560 = ~pi0789 & ~n30454;
  assign n30561 = ~n30457 & ~n30544;
  assign n30562 = pi0789 & ~n30561;
  assign n30563 = ~n30560 & ~n30562;
  assign n30564 = ~pi0626 & ~n30563;
  assign n30565 = pi0626 & n30345;
  assign n30566 = pi0641 & ~n30565;
  assign n30567 = ~n30564 & n30566;
  assign n30568 = ~pi1158 & ~n30567;
  assign n30569 = ~n30559 & n30568;
  assign n30570 = pi0626 & n30554;
  assign n30571 = ~pi0626 & n30377;
  assign n30572 = pi0641 & ~n30571;
  assign n30573 = ~n30570 & n30572;
  assign n30574 = pi0626 & ~n30563;
  assign n30575 = ~pi0626 & n30345;
  assign n30576 = ~pi0641 & ~n30575;
  assign n30577 = ~n30574 & n30576;
  assign n30578 = pi1158 & ~n30577;
  assign n30579 = ~n30573 & n30578;
  assign n30580 = ~n30569 & ~n30579;
  assign n30581 = pi0788 & ~n30580;
  assign n30582 = ~n30555 & ~n30581;
  assign n30583 = ~pi0628 & n30582;
  assign n30584 = ~n17969 & ~n30563;
  assign n30585 = n17969 & n30345;
  assign n30586 = ~n30584 & ~n30585;
  assign n30587 = pi0628 & n30586;
  assign n30588 = ~pi1156 & ~n30587;
  assign n30589 = ~n30583 & n30588;
  assign n30590 = ~pi0629 & ~n30385;
  assign n30591 = ~n30589 & n30590;
  assign n30592 = pi0628 & n30582;
  assign n30593 = ~pi0628 & n30586;
  assign n30594 = pi1156 & ~n30593;
  assign n30595 = ~n30592 & n30594;
  assign n30596 = pi0629 & ~n30389;
  assign n30597 = ~n30595 & n30596;
  assign n30598 = ~n30591 & ~n30597;
  assign n30599 = pi0792 & ~n30598;
  assign n30600 = ~pi0792 & n30582;
  assign n30601 = ~n30599 & ~n30600;
  assign n30602 = ~pi0647 & ~n30601;
  assign n30603 = ~n17779 & ~n30586;
  assign n30604 = n17779 & n30345;
  assign n30605 = ~n30603 & ~n30604;
  assign n30606 = pi0647 & n30605;
  assign n30607 = ~pi1157 & ~n30606;
  assign n30608 = ~n30602 & n30607;
  assign n30609 = ~pi0630 & ~n30397;
  assign n30610 = ~n30608 & n30609;
  assign n30611 = pi0647 & ~n30601;
  assign n30612 = ~pi0647 & n30605;
  assign n30613 = pi1157 & ~n30612;
  assign n30614 = ~n30611 & n30613;
  assign n30615 = pi0630 & ~n30401;
  assign n30616 = ~n30614 & n30615;
  assign n30617 = ~n30610 & ~n30616;
  assign n30618 = pi0787 & ~n30617;
  assign n30619 = ~pi0787 & ~n30601;
  assign n30620 = ~n30618 & ~n30619;
  assign n30621 = pi0644 & ~n30620;
  assign n30622 = pi0715 & ~n30405;
  assign n30623 = ~n30621 & n30622;
  assign n30624 = n17804 & ~n30345;
  assign n30625 = ~n17804 & n30605;
  assign n30626 = ~n30624 & ~n30625;
  assign n30627 = pi0644 & ~n30626;
  assign n30628 = ~pi0644 & ~n30345;
  assign n30629 = ~pi0715 & ~n30628;
  assign n30630 = ~n30627 & n30629;
  assign n30631 = pi1160 & ~n30630;
  assign n30632 = ~n30623 & n30631;
  assign n30633 = ~pi0644 & ~n30620;
  assign n30634 = pi0644 & n30404;
  assign n30635 = ~pi0715 & ~n30634;
  assign n30636 = ~n30633 & n30635;
  assign n30637 = ~pi0644 & ~n30626;
  assign n30638 = pi0644 & ~n30345;
  assign n30639 = pi0715 & ~n30638;
  assign n30640 = ~n30637 & n30639;
  assign n30641 = ~pi1160 & ~n30640;
  assign n30642 = ~n30636 & n30641;
  assign n30643 = pi0790 & ~n30632;
  assign n30644 = ~n30642 & n30643;
  assign n30645 = ~pi0790 & n30620;
  assign n30646 = n6305 & ~n30645;
  assign n30647 = ~n30644 & n30646;
  assign n30648 = ~pi0189 & ~n6305;
  assign n30649 = ~pi0057 & ~n30648;
  assign n30650 = ~n30647 & n30649;
  assign n30651 = pi0057 & pi0189;
  assign n30652 = ~pi0832 & ~n30651;
  assign n30653 = ~n30650 & n30652;
  assign n30654 = pi0189 & ~n2926;
  assign n30655 = pi0772 & n17244;
  assign n30656 = n17291 & n30655;
  assign n30657 = pi1155 & ~n30654;
  assign n30658 = ~n30656 & n30657;
  assign n30659 = pi0727 & n16645;
  assign n30660 = ~n30654 & ~n30659;
  assign n30661 = ~pi0778 & n30660;
  assign n30662 = pi0625 & n30659;
  assign n30663 = ~n30660 & ~n30662;
  assign n30664 = ~pi1153 & ~n30663;
  assign n30665 = pi1153 & ~n30654;
  assign n30666 = ~n30662 & n30665;
  assign n30667 = ~n30664 & ~n30666;
  assign n30668 = pi0778 & ~n30667;
  assign n30669 = ~n30661 & ~n30668;
  assign n30670 = pi0609 & n30669;
  assign n30671 = ~n30654 & ~n30655;
  assign n30672 = pi0727 & n17469;
  assign n30673 = n30671 & ~n30672;
  assign n30674 = pi0625 & n30672;
  assign n30675 = ~n30673 & ~n30674;
  assign n30676 = ~pi1153 & ~n30675;
  assign n30677 = ~pi0608 & ~n30666;
  assign n30678 = ~n30676 & n30677;
  assign n30679 = pi1153 & n30671;
  assign n30680 = ~n30674 & n30679;
  assign n30681 = pi0608 & ~n30664;
  assign n30682 = ~n30680 & n30681;
  assign n30683 = ~n30678 & ~n30682;
  assign n30684 = pi0778 & ~n30683;
  assign n30685 = ~pi0778 & ~n30673;
  assign n30686 = ~n30684 & ~n30685;
  assign n30687 = ~pi0609 & ~n30686;
  assign n30688 = ~pi1155 & ~n30670;
  assign n30689 = ~n30687 & n30688;
  assign n30690 = ~pi0660 & ~n30658;
  assign n30691 = ~n30689 & n30690;
  assign n30692 = n17296 & n30655;
  assign n30693 = ~pi1155 & ~n30654;
  assign n30694 = ~n30692 & n30693;
  assign n30695 = ~pi0609 & n30669;
  assign n30696 = pi0609 & ~n30686;
  assign n30697 = pi1155 & ~n30695;
  assign n30698 = ~n30696 & n30697;
  assign n30699 = pi0660 & ~n30694;
  assign n30700 = ~n30698 & n30699;
  assign n30701 = ~n30691 & ~n30700;
  assign n30702 = pi0785 & ~n30701;
  assign n30703 = ~pi0785 & ~n30686;
  assign n30704 = ~n30702 & ~n30703;
  assign n30705 = ~pi0781 & ~n30704;
  assign n30706 = ~n20225 & n30655;
  assign n30707 = n20319 & n30706;
  assign n30708 = ~pi1154 & ~n30654;
  assign n30709 = ~n30707 & n30708;
  assign n30710 = ~n17075 & n30669;
  assign n30711 = ~n30654 & ~n30710;
  assign n30712 = ~pi0618 & ~n30711;
  assign n30713 = pi0618 & ~n30704;
  assign n30714 = pi1154 & ~n30712;
  assign n30715 = ~n30713 & n30714;
  assign n30716 = pi0627 & ~n30709;
  assign n30717 = ~n30715 & n30716;
  assign n30718 = n20270 & n30706;
  assign n30719 = pi1154 & ~n30654;
  assign n30720 = ~n30718 & n30719;
  assign n30721 = pi0618 & ~n30711;
  assign n30722 = ~pi0618 & ~n30704;
  assign n30723 = ~pi1154 & ~n30721;
  assign n30724 = ~n30722 & n30723;
  assign n30725 = ~pi0627 & ~n30720;
  assign n30726 = ~n30724 & n30725;
  assign n30727 = ~n30717 & ~n30726;
  assign n30728 = pi0781 & ~n30727;
  assign n30729 = ~n23615 & ~n30705;
  assign n30730 = ~n30728 & n30729;
  assign n30731 = ~n20235 & n30706;
  assign n30732 = n20345 & n30731;
  assign n30733 = n16633 & ~n30732;
  assign n30734 = n19150 & n30669;
  assign n30735 = ~n23613 & ~n30734;
  assign n30736 = n20335 & n30731;
  assign n30737 = n16632 & ~n30736;
  assign n30738 = ~n30733 & ~n30737;
  assign n30739 = ~n30735 & n30738;
  assign n30740 = pi0789 & ~n30654;
  assign n30741 = ~n30739 & n30740;
  assign n30742 = n17970 & ~n30741;
  assign n30743 = ~n30730 & n30742;
  assign n30744 = ~n16635 & n30734;
  assign n30745 = ~n30654 & ~n30744;
  assign n30746 = n17865 & ~n30745;
  assign n30747 = n20237 & n30706;
  assign n30748 = ~pi0626 & n30747;
  assign n30749 = ~n30654 & ~n30748;
  assign n30750 = ~pi1158 & ~n30749;
  assign n30751 = pi0641 & ~n30750;
  assign n30752 = ~n30746 & n30751;
  assign n30753 = pi0626 & n30747;
  assign n30754 = ~n30654 & ~n30753;
  assign n30755 = pi1158 & ~n30754;
  assign n30756 = n17866 & ~n30745;
  assign n30757 = ~pi0641 & ~n30755;
  assign n30758 = ~n30756 & n30757;
  assign n30759 = pi0788 & ~n30752;
  assign n30760 = ~n30758 & n30759;
  assign n30761 = ~n20364 & ~n30760;
  assign n30762 = ~n30743 & n30761;
  assign n30763 = ~n17969 & n30747;
  assign n30764 = ~pi0629 & n30763;
  assign n30765 = pi0628 & ~n30764;
  assign n30766 = n19151 & n30669;
  assign n30767 = pi0629 & ~n30766;
  assign n30768 = ~n30765 & ~n30767;
  assign n30769 = ~pi1156 & ~n30768;
  assign n30770 = ~pi0628 & ~n30763;
  assign n30771 = pi0629 & ~n30770;
  assign n30772 = pi0628 & n30766;
  assign n30773 = pi1156 & ~n30771;
  assign n30774 = ~n30772 & n30773;
  assign n30775 = ~n30769 & ~n30774;
  assign n30776 = pi0792 & ~n30654;
  assign n30777 = ~n30775 & n30776;
  assign n30778 = ~n30762 & ~n30777;
  assign n30779 = ~n20206 & ~n30778;
  assign n30780 = ~n17779 & n30763;
  assign n30781 = ~pi0630 & n30780;
  assign n30782 = pi0647 & ~n30781;
  assign n30783 = ~n19142 & n30766;
  assign n30784 = pi0630 & ~n30783;
  assign n30785 = ~n30782 & ~n30784;
  assign n30786 = ~pi1157 & ~n30785;
  assign n30787 = pi0630 & n30780;
  assign n30788 = ~pi0630 & ~n30783;
  assign n30789 = pi0647 & ~n30788;
  assign n30790 = pi1157 & ~n30787;
  assign n30791 = ~n30789 & n30790;
  assign n30792 = ~n30786 & ~n30791;
  assign n30793 = pi0787 & ~n30654;
  assign n30794 = ~n30792 & n30793;
  assign n30795 = ~n30779 & ~n30794;
  assign n30796 = ~pi0790 & n30795;
  assign n30797 = ~n17969 & n23684;
  assign n30798 = n30747 & n30797;
  assign n30799 = pi0644 & n30798;
  assign n30800 = ~pi0715 & ~n30654;
  assign n30801 = ~n30799 & n30800;
  assign n30802 = ~n19342 & n30783;
  assign n30803 = ~n30654 & ~n30802;
  assign n30804 = ~pi0644 & ~n30803;
  assign n30805 = pi0644 & n30795;
  assign n30806 = pi0715 & ~n30804;
  assign n30807 = ~n30805 & n30806;
  assign n30808 = pi1160 & ~n30801;
  assign n30809 = ~n30807 & n30808;
  assign n30810 = ~pi0644 & n30798;
  assign n30811 = pi0715 & ~n30654;
  assign n30812 = ~n30810 & n30811;
  assign n30813 = ~pi0644 & n30795;
  assign n30814 = pi0644 & ~n30803;
  assign n30815 = ~pi0715 & ~n30814;
  assign n30816 = ~n30813 & n30815;
  assign n30817 = ~pi1160 & ~n30812;
  assign n30818 = ~n30816 & n30817;
  assign n30819 = ~n30809 & ~n30818;
  assign n30820 = pi0790 & ~n30819;
  assign n30821 = pi0832 & ~n30796;
  assign n30822 = ~n30820 & n30821;
  assign po0346 = ~n30653 & ~n30822;
  assign n30824 = ~pi0190 & ~n2926;
  assign n30825 = pi0699 & n16645;
  assign n30826 = ~n30824 & ~n30825;
  assign n30827 = ~pi0778 & ~n30826;
  assign n30828 = ~pi0625 & n30825;
  assign n30829 = ~n30826 & ~n30828;
  assign n30830 = pi1153 & ~n30829;
  assign n30831 = ~pi1153 & ~n30824;
  assign n30832 = ~n30828 & n30831;
  assign n30833 = pi0778 & ~n30832;
  assign n30834 = ~n30830 & n30833;
  assign n30835 = ~n30827 & ~n30834;
  assign n30836 = ~n17845 & ~n30835;
  assign n30837 = ~n17847 & n30836;
  assign n30838 = ~n17849 & n30837;
  assign n30839 = ~n17851 & n30838;
  assign n30840 = ~n17857 & n30839;
  assign n30841 = ~pi0647 & n30840;
  assign n30842 = pi0647 & n30824;
  assign n30843 = ~pi1157 & ~n30842;
  assign n30844 = ~n30841 & n30843;
  assign n30845 = pi0630 & n30844;
  assign n30846 = pi0763 & n17244;
  assign n30847 = ~n30824 & ~n30846;
  assign n30848 = ~n17874 & ~n30847;
  assign n30849 = ~pi0785 & ~n30848;
  assign n30850 = n17296 & n30846;
  assign n30851 = n30848 & ~n30850;
  assign n30852 = pi1155 & ~n30851;
  assign n30853 = ~pi1155 & ~n30824;
  assign n30854 = ~n30850 & n30853;
  assign n30855 = ~n30852 & ~n30854;
  assign n30856 = pi0785 & ~n30855;
  assign n30857 = ~n30849 & ~n30856;
  assign n30858 = ~pi0781 & ~n30857;
  assign n30859 = ~n17889 & n30857;
  assign n30860 = pi1154 & ~n30859;
  assign n30861 = ~n17892 & n30857;
  assign n30862 = ~pi1154 & ~n30861;
  assign n30863 = ~n30860 & ~n30862;
  assign n30864 = pi0781 & ~n30863;
  assign n30865 = ~n30858 & ~n30864;
  assign n30866 = ~pi0789 & ~n30865;
  assign n30867 = ~n23078 & n30865;
  assign n30868 = pi1159 & ~n30867;
  assign n30869 = ~n23081 & n30865;
  assign n30870 = ~pi1159 & ~n30869;
  assign n30871 = ~n30868 & ~n30870;
  assign n30872 = pi0789 & ~n30871;
  assign n30873 = ~n30866 & ~n30872;
  assign n30874 = ~n17969 & n30873;
  assign n30875 = n17969 & n30824;
  assign n30876 = ~n30874 & ~n30875;
  assign n30877 = ~n17779 & ~n30876;
  assign n30878 = n17779 & n30824;
  assign n30879 = ~n30877 & ~n30878;
  assign n30880 = ~n20559 & n30879;
  assign n30881 = pi0647 & ~n30840;
  assign n30882 = ~pi0647 & ~n30824;
  assign n30883 = ~n30881 & ~n30882;
  assign n30884 = n17801 & ~n30883;
  assign n30885 = ~n30845 & ~n30884;
  assign n30886 = ~n30880 & n30885;
  assign n30887 = pi0787 & ~n30886;
  assign n30888 = n17871 & n30838;
  assign n30889 = ~pi0626 & ~n30873;
  assign n30890 = pi0626 & ~n30824;
  assign n30891 = n16629 & ~n30890;
  assign n30892 = ~n30889 & n30891;
  assign n30893 = pi0626 & ~n30873;
  assign n30894 = ~pi0626 & ~n30824;
  assign n30895 = n16628 & ~n30894;
  assign n30896 = ~n30893 & n30895;
  assign n30897 = ~n30888 & ~n30892;
  assign n30898 = ~n30896 & n30897;
  assign n30899 = pi0788 & ~n30898;
  assign n30900 = pi0618 & n30836;
  assign n30901 = ~n17168 & ~n30826;
  assign n30902 = pi0625 & n30901;
  assign n30903 = n30847 & ~n30901;
  assign n30904 = ~n30902 & ~n30903;
  assign n30905 = n30831 & ~n30904;
  assign n30906 = ~pi0608 & ~n30830;
  assign n30907 = ~n30905 & n30906;
  assign n30908 = pi1153 & n30847;
  assign n30909 = ~n30902 & n30908;
  assign n30910 = pi0608 & ~n30832;
  assign n30911 = ~n30909 & n30910;
  assign n30912 = ~n30907 & ~n30911;
  assign n30913 = pi0778 & ~n30912;
  assign n30914 = ~pi0778 & ~n30903;
  assign n30915 = ~n30913 & ~n30914;
  assign n30916 = ~pi0609 & ~n30915;
  assign n30917 = pi0609 & ~n30835;
  assign n30918 = ~pi1155 & ~n30917;
  assign n30919 = ~n30916 & n30918;
  assign n30920 = ~pi0660 & ~n30852;
  assign n30921 = ~n30919 & n30920;
  assign n30922 = pi0609 & ~n30915;
  assign n30923 = ~pi0609 & ~n30835;
  assign n30924 = pi1155 & ~n30923;
  assign n30925 = ~n30922 & n30924;
  assign n30926 = pi0660 & ~n30854;
  assign n30927 = ~n30925 & n30926;
  assign n30928 = ~n30921 & ~n30927;
  assign n30929 = pi0785 & ~n30928;
  assign n30930 = ~pi0785 & ~n30915;
  assign n30931 = ~n30929 & ~n30930;
  assign n30932 = ~pi0618 & ~n30931;
  assign n30933 = ~pi1154 & ~n30900;
  assign n30934 = ~n30932 & n30933;
  assign n30935 = ~pi0627 & ~n30860;
  assign n30936 = ~n30934 & n30935;
  assign n30937 = ~pi0618 & n30836;
  assign n30938 = pi0618 & ~n30931;
  assign n30939 = pi1154 & ~n30937;
  assign n30940 = ~n30938 & n30939;
  assign n30941 = pi0627 & ~n30862;
  assign n30942 = ~n30940 & n30941;
  assign n30943 = ~n30936 & ~n30942;
  assign n30944 = pi0781 & ~n30943;
  assign n30945 = ~pi0781 & ~n30931;
  assign n30946 = ~n30944 & ~n30945;
  assign n30947 = ~pi0789 & n30946;
  assign n30948 = ~pi0619 & ~n30946;
  assign n30949 = pi0619 & n30837;
  assign n30950 = ~pi1159 & ~n30949;
  assign n30951 = ~n30948 & n30950;
  assign n30952 = ~pi0648 & ~n30868;
  assign n30953 = ~n30951 & n30952;
  assign n30954 = pi0619 & ~n30946;
  assign n30955 = ~pi0619 & n30837;
  assign n30956 = pi1159 & ~n30955;
  assign n30957 = ~n30954 & n30956;
  assign n30958 = pi0648 & ~n30870;
  assign n30959 = ~n30957 & n30958;
  assign n30960 = pi0789 & ~n30953;
  assign n30961 = ~n30959 & n30960;
  assign n30962 = n17970 & ~n30947;
  assign n30963 = ~n30961 & n30962;
  assign n30964 = ~n30899 & ~n30963;
  assign n30965 = ~n20364 & ~n30964;
  assign n30966 = n17854 & ~n30876;
  assign n30967 = n20851 & n30839;
  assign n30968 = ~n30966 & ~n30967;
  assign n30969 = ~pi0629 & ~n30968;
  assign n30970 = n20855 & n30839;
  assign n30971 = n17853 & ~n30876;
  assign n30972 = ~n30970 & ~n30971;
  assign n30973 = pi0629 & ~n30972;
  assign n30974 = ~n30969 & ~n30973;
  assign n30975 = pi0792 & ~n30974;
  assign n30976 = ~n20206 & ~n30975;
  assign n30977 = ~n30965 & n30976;
  assign n30978 = ~n30887 & ~n30977;
  assign n30979 = ~pi0790 & n30978;
  assign n30980 = ~pi0787 & ~n30840;
  assign n30981 = pi1157 & ~n30883;
  assign n30982 = ~n30844 & ~n30981;
  assign n30983 = pi0787 & ~n30982;
  assign n30984 = ~n30980 & ~n30983;
  assign n30985 = ~pi0644 & n30984;
  assign n30986 = pi0644 & n30978;
  assign n30987 = pi0715 & ~n30985;
  assign n30988 = ~n30986 & n30987;
  assign n30989 = ~n17804 & ~n30879;
  assign n30990 = n17804 & n30824;
  assign n30991 = ~n30989 & ~n30990;
  assign n30992 = pi0644 & ~n30991;
  assign n30993 = ~pi0644 & n30824;
  assign n30994 = ~pi0715 & ~n30993;
  assign n30995 = ~n30992 & n30994;
  assign n30996 = pi1160 & ~n30995;
  assign n30997 = ~n30988 & n30996;
  assign n30998 = ~pi0644 & ~n30991;
  assign n30999 = pi0644 & n30824;
  assign n31000 = pi0715 & ~n30999;
  assign n31001 = ~n30998 & n31000;
  assign n31002 = pi0644 & n30984;
  assign n31003 = ~pi0644 & n30978;
  assign n31004 = ~pi0715 & ~n31002;
  assign n31005 = ~n31003 & n31004;
  assign n31006 = ~pi1160 & ~n31001;
  assign n31007 = ~n31005 & n31006;
  assign n31008 = ~n30997 & ~n31007;
  assign n31009 = pi0790 & ~n31008;
  assign n31010 = pi0832 & ~n30979;
  assign n31011 = ~n31009 & n31010;
  assign n31012 = ~pi0190 & po1038;
  assign n31013 = ~pi0190 & ~n17059;
  assign n31014 = n16635 & ~n31013;
  assign n31015 = pi0190 & ~n2571;
  assign n31016 = ~pi0190 & ~n16641;
  assign n31017 = n16647 & ~n31016;
  assign n31018 = ~pi0190 & n18072;
  assign n31019 = pi0190 & ~n18076;
  assign n31020 = ~pi0038 & ~n31019;
  assign n31021 = ~n31018 & n31020;
  assign n31022 = pi0699 & ~n31017;
  assign n31023 = ~n31021 & n31022;
  assign n31024 = ~pi0190 & ~pi0699;
  assign n31025 = ~n17052 & n31024;
  assign n31026 = n2571 & ~n31025;
  assign n31027 = ~n31023 & n31026;
  assign n31028 = ~n31015 & ~n31027;
  assign n31029 = ~pi0778 & ~n31028;
  assign n31030 = ~pi0625 & n31013;
  assign n31031 = pi0625 & n31028;
  assign n31032 = pi1153 & ~n31030;
  assign n31033 = ~n31031 & n31032;
  assign n31034 = ~pi0625 & n31028;
  assign n31035 = pi0625 & n31013;
  assign n31036 = ~pi1153 & ~n31035;
  assign n31037 = ~n31034 & n31036;
  assign n31038 = ~n31033 & ~n31037;
  assign n31039 = pi0778 & ~n31038;
  assign n31040 = ~n31029 & ~n31039;
  assign n31041 = ~n17075 & ~n31040;
  assign n31042 = n17075 & ~n31013;
  assign n31043 = ~n31041 & ~n31042;
  assign n31044 = ~n16639 & n31043;
  assign n31045 = n16639 & n31013;
  assign n31046 = ~n31044 & ~n31045;
  assign n31047 = ~n16635 & n31046;
  assign n31048 = ~n31014 & ~n31047;
  assign n31049 = ~n16631 & n31048;
  assign n31050 = n16631 & n31013;
  assign n31051 = ~n31049 & ~n31050;
  assign n31052 = ~pi0628 & ~n31051;
  assign n31053 = pi0628 & n31013;
  assign n31054 = ~n31052 & ~n31053;
  assign n31055 = ~pi1156 & ~n31054;
  assign n31056 = pi0628 & ~n31051;
  assign n31057 = ~pi0628 & n31013;
  assign n31058 = ~n31056 & ~n31057;
  assign n31059 = pi1156 & ~n31058;
  assign n31060 = ~n31055 & ~n31059;
  assign n31061 = pi0792 & ~n31060;
  assign n31062 = ~pi0792 & ~n31051;
  assign n31063 = ~n31061 & ~n31062;
  assign n31064 = ~pi0647 & ~n31063;
  assign n31065 = pi0647 & n31013;
  assign n31066 = ~n31064 & ~n31065;
  assign n31067 = ~pi1157 & ~n31066;
  assign n31068 = pi0647 & ~n31063;
  assign n31069 = ~pi0647 & n31013;
  assign n31070 = ~n31068 & ~n31069;
  assign n31071 = pi1157 & ~n31070;
  assign n31072 = ~n31067 & ~n31071;
  assign n31073 = pi0787 & ~n31072;
  assign n31074 = ~pi0787 & ~n31063;
  assign n31075 = ~n31073 & ~n31074;
  assign n31076 = ~pi0644 & ~n31075;
  assign n31077 = pi0715 & ~n31076;
  assign n31078 = ~pi0763 & n17046;
  assign n31079 = pi0190 & n17273;
  assign n31080 = ~n31078 & ~n31079;
  assign n31081 = pi0039 & ~n31080;
  assign n31082 = pi0763 & ~n17234;
  assign n31083 = pi0190 & ~n31082;
  assign n31084 = ~pi0190 & pi0763;
  assign n31085 = n17221 & n31084;
  assign n31086 = ~n22358 & ~n31083;
  assign n31087 = ~n31085 & n31086;
  assign n31088 = ~n31081 & n31087;
  assign n31089 = ~pi0038 & ~n31088;
  assign n31090 = pi0763 & n17280;
  assign n31091 = pi0038 & ~n31016;
  assign n31092 = ~n31090 & n31091;
  assign n31093 = ~n31089 & ~n31092;
  assign n31094 = n2571 & ~n31093;
  assign n31095 = ~n31015 & ~n31094;
  assign n31096 = ~n17117 & ~n31095;
  assign n31097 = n17117 & ~n31013;
  assign n31098 = ~n31096 & ~n31097;
  assign n31099 = ~pi0785 & ~n31098;
  assign n31100 = ~n17291 & ~n31013;
  assign n31101 = pi0609 & n31096;
  assign n31102 = ~n31100 & ~n31101;
  assign n31103 = pi1155 & ~n31102;
  assign n31104 = ~n17296 & ~n31013;
  assign n31105 = ~pi0609 & n31096;
  assign n31106 = ~n31104 & ~n31105;
  assign n31107 = ~pi1155 & ~n31106;
  assign n31108 = ~n31103 & ~n31107;
  assign n31109 = pi0785 & ~n31108;
  assign n31110 = ~n31099 & ~n31109;
  assign n31111 = ~pi0781 & ~n31110;
  assign n31112 = ~pi0618 & n31013;
  assign n31113 = pi0618 & n31110;
  assign n31114 = pi1154 & ~n31112;
  assign n31115 = ~n31113 & n31114;
  assign n31116 = ~pi0618 & n31110;
  assign n31117 = pi0618 & n31013;
  assign n31118 = ~pi1154 & ~n31117;
  assign n31119 = ~n31116 & n31118;
  assign n31120 = ~n31115 & ~n31119;
  assign n31121 = pi0781 & ~n31120;
  assign n31122 = ~n31111 & ~n31121;
  assign n31123 = ~pi0789 & ~n31122;
  assign n31124 = ~pi0619 & n31013;
  assign n31125 = pi0619 & n31122;
  assign n31126 = pi1159 & ~n31124;
  assign n31127 = ~n31125 & n31126;
  assign n31128 = ~pi0619 & n31122;
  assign n31129 = pi0619 & n31013;
  assign n31130 = ~pi1159 & ~n31129;
  assign n31131 = ~n31128 & n31130;
  assign n31132 = ~n31127 & ~n31131;
  assign n31133 = pi0789 & ~n31132;
  assign n31134 = ~n31123 & ~n31133;
  assign n31135 = ~n17969 & n31134;
  assign n31136 = n17969 & n31013;
  assign n31137 = ~n31135 & ~n31136;
  assign n31138 = ~n17779 & ~n31137;
  assign n31139 = n17779 & n31013;
  assign n31140 = ~n31138 & ~n31139;
  assign n31141 = ~n17804 & ~n31140;
  assign n31142 = n17804 & n31013;
  assign n31143 = ~n31141 & ~n31142;
  assign n31144 = pi0644 & ~n31143;
  assign n31145 = ~pi0644 & n31013;
  assign n31146 = ~pi0715 & ~n31145;
  assign n31147 = ~n31144 & n31146;
  assign n31148 = pi1160 & ~n31147;
  assign n31149 = ~n31077 & n31148;
  assign n31150 = pi0644 & ~n31075;
  assign n31151 = ~pi0715 & ~n31150;
  assign n31152 = ~pi0644 & ~n31143;
  assign n31153 = pi0644 & n31013;
  assign n31154 = pi0715 & ~n31153;
  assign n31155 = ~n31152 & n31154;
  assign n31156 = ~pi1160 & ~n31155;
  assign n31157 = ~n31151 & n31156;
  assign n31158 = ~n31149 & ~n31157;
  assign n31159 = pi0790 & ~n31158;
  assign n31160 = n17777 & n31054;
  assign n31161 = ~n20570 & n31137;
  assign n31162 = n17776 & n31058;
  assign n31163 = ~n31160 & ~n31162;
  assign n31164 = ~n31161 & n31163;
  assign n31165 = pi0792 & ~n31164;
  assign n31166 = pi0609 & n31040;
  assign n31167 = ~pi0699 & n31093;
  assign n31168 = ~pi0763 & n24055;
  assign n31169 = ~n17490 & ~n31168;
  assign n31170 = ~pi0039 & ~n31169;
  assign n31171 = ~pi0190 & ~n31170;
  assign n31172 = ~n17469 & ~n30846;
  assign n31173 = pi0190 & ~n31172;
  assign n31174 = n6284 & n31173;
  assign n31175 = pi0038 & ~n31174;
  assign n31176 = ~n31171 & n31175;
  assign n31177 = ~pi0190 & ~n17629;
  assign n31178 = pi0190 & ~n17631;
  assign n31179 = pi0763 & ~n31178;
  assign n31180 = ~n31177 & n31179;
  assign n31181 = ~pi0190 & n17612;
  assign n31182 = pi0190 & n17625;
  assign n31183 = ~pi0763 & ~n31181;
  assign n31184 = ~n31182 & n31183;
  assign n31185 = ~pi0039 & ~n31180;
  assign n31186 = ~n31184 & n31185;
  assign n31187 = pi0190 & n17605;
  assign n31188 = ~pi0190 & ~n17546;
  assign n31189 = pi0763 & ~n31188;
  assign n31190 = ~n31187 & n31189;
  assign n31191 = ~pi0190 & n17404;
  assign n31192 = pi0190 & n17485;
  assign n31193 = ~pi0763 & ~n31192;
  assign n31194 = ~n31191 & n31193;
  assign n31195 = pi0039 & ~n31190;
  assign n31196 = ~n31194 & n31195;
  assign n31197 = ~pi0038 & ~n31186;
  assign n31198 = ~n31196 & n31197;
  assign n31199 = pi0699 & ~n31176;
  assign n31200 = ~n31198 & n31199;
  assign n31201 = n2571 & ~n31200;
  assign n31202 = ~n31167 & n31201;
  assign n31203 = ~n31015 & ~n31202;
  assign n31204 = ~pi0625 & n31203;
  assign n31205 = pi0625 & n31095;
  assign n31206 = ~pi1153 & ~n31205;
  assign n31207 = ~n31204 & n31206;
  assign n31208 = ~pi0608 & ~n31033;
  assign n31209 = ~n31207 & n31208;
  assign n31210 = ~pi0625 & n31095;
  assign n31211 = pi0625 & n31203;
  assign n31212 = pi1153 & ~n31210;
  assign n31213 = ~n31211 & n31212;
  assign n31214 = pi0608 & ~n31037;
  assign n31215 = ~n31213 & n31214;
  assign n31216 = ~n31209 & ~n31215;
  assign n31217 = pi0778 & ~n31216;
  assign n31218 = ~pi0778 & n31203;
  assign n31219 = ~n31217 & ~n31218;
  assign n31220 = ~pi0609 & ~n31219;
  assign n31221 = ~pi1155 & ~n31166;
  assign n31222 = ~n31220 & n31221;
  assign n31223 = ~pi0660 & ~n31103;
  assign n31224 = ~n31222 & n31223;
  assign n31225 = ~pi0609 & n31040;
  assign n31226 = pi0609 & ~n31219;
  assign n31227 = pi1155 & ~n31225;
  assign n31228 = ~n31226 & n31227;
  assign n31229 = pi0660 & ~n31107;
  assign n31230 = ~n31228 & n31229;
  assign n31231 = ~n31224 & ~n31230;
  assign n31232 = pi0785 & ~n31231;
  assign n31233 = ~pi0785 & ~n31219;
  assign n31234 = ~n31232 & ~n31233;
  assign n31235 = ~pi0618 & ~n31234;
  assign n31236 = pi0618 & n31043;
  assign n31237 = ~pi1154 & ~n31236;
  assign n31238 = ~n31235 & n31237;
  assign n31239 = ~pi0627 & ~n31115;
  assign n31240 = ~n31238 & n31239;
  assign n31241 = ~pi0618 & n31043;
  assign n31242 = pi0618 & ~n31234;
  assign n31243 = pi1154 & ~n31241;
  assign n31244 = ~n31242 & n31243;
  assign n31245 = pi0627 & ~n31119;
  assign n31246 = ~n31244 & n31245;
  assign n31247 = ~n31240 & ~n31246;
  assign n31248 = pi0781 & ~n31247;
  assign n31249 = ~pi0781 & ~n31234;
  assign n31250 = ~n31248 & ~n31249;
  assign n31251 = ~pi0789 & n31250;
  assign n31252 = pi0619 & ~n31046;
  assign n31253 = ~pi0619 & ~n31250;
  assign n31254 = ~pi1159 & ~n31252;
  assign n31255 = ~n31253 & n31254;
  assign n31256 = ~pi0648 & ~n31127;
  assign n31257 = ~n31255 & n31256;
  assign n31258 = ~pi0619 & ~n31046;
  assign n31259 = pi0619 & ~n31250;
  assign n31260 = pi1159 & ~n31258;
  assign n31261 = ~n31259 & n31260;
  assign n31262 = pi0648 & ~n31131;
  assign n31263 = ~n31261 & n31262;
  assign n31264 = pi0789 & ~n31257;
  assign n31265 = ~n31263 & n31264;
  assign n31266 = n17970 & ~n31251;
  assign n31267 = ~n31265 & n31266;
  assign n31268 = n17871 & n31048;
  assign n31269 = ~pi0626 & ~n31134;
  assign n31270 = pi0626 & ~n31013;
  assign n31271 = n16629 & ~n31270;
  assign n31272 = ~n31269 & n31271;
  assign n31273 = pi0626 & ~n31134;
  assign n31274 = ~pi0626 & ~n31013;
  assign n31275 = n16628 & ~n31274;
  assign n31276 = ~n31273 & n31275;
  assign n31277 = ~n31268 & ~n31272;
  assign n31278 = ~n31276 & n31277;
  assign n31279 = pi0788 & ~n31278;
  assign n31280 = ~n20364 & ~n31279;
  assign n31281 = ~n31267 & n31280;
  assign n31282 = ~n31165 & ~n31281;
  assign n31283 = ~n20206 & ~n31282;
  assign n31284 = n17802 & n31066;
  assign n31285 = ~n20559 & n31140;
  assign n31286 = n17801 & n31070;
  assign n31287 = ~n31284 & ~n31285;
  assign n31288 = ~n31286 & n31287;
  assign n31289 = pi0787 & ~n31288;
  assign n31290 = ~pi0644 & n31156;
  assign n31291 = pi0644 & n31148;
  assign n31292 = pi0790 & ~n31290;
  assign n31293 = ~n31291 & n31292;
  assign n31294 = ~n31283 & ~n31289;
  assign n31295 = ~n31293 & n31294;
  assign n31296 = ~n31159 & ~n31295;
  assign n31297 = ~po1038 & ~n31296;
  assign n31298 = ~pi0832 & ~n31012;
  assign n31299 = ~n31297 & n31298;
  assign po0347 = ~n31011 & ~n31299;
  assign n31301 = ~pi0191 & ~n2926;
  assign n31302 = pi0729 & n16645;
  assign n31303 = ~n31301 & ~n31302;
  assign n31304 = ~pi0778 & ~n31303;
  assign n31305 = ~pi0625 & n31302;
  assign n31306 = ~n31303 & ~n31305;
  assign n31307 = pi1153 & ~n31306;
  assign n31308 = ~pi1153 & ~n31301;
  assign n31309 = ~n31305 & n31308;
  assign n31310 = pi0778 & ~n31309;
  assign n31311 = ~n31307 & n31310;
  assign n31312 = ~n31304 & ~n31311;
  assign n31313 = ~n17845 & ~n31312;
  assign n31314 = ~n17847 & n31313;
  assign n31315 = ~n17849 & n31314;
  assign n31316 = ~n17851 & n31315;
  assign n31317 = ~n17857 & n31316;
  assign n31318 = ~pi0647 & n31317;
  assign n31319 = pi0647 & n31301;
  assign n31320 = ~pi1157 & ~n31319;
  assign n31321 = ~n31318 & n31320;
  assign n31322 = pi0630 & n31321;
  assign n31323 = pi0746 & n17244;
  assign n31324 = ~n31301 & ~n31323;
  assign n31325 = ~n17874 & ~n31324;
  assign n31326 = ~pi0785 & ~n31325;
  assign n31327 = n17296 & n31323;
  assign n31328 = n31325 & ~n31327;
  assign n31329 = pi1155 & ~n31328;
  assign n31330 = ~pi1155 & ~n31301;
  assign n31331 = ~n31327 & n31330;
  assign n31332 = ~n31329 & ~n31331;
  assign n31333 = pi0785 & ~n31332;
  assign n31334 = ~n31326 & ~n31333;
  assign n31335 = ~pi0781 & ~n31334;
  assign n31336 = ~n17889 & n31334;
  assign n31337 = pi1154 & ~n31336;
  assign n31338 = ~n17892 & n31334;
  assign n31339 = ~pi1154 & ~n31338;
  assign n31340 = ~n31337 & ~n31339;
  assign n31341 = pi0781 & ~n31340;
  assign n31342 = ~n31335 & ~n31341;
  assign n31343 = ~pi0789 & ~n31342;
  assign n31344 = ~n23078 & n31342;
  assign n31345 = pi1159 & ~n31344;
  assign n31346 = ~n23081 & n31342;
  assign n31347 = ~pi1159 & ~n31346;
  assign n31348 = ~n31345 & ~n31347;
  assign n31349 = pi0789 & ~n31348;
  assign n31350 = ~n31343 & ~n31349;
  assign n31351 = ~n17969 & n31350;
  assign n31352 = n17969 & n31301;
  assign n31353 = ~n31351 & ~n31352;
  assign n31354 = ~n17779 & ~n31353;
  assign n31355 = n17779 & n31301;
  assign n31356 = ~n31354 & ~n31355;
  assign n31357 = ~n20559 & n31356;
  assign n31358 = pi0647 & ~n31317;
  assign n31359 = ~pi0647 & ~n31301;
  assign n31360 = ~n31358 & ~n31359;
  assign n31361 = n17801 & ~n31360;
  assign n31362 = ~n31322 & ~n31361;
  assign n31363 = ~n31357 & n31362;
  assign n31364 = pi0787 & ~n31363;
  assign n31365 = n17871 & n31315;
  assign n31366 = ~pi0626 & ~n31350;
  assign n31367 = pi0626 & ~n31301;
  assign n31368 = n16629 & ~n31367;
  assign n31369 = ~n31366 & n31368;
  assign n31370 = pi0626 & ~n31350;
  assign n31371 = ~pi0626 & ~n31301;
  assign n31372 = n16628 & ~n31371;
  assign n31373 = ~n31370 & n31372;
  assign n31374 = ~n31365 & ~n31369;
  assign n31375 = ~n31373 & n31374;
  assign n31376 = pi0788 & ~n31375;
  assign n31377 = pi0618 & n31313;
  assign n31378 = ~n17168 & ~n31303;
  assign n31379 = pi0625 & n31378;
  assign n31380 = n31324 & ~n31378;
  assign n31381 = ~n31379 & ~n31380;
  assign n31382 = n31308 & ~n31381;
  assign n31383 = ~pi0608 & ~n31307;
  assign n31384 = ~n31382 & n31383;
  assign n31385 = pi1153 & n31324;
  assign n31386 = ~n31379 & n31385;
  assign n31387 = pi0608 & ~n31309;
  assign n31388 = ~n31386 & n31387;
  assign n31389 = ~n31384 & ~n31388;
  assign n31390 = pi0778 & ~n31389;
  assign n31391 = ~pi0778 & ~n31380;
  assign n31392 = ~n31390 & ~n31391;
  assign n31393 = ~pi0609 & ~n31392;
  assign n31394 = pi0609 & ~n31312;
  assign n31395 = ~pi1155 & ~n31394;
  assign n31396 = ~n31393 & n31395;
  assign n31397 = ~pi0660 & ~n31329;
  assign n31398 = ~n31396 & n31397;
  assign n31399 = pi0609 & ~n31392;
  assign n31400 = ~pi0609 & ~n31312;
  assign n31401 = pi1155 & ~n31400;
  assign n31402 = ~n31399 & n31401;
  assign n31403 = pi0660 & ~n31331;
  assign n31404 = ~n31402 & n31403;
  assign n31405 = ~n31398 & ~n31404;
  assign n31406 = pi0785 & ~n31405;
  assign n31407 = ~pi0785 & ~n31392;
  assign n31408 = ~n31406 & ~n31407;
  assign n31409 = ~pi0618 & ~n31408;
  assign n31410 = ~pi1154 & ~n31377;
  assign n31411 = ~n31409 & n31410;
  assign n31412 = ~pi0627 & ~n31337;
  assign n31413 = ~n31411 & n31412;
  assign n31414 = ~pi0618 & n31313;
  assign n31415 = pi0618 & ~n31408;
  assign n31416 = pi1154 & ~n31414;
  assign n31417 = ~n31415 & n31416;
  assign n31418 = pi0627 & ~n31339;
  assign n31419 = ~n31417 & n31418;
  assign n31420 = ~n31413 & ~n31419;
  assign n31421 = pi0781 & ~n31420;
  assign n31422 = ~pi0781 & ~n31408;
  assign n31423 = ~n31421 & ~n31422;
  assign n31424 = ~pi0789 & n31423;
  assign n31425 = ~pi0619 & ~n31423;
  assign n31426 = pi0619 & n31314;
  assign n31427 = ~pi1159 & ~n31426;
  assign n31428 = ~n31425 & n31427;
  assign n31429 = ~pi0648 & ~n31345;
  assign n31430 = ~n31428 & n31429;
  assign n31431 = pi0619 & ~n31423;
  assign n31432 = ~pi0619 & n31314;
  assign n31433 = pi1159 & ~n31432;
  assign n31434 = ~n31431 & n31433;
  assign n31435 = pi0648 & ~n31347;
  assign n31436 = ~n31434 & n31435;
  assign n31437 = pi0789 & ~n31430;
  assign n31438 = ~n31436 & n31437;
  assign n31439 = n17970 & ~n31424;
  assign n31440 = ~n31438 & n31439;
  assign n31441 = ~n31376 & ~n31440;
  assign n31442 = ~n20364 & ~n31441;
  assign n31443 = n17854 & ~n31353;
  assign n31444 = n20851 & n31316;
  assign n31445 = ~n31443 & ~n31444;
  assign n31446 = ~pi0629 & ~n31445;
  assign n31447 = n20855 & n31316;
  assign n31448 = n17853 & ~n31353;
  assign n31449 = ~n31447 & ~n31448;
  assign n31450 = pi0629 & ~n31449;
  assign n31451 = ~n31446 & ~n31450;
  assign n31452 = pi0792 & ~n31451;
  assign n31453 = ~n20206 & ~n31452;
  assign n31454 = ~n31442 & n31453;
  assign n31455 = ~n31364 & ~n31454;
  assign n31456 = ~pi0790 & n31455;
  assign n31457 = ~pi0787 & ~n31317;
  assign n31458 = pi1157 & ~n31360;
  assign n31459 = ~n31321 & ~n31458;
  assign n31460 = pi0787 & ~n31459;
  assign n31461 = ~n31457 & ~n31460;
  assign n31462 = ~pi0644 & n31461;
  assign n31463 = pi0644 & n31455;
  assign n31464 = pi0715 & ~n31462;
  assign n31465 = ~n31463 & n31464;
  assign n31466 = ~n17804 & ~n31356;
  assign n31467 = n17804 & n31301;
  assign n31468 = ~n31466 & ~n31467;
  assign n31469 = pi0644 & ~n31468;
  assign n31470 = ~pi0644 & n31301;
  assign n31471 = ~pi0715 & ~n31470;
  assign n31472 = ~n31469 & n31471;
  assign n31473 = pi1160 & ~n31472;
  assign n31474 = ~n31465 & n31473;
  assign n31475 = ~pi0644 & ~n31468;
  assign n31476 = pi0644 & n31301;
  assign n31477 = pi0715 & ~n31476;
  assign n31478 = ~n31475 & n31477;
  assign n31479 = pi0644 & n31461;
  assign n31480 = ~pi0644 & n31455;
  assign n31481 = ~pi0715 & ~n31479;
  assign n31482 = ~n31480 & n31481;
  assign n31483 = ~pi1160 & ~n31478;
  assign n31484 = ~n31482 & n31483;
  assign n31485 = ~n31474 & ~n31484;
  assign n31486 = pi0790 & ~n31485;
  assign n31487 = pi0832 & ~n31456;
  assign n31488 = ~n31486 & n31487;
  assign n31489 = ~pi0191 & po1038;
  assign n31490 = ~pi0191 & ~n17059;
  assign n31491 = n16635 & ~n31490;
  assign n31492 = pi0191 & ~n2571;
  assign n31493 = ~pi0191 & ~n16641;
  assign n31494 = n16647 & ~n31493;
  assign n31495 = ~pi0191 & n18072;
  assign n31496 = pi0191 & ~n18076;
  assign n31497 = ~pi0038 & ~n31496;
  assign n31498 = ~n31495 & n31497;
  assign n31499 = pi0729 & ~n31494;
  assign n31500 = ~n31498 & n31499;
  assign n31501 = ~pi0191 & ~pi0729;
  assign n31502 = ~n17052 & n31501;
  assign n31503 = n2571 & ~n31502;
  assign n31504 = ~n31500 & n31503;
  assign n31505 = ~n31492 & ~n31504;
  assign n31506 = ~pi0778 & ~n31505;
  assign n31507 = ~pi0625 & n31490;
  assign n31508 = pi0625 & n31505;
  assign n31509 = pi1153 & ~n31507;
  assign n31510 = ~n31508 & n31509;
  assign n31511 = ~pi0625 & n31505;
  assign n31512 = pi0625 & n31490;
  assign n31513 = ~pi1153 & ~n31512;
  assign n31514 = ~n31511 & n31513;
  assign n31515 = ~n31510 & ~n31514;
  assign n31516 = pi0778 & ~n31515;
  assign n31517 = ~n31506 & ~n31516;
  assign n31518 = ~n17075 & ~n31517;
  assign n31519 = n17075 & ~n31490;
  assign n31520 = ~n31518 & ~n31519;
  assign n31521 = ~n16639 & n31520;
  assign n31522 = n16639 & n31490;
  assign n31523 = ~n31521 & ~n31522;
  assign n31524 = ~n16635 & n31523;
  assign n31525 = ~n31491 & ~n31524;
  assign n31526 = ~n16631 & n31525;
  assign n31527 = n16631 & n31490;
  assign n31528 = ~n31526 & ~n31527;
  assign n31529 = ~pi0628 & ~n31528;
  assign n31530 = pi0628 & n31490;
  assign n31531 = ~n31529 & ~n31530;
  assign n31532 = ~pi1156 & ~n31531;
  assign n31533 = pi0628 & ~n31528;
  assign n31534 = ~pi0628 & n31490;
  assign n31535 = ~n31533 & ~n31534;
  assign n31536 = pi1156 & ~n31535;
  assign n31537 = ~n31532 & ~n31536;
  assign n31538 = pi0792 & ~n31537;
  assign n31539 = ~pi0792 & ~n31528;
  assign n31540 = ~n31538 & ~n31539;
  assign n31541 = ~pi0647 & ~n31540;
  assign n31542 = pi0647 & n31490;
  assign n31543 = ~n31541 & ~n31542;
  assign n31544 = ~pi1157 & ~n31543;
  assign n31545 = pi0647 & ~n31540;
  assign n31546 = ~pi0647 & n31490;
  assign n31547 = ~n31545 & ~n31546;
  assign n31548 = pi1157 & ~n31547;
  assign n31549 = ~n31544 & ~n31548;
  assign n31550 = pi0787 & ~n31549;
  assign n31551 = ~pi0787 & ~n31540;
  assign n31552 = ~n31550 & ~n31551;
  assign n31553 = ~pi0644 & ~n31552;
  assign n31554 = pi0715 & ~n31553;
  assign n31555 = ~pi0746 & n17046;
  assign n31556 = pi0191 & n17273;
  assign n31557 = ~n31555 & ~n31556;
  assign n31558 = pi0039 & ~n31557;
  assign n31559 = pi0746 & ~n17234;
  assign n31560 = pi0191 & ~n31559;
  assign n31561 = ~pi0191 & pi0746;
  assign n31562 = n17221 & n31561;
  assign n31563 = ~n22439 & ~n31560;
  assign n31564 = ~n31562 & n31563;
  assign n31565 = ~n31558 & n31564;
  assign n31566 = ~pi0038 & ~n31565;
  assign n31567 = pi0746 & n17280;
  assign n31568 = pi0038 & ~n31493;
  assign n31569 = ~n31567 & n31568;
  assign n31570 = ~n31566 & ~n31569;
  assign n31571 = n2571 & ~n31570;
  assign n31572 = ~n31492 & ~n31571;
  assign n31573 = ~n17117 & ~n31572;
  assign n31574 = n17117 & ~n31490;
  assign n31575 = ~n31573 & ~n31574;
  assign n31576 = ~pi0785 & ~n31575;
  assign n31577 = ~n17291 & ~n31490;
  assign n31578 = pi0609 & n31573;
  assign n31579 = ~n31577 & ~n31578;
  assign n31580 = pi1155 & ~n31579;
  assign n31581 = ~n17296 & ~n31490;
  assign n31582 = ~pi0609 & n31573;
  assign n31583 = ~n31581 & ~n31582;
  assign n31584 = ~pi1155 & ~n31583;
  assign n31585 = ~n31580 & ~n31584;
  assign n31586 = pi0785 & ~n31585;
  assign n31587 = ~n31576 & ~n31586;
  assign n31588 = ~pi0781 & ~n31587;
  assign n31589 = ~pi0618 & n31490;
  assign n31590 = pi0618 & n31587;
  assign n31591 = pi1154 & ~n31589;
  assign n31592 = ~n31590 & n31591;
  assign n31593 = ~pi0618 & n31587;
  assign n31594 = pi0618 & n31490;
  assign n31595 = ~pi1154 & ~n31594;
  assign n31596 = ~n31593 & n31595;
  assign n31597 = ~n31592 & ~n31596;
  assign n31598 = pi0781 & ~n31597;
  assign n31599 = ~n31588 & ~n31598;
  assign n31600 = ~pi0789 & ~n31599;
  assign n31601 = ~pi0619 & n31490;
  assign n31602 = pi0619 & n31599;
  assign n31603 = pi1159 & ~n31601;
  assign n31604 = ~n31602 & n31603;
  assign n31605 = ~pi0619 & n31599;
  assign n31606 = pi0619 & n31490;
  assign n31607 = ~pi1159 & ~n31606;
  assign n31608 = ~n31605 & n31607;
  assign n31609 = ~n31604 & ~n31608;
  assign n31610 = pi0789 & ~n31609;
  assign n31611 = ~n31600 & ~n31610;
  assign n31612 = ~n17969 & n31611;
  assign n31613 = n17969 & n31490;
  assign n31614 = ~n31612 & ~n31613;
  assign n31615 = ~n17779 & ~n31614;
  assign n31616 = n17779 & n31490;
  assign n31617 = ~n31615 & ~n31616;
  assign n31618 = ~n17804 & ~n31617;
  assign n31619 = n17804 & n31490;
  assign n31620 = ~n31618 & ~n31619;
  assign n31621 = pi0644 & ~n31620;
  assign n31622 = ~pi0644 & n31490;
  assign n31623 = ~pi0715 & ~n31622;
  assign n31624 = ~n31621 & n31623;
  assign n31625 = pi1160 & ~n31624;
  assign n31626 = ~n31554 & n31625;
  assign n31627 = pi0644 & ~n31552;
  assign n31628 = ~pi0715 & ~n31627;
  assign n31629 = ~pi0644 & ~n31620;
  assign n31630 = pi0644 & n31490;
  assign n31631 = pi0715 & ~n31630;
  assign n31632 = ~n31629 & n31631;
  assign n31633 = ~pi1160 & ~n31632;
  assign n31634 = ~n31628 & n31633;
  assign n31635 = ~n31626 & ~n31634;
  assign n31636 = pi0790 & ~n31635;
  assign n31637 = n17777 & n31531;
  assign n31638 = ~n20570 & n31614;
  assign n31639 = n17776 & n31535;
  assign n31640 = ~n31637 & ~n31639;
  assign n31641 = ~n31638 & n31640;
  assign n31642 = pi0792 & ~n31641;
  assign n31643 = pi0609 & n31517;
  assign n31644 = ~pi0729 & n31570;
  assign n31645 = ~pi0746 & n24055;
  assign n31646 = ~n17490 & ~n31645;
  assign n31647 = ~pi0039 & ~n31646;
  assign n31648 = ~pi0191 & ~n31647;
  assign n31649 = ~n17469 & ~n31323;
  assign n31650 = pi0191 & ~n31649;
  assign n31651 = n6284 & n31650;
  assign n31652 = pi0038 & ~n31651;
  assign n31653 = ~n31648 & n31652;
  assign n31654 = ~pi0191 & ~n17629;
  assign n31655 = pi0191 & ~n17631;
  assign n31656 = pi0746 & ~n31655;
  assign n31657 = ~n31654 & n31656;
  assign n31658 = ~pi0191 & n17612;
  assign n31659 = pi0191 & n17625;
  assign n31660 = ~pi0746 & ~n31658;
  assign n31661 = ~n31659 & n31660;
  assign n31662 = ~pi0039 & ~n31657;
  assign n31663 = ~n31661 & n31662;
  assign n31664 = pi0191 & n17605;
  assign n31665 = ~pi0191 & ~n17546;
  assign n31666 = pi0746 & ~n31665;
  assign n31667 = ~n31664 & n31666;
  assign n31668 = ~pi0191 & n17404;
  assign n31669 = pi0191 & n17485;
  assign n31670 = ~pi0746 & ~n31669;
  assign n31671 = ~n31668 & n31670;
  assign n31672 = pi0039 & ~n31667;
  assign n31673 = ~n31671 & n31672;
  assign n31674 = ~pi0038 & ~n31663;
  assign n31675 = ~n31673 & n31674;
  assign n31676 = pi0729 & ~n31653;
  assign n31677 = ~n31675 & n31676;
  assign n31678 = n2571 & ~n31677;
  assign n31679 = ~n31644 & n31678;
  assign n31680 = ~n31492 & ~n31679;
  assign n31681 = ~pi0625 & n31680;
  assign n31682 = pi0625 & n31572;
  assign n31683 = ~pi1153 & ~n31682;
  assign n31684 = ~n31681 & n31683;
  assign n31685 = ~pi0608 & ~n31510;
  assign n31686 = ~n31684 & n31685;
  assign n31687 = ~pi0625 & n31572;
  assign n31688 = pi0625 & n31680;
  assign n31689 = pi1153 & ~n31687;
  assign n31690 = ~n31688 & n31689;
  assign n31691 = pi0608 & ~n31514;
  assign n31692 = ~n31690 & n31691;
  assign n31693 = ~n31686 & ~n31692;
  assign n31694 = pi0778 & ~n31693;
  assign n31695 = ~pi0778 & n31680;
  assign n31696 = ~n31694 & ~n31695;
  assign n31697 = ~pi0609 & ~n31696;
  assign n31698 = ~pi1155 & ~n31643;
  assign n31699 = ~n31697 & n31698;
  assign n31700 = ~pi0660 & ~n31580;
  assign n31701 = ~n31699 & n31700;
  assign n31702 = ~pi0609 & n31517;
  assign n31703 = pi0609 & ~n31696;
  assign n31704 = pi1155 & ~n31702;
  assign n31705 = ~n31703 & n31704;
  assign n31706 = pi0660 & ~n31584;
  assign n31707 = ~n31705 & n31706;
  assign n31708 = ~n31701 & ~n31707;
  assign n31709 = pi0785 & ~n31708;
  assign n31710 = ~pi0785 & ~n31696;
  assign n31711 = ~n31709 & ~n31710;
  assign n31712 = ~pi0618 & ~n31711;
  assign n31713 = pi0618 & n31520;
  assign n31714 = ~pi1154 & ~n31713;
  assign n31715 = ~n31712 & n31714;
  assign n31716 = ~pi0627 & ~n31592;
  assign n31717 = ~n31715 & n31716;
  assign n31718 = ~pi0618 & n31520;
  assign n31719 = pi0618 & ~n31711;
  assign n31720 = pi1154 & ~n31718;
  assign n31721 = ~n31719 & n31720;
  assign n31722 = pi0627 & ~n31596;
  assign n31723 = ~n31721 & n31722;
  assign n31724 = ~n31717 & ~n31723;
  assign n31725 = pi0781 & ~n31724;
  assign n31726 = ~pi0781 & ~n31711;
  assign n31727 = ~n31725 & ~n31726;
  assign n31728 = ~pi0789 & n31727;
  assign n31729 = pi0619 & ~n31523;
  assign n31730 = ~pi0619 & ~n31727;
  assign n31731 = ~pi1159 & ~n31729;
  assign n31732 = ~n31730 & n31731;
  assign n31733 = ~pi0648 & ~n31604;
  assign n31734 = ~n31732 & n31733;
  assign n31735 = ~pi0619 & ~n31523;
  assign n31736 = pi0619 & ~n31727;
  assign n31737 = pi1159 & ~n31735;
  assign n31738 = ~n31736 & n31737;
  assign n31739 = pi0648 & ~n31608;
  assign n31740 = ~n31738 & n31739;
  assign n31741 = pi0789 & ~n31734;
  assign n31742 = ~n31740 & n31741;
  assign n31743 = n17970 & ~n31728;
  assign n31744 = ~n31742 & n31743;
  assign n31745 = n17871 & n31525;
  assign n31746 = ~pi0626 & ~n31611;
  assign n31747 = pi0626 & ~n31490;
  assign n31748 = n16629 & ~n31747;
  assign n31749 = ~n31746 & n31748;
  assign n31750 = pi0626 & ~n31611;
  assign n31751 = ~pi0626 & ~n31490;
  assign n31752 = n16628 & ~n31751;
  assign n31753 = ~n31750 & n31752;
  assign n31754 = ~n31745 & ~n31749;
  assign n31755 = ~n31753 & n31754;
  assign n31756 = pi0788 & ~n31755;
  assign n31757 = ~n20364 & ~n31756;
  assign n31758 = ~n31744 & n31757;
  assign n31759 = ~n31642 & ~n31758;
  assign n31760 = ~n20206 & ~n31759;
  assign n31761 = n17802 & n31543;
  assign n31762 = ~n20559 & n31617;
  assign n31763 = n17801 & n31547;
  assign n31764 = ~n31761 & ~n31762;
  assign n31765 = ~n31763 & n31764;
  assign n31766 = pi0787 & ~n31765;
  assign n31767 = ~pi0644 & n31633;
  assign n31768 = pi0644 & n31625;
  assign n31769 = pi0790 & ~n31767;
  assign n31770 = ~n31768 & n31769;
  assign n31771 = ~n31760 & ~n31766;
  assign n31772 = ~n31770 & n31771;
  assign n31773 = ~n31636 & ~n31772;
  assign n31774 = ~po1038 & ~n31773;
  assign n31775 = ~pi0832 & ~n31489;
  assign n31776 = ~n31774 & n31775;
  assign po0348 = ~n31488 & ~n31776;
  assign n31778 = ~pi0192 & ~n2926;
  assign n31779 = pi0691 & n16645;
  assign n31780 = ~n31778 & ~n31779;
  assign n31781 = ~pi0778 & ~n31780;
  assign n31782 = ~pi0625 & n31779;
  assign n31783 = ~n31780 & ~n31782;
  assign n31784 = pi1153 & ~n31783;
  assign n31785 = ~pi1153 & ~n31778;
  assign n31786 = ~n31782 & n31785;
  assign n31787 = pi0778 & ~n31786;
  assign n31788 = ~n31784 & n31787;
  assign n31789 = ~n31781 & ~n31788;
  assign n31790 = ~n17845 & ~n31789;
  assign n31791 = ~n17847 & n31790;
  assign n31792 = ~n17849 & n31791;
  assign n31793 = ~n17851 & n31792;
  assign n31794 = ~n17857 & n31793;
  assign n31795 = ~pi0647 & n31794;
  assign n31796 = pi0647 & n31778;
  assign n31797 = ~pi1157 & ~n31796;
  assign n31798 = ~n31795 & n31797;
  assign n31799 = pi0630 & n31798;
  assign n31800 = pi0764 & n17244;
  assign n31801 = ~n31778 & ~n31800;
  assign n31802 = ~n17874 & ~n31801;
  assign n31803 = ~pi0785 & ~n31802;
  assign n31804 = n17296 & n31800;
  assign n31805 = n31802 & ~n31804;
  assign n31806 = pi1155 & ~n31805;
  assign n31807 = ~pi1155 & ~n31778;
  assign n31808 = ~n31804 & n31807;
  assign n31809 = ~n31806 & ~n31808;
  assign n31810 = pi0785 & ~n31809;
  assign n31811 = ~n31803 & ~n31810;
  assign n31812 = ~pi0781 & ~n31811;
  assign n31813 = ~n17889 & n31811;
  assign n31814 = pi1154 & ~n31813;
  assign n31815 = ~n17892 & n31811;
  assign n31816 = ~pi1154 & ~n31815;
  assign n31817 = ~n31814 & ~n31816;
  assign n31818 = pi0781 & ~n31817;
  assign n31819 = ~n31812 & ~n31818;
  assign n31820 = ~pi0789 & ~n31819;
  assign n31821 = ~n23078 & n31819;
  assign n31822 = pi1159 & ~n31821;
  assign n31823 = ~n23081 & n31819;
  assign n31824 = ~pi1159 & ~n31823;
  assign n31825 = ~n31822 & ~n31824;
  assign n31826 = pi0789 & ~n31825;
  assign n31827 = ~n31820 & ~n31826;
  assign n31828 = ~n17969 & n31827;
  assign n31829 = n17969 & n31778;
  assign n31830 = ~n31828 & ~n31829;
  assign n31831 = ~n17779 & ~n31830;
  assign n31832 = n17779 & n31778;
  assign n31833 = ~n31831 & ~n31832;
  assign n31834 = ~n20559 & n31833;
  assign n31835 = pi0647 & ~n31794;
  assign n31836 = ~pi0647 & ~n31778;
  assign n31837 = ~n31835 & ~n31836;
  assign n31838 = n17801 & ~n31837;
  assign n31839 = ~n31799 & ~n31838;
  assign n31840 = ~n31834 & n31839;
  assign n31841 = pi0787 & ~n31840;
  assign n31842 = n17871 & n31792;
  assign n31843 = ~pi0626 & ~n31827;
  assign n31844 = pi0626 & ~n31778;
  assign n31845 = n16629 & ~n31844;
  assign n31846 = ~n31843 & n31845;
  assign n31847 = pi0626 & ~n31827;
  assign n31848 = ~pi0626 & ~n31778;
  assign n31849 = n16628 & ~n31848;
  assign n31850 = ~n31847 & n31849;
  assign n31851 = ~n31842 & ~n31846;
  assign n31852 = ~n31850 & n31851;
  assign n31853 = pi0788 & ~n31852;
  assign n31854 = pi0618 & n31790;
  assign n31855 = ~n17168 & ~n31780;
  assign n31856 = pi0625 & n31855;
  assign n31857 = n31801 & ~n31855;
  assign n31858 = ~n31856 & ~n31857;
  assign n31859 = n31785 & ~n31858;
  assign n31860 = ~pi0608 & ~n31784;
  assign n31861 = ~n31859 & n31860;
  assign n31862 = pi1153 & n31801;
  assign n31863 = ~n31856 & n31862;
  assign n31864 = pi0608 & ~n31786;
  assign n31865 = ~n31863 & n31864;
  assign n31866 = ~n31861 & ~n31865;
  assign n31867 = pi0778 & ~n31866;
  assign n31868 = ~pi0778 & ~n31857;
  assign n31869 = ~n31867 & ~n31868;
  assign n31870 = ~pi0609 & ~n31869;
  assign n31871 = pi0609 & ~n31789;
  assign n31872 = ~pi1155 & ~n31871;
  assign n31873 = ~n31870 & n31872;
  assign n31874 = ~pi0660 & ~n31806;
  assign n31875 = ~n31873 & n31874;
  assign n31876 = pi0609 & ~n31869;
  assign n31877 = ~pi0609 & ~n31789;
  assign n31878 = pi1155 & ~n31877;
  assign n31879 = ~n31876 & n31878;
  assign n31880 = pi0660 & ~n31808;
  assign n31881 = ~n31879 & n31880;
  assign n31882 = ~n31875 & ~n31881;
  assign n31883 = pi0785 & ~n31882;
  assign n31884 = ~pi0785 & ~n31869;
  assign n31885 = ~n31883 & ~n31884;
  assign n31886 = ~pi0618 & ~n31885;
  assign n31887 = ~pi1154 & ~n31854;
  assign n31888 = ~n31886 & n31887;
  assign n31889 = ~pi0627 & ~n31814;
  assign n31890 = ~n31888 & n31889;
  assign n31891 = ~pi0618 & n31790;
  assign n31892 = pi0618 & ~n31885;
  assign n31893 = pi1154 & ~n31891;
  assign n31894 = ~n31892 & n31893;
  assign n31895 = pi0627 & ~n31816;
  assign n31896 = ~n31894 & n31895;
  assign n31897 = ~n31890 & ~n31896;
  assign n31898 = pi0781 & ~n31897;
  assign n31899 = ~pi0781 & ~n31885;
  assign n31900 = ~n31898 & ~n31899;
  assign n31901 = ~pi0789 & n31900;
  assign n31902 = ~pi0619 & ~n31900;
  assign n31903 = pi0619 & n31791;
  assign n31904 = ~pi1159 & ~n31903;
  assign n31905 = ~n31902 & n31904;
  assign n31906 = ~pi0648 & ~n31822;
  assign n31907 = ~n31905 & n31906;
  assign n31908 = pi0619 & ~n31900;
  assign n31909 = ~pi0619 & n31791;
  assign n31910 = pi1159 & ~n31909;
  assign n31911 = ~n31908 & n31910;
  assign n31912 = pi0648 & ~n31824;
  assign n31913 = ~n31911 & n31912;
  assign n31914 = pi0789 & ~n31907;
  assign n31915 = ~n31913 & n31914;
  assign n31916 = n17970 & ~n31901;
  assign n31917 = ~n31915 & n31916;
  assign n31918 = ~n31853 & ~n31917;
  assign n31919 = ~n20364 & ~n31918;
  assign n31920 = n17854 & ~n31830;
  assign n31921 = n20851 & n31793;
  assign n31922 = ~n31920 & ~n31921;
  assign n31923 = ~pi0629 & ~n31922;
  assign n31924 = n20855 & n31793;
  assign n31925 = n17853 & ~n31830;
  assign n31926 = ~n31924 & ~n31925;
  assign n31927 = pi0629 & ~n31926;
  assign n31928 = ~n31923 & ~n31927;
  assign n31929 = pi0792 & ~n31928;
  assign n31930 = ~n20206 & ~n31929;
  assign n31931 = ~n31919 & n31930;
  assign n31932 = ~n31841 & ~n31931;
  assign n31933 = ~pi0790 & n31932;
  assign n31934 = ~pi0787 & ~n31794;
  assign n31935 = pi1157 & ~n31837;
  assign n31936 = ~n31798 & ~n31935;
  assign n31937 = pi0787 & ~n31936;
  assign n31938 = ~n31934 & ~n31937;
  assign n31939 = ~pi0644 & n31938;
  assign n31940 = pi0644 & n31932;
  assign n31941 = pi0715 & ~n31939;
  assign n31942 = ~n31940 & n31941;
  assign n31943 = ~n17804 & ~n31833;
  assign n31944 = n17804 & n31778;
  assign n31945 = ~n31943 & ~n31944;
  assign n31946 = pi0644 & ~n31945;
  assign n31947 = ~pi0644 & n31778;
  assign n31948 = ~pi0715 & ~n31947;
  assign n31949 = ~n31946 & n31948;
  assign n31950 = pi1160 & ~n31949;
  assign n31951 = ~n31942 & n31950;
  assign n31952 = ~pi0644 & ~n31945;
  assign n31953 = pi0644 & n31778;
  assign n31954 = pi0715 & ~n31953;
  assign n31955 = ~n31952 & n31954;
  assign n31956 = pi0644 & n31938;
  assign n31957 = ~pi0644 & n31932;
  assign n31958 = ~pi0715 & ~n31956;
  assign n31959 = ~n31957 & n31958;
  assign n31960 = ~pi1160 & ~n31955;
  assign n31961 = ~n31959 & n31960;
  assign n31962 = ~n31951 & ~n31961;
  assign n31963 = pi0790 & ~n31962;
  assign n31964 = pi0832 & ~n31933;
  assign n31965 = ~n31963 & n31964;
  assign n31966 = ~pi0192 & po1038;
  assign n31967 = ~pi0192 & ~n17059;
  assign n31968 = n16635 & ~n31967;
  assign n31969 = pi0192 & ~n2571;
  assign n31970 = ~pi0192 & ~n16641;
  assign n31971 = n16647 & ~n31970;
  assign n31972 = ~pi0192 & n18072;
  assign n31973 = pi0192 & ~n18076;
  assign n31974 = ~pi0038 & ~n31973;
  assign n31975 = ~n31972 & n31974;
  assign n31976 = pi0691 & ~n31971;
  assign n31977 = ~n31975 & n31976;
  assign n31978 = ~pi0192 & ~pi0691;
  assign n31979 = ~n17052 & n31978;
  assign n31980 = n2571 & ~n31979;
  assign n31981 = ~n31977 & n31980;
  assign n31982 = ~n31969 & ~n31981;
  assign n31983 = ~pi0778 & ~n31982;
  assign n31984 = ~pi0625 & n31967;
  assign n31985 = pi0625 & n31982;
  assign n31986 = pi1153 & ~n31984;
  assign n31987 = ~n31985 & n31986;
  assign n31988 = ~pi0625 & n31982;
  assign n31989 = pi0625 & n31967;
  assign n31990 = ~pi1153 & ~n31989;
  assign n31991 = ~n31988 & n31990;
  assign n31992 = ~n31987 & ~n31991;
  assign n31993 = pi0778 & ~n31992;
  assign n31994 = ~n31983 & ~n31993;
  assign n31995 = ~n17075 & ~n31994;
  assign n31996 = n17075 & ~n31967;
  assign n31997 = ~n31995 & ~n31996;
  assign n31998 = ~n16639 & n31997;
  assign n31999 = n16639 & n31967;
  assign n32000 = ~n31998 & ~n31999;
  assign n32001 = ~n16635 & n32000;
  assign n32002 = ~n31968 & ~n32001;
  assign n32003 = ~n16631 & n32002;
  assign n32004 = n16631 & n31967;
  assign n32005 = ~n32003 & ~n32004;
  assign n32006 = ~pi0628 & ~n32005;
  assign n32007 = pi0628 & n31967;
  assign n32008 = ~n32006 & ~n32007;
  assign n32009 = ~pi1156 & ~n32008;
  assign n32010 = pi0628 & ~n32005;
  assign n32011 = ~pi0628 & n31967;
  assign n32012 = ~n32010 & ~n32011;
  assign n32013 = pi1156 & ~n32012;
  assign n32014 = ~n32009 & ~n32013;
  assign n32015 = pi0792 & ~n32014;
  assign n32016 = ~pi0792 & ~n32005;
  assign n32017 = ~n32015 & ~n32016;
  assign n32018 = ~pi0647 & ~n32017;
  assign n32019 = pi0647 & n31967;
  assign n32020 = ~n32018 & ~n32019;
  assign n32021 = ~pi1157 & ~n32020;
  assign n32022 = pi0647 & ~n32017;
  assign n32023 = ~pi0647 & n31967;
  assign n32024 = ~n32022 & ~n32023;
  assign n32025 = pi1157 & ~n32024;
  assign n32026 = ~n32021 & ~n32025;
  assign n32027 = pi0787 & ~n32026;
  assign n32028 = ~pi0787 & ~n32017;
  assign n32029 = ~n32027 & ~n32028;
  assign n32030 = ~pi0644 & ~n32029;
  assign n32031 = pi0715 & ~n32030;
  assign n32032 = ~pi0764 & n17046;
  assign n32033 = pi0192 & n17273;
  assign n32034 = ~n32032 & ~n32033;
  assign n32035 = pi0039 & ~n32034;
  assign n32036 = pi0764 & ~n17234;
  assign n32037 = pi0192 & ~n32036;
  assign n32038 = ~pi0192 & pi0764;
  assign n32039 = n17221 & n32038;
  assign n32040 = ~n22600 & ~n32037;
  assign n32041 = ~n32039 & n32040;
  assign n32042 = ~n32035 & n32041;
  assign n32043 = ~pi0038 & ~n32042;
  assign n32044 = pi0764 & n17280;
  assign n32045 = pi0038 & ~n31970;
  assign n32046 = ~n32044 & n32045;
  assign n32047 = ~n32043 & ~n32046;
  assign n32048 = n2571 & ~n32047;
  assign n32049 = ~n31969 & ~n32048;
  assign n32050 = ~n17117 & ~n32049;
  assign n32051 = n17117 & ~n31967;
  assign n32052 = ~n32050 & ~n32051;
  assign n32053 = ~pi0785 & ~n32052;
  assign n32054 = ~n17291 & ~n31967;
  assign n32055 = pi0609 & n32050;
  assign n32056 = ~n32054 & ~n32055;
  assign n32057 = pi1155 & ~n32056;
  assign n32058 = ~n17296 & ~n31967;
  assign n32059 = ~pi0609 & n32050;
  assign n32060 = ~n32058 & ~n32059;
  assign n32061 = ~pi1155 & ~n32060;
  assign n32062 = ~n32057 & ~n32061;
  assign n32063 = pi0785 & ~n32062;
  assign n32064 = ~n32053 & ~n32063;
  assign n32065 = ~pi0781 & ~n32064;
  assign n32066 = ~pi0618 & n31967;
  assign n32067 = pi0618 & n32064;
  assign n32068 = pi1154 & ~n32066;
  assign n32069 = ~n32067 & n32068;
  assign n32070 = ~pi0618 & n32064;
  assign n32071 = pi0618 & n31967;
  assign n32072 = ~pi1154 & ~n32071;
  assign n32073 = ~n32070 & n32072;
  assign n32074 = ~n32069 & ~n32073;
  assign n32075 = pi0781 & ~n32074;
  assign n32076 = ~n32065 & ~n32075;
  assign n32077 = ~pi0789 & ~n32076;
  assign n32078 = ~pi0619 & n31967;
  assign n32079 = pi0619 & n32076;
  assign n32080 = pi1159 & ~n32078;
  assign n32081 = ~n32079 & n32080;
  assign n32082 = ~pi0619 & n32076;
  assign n32083 = pi0619 & n31967;
  assign n32084 = ~pi1159 & ~n32083;
  assign n32085 = ~n32082 & n32084;
  assign n32086 = ~n32081 & ~n32085;
  assign n32087 = pi0789 & ~n32086;
  assign n32088 = ~n32077 & ~n32087;
  assign n32089 = ~n17969 & n32088;
  assign n32090 = n17969 & n31967;
  assign n32091 = ~n32089 & ~n32090;
  assign n32092 = ~n17779 & ~n32091;
  assign n32093 = n17779 & n31967;
  assign n32094 = ~n32092 & ~n32093;
  assign n32095 = ~n17804 & ~n32094;
  assign n32096 = n17804 & n31967;
  assign n32097 = ~n32095 & ~n32096;
  assign n32098 = pi0644 & ~n32097;
  assign n32099 = ~pi0644 & n31967;
  assign n32100 = ~pi0715 & ~n32099;
  assign n32101 = ~n32098 & n32100;
  assign n32102 = pi1160 & ~n32101;
  assign n32103 = ~n32031 & n32102;
  assign n32104 = pi0644 & ~n32029;
  assign n32105 = ~pi0715 & ~n32104;
  assign n32106 = ~pi0644 & ~n32097;
  assign n32107 = pi0644 & n31967;
  assign n32108 = pi0715 & ~n32107;
  assign n32109 = ~n32106 & n32108;
  assign n32110 = ~pi1160 & ~n32109;
  assign n32111 = ~n32105 & n32110;
  assign n32112 = ~n32103 & ~n32111;
  assign n32113 = pi0790 & ~n32112;
  assign n32114 = n17777 & n32008;
  assign n32115 = ~n20570 & n32091;
  assign n32116 = n17776 & n32012;
  assign n32117 = ~n32114 & ~n32116;
  assign n32118 = ~n32115 & n32117;
  assign n32119 = pi0792 & ~n32118;
  assign n32120 = pi0609 & n31994;
  assign n32121 = ~pi0691 & n32047;
  assign n32122 = ~pi0764 & n24055;
  assign n32123 = ~n17490 & ~n32122;
  assign n32124 = ~pi0039 & ~n32123;
  assign n32125 = ~pi0192 & ~n32124;
  assign n32126 = ~n17469 & ~n31800;
  assign n32127 = pi0192 & ~n32126;
  assign n32128 = n6284 & n32127;
  assign n32129 = pi0038 & ~n32128;
  assign n32130 = ~n32125 & n32129;
  assign n32131 = ~pi0192 & ~n17629;
  assign n32132 = pi0192 & ~n17631;
  assign n32133 = pi0764 & ~n32132;
  assign n32134 = ~n32131 & n32133;
  assign n32135 = ~pi0192 & n17612;
  assign n32136 = pi0192 & n17625;
  assign n32137 = ~pi0764 & ~n32135;
  assign n32138 = ~n32136 & n32137;
  assign n32139 = ~pi0039 & ~n32134;
  assign n32140 = ~n32138 & n32139;
  assign n32141 = pi0192 & n17605;
  assign n32142 = ~pi0192 & ~n17546;
  assign n32143 = pi0764 & ~n32142;
  assign n32144 = ~n32141 & n32143;
  assign n32145 = ~pi0192 & n17404;
  assign n32146 = pi0192 & n17485;
  assign n32147 = ~pi0764 & ~n32146;
  assign n32148 = ~n32145 & n32147;
  assign n32149 = pi0039 & ~n32144;
  assign n32150 = ~n32148 & n32149;
  assign n32151 = ~pi0038 & ~n32140;
  assign n32152 = ~n32150 & n32151;
  assign n32153 = pi0691 & ~n32130;
  assign n32154 = ~n32152 & n32153;
  assign n32155 = n2571 & ~n32154;
  assign n32156 = ~n32121 & n32155;
  assign n32157 = ~n31969 & ~n32156;
  assign n32158 = ~pi0625 & n32157;
  assign n32159 = pi0625 & n32049;
  assign n32160 = ~pi1153 & ~n32159;
  assign n32161 = ~n32158 & n32160;
  assign n32162 = ~pi0608 & ~n31987;
  assign n32163 = ~n32161 & n32162;
  assign n32164 = ~pi0625 & n32049;
  assign n32165 = pi0625 & n32157;
  assign n32166 = pi1153 & ~n32164;
  assign n32167 = ~n32165 & n32166;
  assign n32168 = pi0608 & ~n31991;
  assign n32169 = ~n32167 & n32168;
  assign n32170 = ~n32163 & ~n32169;
  assign n32171 = pi0778 & ~n32170;
  assign n32172 = ~pi0778 & n32157;
  assign n32173 = ~n32171 & ~n32172;
  assign n32174 = ~pi0609 & ~n32173;
  assign n32175 = ~pi1155 & ~n32120;
  assign n32176 = ~n32174 & n32175;
  assign n32177 = ~pi0660 & ~n32057;
  assign n32178 = ~n32176 & n32177;
  assign n32179 = ~pi0609 & n31994;
  assign n32180 = pi0609 & ~n32173;
  assign n32181 = pi1155 & ~n32179;
  assign n32182 = ~n32180 & n32181;
  assign n32183 = pi0660 & ~n32061;
  assign n32184 = ~n32182 & n32183;
  assign n32185 = ~n32178 & ~n32184;
  assign n32186 = pi0785 & ~n32185;
  assign n32187 = ~pi0785 & ~n32173;
  assign n32188 = ~n32186 & ~n32187;
  assign n32189 = ~pi0618 & ~n32188;
  assign n32190 = pi0618 & n31997;
  assign n32191 = ~pi1154 & ~n32190;
  assign n32192 = ~n32189 & n32191;
  assign n32193 = ~pi0627 & ~n32069;
  assign n32194 = ~n32192 & n32193;
  assign n32195 = ~pi0618 & n31997;
  assign n32196 = pi0618 & ~n32188;
  assign n32197 = pi1154 & ~n32195;
  assign n32198 = ~n32196 & n32197;
  assign n32199 = pi0627 & ~n32073;
  assign n32200 = ~n32198 & n32199;
  assign n32201 = ~n32194 & ~n32200;
  assign n32202 = pi0781 & ~n32201;
  assign n32203 = ~pi0781 & ~n32188;
  assign n32204 = ~n32202 & ~n32203;
  assign n32205 = ~pi0789 & n32204;
  assign n32206 = pi0619 & ~n32000;
  assign n32207 = ~pi0619 & ~n32204;
  assign n32208 = ~pi1159 & ~n32206;
  assign n32209 = ~n32207 & n32208;
  assign n32210 = ~pi0648 & ~n32081;
  assign n32211 = ~n32209 & n32210;
  assign n32212 = ~pi0619 & ~n32000;
  assign n32213 = pi0619 & ~n32204;
  assign n32214 = pi1159 & ~n32212;
  assign n32215 = ~n32213 & n32214;
  assign n32216 = pi0648 & ~n32085;
  assign n32217 = ~n32215 & n32216;
  assign n32218 = pi0789 & ~n32211;
  assign n32219 = ~n32217 & n32218;
  assign n32220 = n17970 & ~n32205;
  assign n32221 = ~n32219 & n32220;
  assign n32222 = n17871 & n32002;
  assign n32223 = ~pi0626 & ~n32088;
  assign n32224 = pi0626 & ~n31967;
  assign n32225 = n16629 & ~n32224;
  assign n32226 = ~n32223 & n32225;
  assign n32227 = pi0626 & ~n32088;
  assign n32228 = ~pi0626 & ~n31967;
  assign n32229 = n16628 & ~n32228;
  assign n32230 = ~n32227 & n32229;
  assign n32231 = ~n32222 & ~n32226;
  assign n32232 = ~n32230 & n32231;
  assign n32233 = pi0788 & ~n32232;
  assign n32234 = ~n20364 & ~n32233;
  assign n32235 = ~n32221 & n32234;
  assign n32236 = ~n32119 & ~n32235;
  assign n32237 = ~n20206 & ~n32236;
  assign n32238 = n17802 & n32020;
  assign n32239 = ~n20559 & n32094;
  assign n32240 = n17801 & n32024;
  assign n32241 = ~n32238 & ~n32239;
  assign n32242 = ~n32240 & n32241;
  assign n32243 = pi0787 & ~n32242;
  assign n32244 = ~pi0644 & n32110;
  assign n32245 = pi0644 & n32102;
  assign n32246 = pi0790 & ~n32244;
  assign n32247 = ~n32245 & n32246;
  assign n32248 = ~n32237 & ~n32243;
  assign n32249 = ~n32247 & n32248;
  assign n32250 = ~n32113 & ~n32249;
  assign n32251 = ~po1038 & ~n32250;
  assign n32252 = ~pi0832 & ~n31966;
  assign n32253 = ~n32251 & n32252;
  assign po0349 = ~n31965 & ~n32253;
  assign n32255 = ~pi0193 & ~n2926;
  assign n32256 = pi0690 & n16645;
  assign n32257 = ~n32255 & ~n32256;
  assign n32258 = ~pi0778 & ~n32257;
  assign n32259 = ~pi0625 & n32256;
  assign n32260 = ~n32257 & ~n32259;
  assign n32261 = pi1153 & ~n32260;
  assign n32262 = ~pi1153 & ~n32255;
  assign n32263 = ~n32259 & n32262;
  assign n32264 = pi0778 & ~n32263;
  assign n32265 = ~n32261 & n32264;
  assign n32266 = ~n32258 & ~n32265;
  assign n32267 = ~n17845 & ~n32266;
  assign n32268 = ~n17847 & n32267;
  assign n32269 = ~n17849 & n32268;
  assign n32270 = ~n17851 & n32269;
  assign n32271 = ~n17857 & n32270;
  assign n32272 = ~pi0647 & n32271;
  assign n32273 = pi0647 & n32255;
  assign n32274 = ~pi1157 & ~n32273;
  assign n32275 = ~n32272 & n32274;
  assign n32276 = pi0630 & n32275;
  assign n32277 = pi0739 & n17244;
  assign n32278 = ~n32255 & ~n32277;
  assign n32279 = ~n17874 & ~n32278;
  assign n32280 = ~pi0785 & ~n32279;
  assign n32281 = n17296 & n32277;
  assign n32282 = n32279 & ~n32281;
  assign n32283 = pi1155 & ~n32282;
  assign n32284 = ~pi1155 & ~n32255;
  assign n32285 = ~n32281 & n32284;
  assign n32286 = ~n32283 & ~n32285;
  assign n32287 = pi0785 & ~n32286;
  assign n32288 = ~n32280 & ~n32287;
  assign n32289 = ~pi0781 & ~n32288;
  assign n32290 = ~n17889 & n32288;
  assign n32291 = pi1154 & ~n32290;
  assign n32292 = ~n17892 & n32288;
  assign n32293 = ~pi1154 & ~n32292;
  assign n32294 = ~n32291 & ~n32293;
  assign n32295 = pi0781 & ~n32294;
  assign n32296 = ~n32289 & ~n32295;
  assign n32297 = ~pi0789 & ~n32296;
  assign n32298 = ~n23078 & n32296;
  assign n32299 = pi1159 & ~n32298;
  assign n32300 = ~n23081 & n32296;
  assign n32301 = ~pi1159 & ~n32300;
  assign n32302 = ~n32299 & ~n32301;
  assign n32303 = pi0789 & ~n32302;
  assign n32304 = ~n32297 & ~n32303;
  assign n32305 = ~n17969 & n32304;
  assign n32306 = n17969 & n32255;
  assign n32307 = ~n32305 & ~n32306;
  assign n32308 = ~n17779 & ~n32307;
  assign n32309 = n17779 & n32255;
  assign n32310 = ~n32308 & ~n32309;
  assign n32311 = ~n20559 & n32310;
  assign n32312 = pi0647 & ~n32271;
  assign n32313 = ~pi0647 & ~n32255;
  assign n32314 = ~n32312 & ~n32313;
  assign n32315 = n17801 & ~n32314;
  assign n32316 = ~n32276 & ~n32315;
  assign n32317 = ~n32311 & n32316;
  assign n32318 = pi0787 & ~n32317;
  assign n32319 = n17871 & n32269;
  assign n32320 = ~pi0626 & ~n32304;
  assign n32321 = pi0626 & ~n32255;
  assign n32322 = n16629 & ~n32321;
  assign n32323 = ~n32320 & n32322;
  assign n32324 = pi0626 & ~n32304;
  assign n32325 = ~pi0626 & ~n32255;
  assign n32326 = n16628 & ~n32325;
  assign n32327 = ~n32324 & n32326;
  assign n32328 = ~n32319 & ~n32323;
  assign n32329 = ~n32327 & n32328;
  assign n32330 = pi0788 & ~n32329;
  assign n32331 = pi0618 & n32267;
  assign n32332 = ~n17168 & ~n32257;
  assign n32333 = pi0625 & n32332;
  assign n32334 = n32278 & ~n32332;
  assign n32335 = ~n32333 & ~n32334;
  assign n32336 = n32262 & ~n32335;
  assign n32337 = ~pi0608 & ~n32261;
  assign n32338 = ~n32336 & n32337;
  assign n32339 = pi1153 & n32278;
  assign n32340 = ~n32333 & n32339;
  assign n32341 = pi0608 & ~n32263;
  assign n32342 = ~n32340 & n32341;
  assign n32343 = ~n32338 & ~n32342;
  assign n32344 = pi0778 & ~n32343;
  assign n32345 = ~pi0778 & ~n32334;
  assign n32346 = ~n32344 & ~n32345;
  assign n32347 = ~pi0609 & ~n32346;
  assign n32348 = pi0609 & ~n32266;
  assign n32349 = ~pi1155 & ~n32348;
  assign n32350 = ~n32347 & n32349;
  assign n32351 = ~pi0660 & ~n32283;
  assign n32352 = ~n32350 & n32351;
  assign n32353 = pi0609 & ~n32346;
  assign n32354 = ~pi0609 & ~n32266;
  assign n32355 = pi1155 & ~n32354;
  assign n32356 = ~n32353 & n32355;
  assign n32357 = pi0660 & ~n32285;
  assign n32358 = ~n32356 & n32357;
  assign n32359 = ~n32352 & ~n32358;
  assign n32360 = pi0785 & ~n32359;
  assign n32361 = ~pi0785 & ~n32346;
  assign n32362 = ~n32360 & ~n32361;
  assign n32363 = ~pi0618 & ~n32362;
  assign n32364 = ~pi1154 & ~n32331;
  assign n32365 = ~n32363 & n32364;
  assign n32366 = ~pi0627 & ~n32291;
  assign n32367 = ~n32365 & n32366;
  assign n32368 = ~pi0618 & n32267;
  assign n32369 = pi0618 & ~n32362;
  assign n32370 = pi1154 & ~n32368;
  assign n32371 = ~n32369 & n32370;
  assign n32372 = pi0627 & ~n32293;
  assign n32373 = ~n32371 & n32372;
  assign n32374 = ~n32367 & ~n32373;
  assign n32375 = pi0781 & ~n32374;
  assign n32376 = ~pi0781 & ~n32362;
  assign n32377 = ~n32375 & ~n32376;
  assign n32378 = ~pi0789 & n32377;
  assign n32379 = ~pi0619 & ~n32377;
  assign n32380 = pi0619 & n32268;
  assign n32381 = ~pi1159 & ~n32380;
  assign n32382 = ~n32379 & n32381;
  assign n32383 = ~pi0648 & ~n32299;
  assign n32384 = ~n32382 & n32383;
  assign n32385 = pi0619 & ~n32377;
  assign n32386 = ~pi0619 & n32268;
  assign n32387 = pi1159 & ~n32386;
  assign n32388 = ~n32385 & n32387;
  assign n32389 = pi0648 & ~n32301;
  assign n32390 = ~n32388 & n32389;
  assign n32391 = pi0789 & ~n32384;
  assign n32392 = ~n32390 & n32391;
  assign n32393 = n17970 & ~n32378;
  assign n32394 = ~n32392 & n32393;
  assign n32395 = ~n32330 & ~n32394;
  assign n32396 = ~n20364 & ~n32395;
  assign n32397 = n17854 & ~n32307;
  assign n32398 = n20851 & n32270;
  assign n32399 = ~n32397 & ~n32398;
  assign n32400 = ~pi0629 & ~n32399;
  assign n32401 = n20855 & n32270;
  assign n32402 = n17853 & ~n32307;
  assign n32403 = ~n32401 & ~n32402;
  assign n32404 = pi0629 & ~n32403;
  assign n32405 = ~n32400 & ~n32404;
  assign n32406 = pi0792 & ~n32405;
  assign n32407 = ~n20206 & ~n32406;
  assign n32408 = ~n32396 & n32407;
  assign n32409 = ~n32318 & ~n32408;
  assign n32410 = ~pi0790 & n32409;
  assign n32411 = ~pi0787 & ~n32271;
  assign n32412 = pi1157 & ~n32314;
  assign n32413 = ~n32275 & ~n32412;
  assign n32414 = pi0787 & ~n32413;
  assign n32415 = ~n32411 & ~n32414;
  assign n32416 = ~pi0644 & n32415;
  assign n32417 = pi0644 & n32409;
  assign n32418 = pi0715 & ~n32416;
  assign n32419 = ~n32417 & n32418;
  assign n32420 = ~n17804 & ~n32310;
  assign n32421 = n17804 & n32255;
  assign n32422 = ~n32420 & ~n32421;
  assign n32423 = pi0644 & ~n32422;
  assign n32424 = ~pi0644 & n32255;
  assign n32425 = ~pi0715 & ~n32424;
  assign n32426 = ~n32423 & n32425;
  assign n32427 = pi1160 & ~n32426;
  assign n32428 = ~n32419 & n32427;
  assign n32429 = ~pi0644 & ~n32422;
  assign n32430 = pi0644 & n32255;
  assign n32431 = pi0715 & ~n32430;
  assign n32432 = ~n32429 & n32431;
  assign n32433 = pi0644 & n32415;
  assign n32434 = ~pi0644 & n32409;
  assign n32435 = ~pi0715 & ~n32433;
  assign n32436 = ~n32434 & n32435;
  assign n32437 = ~pi1160 & ~n32432;
  assign n32438 = ~n32436 & n32437;
  assign n32439 = ~n32428 & ~n32438;
  assign n32440 = pi0790 & ~n32439;
  assign n32441 = pi0832 & ~n32410;
  assign n32442 = ~n32440 & n32441;
  assign n32443 = ~pi0193 & po1038;
  assign n32444 = ~pi0193 & ~n17059;
  assign n32445 = n16635 & ~n32444;
  assign n32446 = pi0690 & n2571;
  assign n32447 = n32444 & ~n32446;
  assign n32448 = ~pi0193 & ~n16641;
  assign n32449 = n16647 & ~n32448;
  assign n32450 = pi0193 & ~n18076;
  assign n32451 = ~pi0038 & ~n32450;
  assign n32452 = n2571 & ~n32451;
  assign n32453 = ~pi0193 & n18072;
  assign n32454 = ~n32452 & ~n32453;
  assign n32455 = pi0690 & ~n32449;
  assign n32456 = ~n32454 & n32455;
  assign n32457 = ~n32447 & ~n32456;
  assign n32458 = ~pi0778 & n32457;
  assign n32459 = ~pi0625 & n32444;
  assign n32460 = pi0625 & ~n32457;
  assign n32461 = pi1153 & ~n32459;
  assign n32462 = ~n32460 & n32461;
  assign n32463 = pi0625 & n32444;
  assign n32464 = ~pi0625 & ~n32457;
  assign n32465 = ~pi1153 & ~n32463;
  assign n32466 = ~n32464 & n32465;
  assign n32467 = ~n32462 & ~n32466;
  assign n32468 = pi0778 & ~n32467;
  assign n32469 = ~n32458 & ~n32468;
  assign n32470 = ~n17075 & ~n32469;
  assign n32471 = n17075 & ~n32444;
  assign n32472 = ~n32470 & ~n32471;
  assign n32473 = ~n16639 & n32472;
  assign n32474 = n16639 & n32444;
  assign n32475 = ~n32473 & ~n32474;
  assign n32476 = ~n16635 & n32475;
  assign n32477 = ~n32445 & ~n32476;
  assign n32478 = ~n16631 & n32477;
  assign n32479 = n16631 & n32444;
  assign n32480 = ~n32478 & ~n32479;
  assign n32481 = ~pi0792 & n32480;
  assign n32482 = pi0628 & ~n32480;
  assign n32483 = ~pi0628 & n32444;
  assign n32484 = pi1156 & ~n32483;
  assign n32485 = ~n32482 & n32484;
  assign n32486 = pi0628 & n32444;
  assign n32487 = ~pi0628 & ~n32480;
  assign n32488 = ~pi1156 & ~n32486;
  assign n32489 = ~n32487 & n32488;
  assign n32490 = ~n32485 & ~n32489;
  assign n32491 = pi0792 & ~n32490;
  assign n32492 = ~n32481 & ~n32491;
  assign n32493 = ~pi0647 & ~n32492;
  assign n32494 = pi0647 & ~n32444;
  assign n32495 = ~n32493 & ~n32494;
  assign n32496 = ~pi1157 & n32495;
  assign n32497 = pi0647 & ~n32492;
  assign n32498 = ~pi0647 & ~n32444;
  assign n32499 = ~n32497 & ~n32498;
  assign n32500 = pi1157 & n32499;
  assign n32501 = ~n32496 & ~n32500;
  assign n32502 = pi0787 & ~n32501;
  assign n32503 = ~pi0787 & n32492;
  assign n32504 = ~n32502 & ~n32503;
  assign n32505 = ~pi0644 & ~n32504;
  assign n32506 = pi0715 & ~n32505;
  assign n32507 = pi0193 & ~n2571;
  assign n32508 = pi0739 & n17280;
  assign n32509 = ~n32448 & ~n32508;
  assign n32510 = pi0038 & ~n32509;
  assign n32511 = ~pi0193 & n17221;
  assign n32512 = pi0193 & ~n17275;
  assign n32513 = pi0739 & ~n32512;
  assign n32514 = ~n32511 & n32513;
  assign n32515 = ~pi0193 & ~pi0739;
  assign n32516 = ~n17048 & n32515;
  assign n32517 = ~n32514 & ~n32516;
  assign n32518 = ~pi0038 & ~n32517;
  assign n32519 = ~n32510 & ~n32518;
  assign n32520 = n2571 & n32519;
  assign n32521 = ~n32507 & ~n32520;
  assign n32522 = ~n17117 & ~n32521;
  assign n32523 = n17117 & ~n32444;
  assign n32524 = ~n32522 & ~n32523;
  assign n32525 = ~pi0785 & ~n32524;
  assign n32526 = ~n17291 & ~n32444;
  assign n32527 = pi0609 & n32522;
  assign n32528 = ~n32526 & ~n32527;
  assign n32529 = pi1155 & ~n32528;
  assign n32530 = ~n17296 & ~n32444;
  assign n32531 = ~pi0609 & n32522;
  assign n32532 = ~n32530 & ~n32531;
  assign n32533 = ~pi1155 & ~n32532;
  assign n32534 = ~n32529 & ~n32533;
  assign n32535 = pi0785 & ~n32534;
  assign n32536 = ~n32525 & ~n32535;
  assign n32537 = ~pi0781 & ~n32536;
  assign n32538 = ~pi0618 & n32444;
  assign n32539 = pi0618 & n32536;
  assign n32540 = pi1154 & ~n32538;
  assign n32541 = ~n32539 & n32540;
  assign n32542 = ~pi0618 & n32536;
  assign n32543 = pi0618 & n32444;
  assign n32544 = ~pi1154 & ~n32543;
  assign n32545 = ~n32542 & n32544;
  assign n32546 = ~n32541 & ~n32545;
  assign n32547 = pi0781 & ~n32546;
  assign n32548 = ~n32537 & ~n32547;
  assign n32549 = ~pi0789 & ~n32548;
  assign n32550 = ~pi0619 & n32444;
  assign n32551 = pi0619 & n32548;
  assign n32552 = pi1159 & ~n32550;
  assign n32553 = ~n32551 & n32552;
  assign n32554 = ~pi0619 & n32548;
  assign n32555 = pi0619 & n32444;
  assign n32556 = ~pi1159 & ~n32555;
  assign n32557 = ~n32554 & n32556;
  assign n32558 = ~n32553 & ~n32557;
  assign n32559 = pi0789 & ~n32558;
  assign n32560 = ~n32549 & ~n32559;
  assign n32561 = ~n17969 & n32560;
  assign n32562 = n17969 & n32444;
  assign n32563 = ~n32561 & ~n32562;
  assign n32564 = ~n17779 & ~n32563;
  assign n32565 = n17779 & n32444;
  assign n32566 = ~n32564 & ~n32565;
  assign n32567 = ~n17804 & ~n32566;
  assign n32568 = n17804 & n32444;
  assign n32569 = ~n32567 & ~n32568;
  assign n32570 = pi0644 & ~n32569;
  assign n32571 = ~pi0644 & n32444;
  assign n32572 = ~pi0715 & ~n32571;
  assign n32573 = ~n32570 & n32572;
  assign n32574 = pi1160 & ~n32573;
  assign n32575 = ~n32506 & n32574;
  assign n32576 = pi0644 & ~n32504;
  assign n32577 = ~pi0715 & ~n32576;
  assign n32578 = ~pi0644 & ~n32569;
  assign n32579 = pi0644 & n32444;
  assign n32580 = pi0715 & ~n32579;
  assign n32581 = ~n32578 & n32580;
  assign n32582 = ~pi1160 & ~n32581;
  assign n32583 = ~n32577 & n32582;
  assign n32584 = ~n32575 & ~n32583;
  assign n32585 = pi0790 & ~n32584;
  assign n32586 = ~pi0629 & n32485;
  assign n32587 = ~n20570 & n32563;
  assign n32588 = pi0629 & n32489;
  assign n32589 = ~n32586 & ~n32588;
  assign n32590 = ~n32587 & n32589;
  assign n32591 = pi0792 & ~n32590;
  assign n32592 = pi0609 & n32469;
  assign n32593 = ~pi0690 & ~n32519;
  assign n32594 = ~pi0193 & n17629;
  assign n32595 = pi0193 & n17631;
  assign n32596 = pi0739 & ~n32595;
  assign n32597 = ~n32594 & n32596;
  assign n32598 = pi0193 & ~n17625;
  assign n32599 = ~pi0193 & ~n17612;
  assign n32600 = ~pi0739 & ~n32598;
  assign n32601 = ~n32599 & n32600;
  assign n32602 = ~n32597 & ~n32601;
  assign n32603 = ~pi0039 & ~n32602;
  assign n32604 = pi0193 & n17605;
  assign n32605 = ~pi0193 & ~n17546;
  assign n32606 = pi0739 & ~n32605;
  assign n32607 = ~n32604 & n32606;
  assign n32608 = ~pi0193 & n17404;
  assign n32609 = pi0193 & n17485;
  assign n32610 = ~pi0739 & ~n32609;
  assign n32611 = ~n32608 & n32610;
  assign n32612 = pi0039 & ~n32607;
  assign n32613 = ~n32611 & n32612;
  assign n32614 = ~pi0038 & ~n32603;
  assign n32615 = ~n32613 & n32614;
  assign n32616 = ~pi0739 & n24055;
  assign n32617 = ~n17490 & ~n32616;
  assign n32618 = ~pi0039 & ~n32617;
  assign n32619 = ~pi0193 & ~n32618;
  assign n32620 = ~n17469 & ~n32277;
  assign n32621 = pi0193 & ~n32620;
  assign n32622 = n6284 & n32621;
  assign n32623 = pi0038 & ~n32622;
  assign n32624 = ~n32619 & n32623;
  assign n32625 = pi0690 & ~n32624;
  assign n32626 = ~n32615 & n32625;
  assign n32627 = n2571 & ~n32626;
  assign n32628 = ~n32593 & n32627;
  assign n32629 = ~n32507 & ~n32628;
  assign n32630 = ~pi0625 & n32629;
  assign n32631 = pi0625 & n32521;
  assign n32632 = ~pi1153 & ~n32631;
  assign n32633 = ~n32630 & n32632;
  assign n32634 = ~pi0608 & ~n32462;
  assign n32635 = ~n32633 & n32634;
  assign n32636 = ~pi0625 & n32521;
  assign n32637 = pi0625 & n32629;
  assign n32638 = pi1153 & ~n32636;
  assign n32639 = ~n32637 & n32638;
  assign n32640 = pi0608 & ~n32466;
  assign n32641 = ~n32639 & n32640;
  assign n32642 = ~n32635 & ~n32641;
  assign n32643 = pi0778 & ~n32642;
  assign n32644 = ~pi0778 & n32629;
  assign n32645 = ~n32643 & ~n32644;
  assign n32646 = ~pi0609 & ~n32645;
  assign n32647 = ~pi1155 & ~n32592;
  assign n32648 = ~n32646 & n32647;
  assign n32649 = ~pi0660 & ~n32529;
  assign n32650 = ~n32648 & n32649;
  assign n32651 = ~pi0609 & n32469;
  assign n32652 = pi0609 & ~n32645;
  assign n32653 = pi1155 & ~n32651;
  assign n32654 = ~n32652 & n32653;
  assign n32655 = pi0660 & ~n32533;
  assign n32656 = ~n32654 & n32655;
  assign n32657 = ~n32650 & ~n32656;
  assign n32658 = pi0785 & ~n32657;
  assign n32659 = ~pi0785 & ~n32645;
  assign n32660 = ~n32658 & ~n32659;
  assign n32661 = ~pi0618 & ~n32660;
  assign n32662 = pi0618 & n32472;
  assign n32663 = ~pi1154 & ~n32662;
  assign n32664 = ~n32661 & n32663;
  assign n32665 = ~pi0627 & ~n32541;
  assign n32666 = ~n32664 & n32665;
  assign n32667 = ~pi0618 & n32472;
  assign n32668 = pi0618 & ~n32660;
  assign n32669 = pi1154 & ~n32667;
  assign n32670 = ~n32668 & n32669;
  assign n32671 = pi0627 & ~n32545;
  assign n32672 = ~n32670 & n32671;
  assign n32673 = ~n32666 & ~n32672;
  assign n32674 = pi0781 & ~n32673;
  assign n32675 = ~pi0781 & ~n32660;
  assign n32676 = ~n32674 & ~n32675;
  assign n32677 = ~pi0789 & n32676;
  assign n32678 = pi0619 & ~n32475;
  assign n32679 = ~pi0619 & ~n32676;
  assign n32680 = ~pi1159 & ~n32678;
  assign n32681 = ~n32679 & n32680;
  assign n32682 = ~pi0648 & ~n32553;
  assign n32683 = ~n32681 & n32682;
  assign n32684 = ~pi0619 & ~n32475;
  assign n32685 = pi0619 & ~n32676;
  assign n32686 = pi1159 & ~n32684;
  assign n32687 = ~n32685 & n32686;
  assign n32688 = pi0648 & ~n32557;
  assign n32689 = ~n32687 & n32688;
  assign n32690 = pi0789 & ~n32683;
  assign n32691 = ~n32689 & n32690;
  assign n32692 = n17970 & ~n32677;
  assign n32693 = ~n32691 & n32692;
  assign n32694 = n17871 & n32477;
  assign n32695 = ~pi0626 & ~n32560;
  assign n32696 = pi0626 & ~n32444;
  assign n32697 = n16629 & ~n32696;
  assign n32698 = ~n32695 & n32697;
  assign n32699 = pi0626 & ~n32560;
  assign n32700 = ~pi0626 & ~n32444;
  assign n32701 = n16628 & ~n32700;
  assign n32702 = ~n32699 & n32701;
  assign n32703 = ~n32694 & ~n32698;
  assign n32704 = ~n32702 & n32703;
  assign n32705 = pi0788 & ~n32704;
  assign n32706 = ~n20364 & ~n32705;
  assign n32707 = ~n32693 & n32706;
  assign n32708 = ~n32591 & ~n32707;
  assign n32709 = ~n20206 & ~n32708;
  assign n32710 = n17802 & ~n32495;
  assign n32711 = ~n20559 & n32566;
  assign n32712 = n17801 & ~n32499;
  assign n32713 = ~n32710 & ~n32712;
  assign n32714 = ~n32711 & n32713;
  assign n32715 = pi0787 & ~n32714;
  assign n32716 = ~pi0644 & n32582;
  assign n32717 = pi0644 & n32574;
  assign n32718 = pi0790 & ~n32716;
  assign n32719 = ~n32717 & n32718;
  assign n32720 = ~n32709 & ~n32715;
  assign n32721 = ~n32719 & n32720;
  assign n32722 = ~n32585 & ~n32721;
  assign n32723 = ~po1038 & ~n32722;
  assign n32724 = ~pi0832 & ~n32443;
  assign n32725 = ~n32723 & n32724;
  assign po0350 = ~n32442 & ~n32725;
  assign n32727 = ~pi0194 & ~n17059;
  assign n32728 = n16635 & ~n32727;
  assign n32729 = pi0194 & ~n24385;
  assign n32730 = ~pi0194 & n24388;
  assign n32731 = pi0730 & ~n32730;
  assign n32732 = ~pi0194 & ~n17052;
  assign n32733 = ~pi0730 & n32732;
  assign n32734 = n2571 & ~n32733;
  assign n32735 = ~n32731 & n32734;
  assign n32736 = ~n32729 & ~n32735;
  assign n32737 = ~pi0778 & ~n32736;
  assign n32738 = ~pi0625 & n32727;
  assign n32739 = pi0625 & n32736;
  assign n32740 = pi1153 & ~n32738;
  assign n32741 = ~n32739 & n32740;
  assign n32742 = ~pi0625 & n32736;
  assign n32743 = pi0625 & n32727;
  assign n32744 = ~pi1153 & ~n32743;
  assign n32745 = ~n32742 & n32744;
  assign n32746 = ~n32741 & ~n32745;
  assign n32747 = pi0778 & ~n32746;
  assign n32748 = ~n32737 & ~n32747;
  assign n32749 = ~n17075 & ~n32748;
  assign n32750 = n17075 & ~n32727;
  assign n32751 = ~n32749 & ~n32750;
  assign n32752 = ~n16639 & n32751;
  assign n32753 = n16639 & n32727;
  assign n32754 = ~n32752 & ~n32753;
  assign n32755 = ~n16635 & n32754;
  assign n32756 = ~n32728 & ~n32755;
  assign n32757 = ~n16631 & n32756;
  assign n32758 = n16631 & n32727;
  assign n32759 = ~n32757 & ~n32758;
  assign n32760 = ~pi0792 & n32759;
  assign n32761 = ~pi0628 & n32727;
  assign n32762 = pi0628 & ~n32759;
  assign n32763 = pi1156 & ~n32761;
  assign n32764 = ~n32762 & n32763;
  assign n32765 = pi0628 & n32727;
  assign n32766 = ~pi0628 & ~n32759;
  assign n32767 = ~pi1156 & ~n32765;
  assign n32768 = ~n32766 & n32767;
  assign n32769 = ~n32764 & ~n32768;
  assign n32770 = pi0792 & ~n32769;
  assign n32771 = ~n32760 & ~n32770;
  assign n32772 = ~pi0787 & ~n32771;
  assign n32773 = ~pi0647 & n32727;
  assign n32774 = pi0647 & n32771;
  assign n32775 = pi1157 & ~n32773;
  assign n32776 = ~n32774 & n32775;
  assign n32777 = ~pi0647 & n32771;
  assign n32778 = pi0647 & n32727;
  assign n32779 = ~pi1157 & ~n32778;
  assign n32780 = ~n32777 & n32779;
  assign n32781 = ~n32776 & ~n32780;
  assign n32782 = pi0787 & ~n32781;
  assign n32783 = ~n32772 & ~n32782;
  assign n32784 = ~pi0644 & n32783;
  assign n32785 = ~pi0618 & n32727;
  assign n32786 = pi0194 & ~n2571;
  assign n32787 = ~pi0194 & n19439;
  assign n32788 = pi0194 & n24447;
  assign n32789 = ~n32787 & ~n32788;
  assign n32790 = pi0748 & ~n32789;
  assign n32791 = ~pi0748 & ~n32732;
  assign n32792 = ~n32790 & ~n32791;
  assign n32793 = n2571 & ~n32792;
  assign n32794 = ~n32786 & ~n32793;
  assign n32795 = ~n17117 & ~n32794;
  assign n32796 = n17117 & ~n32727;
  assign n32797 = ~n32795 & ~n32796;
  assign n32798 = ~pi0785 & ~n32797;
  assign n32799 = ~n17291 & ~n32727;
  assign n32800 = pi0609 & n32795;
  assign n32801 = ~n32799 & ~n32800;
  assign n32802 = pi1155 & ~n32801;
  assign n32803 = ~n17296 & ~n32727;
  assign n32804 = ~pi0609 & n32795;
  assign n32805 = ~n32803 & ~n32804;
  assign n32806 = ~pi1155 & ~n32805;
  assign n32807 = ~n32802 & ~n32806;
  assign n32808 = pi0785 & ~n32807;
  assign n32809 = ~n32798 & ~n32808;
  assign n32810 = pi0618 & n32809;
  assign n32811 = pi1154 & ~n32785;
  assign n32812 = ~n32810 & n32811;
  assign n32813 = ~pi0730 & n32792;
  assign n32814 = pi0194 & n19496;
  assign n32815 = ~pi0194 & ~n19488;
  assign n32816 = pi0748 & ~n32815;
  assign n32817 = ~n32814 & n32816;
  assign n32818 = pi0194 & ~n24549;
  assign n32819 = ~pi0194 & n19477;
  assign n32820 = ~pi0748 & ~n32818;
  assign n32821 = ~n32819 & n32820;
  assign n32822 = pi0730 & ~n32817;
  assign n32823 = ~n32821 & n32822;
  assign n32824 = n2571 & ~n32813;
  assign n32825 = ~n32823 & n32824;
  assign n32826 = ~n32786 & ~n32825;
  assign n32827 = ~pi0625 & n32826;
  assign n32828 = pi0625 & n32794;
  assign n32829 = ~pi1153 & ~n32828;
  assign n32830 = ~n32827 & n32829;
  assign n32831 = ~pi0608 & ~n32741;
  assign n32832 = ~n32830 & n32831;
  assign n32833 = ~pi0625 & n32794;
  assign n32834 = pi0625 & n32826;
  assign n32835 = pi1153 & ~n32833;
  assign n32836 = ~n32834 & n32835;
  assign n32837 = pi0608 & ~n32745;
  assign n32838 = ~n32836 & n32837;
  assign n32839 = ~n32832 & ~n32838;
  assign n32840 = pi0778 & ~n32839;
  assign n32841 = ~pi0778 & n32826;
  assign n32842 = ~n32840 & ~n32841;
  assign n32843 = ~pi0609 & ~n32842;
  assign n32844 = pi0609 & n32748;
  assign n32845 = ~pi1155 & ~n32844;
  assign n32846 = ~n32843 & n32845;
  assign n32847 = ~pi0660 & ~n32802;
  assign n32848 = ~n32846 & n32847;
  assign n32849 = ~pi0609 & n32748;
  assign n32850 = pi0609 & ~n32842;
  assign n32851 = pi1155 & ~n32849;
  assign n32852 = ~n32850 & n32851;
  assign n32853 = pi0660 & ~n32806;
  assign n32854 = ~n32852 & n32853;
  assign n32855 = ~n32848 & ~n32854;
  assign n32856 = pi0785 & ~n32855;
  assign n32857 = ~pi0785 & ~n32842;
  assign n32858 = ~n32856 & ~n32857;
  assign n32859 = ~pi0618 & ~n32858;
  assign n32860 = pi0618 & n32751;
  assign n32861 = ~pi1154 & ~n32860;
  assign n32862 = ~n32859 & n32861;
  assign n32863 = ~pi0627 & ~n32812;
  assign n32864 = ~n32862 & n32863;
  assign n32865 = ~pi0618 & n32809;
  assign n32866 = pi0618 & n32727;
  assign n32867 = ~pi1154 & ~n32866;
  assign n32868 = ~n32865 & n32867;
  assign n32869 = ~pi0618 & n32751;
  assign n32870 = pi0618 & ~n32858;
  assign n32871 = pi1154 & ~n32869;
  assign n32872 = ~n32870 & n32871;
  assign n32873 = pi0627 & ~n32868;
  assign n32874 = ~n32872 & n32873;
  assign n32875 = ~n32864 & ~n32874;
  assign n32876 = pi0781 & ~n32875;
  assign n32877 = ~pi0781 & ~n32858;
  assign n32878 = ~n32876 & ~n32877;
  assign n32879 = ~pi0619 & ~n32878;
  assign n32880 = pi0619 & ~n32754;
  assign n32881 = ~pi1159 & ~n32880;
  assign n32882 = ~n32879 & n32881;
  assign n32883 = ~pi0619 & n32727;
  assign n32884 = ~pi0781 & ~n32809;
  assign n32885 = ~n32812 & ~n32868;
  assign n32886 = pi0781 & ~n32885;
  assign n32887 = ~n32884 & ~n32886;
  assign n32888 = pi0619 & n32887;
  assign n32889 = pi1159 & ~n32883;
  assign n32890 = ~n32888 & n32889;
  assign n32891 = ~pi0648 & ~n32890;
  assign n32892 = ~n32882 & n32891;
  assign n32893 = pi0619 & ~n32878;
  assign n32894 = ~pi0619 & ~n32754;
  assign n32895 = pi1159 & ~n32894;
  assign n32896 = ~n32893 & n32895;
  assign n32897 = ~pi0619 & n32887;
  assign n32898 = pi0619 & n32727;
  assign n32899 = ~pi1159 & ~n32898;
  assign n32900 = ~n32897 & n32899;
  assign n32901 = pi0648 & ~n32900;
  assign n32902 = ~n32896 & n32901;
  assign n32903 = ~n32892 & ~n32902;
  assign n32904 = pi0789 & ~n32903;
  assign n32905 = ~pi0789 & ~n32878;
  assign n32906 = ~n32904 & ~n32905;
  assign n32907 = ~pi0788 & n32906;
  assign n32908 = ~pi0626 & n32906;
  assign n32909 = pi0626 & ~n32756;
  assign n32910 = ~pi0641 & ~n32909;
  assign n32911 = ~n32908 & n32910;
  assign n32912 = ~pi0789 & ~n32887;
  assign n32913 = ~n32890 & ~n32900;
  assign n32914 = pi0789 & ~n32913;
  assign n32915 = ~n32912 & ~n32914;
  assign n32916 = ~pi0626 & ~n32915;
  assign n32917 = pi0626 & ~n32727;
  assign n32918 = pi0641 & ~n32917;
  assign n32919 = ~n32916 & n32918;
  assign n32920 = ~pi1158 & ~n32919;
  assign n32921 = ~n32911 & n32920;
  assign n32922 = pi0626 & n32906;
  assign n32923 = ~pi0626 & ~n32756;
  assign n32924 = pi0641 & ~n32923;
  assign n32925 = ~n32922 & n32924;
  assign n32926 = pi0626 & ~n32915;
  assign n32927 = ~pi0626 & ~n32727;
  assign n32928 = ~pi0641 & ~n32927;
  assign n32929 = ~n32926 & n32928;
  assign n32930 = pi1158 & ~n32929;
  assign n32931 = ~n32925 & n32930;
  assign n32932 = ~n32921 & ~n32931;
  assign n32933 = pi0788 & ~n32932;
  assign n32934 = ~n32907 & ~n32933;
  assign n32935 = ~pi0628 & n32934;
  assign n32936 = ~n17969 & n32915;
  assign n32937 = n17969 & n32727;
  assign n32938 = ~n32936 & ~n32937;
  assign n32939 = pi0628 & ~n32938;
  assign n32940 = ~pi1156 & ~n32939;
  assign n32941 = ~n32935 & n32940;
  assign n32942 = ~pi0629 & ~n32764;
  assign n32943 = ~n32941 & n32942;
  assign n32944 = pi0628 & n32934;
  assign n32945 = ~pi0628 & ~n32938;
  assign n32946 = pi1156 & ~n32945;
  assign n32947 = ~n32944 & n32946;
  assign n32948 = pi0629 & ~n32768;
  assign n32949 = ~n32947 & n32948;
  assign n32950 = ~n32943 & ~n32949;
  assign n32951 = pi0792 & ~n32950;
  assign n32952 = ~pi0792 & n32934;
  assign n32953 = ~n32951 & ~n32952;
  assign n32954 = ~pi0647 & ~n32953;
  assign n32955 = ~n17779 & ~n32938;
  assign n32956 = n17779 & n32727;
  assign n32957 = ~n32955 & ~n32956;
  assign n32958 = pi0647 & ~n32957;
  assign n32959 = ~pi1157 & ~n32958;
  assign n32960 = ~n32954 & n32959;
  assign n32961 = ~pi0630 & ~n32776;
  assign n32962 = ~n32960 & n32961;
  assign n32963 = pi0647 & ~n32953;
  assign n32964 = ~pi0647 & ~n32957;
  assign n32965 = pi1157 & ~n32964;
  assign n32966 = ~n32963 & n32965;
  assign n32967 = pi0630 & ~n32780;
  assign n32968 = ~n32966 & n32967;
  assign n32969 = ~n32962 & ~n32968;
  assign n32970 = pi0787 & ~n32969;
  assign n32971 = ~pi0787 & ~n32953;
  assign n32972 = ~n32970 & ~n32971;
  assign n32973 = pi0644 & ~n32972;
  assign n32974 = pi0715 & ~n32784;
  assign n32975 = ~n32973 & n32974;
  assign n32976 = n17804 & ~n32727;
  assign n32977 = ~n17804 & n32957;
  assign n32978 = ~n32976 & ~n32977;
  assign n32979 = pi0644 & n32978;
  assign n32980 = ~pi0644 & n32727;
  assign n32981 = ~pi0715 & ~n32980;
  assign n32982 = ~n32979 & n32981;
  assign n32983 = pi1160 & ~n32982;
  assign n32984 = ~n32975 & n32983;
  assign n32985 = ~pi0644 & ~n32972;
  assign n32986 = pi0644 & n32783;
  assign n32987 = ~pi0715 & ~n32986;
  assign n32988 = ~n32985 & n32987;
  assign n32989 = ~pi0644 & n32978;
  assign n32990 = pi0644 & n32727;
  assign n32991 = pi0715 & ~n32990;
  assign n32992 = ~n32989 & n32991;
  assign n32993 = ~pi1160 & ~n32992;
  assign n32994 = ~n32988 & n32993;
  assign n32995 = pi0790 & ~n32984;
  assign n32996 = ~n32994 & n32995;
  assign n32997 = ~pi0790 & n32972;
  assign n32998 = ~po1038 & ~n32997;
  assign n32999 = ~n32996 & n32998;
  assign n33000 = ~pi0194 & po1038;
  assign n33001 = ~pi0832 & ~n33000;
  assign n33002 = ~n32999 & n33001;
  assign n33003 = ~pi0194 & ~n2926;
  assign n33004 = pi0730 & n16645;
  assign n33005 = ~n33003 & ~n33004;
  assign n33006 = ~pi0778 & n33005;
  assign n33007 = ~pi0625 & n33004;
  assign n33008 = ~n33005 & ~n33007;
  assign n33009 = pi1153 & ~n33008;
  assign n33010 = ~pi1153 & ~n33003;
  assign n33011 = ~n33007 & n33010;
  assign n33012 = ~n33009 & ~n33011;
  assign n33013 = pi0778 & ~n33012;
  assign n33014 = ~n33006 & ~n33013;
  assign n33015 = ~n17845 & n33014;
  assign n33016 = ~n17847 & n33015;
  assign n33017 = ~n17849 & n33016;
  assign n33018 = ~n17851 & n33017;
  assign n33019 = ~n17857 & n33018;
  assign n33020 = ~pi0647 & n33019;
  assign n33021 = pi0647 & n33003;
  assign n33022 = ~pi1157 & ~n33021;
  assign n33023 = ~n33020 & n33022;
  assign n33024 = pi0630 & n33023;
  assign n33025 = pi0748 & n17244;
  assign n33026 = ~n33003 & ~n33025;
  assign n33027 = ~n17874 & ~n33026;
  assign n33028 = ~pi0785 & ~n33027;
  assign n33029 = ~n17879 & ~n33026;
  assign n33030 = pi1155 & ~n33029;
  assign n33031 = ~n17882 & n33027;
  assign n33032 = ~pi1155 & ~n33031;
  assign n33033 = ~n33030 & ~n33032;
  assign n33034 = pi0785 & ~n33033;
  assign n33035 = ~n33028 & ~n33034;
  assign n33036 = ~pi0781 & ~n33035;
  assign n33037 = ~n17889 & n33035;
  assign n33038 = pi1154 & ~n33037;
  assign n33039 = ~n17892 & n33035;
  assign n33040 = ~pi1154 & ~n33039;
  assign n33041 = ~n33038 & ~n33040;
  assign n33042 = pi0781 & ~n33041;
  assign n33043 = ~n33036 & ~n33042;
  assign n33044 = ~pi0789 & ~n33043;
  assign n33045 = ~pi0619 & n33003;
  assign n33046 = pi0619 & n33043;
  assign n33047 = pi1159 & ~n33045;
  assign n33048 = ~n33046 & n33047;
  assign n33049 = ~pi0619 & n33043;
  assign n33050 = pi0619 & n33003;
  assign n33051 = ~pi1159 & ~n33050;
  assign n33052 = ~n33049 & n33051;
  assign n33053 = ~n33048 & ~n33052;
  assign n33054 = pi0789 & ~n33053;
  assign n33055 = ~n33044 & ~n33054;
  assign n33056 = ~n17969 & n33055;
  assign n33057 = n17969 & n33003;
  assign n33058 = ~n33056 & ~n33057;
  assign n33059 = ~n17779 & ~n33058;
  assign n33060 = n17779 & n33003;
  assign n33061 = ~n33059 & ~n33060;
  assign n33062 = ~n20559 & n33061;
  assign n33063 = pi0647 & ~n33019;
  assign n33064 = ~pi0647 & ~n33003;
  assign n33065 = ~n33063 & ~n33064;
  assign n33066 = n17801 & ~n33065;
  assign n33067 = ~n33024 & ~n33066;
  assign n33068 = ~n33062 & n33067;
  assign n33069 = pi0787 & ~n33068;
  assign n33070 = n17871 & n33017;
  assign n33071 = ~pi0626 & ~n33055;
  assign n33072 = pi0626 & ~n33003;
  assign n33073 = n16629 & ~n33072;
  assign n33074 = ~n33071 & n33073;
  assign n33075 = pi0626 & ~n33055;
  assign n33076 = ~pi0626 & ~n33003;
  assign n33077 = n16628 & ~n33076;
  assign n33078 = ~n33075 & n33077;
  assign n33079 = ~n33070 & ~n33074;
  assign n33080 = ~n33078 & n33079;
  assign n33081 = pi0788 & ~n33080;
  assign n33082 = pi0618 & n33015;
  assign n33083 = pi0609 & n33014;
  assign n33084 = ~n17168 & ~n33005;
  assign n33085 = pi0625 & n33084;
  assign n33086 = n33026 & ~n33084;
  assign n33087 = ~n33085 & ~n33086;
  assign n33088 = n33010 & ~n33087;
  assign n33089 = ~pi0608 & ~n33009;
  assign n33090 = ~n33088 & n33089;
  assign n33091 = pi1153 & n33026;
  assign n33092 = ~n33085 & n33091;
  assign n33093 = pi0608 & ~n33011;
  assign n33094 = ~n33092 & n33093;
  assign n33095 = ~n33090 & ~n33094;
  assign n33096 = pi0778 & ~n33095;
  assign n33097 = ~pi0778 & ~n33086;
  assign n33098 = ~n33096 & ~n33097;
  assign n33099 = ~pi0609 & ~n33098;
  assign n33100 = ~pi1155 & ~n33083;
  assign n33101 = ~n33099 & n33100;
  assign n33102 = ~pi0660 & ~n33030;
  assign n33103 = ~n33101 & n33102;
  assign n33104 = ~pi0609 & n33014;
  assign n33105 = pi0609 & ~n33098;
  assign n33106 = pi1155 & ~n33104;
  assign n33107 = ~n33105 & n33106;
  assign n33108 = pi0660 & ~n33032;
  assign n33109 = ~n33107 & n33108;
  assign n33110 = ~n33103 & ~n33109;
  assign n33111 = pi0785 & ~n33110;
  assign n33112 = ~pi0785 & ~n33098;
  assign n33113 = ~n33111 & ~n33112;
  assign n33114 = ~pi0618 & ~n33113;
  assign n33115 = ~pi1154 & ~n33082;
  assign n33116 = ~n33114 & n33115;
  assign n33117 = ~pi0627 & ~n33038;
  assign n33118 = ~n33116 & n33117;
  assign n33119 = ~pi0618 & n33015;
  assign n33120 = pi0618 & ~n33113;
  assign n33121 = pi1154 & ~n33119;
  assign n33122 = ~n33120 & n33121;
  assign n33123 = pi0627 & ~n33040;
  assign n33124 = ~n33122 & n33123;
  assign n33125 = ~n33118 & ~n33124;
  assign n33126 = pi0781 & ~n33125;
  assign n33127 = ~pi0781 & ~n33113;
  assign n33128 = ~n33126 & ~n33127;
  assign n33129 = ~pi0789 & n33128;
  assign n33130 = ~pi0619 & ~n33128;
  assign n33131 = pi0619 & n33016;
  assign n33132 = ~pi1159 & ~n33131;
  assign n33133 = ~n33130 & n33132;
  assign n33134 = ~pi0648 & ~n33048;
  assign n33135 = ~n33133 & n33134;
  assign n33136 = pi0619 & ~n33128;
  assign n33137 = ~pi0619 & n33016;
  assign n33138 = pi1159 & ~n33137;
  assign n33139 = ~n33136 & n33138;
  assign n33140 = pi0648 & ~n33052;
  assign n33141 = ~n33139 & n33140;
  assign n33142 = pi0789 & ~n33135;
  assign n33143 = ~n33141 & n33142;
  assign n33144 = n17970 & ~n33129;
  assign n33145 = ~n33143 & n33144;
  assign n33146 = ~n33081 & ~n33145;
  assign n33147 = ~n20364 & ~n33146;
  assign n33148 = n17854 & ~n33058;
  assign n33149 = n20851 & n33018;
  assign n33150 = ~n33148 & ~n33149;
  assign n33151 = ~pi0629 & ~n33150;
  assign n33152 = n20855 & n33018;
  assign n33153 = n17853 & ~n33058;
  assign n33154 = ~n33152 & ~n33153;
  assign n33155 = pi0629 & ~n33154;
  assign n33156 = ~n33151 & ~n33155;
  assign n33157 = pi0792 & ~n33156;
  assign n33158 = ~n20206 & ~n33157;
  assign n33159 = ~n33147 & n33158;
  assign n33160 = ~n33069 & ~n33159;
  assign n33161 = ~pi0790 & n33160;
  assign n33162 = ~pi0787 & ~n33019;
  assign n33163 = pi1157 & ~n33065;
  assign n33164 = ~n33023 & ~n33163;
  assign n33165 = pi0787 & ~n33164;
  assign n33166 = ~n33162 & ~n33165;
  assign n33167 = ~pi0644 & n33166;
  assign n33168 = pi0644 & n33160;
  assign n33169 = pi0715 & ~n33167;
  assign n33170 = ~n33168 & n33169;
  assign n33171 = ~n17804 & ~n33061;
  assign n33172 = n17804 & n33003;
  assign n33173 = ~n33171 & ~n33172;
  assign n33174 = pi0644 & ~n33173;
  assign n33175 = ~pi0644 & n33003;
  assign n33176 = ~pi0715 & ~n33175;
  assign n33177 = ~n33174 & n33176;
  assign n33178 = pi1160 & ~n33177;
  assign n33179 = ~n33170 & n33178;
  assign n33180 = ~pi0644 & ~n33173;
  assign n33181 = pi0644 & n33003;
  assign n33182 = pi0715 & ~n33181;
  assign n33183 = ~n33180 & n33182;
  assign n33184 = pi0644 & n33166;
  assign n33185 = ~pi0644 & n33160;
  assign n33186 = ~pi0715 & ~n33184;
  assign n33187 = ~n33185 & n33186;
  assign n33188 = ~pi1160 & ~n33183;
  assign n33189 = ~n33187 & n33188;
  assign n33190 = ~n33179 & ~n33189;
  assign n33191 = pi0790 & ~n33190;
  assign n33192 = pi0832 & ~n33161;
  assign n33193 = ~n33191 & n33192;
  assign po0351 = ~n33002 & ~n33193;
  assign n33195 = ~pi0138 & n16565;
  assign n33196 = ~pi0196 & n33195;
  assign n33197 = pi0195 & ~n33196;
  assign n33198 = ~n11477 & n16193;
  assign n33199 = ~n6198 & n16168;
  assign n33200 = n16167 & ~n16493;
  assign n33201 = ~n11480 & ~n33199;
  assign n33202 = ~n33198 & ~n33200;
  assign n33203 = n33201 & n33202;
  assign n33204 = pi0232 & ~n33203;
  assign n33205 = ~n16491 & ~n33204;
  assign n33206 = pi0039 & ~n33205;
  assign n33207 = n13910 & ~n16170;
  assign n33208 = ~pi0039 & ~n33207;
  assign n33209 = n10200 & ~n33197;
  assign n33210 = ~n33208 & n33209;
  assign n33211 = ~n33206 & n33210;
  assign n33212 = ~pi0171 & n9326;
  assign n33213 = ~n16522 & ~n33212;
  assign n33214 = n9036 & ~n33213;
  assign n33215 = n9291 & ~n33214;
  assign n33216 = ~pi0192 & n16511;
  assign n33217 = pi0192 & n16520;
  assign n33218 = ~n33215 & ~n33216;
  assign n33219 = ~n33217 & n33218;
  assign n33220 = pi0232 & ~n33219;
  assign n33221 = ~n16517 & ~n33220;
  assign n33222 = pi0039 & ~n33221;
  assign n33223 = pi0192 & n16539;
  assign n33224 = ~n9605 & ~n16162;
  assign n33225 = pi0171 & n13737;
  assign n33226 = ~n33224 & ~n33225;
  assign n33227 = pi0299 & ~n33226;
  assign n33228 = ~pi0192 & n16533;
  assign n33229 = pi0232 & ~n33228;
  assign n33230 = ~n33223 & n33229;
  assign n33231 = ~n33227 & n33230;
  assign n33232 = n16536 & ~n33231;
  assign n33233 = n2608 & ~n33222;
  assign n33234 = ~n33232 & n33233;
  assign n33235 = ~pi0087 & ~n33234;
  assign n33236 = n16508 & ~n33235;
  assign n33237 = ~pi0092 & ~n33236;
  assign n33238 = n16507 & ~n33237;
  assign n33239 = ~pi0055 & ~n33238;
  assign n33240 = ~n16559 & ~n33239;
  assign n33241 = n2529 & ~n33240;
  assign n33242 = n9883 & n33197;
  assign n33243 = ~n33241 & n33242;
  assign po0352 = n33211 | n33243;
  assign n33245 = n13132 & n16492;
  assign n33246 = ~pi0170 & n9039;
  assign n33247 = ~n16492 & ~n33246;
  assign n33248 = n13130 & ~n33247;
  assign n33249 = pi0232 & ~n33245;
  assign n33250 = ~n33248 & n33249;
  assign n33251 = ~n16491 & ~n33250;
  assign n33252 = pi0039 & ~n33251;
  assign n33253 = n13910 & n16287;
  assign n33254 = ~pi0039 & ~n33253;
  assign n33255 = ~pi0038 & ~n33254;
  assign n33256 = ~n33252 & n33255;
  assign n33257 = pi0194 & ~n33256;
  assign n33258 = pi0299 & ~n33251;
  assign n33259 = ~n11478 & ~n33258;
  assign n33260 = pi0039 & ~n33259;
  assign n33261 = n13910 & ~n16275;
  assign n33262 = ~pi0039 & ~n33261;
  assign n33263 = ~pi0038 & ~n33262;
  assign n33264 = ~n33260 & n33263;
  assign n33265 = ~pi0194 & ~n33264;
  assign n33266 = n10197 & ~n33257;
  assign n33267 = ~n33265 & n33266;
  assign n33268 = ~pi0196 & ~n33267;
  assign n33269 = ~pi0170 & n9326;
  assign n33270 = ~n16522 & ~n33269;
  assign n33271 = n9036 & ~n33270;
  assign n33272 = n9291 & ~n33271;
  assign n33273 = ~n16511 & ~n33272;
  assign n33274 = pi0232 & ~n33273;
  assign n33275 = ~n16517 & ~n33274;
  assign n33276 = pi0232 & n16520;
  assign n33277 = n33275 & ~n33276;
  assign n33278 = pi0039 & ~n33277;
  assign n33279 = ~pi0038 & pi0194;
  assign n33280 = ~n33278 & n33279;
  assign n33281 = pi0039 & ~n33275;
  assign n33282 = ~pi0038 & ~pi0194;
  assign n33283 = ~n33281 & n33282;
  assign n33284 = ~n33280 & ~n33283;
  assign n33285 = ~n16536 & ~n33284;
  assign n33286 = ~n9605 & ~n16274;
  assign n33287 = pi0170 & n13737;
  assign n33288 = ~n33286 & ~n33287;
  assign n33289 = pi0299 & ~n33288;
  assign n33290 = ~n16539 & n33280;
  assign n33291 = ~n16533 & n33283;
  assign n33292 = ~n33290 & ~n33291;
  assign n33293 = pi0232 & ~n33289;
  assign n33294 = ~n33292 & n33293;
  assign n33295 = ~n33285 & ~n33294;
  assign n33296 = ~pi0100 & ~n33295;
  assign n33297 = ~pi0087 & ~n33296;
  assign n33298 = n16508 & ~n33297;
  assign n33299 = ~pi0092 & ~n33298;
  assign n33300 = n16507 & ~n33299;
  assign n33301 = ~pi0055 & ~n33300;
  assign n33302 = ~n16559 & ~n33301;
  assign n33303 = n2529 & ~n33302;
  assign n33304 = n9883 & ~n33303;
  assign n33305 = pi0196 & ~n33304;
  assign n33306 = ~n33195 & ~n33268;
  assign n33307 = ~n33305 & n33306;
  assign n33308 = pi0195 & ~pi0196;
  assign n33309 = ~n33267 & ~n33308;
  assign n33310 = ~n33304 & n33308;
  assign n33311 = n33195 & ~n33309;
  assign n33312 = ~n33310 & n33311;
  assign po0353 = n33307 | n33312;
  assign n33314 = ~pi0197 & ~n2926;
  assign n33315 = ~pi0767 & pi0947;
  assign n33316 = ~pi0698 & n20902;
  assign n33317 = ~n33315 & ~n33316;
  assign n33318 = n2926 & ~n33317;
  assign n33319 = pi0832 & ~n33314;
  assign n33320 = ~n33318 & n33319;
  assign n33321 = ~pi0197 & ~n10197;
  assign n33322 = n16641 & ~n33315;
  assign n33323 = pi0197 & ~n17050;
  assign n33324 = pi0038 & ~n33322;
  assign n33325 = ~n33323 & n33324;
  assign n33326 = ~pi0197 & ~n16958;
  assign n33327 = n16958 & n33315;
  assign n33328 = ~pi0039 & ~n33326;
  assign n33329 = ~n33327 & n33328;
  assign n33330 = ~pi0197 & ~n21001;
  assign n33331 = pi0197 & ~n21162;
  assign n33332 = pi0299 & ~n33331;
  assign n33333 = ~n33330 & n33332;
  assign n33334 = ~pi0197 & ~n17024;
  assign n33335 = n21019 & ~n33334;
  assign n33336 = ~pi0767 & ~n33335;
  assign n33337 = ~n33333 & n33336;
  assign n33338 = ~pi0197 & pi0767;
  assign n33339 = ~n17046 & n33338;
  assign n33340 = pi0039 & ~n33339;
  assign n33341 = ~n33337 & n33340;
  assign n33342 = ~pi0038 & ~n33329;
  assign n33343 = ~n33341 & n33342;
  assign n33344 = ~n33325 & ~n33343;
  assign n33345 = pi0698 & ~n33344;
  assign n33346 = ~n21114 & n33329;
  assign n33347 = n21111 & ~n33334;
  assign n33348 = pi0197 & n21108;
  assign n33349 = ~pi0197 & n21092;
  assign n33350 = pi0299 & ~n33348;
  assign n33351 = ~n33349 & n33350;
  assign n33352 = pi0767 & ~n33347;
  assign n33353 = ~n33351 & n33352;
  assign n33354 = ~pi0197 & n21064;
  assign n33355 = pi0197 & n21080;
  assign n33356 = ~pi0767 & ~n33355;
  assign n33357 = ~n33354 & n33356;
  assign n33358 = pi0039 & ~n33353;
  assign n33359 = ~n33357 & n33358;
  assign n33360 = ~n33346 & ~n33359;
  assign n33361 = ~pi0038 & ~n33360;
  assign n33362 = ~pi0197 & ~n16641;
  assign n33363 = pi0767 & pi0947;
  assign n33364 = ~pi0039 & ~n33363;
  assign n33365 = n21239 & n33364;
  assign n33366 = pi0038 & ~n33362;
  assign n33367 = ~n33365 & n33366;
  assign n33368 = ~pi0698 & ~n33367;
  assign n33369 = ~n33361 & n33368;
  assign n33370 = ~n33345 & ~n33369;
  assign n33371 = n10197 & ~n33370;
  assign n33372 = ~pi0832 & ~n33321;
  assign n33373 = ~n33371 & n33372;
  assign po0354 = ~n33320 & ~n33373;
  assign n33375 = n2530 & ~n16958;
  assign n33376 = n18591 & ~n33375;
  assign n33377 = pi0198 & ~n33376;
  assign n33378 = pi0198 & ~n16797;
  assign n33379 = pi0198 & ~n16653;
  assign n33380 = ~po1101 & ~n33379;
  assign n33381 = n33378 & ~n33380;
  assign n33382 = n6192 & ~n16721;
  assign n33383 = ~n6192 & ~n16723;
  assign n33384 = pi0198 & ~n33382;
  assign n33385 = ~n33383 & n33384;
  assign n33386 = ~n6242 & n33385;
  assign n33387 = ~n33381 & ~n33386;
  assign n33388 = pi0215 & ~n33387;
  assign n33389 = n3448 & ~n33379;
  assign n33390 = pi0198 & ~n16684;
  assign n33391 = po1101 & ~n33390;
  assign n33392 = ~n33380 & ~n33391;
  assign n33393 = n6242 & n33392;
  assign n33394 = pi0198 & ~n17143;
  assign n33395 = ~n6242 & n33394;
  assign n33396 = ~n3448 & ~n33393;
  assign n33397 = ~n33395 & n33396;
  assign n33398 = ~pi0215 & ~n33389;
  assign n33399 = ~n33397 & n33398;
  assign n33400 = pi0299 & ~n33388;
  assign n33401 = ~n33399 & n33400;
  assign n33402 = ~n6205 & n33385;
  assign n33403 = ~n33381 & ~n33402;
  assign n33404 = pi0223 & ~n33403;
  assign n33405 = n2603 & ~n33379;
  assign n33406 = ~n6205 & n33394;
  assign n33407 = n6205 & n33392;
  assign n33408 = ~n2603 & ~n33407;
  assign n33409 = ~n33406 & n33408;
  assign n33410 = ~pi0223 & ~n33405;
  assign n33411 = ~n33409 & n33410;
  assign n33412 = ~pi0299 & ~n33404;
  assign n33413 = ~n33411 & n33412;
  assign n33414 = n2571 & n10982;
  assign n33415 = ~n33401 & n33414;
  assign n33416 = ~n33413 & n33415;
  assign n33417 = ~n33377 & ~n33416;
  assign n33418 = ~n19149 & n33417;
  assign n33419 = n16639 & ~n33417;
  assign n33420 = pi0198 & ~n2571;
  assign n33421 = pi0039 & pi0198;
  assign n33422 = pi0038 & ~n33421;
  assign n33423 = pi0198 & ~n16667;
  assign n33424 = pi0634 & n16644;
  assign n33425 = n16667 & n33424;
  assign n33426 = ~n33423 & ~n33425;
  assign n33427 = ~pi0039 & ~n33426;
  assign n33428 = n33422 & ~n33427;
  assign n33429 = pi0198 & n16721;
  assign n33430 = pi0634 & ~n16721;
  assign n33431 = n16658 & n33430;
  assign n33432 = ~n33429 & ~n33431;
  assign n33433 = n6195 & ~n33432;
  assign n33434 = ~pi0680 & n33385;
  assign n33435 = n6192 & n33432;
  assign n33436 = ~n16658 & ~n33379;
  assign n33437 = pi0634 & ~n33436;
  assign n33438 = ~n33379 & ~n33437;
  assign n33439 = ~n6197 & n33438;
  assign n33440 = n6197 & n33432;
  assign n33441 = ~n33439 & ~n33440;
  assign n33442 = ~n6192 & ~n33441;
  assign n33443 = n17323 & ~n33435;
  assign n33444 = ~n33442 & n33443;
  assign n33445 = ~n33433 & ~n33434;
  assign n33446 = ~n33444 & n33445;
  assign n33447 = ~n6205 & n33446;
  assign n33448 = n33378 & n33434;
  assign n33449 = n6197 & ~n33438;
  assign n33450 = ~n6197 & ~n33432;
  assign n33451 = ~n33449 & ~n33450;
  assign n33452 = n6192 & n33451;
  assign n33453 = ~n6192 & n33438;
  assign n33454 = n17323 & ~n33453;
  assign n33455 = ~n33452 & n33454;
  assign n33456 = n6195 & ~n33451;
  assign n33457 = ~n33448 & ~n33456;
  assign n33458 = ~n33455 & n33457;
  assign n33459 = n6205 & n33458;
  assign n33460 = pi0223 & ~n33447;
  assign n33461 = ~n33459 & n33460;
  assign n33462 = pi0680 & n33437;
  assign n33463 = ~n33379 & ~n33462;
  assign n33464 = n2603 & n33463;
  assign n33465 = pi0198 & n16681;
  assign n33466 = pi0634 & n16686;
  assign n33467 = ~n33465 & ~n33466;
  assign n33468 = ~n6197 & ~n33467;
  assign n33469 = ~n33449 & ~n33468;
  assign n33470 = n6195 & ~n33469;
  assign n33471 = n6192 & n33469;
  assign n33472 = n33454 & ~n33471;
  assign n33473 = ~n6192 & ~n33379;
  assign n33474 = n6192 & ~n33390;
  assign n33475 = ~pi0680 & ~n33473;
  assign n33476 = ~n33474 & n33475;
  assign n33477 = ~n33470 & ~n33476;
  assign n33478 = ~n33472 & n33477;
  assign n33479 = n6205 & ~n33478;
  assign n33480 = pi0198 & n16753;
  assign n33481 = n6195 & ~n33467;
  assign n33482 = n6192 & n33467;
  assign n33483 = n6197 & n33467;
  assign n33484 = ~n33439 & ~n33483;
  assign n33485 = ~n6192 & ~n33484;
  assign n33486 = n17323 & ~n33482;
  assign n33487 = ~n33485 & n33486;
  assign n33488 = ~n33480 & ~n33481;
  assign n33489 = ~n33487 & n33488;
  assign n33490 = ~n6205 & ~n33489;
  assign n33491 = ~n2603 & ~n33479;
  assign n33492 = ~n33490 & n33491;
  assign n33493 = ~pi0223 & ~n33464;
  assign n33494 = ~n33492 & n33493;
  assign n33495 = ~pi0299 & ~n33461;
  assign n33496 = ~n33494 & n33495;
  assign n33497 = ~n6242 & n33446;
  assign n33498 = n6242 & n33458;
  assign n33499 = pi0215 & ~n33497;
  assign n33500 = ~n33498 & n33499;
  assign n33501 = n3448 & n33463;
  assign n33502 = ~n6242 & ~n33489;
  assign n33503 = n6242 & ~n33478;
  assign n33504 = ~n3448 & ~n33502;
  assign n33505 = ~n33503 & n33504;
  assign n33506 = ~pi0215 & ~n33501;
  assign n33507 = ~n33505 & n33506;
  assign n33508 = pi0299 & ~n33500;
  assign n33509 = ~n33507 & n33508;
  assign n33510 = ~n33496 & ~n33509;
  assign n33511 = pi0039 & ~n33510;
  assign n33512 = pi0634 & pi0680;
  assign n33513 = pi0198 & n16931;
  assign n33514 = ~n16896 & n33512;
  assign n33515 = ~n33513 & n33514;
  assign n33516 = ~n16929 & ~n33515;
  assign n33517 = ~pi0299 & ~n33516;
  assign n33518 = ~pi0198 & n16923;
  assign n33519 = pi0198 & ~n16944;
  assign n33520 = ~n33518 & ~n33519;
  assign n33521 = n33512 & ~n33520;
  assign n33522 = pi0198 & ~n16941;
  assign n33523 = ~n33512 & n33522;
  assign n33524 = ~n33521 & ~n33523;
  assign n33525 = pi0299 & ~n33524;
  assign n33526 = ~pi0039 & ~n33517;
  assign n33527 = ~n33525 & n33526;
  assign n33528 = ~n33511 & ~n33527;
  assign n33529 = ~pi0038 & ~n33528;
  assign n33530 = n2571 & ~n33428;
  assign n33531 = ~n33529 & n33530;
  assign n33532 = ~n33420 & ~n33531;
  assign n33533 = ~pi0778 & ~n33532;
  assign n33534 = ~pi0625 & n33417;
  assign n33535 = pi0625 & n33532;
  assign n33536 = pi1153 & ~n33534;
  assign n33537 = ~n33535 & n33536;
  assign n33538 = ~pi0625 & n33532;
  assign n33539 = pi0625 & n33417;
  assign n33540 = ~pi1153 & ~n33539;
  assign n33541 = ~n33538 & n33540;
  assign n33542 = ~n33537 & ~n33541;
  assign n33543 = pi0778 & ~n33542;
  assign n33544 = ~n33533 & ~n33543;
  assign n33545 = ~n17075 & n33544;
  assign n33546 = n17075 & n33417;
  assign n33547 = ~n33545 & ~n33546;
  assign n33548 = ~n16639 & n33547;
  assign n33549 = ~n33419 & ~n33548;
  assign n33550 = ~n16635 & n33549;
  assign n33551 = ~n16631 & n33550;
  assign n33552 = ~n33418 & ~n33551;
  assign n33553 = ~pi0792 & n33552;
  assign n33554 = pi0628 & ~n33552;
  assign n33555 = ~pi0628 & n33417;
  assign n33556 = ~n33554 & ~n33555;
  assign n33557 = pi1156 & n33556;
  assign n33558 = pi0628 & n33417;
  assign n33559 = ~pi0628 & ~n33552;
  assign n33560 = ~pi1156 & ~n33558;
  assign n33561 = ~n33559 & n33560;
  assign n33562 = ~n33557 & ~n33561;
  assign n33563 = pi0792 & ~n33562;
  assign n33564 = ~n33553 & ~n33563;
  assign n33565 = ~pi0647 & n33564;
  assign n33566 = pi0647 & n33417;
  assign n33567 = ~pi1157 & ~n33566;
  assign n33568 = ~n33565 & n33567;
  assign n33569 = pi0630 & n33568;
  assign n33570 = n17779 & ~n33417;
  assign n33571 = ~n17127 & ~n17131;
  assign n33572 = pi0633 & ~n33571;
  assign n33573 = ~n16929 & ~n33572;
  assign n33574 = ~n17136 & ~n33573;
  assign n33575 = ~pi0299 & n33574;
  assign n33576 = pi0603 & pi0633;
  assign n33577 = ~n33522 & ~n33576;
  assign n33578 = pi0198 & ~n17122;
  assign n33579 = ~pi0198 & n17230;
  assign n33580 = ~n33578 & ~n33579;
  assign n33581 = n33576 & n33580;
  assign n33582 = ~n33577 & ~n33581;
  assign n33583 = pi0299 & n33582;
  assign n33584 = ~pi0039 & ~n33575;
  assign n33585 = ~n33583 & n33584;
  assign n33586 = pi0633 & n17239;
  assign n33587 = ~n33385 & ~n33586;
  assign n33588 = ~n6195 & ~n33587;
  assign n33589 = pi0633 & n16653;
  assign n33590 = ~n17144 & n33589;
  assign n33591 = ~n16721 & n33590;
  assign n33592 = ~n33429 & ~n33591;
  assign n33593 = n17188 & ~n33592;
  assign n33594 = ~n33588 & ~n33593;
  assign n33595 = ~n6205 & n33594;
  assign n33596 = ~n33379 & ~n33590;
  assign n33597 = pi0603 & ~n33596;
  assign n33598 = ~pi0603 & n33379;
  assign n33599 = ~n33597 & ~n33598;
  assign n33600 = ~n17167 & n33599;
  assign n33601 = n6197 & ~n33596;
  assign n33602 = ~n33378 & ~n33591;
  assign n33603 = ~n33601 & n33602;
  assign n33604 = pi0603 & ~n33603;
  assign n33605 = n17167 & ~n33598;
  assign n33606 = ~n33604 & n33605;
  assign n33607 = ~n33600 & ~n33606;
  assign n33608 = ~n6195 & n33607;
  assign n33609 = ~n33378 & ~n33604;
  assign n33610 = n6195 & ~n33609;
  assign n33611 = ~n33608 & ~n33610;
  assign n33612 = n6205 & n33611;
  assign n33613 = pi0223 & ~n33595;
  assign n33614 = ~n33612 & n33613;
  assign n33615 = n2603 & n33599;
  assign n33616 = pi0642 & ~n33597;
  assign n33617 = pi0633 & n17147;
  assign n33618 = ~n33465 & ~n33617;
  assign n33619 = ~n6197 & ~n33618;
  assign n33620 = ~n33601 & ~n33619;
  assign n33621 = pi0603 & ~n33620;
  assign n33622 = ~pi0642 & ~n33621;
  assign n33623 = n6191 & ~n33616;
  assign n33624 = ~n33622 & n33623;
  assign n33625 = ~n6191 & n33597;
  assign n33626 = ~n33598 & ~n33625;
  assign n33627 = ~n33624 & n33626;
  assign n33628 = ~n6195 & n33627;
  assign n33629 = ~pi0603 & n33390;
  assign n33630 = n6195 & ~n33629;
  assign n33631 = ~n33621 & n33630;
  assign n33632 = ~n33628 & ~n33631;
  assign n33633 = n6205 & n33632;
  assign n33634 = pi0603 & ~n33618;
  assign n33635 = n17167 & n33634;
  assign n33636 = pi0198 & n17149;
  assign n33637 = n6197 & n33618;
  assign n33638 = ~n6197 & n33596;
  assign n33639 = pi0603 & ~n17167;
  assign n33640 = ~n33638 & n33639;
  assign n33641 = ~n33637 & n33640;
  assign n33642 = ~n33635 & ~n33636;
  assign n33643 = ~n33641 & n33642;
  assign n33644 = ~n6195 & n33643;
  assign n33645 = n6195 & ~n33465;
  assign n33646 = ~n33634 & n33645;
  assign n33647 = ~n33644 & ~n33646;
  assign n33648 = ~n6205 & n33647;
  assign n33649 = ~n2603 & ~n33648;
  assign n33650 = ~n33633 & n33649;
  assign n33651 = ~pi0223 & ~n33615;
  assign n33652 = ~n33650 & n33651;
  assign n33653 = ~n33614 & ~n33652;
  assign n33654 = ~pi0299 & ~n33653;
  assign n33655 = ~n6242 & n33594;
  assign n33656 = n6242 & n33611;
  assign n33657 = pi0215 & ~n33655;
  assign n33658 = ~n33656 & n33657;
  assign n33659 = n3448 & n33599;
  assign n33660 = ~n6242 & n33647;
  assign n33661 = n6242 & n33632;
  assign n33662 = ~n3448 & ~n33660;
  assign n33663 = ~n33661 & n33662;
  assign n33664 = ~pi0215 & ~n33659;
  assign n33665 = ~n33663 & n33664;
  assign n33666 = ~n33658 & ~n33665;
  assign n33667 = pi0299 & ~n33666;
  assign n33668 = pi0039 & ~n33654;
  assign n33669 = ~n33667 & n33668;
  assign n33670 = ~n33585 & ~n33669;
  assign n33671 = ~pi0038 & ~n33670;
  assign n33672 = pi0633 & n17168;
  assign n33673 = n16667 & n33672;
  assign n33674 = ~n33423 & ~n33673;
  assign n33675 = ~pi0039 & ~n33674;
  assign n33676 = n33422 & ~n33675;
  assign n33677 = n2571 & ~n33676;
  assign n33678 = ~n33671 & n33677;
  assign n33679 = ~n33420 & ~n33678;
  assign n33680 = ~n17117 & ~n33679;
  assign n33681 = n17117 & ~n33417;
  assign n33682 = ~n33680 & ~n33681;
  assign n33683 = ~pi0785 & ~n33682;
  assign n33684 = ~n17291 & ~n33417;
  assign n33685 = pi0609 & n33680;
  assign n33686 = ~n33684 & ~n33685;
  assign n33687 = pi1155 & ~n33686;
  assign n33688 = ~n17296 & ~n33417;
  assign n33689 = ~pi0609 & n33680;
  assign n33690 = ~n33688 & ~n33689;
  assign n33691 = ~pi1155 & ~n33690;
  assign n33692 = ~n33687 & ~n33691;
  assign n33693 = pi0785 & ~n33692;
  assign n33694 = ~n33683 & ~n33693;
  assign n33695 = ~pi0781 & ~n33694;
  assign n33696 = ~pi0618 & n33417;
  assign n33697 = pi0618 & n33694;
  assign n33698 = pi1154 & ~n33696;
  assign n33699 = ~n33697 & n33698;
  assign n33700 = ~pi0618 & n33694;
  assign n33701 = pi0618 & n33417;
  assign n33702 = ~pi1154 & ~n33701;
  assign n33703 = ~n33700 & n33702;
  assign n33704 = ~n33699 & ~n33703;
  assign n33705 = pi0781 & ~n33704;
  assign n33706 = ~n33695 & ~n33705;
  assign n33707 = ~pi0789 & ~n33706;
  assign n33708 = ~pi0619 & n33417;
  assign n33709 = pi0619 & n33706;
  assign n33710 = pi1159 & ~n33708;
  assign n33711 = ~n33709 & n33710;
  assign n33712 = ~pi0619 & n33706;
  assign n33713 = pi0619 & n33417;
  assign n33714 = ~pi1159 & ~n33713;
  assign n33715 = ~n33712 & n33714;
  assign n33716 = ~n33711 & ~n33715;
  assign n33717 = pi0789 & ~n33716;
  assign n33718 = ~n33707 & ~n33717;
  assign n33719 = ~n17969 & n33718;
  assign n33720 = n17969 & n33417;
  assign n33721 = ~n33719 & ~n33720;
  assign n33722 = ~n17779 & n33721;
  assign n33723 = ~n33570 & ~n33722;
  assign n33724 = ~n20559 & ~n33723;
  assign n33725 = pi0647 & ~n33564;
  assign n33726 = ~pi0647 & ~n33417;
  assign n33727 = ~n33725 & ~n33726;
  assign n33728 = n17801 & ~n33727;
  assign n33729 = ~n33569 & ~n33728;
  assign n33730 = ~n33724 & n33729;
  assign n33731 = pi0787 & ~n33730;
  assign n33732 = pi0629 & n33561;
  assign n33733 = ~n20570 & n33721;
  assign n33734 = n17776 & n33556;
  assign n33735 = ~n33732 & ~n33734;
  assign n33736 = ~n33733 & n33735;
  assign n33737 = pi0792 & ~n33736;
  assign n33738 = n16635 & n33417;
  assign n33739 = ~n33550 & ~n33738;
  assign n33740 = n17871 & ~n33739;
  assign n33741 = ~pi0626 & ~n33718;
  assign n33742 = pi0626 & ~n33417;
  assign n33743 = n16629 & ~n33742;
  assign n33744 = ~n33741 & n33743;
  assign n33745 = pi0626 & ~n33718;
  assign n33746 = ~pi0626 & ~n33417;
  assign n33747 = n16628 & ~n33746;
  assign n33748 = ~n33745 & n33747;
  assign n33749 = ~n33740 & ~n33744;
  assign n33750 = ~n33748 & n33749;
  assign n33751 = pi0788 & ~n33750;
  assign n33752 = pi0609 & n33544;
  assign n33753 = pi0634 & n17645;
  assign n33754 = n33674 & ~n33753;
  assign n33755 = ~pi0039 & ~n33754;
  assign n33756 = n33422 & ~n33755;
  assign n33757 = ~n33512 & n33582;
  assign n33758 = ~pi0603 & ~n33520;
  assign n33759 = ~pi0198 & ~pi0665;
  assign n33760 = n17122 & n33759;
  assign n33761 = ~n17230 & n33519;
  assign n33762 = ~pi0633 & ~n33760;
  assign n33763 = ~n33761 & n33762;
  assign n33764 = pi0198 & ~pi0665;
  assign n33765 = pi0633 & ~n33764;
  assign n33766 = ~n33518 & n33765;
  assign n33767 = n33580 & n33766;
  assign n33768 = pi0603 & ~n33763;
  assign n33769 = ~n33767 & n33768;
  assign n33770 = ~n33758 & ~n33769;
  assign n33771 = n33512 & ~n33770;
  assign n33772 = pi0299 & ~n33757;
  assign n33773 = ~n33771 & n33772;
  assign n33774 = ~pi0680 & n33574;
  assign n33775 = ~pi0603 & n33516;
  assign n33776 = pi0198 & ~pi0633;
  assign n33777 = pi0634 & ~pi0665;
  assign n33778 = ~n33776 & n33777;
  assign n33779 = ~n17126 & n33778;
  assign n33780 = ~pi0634 & n16929;
  assign n33781 = pi0634 & n16932;
  assign n33782 = ~n17133 & n33781;
  assign n33783 = ~n33780 & ~n33782;
  assign n33784 = ~pi0633 & ~n33783;
  assign n33785 = pi0603 & ~n33779;
  assign n33786 = ~n33572 & n33785;
  assign n33787 = ~n33784 & n33786;
  assign n33788 = pi0680 & ~n33775;
  assign n33789 = ~n33787 & n33788;
  assign n33790 = ~pi0299 & ~n33774;
  assign n33791 = ~n33789 & n33790;
  assign n33792 = ~n33773 & ~n33791;
  assign n33793 = ~pi0039 & ~n33792;
  assign n33794 = n17355 & n33437;
  assign n33795 = n33599 & ~n33794;
  assign n33796 = n2603 & n33795;
  assign n33797 = ~pi0680 & n33627;
  assign n33798 = ~pi0603 & ~n33438;
  assign n33799 = n17159 & n33777;
  assign n33800 = n33596 & ~n33799;
  assign n33801 = pi0603 & ~n33800;
  assign n33802 = ~n33798 & ~n33801;
  assign n33803 = ~n6191 & ~n33802;
  assign n33804 = n6197 & ~n33800;
  assign n33805 = pi0634 & n17424;
  assign n33806 = n33618 & ~n33805;
  assign n33807 = ~n6197 & ~n33806;
  assign n33808 = ~n33804 & ~n33807;
  assign n33809 = pi0603 & ~n33808;
  assign n33810 = ~pi0642 & n33809;
  assign n33811 = pi0642 & n33801;
  assign n33812 = ~n33798 & ~n33811;
  assign n33813 = ~n33810 & n33812;
  assign n33814 = n6191 & ~n33813;
  assign n33815 = ~n16657 & ~n33803;
  assign n33816 = ~n33814 & n33815;
  assign n33817 = ~pi0603 & ~n33469;
  assign n33818 = n16657 & ~n33817;
  assign n33819 = ~n33809 & n33818;
  assign n33820 = ~n33816 & ~n33819;
  assign n33821 = pi0680 & ~n33820;
  assign n33822 = ~n33797 & ~n33821;
  assign n33823 = n6205 & n33822;
  assign n33824 = ~pi0680 & ~n33643;
  assign n33825 = ~pi0603 & n33484;
  assign n33826 = ~n17167 & n33801;
  assign n33827 = ~n33640 & ~n33826;
  assign n33828 = ~n6192 & n33827;
  assign n33829 = ~n6197 & ~n33827;
  assign n33830 = n33806 & ~n33829;
  assign n33831 = ~n33828 & ~n33830;
  assign n33832 = ~n33825 & ~n33831;
  assign n33833 = n17323 & ~n33832;
  assign n33834 = ~n17168 & ~n33467;
  assign n33835 = ~n33634 & ~n33834;
  assign n33836 = n6195 & ~n33835;
  assign n33837 = ~n33824 & ~n33836;
  assign n33838 = ~n33833 & n33837;
  assign n33839 = ~n6205 & ~n33838;
  assign n33840 = ~n2603 & ~n33839;
  assign n33841 = ~n33823 & n33840;
  assign n33842 = ~pi0223 & ~n33796;
  assign n33843 = ~n33841 & n33842;
  assign n33844 = ~pi0680 & ~n33587;
  assign n33845 = n17191 & n33759;
  assign n33846 = n17144 & n33764;
  assign n33847 = ~n33429 & ~n33846;
  assign n33848 = ~n33845 & n33847;
  assign n33849 = pi0634 & ~n33848;
  assign n33850 = ~pi0634 & n33429;
  assign n33851 = ~n33591 & ~n33850;
  assign n33852 = ~n33849 & n33851;
  assign n33853 = pi0603 & ~n33852;
  assign n33854 = ~pi0603 & ~n33432;
  assign n33855 = ~n33853 & ~n33854;
  assign n33856 = n6195 & ~n33855;
  assign n33857 = n17167 & n33853;
  assign n33858 = ~pi0603 & n33441;
  assign n33859 = ~n33827 & ~n33852;
  assign n33860 = ~n33829 & ~n33858;
  assign n33861 = ~n33857 & ~n33859;
  assign n33862 = n33860 & n33861;
  assign n33863 = n17323 & ~n33862;
  assign n33864 = ~n33844 & ~n33856;
  assign n33865 = ~n33863 & n33864;
  assign n33866 = ~n6205 & n33865;
  assign n33867 = ~pi0680 & n33607;
  assign n33868 = ~n6197 & ~n33852;
  assign n33869 = ~n33804 & ~n33868;
  assign n33870 = pi0603 & ~n33869;
  assign n33871 = ~pi0603 & ~n33451;
  assign n33872 = ~n33870 & ~n33871;
  assign n33873 = n6195 & ~n33872;
  assign n33874 = ~n17167 & n33802;
  assign n33875 = n17167 & ~n33798;
  assign n33876 = ~n33870 & n33875;
  assign n33877 = n17323 & ~n33874;
  assign n33878 = ~n33876 & n33877;
  assign n33879 = ~n33867 & ~n33873;
  assign n33880 = ~n33878 & n33879;
  assign n33881 = n6205 & n33880;
  assign n33882 = pi0223 & ~n33866;
  assign n33883 = ~n33881 & n33882;
  assign n33884 = ~n33843 & ~n33883;
  assign n33885 = ~pi0299 & ~n33884;
  assign n33886 = n3448 & n33795;
  assign n33887 = n6242 & n33822;
  assign n33888 = ~n6242 & ~n33838;
  assign n33889 = ~n3448 & ~n33888;
  assign n33890 = ~n33887 & n33889;
  assign n33891 = ~pi0215 & ~n33886;
  assign n33892 = ~n33890 & n33891;
  assign n33893 = ~n6242 & n33865;
  assign n33894 = n6242 & n33880;
  assign n33895 = pi0215 & ~n33893;
  assign n33896 = ~n33894 & n33895;
  assign n33897 = ~n33892 & ~n33896;
  assign n33898 = pi0299 & ~n33897;
  assign n33899 = pi0039 & ~n33885;
  assign n33900 = ~n33898 & n33899;
  assign n33901 = ~n33793 & ~n33900;
  assign n33902 = ~pi0038 & ~n33901;
  assign n33903 = n2571 & ~n33756;
  assign n33904 = ~n33902 & n33903;
  assign n33905 = ~n33420 & ~n33904;
  assign n33906 = ~pi0625 & n33905;
  assign n33907 = pi0625 & n33679;
  assign n33908 = ~pi1153 & ~n33907;
  assign n33909 = ~n33906 & n33908;
  assign n33910 = ~pi0608 & ~n33537;
  assign n33911 = ~n33909 & n33910;
  assign n33912 = ~pi0625 & n33679;
  assign n33913 = pi0625 & n33905;
  assign n33914 = pi1153 & ~n33912;
  assign n33915 = ~n33913 & n33914;
  assign n33916 = pi0608 & ~n33541;
  assign n33917 = ~n33915 & n33916;
  assign n33918 = ~n33911 & ~n33917;
  assign n33919 = pi0778 & ~n33918;
  assign n33920 = ~pi0778 & n33905;
  assign n33921 = ~n33919 & ~n33920;
  assign n33922 = ~pi0609 & ~n33921;
  assign n33923 = ~pi1155 & ~n33752;
  assign n33924 = ~n33922 & n33923;
  assign n33925 = ~pi0660 & ~n33687;
  assign n33926 = ~n33924 & n33925;
  assign n33927 = ~pi0609 & n33544;
  assign n33928 = pi0609 & ~n33921;
  assign n33929 = pi1155 & ~n33927;
  assign n33930 = ~n33928 & n33929;
  assign n33931 = pi0660 & ~n33691;
  assign n33932 = ~n33930 & n33931;
  assign n33933 = ~n33926 & ~n33932;
  assign n33934 = pi0785 & ~n33933;
  assign n33935 = ~pi0785 & ~n33921;
  assign n33936 = ~n33934 & ~n33935;
  assign n33937 = ~pi0618 & ~n33936;
  assign n33938 = pi0618 & ~n33547;
  assign n33939 = ~pi1154 & ~n33938;
  assign n33940 = ~n33937 & n33939;
  assign n33941 = ~pi0627 & ~n33699;
  assign n33942 = ~n33940 & n33941;
  assign n33943 = pi0618 & ~n33936;
  assign n33944 = ~pi0618 & ~n33547;
  assign n33945 = pi1154 & ~n33944;
  assign n33946 = ~n33943 & n33945;
  assign n33947 = pi0627 & ~n33703;
  assign n33948 = ~n33946 & n33947;
  assign n33949 = ~n33942 & ~n33948;
  assign n33950 = pi0781 & ~n33949;
  assign n33951 = ~pi0781 & ~n33936;
  assign n33952 = ~n33950 & ~n33951;
  assign n33953 = ~pi0789 & n33952;
  assign n33954 = ~pi0619 & ~n33952;
  assign n33955 = pi0619 & n33549;
  assign n33956 = ~pi1159 & ~n33955;
  assign n33957 = ~n33954 & n33956;
  assign n33958 = ~pi0648 & ~n33711;
  assign n33959 = ~n33957 & n33958;
  assign n33960 = ~pi0619 & n33549;
  assign n33961 = pi0619 & ~n33952;
  assign n33962 = pi1159 & ~n33960;
  assign n33963 = ~n33961 & n33962;
  assign n33964 = pi0648 & ~n33715;
  assign n33965 = ~n33963 & n33964;
  assign n33966 = pi0789 & ~n33959;
  assign n33967 = ~n33965 & n33966;
  assign n33968 = n17970 & ~n33953;
  assign n33969 = ~n33967 & n33968;
  assign n33970 = ~n33751 & ~n33969;
  assign n33971 = ~n33737 & ~n33970;
  assign n33972 = n20364 & n33736;
  assign n33973 = ~n20206 & ~n33972;
  assign n33974 = ~n33971 & n33973;
  assign n33975 = ~n33731 & ~n33974;
  assign n33976 = ~pi0790 & ~n33975;
  assign n33977 = ~pi0787 & ~n33564;
  assign n33978 = pi1157 & ~n33727;
  assign n33979 = ~n33568 & ~n33978;
  assign n33980 = pi0787 & ~n33979;
  assign n33981 = ~n33977 & ~n33980;
  assign n33982 = ~pi0644 & n33981;
  assign n33983 = pi0644 & n33975;
  assign n33984 = pi0715 & ~n33982;
  assign n33985 = ~n33983 & n33984;
  assign n33986 = ~n17804 & n33723;
  assign n33987 = n17804 & n33417;
  assign n33988 = ~n33986 & ~n33987;
  assign n33989 = pi0644 & ~n33988;
  assign n33990 = ~pi0644 & n33417;
  assign n33991 = ~pi0715 & ~n33990;
  assign n33992 = ~n33989 & n33991;
  assign n33993 = pi1160 & ~n33992;
  assign n33994 = ~n33985 & n33993;
  assign n33995 = ~pi0644 & ~n33988;
  assign n33996 = pi0644 & n33417;
  assign n33997 = pi0715 & ~n33996;
  assign n33998 = ~n33995 & n33997;
  assign n33999 = pi0644 & n33981;
  assign n34000 = ~pi0644 & n33975;
  assign n34001 = ~pi0715 & ~n33999;
  assign n34002 = ~n34000 & n34001;
  assign n34003 = ~pi1160 & ~n33998;
  assign n34004 = ~n34002 & n34003;
  assign n34005 = pi0790 & ~n33994;
  assign n34006 = ~n34004 & n34005;
  assign n34007 = ~n33976 & ~n34006;
  assign n34008 = ~po1038 & ~n34007;
  assign n34009 = pi0198 & po1038;
  assign po0355 = n34008 | n34009;
  assign n34011 = pi0199 & ~n17059;
  assign n34012 = ~pi0619 & ~n34011;
  assign n34013 = ~pi0617 & ~n34011;
  assign n34014 = ~pi0199 & ~n19432;
  assign n34015 = n19438 & ~n34014;
  assign n34016 = ~pi0199 & ~n17275;
  assign n34017 = pi0199 & n17221;
  assign n34018 = ~pi0038 & ~n34016;
  assign n34019 = ~n34017 & n34018;
  assign n34020 = ~n34015 & ~n34019;
  assign n34021 = n2571 & ~n34020;
  assign n34022 = pi0199 & ~n2571;
  assign n34023 = pi0617 & ~n34022;
  assign n34024 = ~n34021 & n34023;
  assign n34025 = ~n34013 & ~n34024;
  assign n34026 = ~n17117 & ~n34025;
  assign n34027 = n17117 & ~n34011;
  assign n34028 = ~n34026 & ~n34027;
  assign n34029 = ~pi0785 & n34028;
  assign n34030 = ~pi0609 & ~n34011;
  assign n34031 = pi0609 & ~n34028;
  assign n34032 = pi1155 & ~n34030;
  assign n34033 = ~n34031 & n34032;
  assign n34034 = ~pi0609 & ~n34028;
  assign n34035 = pi0609 & ~n34011;
  assign n34036 = ~pi1155 & ~n34035;
  assign n34037 = ~n34034 & n34036;
  assign n34038 = ~n34033 & ~n34037;
  assign n34039 = pi0785 & ~n34038;
  assign n34040 = ~n34029 & ~n34039;
  assign n34041 = ~pi0781 & ~n34040;
  assign n34042 = ~pi0618 & ~n34011;
  assign n34043 = pi0618 & n34040;
  assign n34044 = pi1154 & ~n34042;
  assign n34045 = ~n34043 & n34044;
  assign n34046 = pi0618 & ~n34011;
  assign n34047 = ~pi0618 & n34040;
  assign n34048 = ~pi1154 & ~n34046;
  assign n34049 = ~n34047 & n34048;
  assign n34050 = ~n34045 & ~n34049;
  assign n34051 = pi0781 & ~n34050;
  assign n34052 = ~n34041 & ~n34051;
  assign n34053 = pi0619 & n34052;
  assign n34054 = pi1159 & ~n34012;
  assign n34055 = ~n34053 & n34054;
  assign n34056 = ~pi0625 & ~n34011;
  assign n34057 = ~pi0637 & ~n34011;
  assign n34058 = ~pi0199 & ~n16641;
  assign n34059 = n19899 & ~n34058;
  assign n34060 = pi0199 & ~n16840;
  assign n34061 = ~pi0199 & ~n16749;
  assign n34062 = pi0039 & ~n34061;
  assign n34063 = ~n34060 & n34062;
  assign n34064 = pi0199 & ~n16948;
  assign n34065 = ~pi0199 & n16926;
  assign n34066 = ~pi0039 & ~n34064;
  assign n34067 = ~n34065 & n34066;
  assign n34068 = ~pi0038 & ~n34067;
  assign n34069 = ~n34063 & n34068;
  assign n34070 = ~n34059 & ~n34069;
  assign n34071 = n2571 & ~n34070;
  assign n34072 = pi0637 & ~n34022;
  assign n34073 = ~n34071 & n34072;
  assign n34074 = ~n34057 & ~n34073;
  assign n34075 = pi0625 & ~n34074;
  assign n34076 = pi1153 & ~n34056;
  assign n34077 = ~n34075 & n34076;
  assign n34078 = ~pi0637 & n34025;
  assign n34079 = pi0199 & n19476;
  assign n34080 = n2571 & ~n24549;
  assign n34081 = ~pi0199 & ~n34080;
  assign n34082 = ~pi0617 & ~n19472;
  assign n34083 = ~n34081 & n34082;
  assign n34084 = ~n34079 & n34083;
  assign n34085 = n2571 & n19496;
  assign n34086 = ~pi0199 & ~n34085;
  assign n34087 = pi0199 & n19488;
  assign n34088 = pi0617 & ~n34087;
  assign n34089 = ~n34086 & n34088;
  assign n34090 = ~n34022 & ~n34089;
  assign n34091 = ~n34084 & n34090;
  assign n34092 = pi0637 & ~n34091;
  assign n34093 = ~n34078 & ~n34092;
  assign n34094 = ~pi0625 & n34093;
  assign n34095 = pi0625 & ~n34025;
  assign n34096 = ~pi1153 & ~n34095;
  assign n34097 = ~n34094 & n34096;
  assign n34098 = ~pi0608 & ~n34077;
  assign n34099 = ~n34097 & n34098;
  assign n34100 = ~pi0625 & ~n34074;
  assign n34101 = pi0625 & ~n34011;
  assign n34102 = ~pi1153 & ~n34101;
  assign n34103 = ~n34100 & n34102;
  assign n34104 = pi0625 & n34093;
  assign n34105 = ~pi0625 & ~n34025;
  assign n34106 = pi1153 & ~n34105;
  assign n34107 = ~n34104 & n34106;
  assign n34108 = pi0608 & ~n34103;
  assign n34109 = ~n34107 & n34108;
  assign n34110 = ~n34099 & ~n34109;
  assign n34111 = pi0778 & ~n34110;
  assign n34112 = ~pi0778 & n34093;
  assign n34113 = ~n34111 & ~n34112;
  assign n34114 = ~pi0609 & ~n34113;
  assign n34115 = ~pi0778 & n34074;
  assign n34116 = ~n34077 & ~n34103;
  assign n34117 = pi0778 & ~n34116;
  assign n34118 = ~n34115 & ~n34117;
  assign n34119 = pi0609 & n34118;
  assign n34120 = ~pi1155 & ~n34119;
  assign n34121 = ~n34114 & n34120;
  assign n34122 = ~pi0660 & ~n34033;
  assign n34123 = ~n34121 & n34122;
  assign n34124 = ~pi0609 & n34118;
  assign n34125 = pi0609 & ~n34113;
  assign n34126 = pi1155 & ~n34124;
  assign n34127 = ~n34125 & n34126;
  assign n34128 = pi0660 & ~n34037;
  assign n34129 = ~n34127 & n34128;
  assign n34130 = ~n34123 & ~n34129;
  assign n34131 = pi0785 & ~n34130;
  assign n34132 = ~pi0785 & ~n34113;
  assign n34133 = ~n34131 & ~n34132;
  assign n34134 = ~pi0618 & ~n34133;
  assign n34135 = n17075 & ~n34011;
  assign n34136 = ~n17075 & n34118;
  assign n34137 = ~n34135 & ~n34136;
  assign n34138 = pi0618 & ~n34137;
  assign n34139 = ~pi1154 & ~n34138;
  assign n34140 = ~n34134 & n34139;
  assign n34141 = ~pi0627 & ~n34045;
  assign n34142 = ~n34140 & n34141;
  assign n34143 = pi0618 & ~n34133;
  assign n34144 = ~pi0618 & ~n34137;
  assign n34145 = pi1154 & ~n34144;
  assign n34146 = ~n34143 & n34145;
  assign n34147 = pi0627 & ~n34049;
  assign n34148 = ~n34146 & n34147;
  assign n34149 = ~n34142 & ~n34148;
  assign n34150 = pi0781 & ~n34149;
  assign n34151 = ~pi0781 & ~n34133;
  assign n34152 = ~n34150 & ~n34151;
  assign n34153 = ~pi0619 & ~n34152;
  assign n34154 = ~n16639 & n34137;
  assign n34155 = n16639 & n34011;
  assign n34156 = ~n34154 & ~n34155;
  assign n34157 = pi0619 & n34156;
  assign n34158 = ~pi1159 & ~n34157;
  assign n34159 = ~n34153 & n34158;
  assign n34160 = ~pi0648 & ~n34055;
  assign n34161 = ~n34159 & n34160;
  assign n34162 = pi0619 & ~n34011;
  assign n34163 = ~pi0619 & n34052;
  assign n34164 = ~pi1159 & ~n34162;
  assign n34165 = ~n34163 & n34164;
  assign n34166 = ~pi0619 & n34156;
  assign n34167 = pi0619 & ~n34152;
  assign n34168 = pi1159 & ~n34166;
  assign n34169 = ~n34167 & n34168;
  assign n34170 = pi0648 & ~n34165;
  assign n34171 = ~n34169 & n34170;
  assign n34172 = ~n34161 & ~n34171;
  assign n34173 = pi0789 & ~n34172;
  assign n34174 = ~pi0789 & ~n34152;
  assign n34175 = ~n34173 & ~n34174;
  assign n34176 = ~pi0788 & n34175;
  assign n34177 = ~pi0626 & n34175;
  assign n34178 = n16635 & ~n34011;
  assign n34179 = ~n16635 & n34156;
  assign n34180 = ~n34178 & ~n34179;
  assign n34181 = pi0626 & n34180;
  assign n34182 = ~pi0641 & ~n34181;
  assign n34183 = ~n34177 & n34182;
  assign n34184 = ~pi0789 & ~n34052;
  assign n34185 = ~n34055 & ~n34165;
  assign n34186 = pi0789 & ~n34185;
  assign n34187 = ~n34184 & ~n34186;
  assign n34188 = ~pi0626 & ~n34187;
  assign n34189 = pi0626 & n34011;
  assign n34190 = pi0641 & ~n34189;
  assign n34191 = ~n34188 & n34190;
  assign n34192 = ~pi1158 & ~n34191;
  assign n34193 = ~n34183 & n34192;
  assign n34194 = ~pi0626 & n34180;
  assign n34195 = pi0626 & n34175;
  assign n34196 = pi0641 & ~n34194;
  assign n34197 = ~n34195 & n34196;
  assign n34198 = pi0626 & ~n34187;
  assign n34199 = ~pi0626 & n34011;
  assign n34200 = ~pi0641 & ~n34199;
  assign n34201 = ~n34198 & n34200;
  assign n34202 = pi1158 & ~n34201;
  assign n34203 = ~n34197 & n34202;
  assign n34204 = ~n34193 & ~n34203;
  assign n34205 = pi0788 & ~n34204;
  assign n34206 = ~n34176 & ~n34205;
  assign n34207 = ~pi0628 & n34206;
  assign n34208 = ~n17969 & ~n34187;
  assign n34209 = n17969 & n34011;
  assign n34210 = ~n34208 & ~n34209;
  assign n34211 = pi0628 & n34210;
  assign n34212 = ~pi1156 & ~n34211;
  assign n34213 = ~n34207 & n34212;
  assign n34214 = ~pi0628 & ~n34011;
  assign n34215 = ~n16631 & n34180;
  assign n34216 = n16631 & n34011;
  assign n34217 = ~n34215 & ~n34216;
  assign n34218 = pi0628 & n34217;
  assign n34219 = pi1156 & ~n34214;
  assign n34220 = ~n34218 & n34219;
  assign n34221 = ~pi0629 & ~n34220;
  assign n34222 = ~n34213 & n34221;
  assign n34223 = pi0628 & n34206;
  assign n34224 = ~pi0628 & n34210;
  assign n34225 = pi1156 & ~n34224;
  assign n34226 = ~n34223 & n34225;
  assign n34227 = pi0628 & ~n34011;
  assign n34228 = ~pi0628 & n34217;
  assign n34229 = ~pi1156 & ~n34227;
  assign n34230 = ~n34228 & n34229;
  assign n34231 = pi0629 & ~n34230;
  assign n34232 = ~n34226 & n34231;
  assign n34233 = ~n34222 & ~n34232;
  assign n34234 = pi0792 & ~n34233;
  assign n34235 = ~pi0792 & n34206;
  assign n34236 = ~n34234 & ~n34235;
  assign n34237 = ~pi0647 & ~n34236;
  assign n34238 = ~n17779 & ~n34210;
  assign n34239 = n17779 & n34011;
  assign n34240 = ~n34238 & ~n34239;
  assign n34241 = pi0647 & n34240;
  assign n34242 = ~pi1157 & ~n34241;
  assign n34243 = ~n34237 & n34242;
  assign n34244 = ~pi0647 & ~n34011;
  assign n34245 = ~pi0792 & ~n34217;
  assign n34246 = ~n34220 & ~n34230;
  assign n34247 = pi0792 & ~n34246;
  assign n34248 = ~n34245 & ~n34247;
  assign n34249 = pi0647 & n34248;
  assign n34250 = pi1157 & ~n34244;
  assign n34251 = ~n34249 & n34250;
  assign n34252 = ~pi0630 & ~n34251;
  assign n34253 = ~n34243 & n34252;
  assign n34254 = pi0647 & ~n34236;
  assign n34255 = ~pi0647 & n34240;
  assign n34256 = pi1157 & ~n34255;
  assign n34257 = ~n34254 & n34256;
  assign n34258 = pi0647 & ~n34011;
  assign n34259 = ~pi0647 & n34248;
  assign n34260 = ~pi1157 & ~n34258;
  assign n34261 = ~n34259 & n34260;
  assign n34262 = pi0630 & ~n34261;
  assign n34263 = ~n34257 & n34262;
  assign n34264 = ~n34253 & ~n34263;
  assign n34265 = pi0787 & ~n34264;
  assign n34266 = ~pi0787 & ~n34236;
  assign n34267 = ~n34265 & ~n34266;
  assign n34268 = ~pi0790 & n34267;
  assign n34269 = ~pi0787 & ~n34248;
  assign n34270 = ~n34251 & ~n34261;
  assign n34271 = pi0787 & ~n34270;
  assign n34272 = ~n34269 & ~n34271;
  assign n34273 = ~pi0644 & n34272;
  assign n34274 = pi0644 & ~n34267;
  assign n34275 = pi0715 & ~n34273;
  assign n34276 = ~n34274 & n34275;
  assign n34277 = n17804 & ~n34011;
  assign n34278 = ~n17804 & n34240;
  assign n34279 = ~n34277 & ~n34278;
  assign n34280 = pi0644 & ~n34279;
  assign n34281 = ~pi0644 & ~n34011;
  assign n34282 = ~pi0715 & ~n34281;
  assign n34283 = ~n34280 & n34282;
  assign n34284 = pi1160 & ~n34283;
  assign n34285 = ~n34276 & n34284;
  assign n34286 = ~pi0644 & ~n34267;
  assign n34287 = pi0644 & n34272;
  assign n34288 = ~pi0715 & ~n34287;
  assign n34289 = ~n34286 & n34288;
  assign n34290 = ~pi0644 & ~n34279;
  assign n34291 = pi0644 & ~n34011;
  assign n34292 = pi0715 & ~n34291;
  assign n34293 = ~n34290 & n34292;
  assign n34294 = ~pi1160 & ~n34293;
  assign n34295 = ~n34289 & n34294;
  assign n34296 = pi0790 & ~n34285;
  assign n34297 = ~n34295 & n34296;
  assign n34298 = ~n34268 & ~n34297;
  assign n34299 = ~po1038 & ~n34298;
  assign n34300 = pi0199 & po1038;
  assign po0356 = n34299 | n34300;
  assign n34302 = pi0200 & ~n17059;
  assign n34303 = ~pi0606 & ~n34302;
  assign n34304 = pi0200 & ~n2571;
  assign n34305 = ~pi0200 & ~n19432;
  assign n34306 = n19438 & ~n34305;
  assign n34307 = ~pi0200 & ~n17275;
  assign n34308 = pi0200 & n17221;
  assign n34309 = ~pi0038 & ~n34307;
  assign n34310 = ~n34308 & n34309;
  assign n34311 = ~n34306 & ~n34310;
  assign n34312 = n2571 & ~n34311;
  assign n34313 = pi0606 & ~n34304;
  assign n34314 = ~n34312 & n34313;
  assign n34315 = ~n34303 & ~n34314;
  assign n34316 = ~n17117 & ~n34315;
  assign n34317 = n17117 & ~n34302;
  assign n34318 = ~n34316 & ~n34317;
  assign n34319 = ~pi0785 & n34318;
  assign n34320 = ~pi0609 & ~n34302;
  assign n34321 = pi0609 & ~n34318;
  assign n34322 = pi1155 & ~n34320;
  assign n34323 = ~n34321 & n34322;
  assign n34324 = ~pi0609 & ~n34318;
  assign n34325 = pi0609 & ~n34302;
  assign n34326 = ~pi1155 & ~n34325;
  assign n34327 = ~n34324 & n34326;
  assign n34328 = ~n34323 & ~n34327;
  assign n34329 = pi0785 & ~n34328;
  assign n34330 = ~n34319 & ~n34329;
  assign n34331 = ~pi0781 & ~n34330;
  assign n34332 = ~pi0618 & ~n34302;
  assign n34333 = pi0618 & n34330;
  assign n34334 = pi1154 & ~n34332;
  assign n34335 = ~n34333 & n34334;
  assign n34336 = pi0618 & ~n34302;
  assign n34337 = ~pi0618 & n34330;
  assign n34338 = ~pi1154 & ~n34336;
  assign n34339 = ~n34337 & n34338;
  assign n34340 = ~n34335 & ~n34339;
  assign n34341 = pi0781 & ~n34340;
  assign n34342 = ~n34331 & ~n34341;
  assign n34343 = ~pi0789 & ~n34342;
  assign n34344 = ~pi0619 & ~n34302;
  assign n34345 = pi0619 & n34342;
  assign n34346 = pi1159 & ~n34344;
  assign n34347 = ~n34345 & n34346;
  assign n34348 = pi0619 & ~n34302;
  assign n34349 = ~pi0619 & n34342;
  assign n34350 = ~pi1159 & ~n34348;
  assign n34351 = ~n34349 & n34350;
  assign n34352 = ~n34347 & ~n34351;
  assign n34353 = pi0789 & ~n34352;
  assign n34354 = ~n34343 & ~n34353;
  assign n34355 = ~n17969 & ~n34354;
  assign n34356 = n17969 & n34302;
  assign n34357 = ~n34355 & ~n34356;
  assign n34358 = ~n17779 & ~n34357;
  assign n34359 = n17779 & n34302;
  assign n34360 = ~n34358 & ~n34359;
  assign n34361 = ~n17804 & ~n34360;
  assign n34362 = n17804 & n34302;
  assign n34363 = ~n34361 & ~n34362;
  assign n34364 = ~pi0644 & n34363;
  assign n34365 = pi0644 & ~n34302;
  assign n34366 = pi0715 & ~n34365;
  assign n34367 = ~n34364 & n34366;
  assign n34368 = n16635 & ~n34302;
  assign n34369 = n17075 & ~n34302;
  assign n34370 = ~pi0643 & ~n34302;
  assign n34371 = ~pi0200 & ~n16641;
  assign n34372 = n19899 & ~n34371;
  assign n34373 = ~pi0200 & n16733;
  assign n34374 = pi0200 & n16823;
  assign n34375 = ~pi0299 & ~n34373;
  assign n34376 = ~n34374 & n34375;
  assign n34377 = ~pi0200 & n16747;
  assign n34378 = pi0200 & n16838;
  assign n34379 = pi0299 & ~n34377;
  assign n34380 = ~n34378 & n34379;
  assign n34381 = ~n34376 & ~n34380;
  assign n34382 = pi0039 & ~n34381;
  assign n34383 = ~pi0200 & ~n16926;
  assign n34384 = pi0200 & n16948;
  assign n34385 = ~pi0039 & ~n34383;
  assign n34386 = ~n34384 & n34385;
  assign n34387 = ~n34382 & ~n34386;
  assign n34388 = ~pi0038 & ~n34387;
  assign n34389 = ~n34372 & ~n34388;
  assign n34390 = n2571 & ~n34389;
  assign n34391 = pi0643 & ~n34304;
  assign n34392 = ~n34390 & n34391;
  assign n34393 = ~n34370 & ~n34392;
  assign n34394 = ~pi0778 & n34393;
  assign n34395 = ~pi0625 & ~n34302;
  assign n34396 = pi0625 & ~n34393;
  assign n34397 = pi1153 & ~n34395;
  assign n34398 = ~n34396 & n34397;
  assign n34399 = ~pi0625 & ~n34393;
  assign n34400 = pi0625 & ~n34302;
  assign n34401 = ~pi1153 & ~n34400;
  assign n34402 = ~n34399 & n34401;
  assign n34403 = ~n34398 & ~n34402;
  assign n34404 = pi0778 & ~n34403;
  assign n34405 = ~n34394 & ~n34404;
  assign n34406 = ~n17075 & n34405;
  assign n34407 = ~n34369 & ~n34406;
  assign n34408 = ~n16639 & n34407;
  assign n34409 = n16639 & n34302;
  assign n34410 = ~n34408 & ~n34409;
  assign n34411 = ~n16635 & n34410;
  assign n34412 = ~n34368 & ~n34411;
  assign n34413 = ~n16631 & n34412;
  assign n34414 = n16631 & n34302;
  assign n34415 = ~n34413 & ~n34414;
  assign n34416 = ~pi0792 & ~n34415;
  assign n34417 = pi0628 & ~n34302;
  assign n34418 = ~pi0628 & n34415;
  assign n34419 = ~pi1156 & ~n34417;
  assign n34420 = ~n34418 & n34419;
  assign n34421 = ~pi0628 & ~n34302;
  assign n34422 = pi0628 & n34415;
  assign n34423 = pi1156 & ~n34421;
  assign n34424 = ~n34422 & n34423;
  assign n34425 = ~n34420 & ~n34424;
  assign n34426 = pi0792 & ~n34425;
  assign n34427 = ~n34416 & ~n34426;
  assign n34428 = ~pi0787 & ~n34427;
  assign n34429 = pi0647 & ~n34427;
  assign n34430 = ~pi0647 & n34302;
  assign n34431 = ~n34429 & ~n34430;
  assign n34432 = pi1157 & ~n34431;
  assign n34433 = pi0647 & ~n34302;
  assign n34434 = ~pi0647 & n34427;
  assign n34435 = ~pi1157 & ~n34433;
  assign n34436 = ~n34434 & n34435;
  assign n34437 = ~n34432 & ~n34436;
  assign n34438 = pi0787 & ~n34437;
  assign n34439 = ~n34428 & ~n34438;
  assign n34440 = pi0644 & n34439;
  assign n34441 = ~pi0629 & n34424;
  assign n34442 = ~n20570 & ~n34357;
  assign n34443 = pi0629 & n34420;
  assign n34444 = ~n34441 & ~n34443;
  assign n34445 = ~n34442 & n34444;
  assign n34446 = pi0792 & ~n34445;
  assign n34447 = pi0609 & n34405;
  assign n34448 = ~pi0643 & n34315;
  assign n34449 = ~n19491 & ~n19492;
  assign n34450 = ~pi0200 & ~n34449;
  assign n34451 = pi0038 & pi0200;
  assign n34452 = n19485 & n34451;
  assign n34453 = ~pi0200 & ~n19493;
  assign n34454 = pi0200 & ~n24754;
  assign n34455 = ~pi0038 & ~n34453;
  assign n34456 = ~n34454 & n34455;
  assign n34457 = pi0606 & n2571;
  assign n34458 = ~n34452 & n34457;
  assign n34459 = ~n34450 & n34458;
  assign n34460 = ~n34456 & n34459;
  assign n34461 = ~n16647 & ~n17355;
  assign n34462 = n34372 & ~n34461;
  assign n34463 = ~pi0200 & ~n19467;
  assign n34464 = pi0200 & ~n19475;
  assign n34465 = ~pi0038 & ~n34463;
  assign n34466 = ~n34464 & n34465;
  assign n34467 = ~n34462 & ~n34466;
  assign n34468 = ~pi0606 & n2571;
  assign n34469 = ~n34467 & n34468;
  assign n34470 = ~n34304 & ~n34460;
  assign n34471 = ~n34469 & n34470;
  assign n34472 = pi0643 & ~n34471;
  assign n34473 = ~n34448 & ~n34472;
  assign n34474 = ~pi0625 & n34473;
  assign n34475 = pi0625 & ~n34315;
  assign n34476 = ~pi1153 & ~n34475;
  assign n34477 = ~n34474 & n34476;
  assign n34478 = ~pi0608 & ~n34398;
  assign n34479 = ~n34477 & n34478;
  assign n34480 = pi0625 & n34473;
  assign n34481 = ~pi0625 & ~n34315;
  assign n34482 = pi1153 & ~n34481;
  assign n34483 = ~n34480 & n34482;
  assign n34484 = pi0608 & ~n34402;
  assign n34485 = ~n34483 & n34484;
  assign n34486 = ~n34479 & ~n34485;
  assign n34487 = pi0778 & ~n34486;
  assign n34488 = ~pi0778 & n34473;
  assign n34489 = ~n34487 & ~n34488;
  assign n34490 = ~pi0609 & ~n34489;
  assign n34491 = ~pi1155 & ~n34447;
  assign n34492 = ~n34490 & n34491;
  assign n34493 = ~pi0660 & ~n34323;
  assign n34494 = ~n34492 & n34493;
  assign n34495 = ~pi0609 & n34405;
  assign n34496 = pi0609 & ~n34489;
  assign n34497 = pi1155 & ~n34495;
  assign n34498 = ~n34496 & n34497;
  assign n34499 = pi0660 & ~n34327;
  assign n34500 = ~n34498 & n34499;
  assign n34501 = ~n34494 & ~n34500;
  assign n34502 = pi0785 & ~n34501;
  assign n34503 = ~pi0785 & ~n34489;
  assign n34504 = ~n34502 & ~n34503;
  assign n34505 = ~pi0618 & ~n34504;
  assign n34506 = pi0618 & ~n34407;
  assign n34507 = ~pi1154 & ~n34506;
  assign n34508 = ~n34505 & n34507;
  assign n34509 = ~pi0627 & ~n34335;
  assign n34510 = ~n34508 & n34509;
  assign n34511 = pi0618 & ~n34504;
  assign n34512 = ~pi0618 & ~n34407;
  assign n34513 = pi1154 & ~n34512;
  assign n34514 = ~n34511 & n34513;
  assign n34515 = pi0627 & ~n34339;
  assign n34516 = ~n34514 & n34515;
  assign n34517 = ~n34510 & ~n34516;
  assign n34518 = pi0781 & ~n34517;
  assign n34519 = ~pi0781 & ~n34504;
  assign n34520 = ~n34518 & ~n34519;
  assign n34521 = ~pi0789 & n34520;
  assign n34522 = ~pi0619 & ~n34520;
  assign n34523 = pi0619 & n34410;
  assign n34524 = ~pi1159 & ~n34523;
  assign n34525 = ~n34522 & n34524;
  assign n34526 = ~pi0648 & ~n34347;
  assign n34527 = ~n34525 & n34526;
  assign n34528 = pi0619 & ~n34520;
  assign n34529 = ~pi0619 & n34410;
  assign n34530 = pi1159 & ~n34529;
  assign n34531 = ~n34528 & n34530;
  assign n34532 = pi0648 & ~n34351;
  assign n34533 = ~n34531 & n34532;
  assign n34534 = pi0789 & ~n34527;
  assign n34535 = ~n34533 & n34534;
  assign n34536 = n17970 & ~n34521;
  assign n34537 = ~n34535 & n34536;
  assign n34538 = n17871 & ~n34412;
  assign n34539 = pi0626 & n34302;
  assign n34540 = ~pi0626 & ~n34354;
  assign n34541 = n16629 & ~n34539;
  assign n34542 = ~n34540 & n34541;
  assign n34543 = ~pi0626 & n34302;
  assign n34544 = pi0626 & ~n34354;
  assign n34545 = n16628 & ~n34543;
  assign n34546 = ~n34544 & n34545;
  assign n34547 = ~n34538 & ~n34542;
  assign n34548 = ~n34546 & n34547;
  assign n34549 = pi0788 & ~n34548;
  assign n34550 = ~n20364 & ~n34549;
  assign n34551 = ~n34537 & n34550;
  assign n34552 = ~n34446 & ~n34551;
  assign n34553 = ~n20206 & ~n34552;
  assign n34554 = pi0630 & n34436;
  assign n34555 = ~n20559 & ~n34360;
  assign n34556 = n17801 & ~n34431;
  assign n34557 = ~n34554 & ~n34555;
  assign n34558 = ~n34556 & n34557;
  assign n34559 = pi0787 & ~n34558;
  assign n34560 = ~n34553 & ~n34559;
  assign n34561 = ~pi0644 & n34560;
  assign n34562 = ~pi0715 & ~n34440;
  assign n34563 = ~n34561 & n34562;
  assign n34564 = ~pi1160 & ~n34367;
  assign n34565 = ~n34563 & n34564;
  assign n34566 = ~pi0644 & n34439;
  assign n34567 = pi0644 & n34560;
  assign n34568 = pi0715 & ~n34566;
  assign n34569 = ~n34567 & n34568;
  assign n34570 = pi0644 & n34363;
  assign n34571 = ~pi0644 & ~n34302;
  assign n34572 = ~pi0715 & ~n34571;
  assign n34573 = ~n34570 & n34572;
  assign n34574 = pi1160 & ~n34573;
  assign n34575 = ~n34569 & n34574;
  assign n34576 = ~n34565 & ~n34575;
  assign n34577 = pi0790 & ~n34576;
  assign n34578 = ~pi0790 & n34560;
  assign n34579 = ~n34577 & ~n34578;
  assign n34580 = ~po1038 & ~n34579;
  assign n34581 = ~pi0200 & po1038;
  assign po0357 = ~n34580 & ~n34581;
  assign n34583 = pi0233 & pi0237;
  assign n34584 = pi0057 & pi0332;
  assign n34585 = n2572 & n6573;
  assign n34586 = n2521 & n34585;
  assign n34587 = ~pi0332 & ~n34586;
  assign n34588 = n6304 & ~n34587;
  assign n34589 = pi0332 & ~n6304;
  assign n34590 = pi0059 & ~n34589;
  assign n34591 = ~n34588 & n34590;
  assign n34592 = pi0332 & ~n2529;
  assign n34593 = ~pi0059 & ~n34592;
  assign n34594 = pi0055 & n34587;
  assign n34595 = pi0074 & pi0332;
  assign n34596 = ~pi0055 & ~n34595;
  assign n34597 = n2726 & n11086;
  assign n34598 = pi0468 & n6192;
  assign n34599 = ~pi0299 & pi0587;
  assign n34600 = ~n21044 & ~n34599;
  assign n34601 = ~pi0468 & ~n34600;
  assign n34602 = ~n34598 & ~n34601;
  assign n34603 = n34597 & ~n34602;
  assign n34604 = ~pi0332 & ~n34603;
  assign n34605 = n7363 & ~n34604;
  assign n34606 = n2521 & n6585;
  assign n34607 = ~pi0332 & ~n34606;
  assign n34608 = n15625 & ~n34607;
  assign n34609 = pi0332 & ~n2611;
  assign n34610 = ~n34608 & ~n34609;
  assign n34611 = ~n34605 & n34610;
  assign n34612 = ~pi0074 & ~n34611;
  assign n34613 = n34596 & ~n34612;
  assign n34614 = n2529 & ~n34594;
  assign n34615 = ~n34613 & n34614;
  assign n34616 = n34593 & ~n34615;
  assign n34617 = ~pi0057 & ~n34591;
  assign n34618 = ~n34616 & n34617;
  assign n34619 = ~n34584 & ~n34618;
  assign n34620 = ~n34583 & ~n34619;
  assign n34621 = ~pi0332 & ~n6192;
  assign n34622 = ~pi0947 & ~n34621;
  assign n34623 = pi0096 & pi0210;
  assign n34624 = pi0332 & n34623;
  assign n34625 = ~pi0032 & pi0070;
  assign n34626 = ~pi0070 & ~pi0841;
  assign n34627 = pi0032 & n34626;
  assign n34628 = ~n34625 & ~n34627;
  assign n34629 = ~pi0210 & ~n34628;
  assign n34630 = ~pi0032 & ~pi0096;
  assign n34631 = pi0070 & n34630;
  assign n34632 = ~pi0332 & ~n34631;
  assign n34633 = ~n34629 & n34632;
  assign n34634 = ~n34624 & ~n34633;
  assign n34635 = ~n6197 & n34634;
  assign n34636 = n6192 & ~n34635;
  assign n34637 = n34622 & ~n34636;
  assign n34638 = n6192 & ~n34634;
  assign n34639 = pi0332 & pi0468;
  assign n34640 = ~pi0468 & ~n34633;
  assign n34641 = ~n34639 & ~n34640;
  assign n34642 = ~n6192 & n34641;
  assign n34643 = pi0947 & ~n34638;
  assign n34644 = ~n34642 & n34643;
  assign n34645 = ~n34637 & ~n34644;
  assign n34646 = pi0057 & ~n34645;
  assign n34647 = ~n6304 & n34645;
  assign n34648 = ~n2572 & n34645;
  assign n34649 = pi0032 & ~n34626;
  assign n34650 = ~pi0095 & n2736;
  assign n34651 = ~n34649 & n34650;
  assign n34652 = n2706 & n34651;
  assign n34653 = n2728 & n34652;
  assign n34654 = n34628 & ~n34653;
  assign n34655 = ~pi0210 & ~n34654;
  assign n34656 = ~pi0095 & n2975;
  assign n34657 = ~pi0070 & ~n34656;
  assign n34658 = n34630 & ~n34657;
  assign n34659 = pi0210 & n34658;
  assign n34660 = ~pi0332 & ~n34655;
  assign n34661 = ~n34659 & n34660;
  assign n34662 = ~n34624 & ~n34661;
  assign n34663 = ~n6197 & n34662;
  assign n34664 = n6192 & ~n34663;
  assign n34665 = n34622 & ~n34664;
  assign n34666 = n6192 & ~n34662;
  assign n34667 = ~pi0468 & ~n34661;
  assign n34668 = ~n34639 & ~n34667;
  assign n34669 = ~n6192 & n34668;
  assign n34670 = pi0947 & ~n34666;
  assign n34671 = ~n34669 & n34670;
  assign n34672 = ~n34665 & ~n34671;
  assign n34673 = n2572 & n34672;
  assign n34674 = ~n34648 & ~n34673;
  assign n34675 = n6304 & ~n34674;
  assign n34676 = pi0059 & ~n34647;
  assign n34677 = ~n34675 & n34676;
  assign n34678 = ~n2529 & n34645;
  assign n34679 = pi0055 & n34674;
  assign n34680 = ~pi0074 & n2611;
  assign n34681 = pi0299 & ~n34645;
  assign n34682 = pi0096 & pi0198;
  assign n34683 = pi0332 & n34682;
  assign n34684 = ~pi0198 & ~n34628;
  assign n34685 = n34632 & ~n34684;
  assign n34686 = ~n34683 & ~n34685;
  assign n34687 = n6192 & ~n34686;
  assign n34688 = n6583 & ~n34685;
  assign n34689 = n34621 & ~n34688;
  assign n34690 = ~pi0299 & ~n6582;
  assign n34691 = ~n34687 & n34690;
  assign n34692 = ~n34689 & n34691;
  assign n34693 = ~n34680 & ~n34692;
  assign n34694 = ~n34681 & n34693;
  assign n34695 = n2726 & n2962;
  assign n34696 = n34651 & n34695;
  assign n34697 = n34628 & ~n34696;
  assign n34698 = ~pi0210 & ~n34697;
  assign n34699 = ~pi0095 & n2517;
  assign n34700 = n34695 & n34699;
  assign n34701 = ~pi0070 & ~n34700;
  assign n34702 = n34630 & ~n34701;
  assign n34703 = pi0210 & n34702;
  assign n34704 = ~pi0332 & ~n34698;
  assign n34705 = ~n34703 & n34704;
  assign n34706 = ~n34624 & ~n34705;
  assign n34707 = ~n6197 & n34706;
  assign n34708 = n6192 & ~n34707;
  assign n34709 = n34622 & ~n34708;
  assign n34710 = n6192 & ~n34706;
  assign n34711 = ~pi0468 & ~n34705;
  assign n34712 = ~n34639 & ~n34711;
  assign n34713 = ~n6192 & n34712;
  assign n34714 = pi0947 & ~n34710;
  assign n34715 = ~n34713 & n34714;
  assign n34716 = pi0299 & ~n34709;
  assign n34717 = ~n34715 & n34716;
  assign n34718 = ~pi0587 & ~n34621;
  assign n34719 = ~pi0198 & ~n34697;
  assign n34720 = pi0198 & n34702;
  assign n34721 = ~pi0332 & ~n34719;
  assign n34722 = ~n34720 & n34721;
  assign n34723 = ~n34683 & ~n34722;
  assign n34724 = ~n6197 & n34723;
  assign n34725 = n6192 & ~n34724;
  assign n34726 = n34718 & ~n34725;
  assign n34727 = n6192 & ~n34723;
  assign n34728 = ~pi0468 & ~n34722;
  assign n34729 = ~n6192 & ~n34639;
  assign n34730 = ~n34728 & n34729;
  assign n34731 = pi0587 & ~n34727;
  assign n34732 = ~n34730 & n34731;
  assign n34733 = ~pi0299 & ~n34726;
  assign n34734 = ~n34732 & n34733;
  assign n34735 = ~n34717 & ~n34734;
  assign n34736 = n7363 & ~n34735;
  assign n34737 = pi0299 & ~n34672;
  assign n34738 = ~pi0198 & ~n34654;
  assign n34739 = pi0198 & n34658;
  assign n34740 = ~pi0332 & ~n34738;
  assign n34741 = ~n34739 & n34740;
  assign n34742 = ~n34683 & ~n34741;
  assign n34743 = ~n6197 & n34742;
  assign n34744 = n6192 & ~n34743;
  assign n34745 = n34718 & ~n34744;
  assign n34746 = n6192 & ~n34742;
  assign n34747 = ~pi0468 & ~n34741;
  assign n34748 = n34729 & ~n34747;
  assign n34749 = pi0587 & ~n34746;
  assign n34750 = ~n34748 & n34749;
  assign n34751 = ~n34745 & ~n34750;
  assign n34752 = ~pi0299 & ~n34751;
  assign n34753 = n15625 & ~n34737;
  assign n34754 = ~n34752 & n34753;
  assign n34755 = ~n34736 & ~n34754;
  assign n34756 = ~pi0074 & ~n34755;
  assign n34757 = ~pi0055 & ~n34694;
  assign n34758 = ~n34756 & n34757;
  assign n34759 = n2529 & ~n34679;
  assign n34760 = ~n34758 & n34759;
  assign n34761 = ~pi0059 & ~n34678;
  assign n34762 = ~n34760 & n34761;
  assign n34763 = ~n34677 & ~n34762;
  assign n34764 = ~pi0057 & ~n34763;
  assign n34765 = ~n34646 & ~n34764;
  assign n34766 = n34583 & ~n34765;
  assign n34767 = ~n34620 & ~n34766;
  assign n34768 = ~pi0201 & ~n34767;
  assign n34769 = ~n6573 & ~n16479;
  assign n34770 = n6583 & n34682;
  assign n34771 = n16479 & ~n34770;
  assign n34772 = ~n16479 & ~n34623;
  assign n34773 = ~n34769 & ~n34771;
  assign n34774 = ~n34772 & n34773;
  assign n34775 = n34583 & n34774;
  assign n34776 = pi0201 & ~n34775;
  assign po0358 = ~n34768 & ~n34776;
  assign n34778 = ~pi0233 & pi0237;
  assign n34779 = ~n34619 & ~n34778;
  assign n34780 = ~n34765 & n34778;
  assign n34781 = ~n34779 & ~n34780;
  assign n34782 = ~pi0202 & ~n34781;
  assign n34783 = n34774 & n34778;
  assign n34784 = pi0202 & ~n34783;
  assign po0359 = ~n34782 & ~n34784;
  assign n34786 = ~pi0233 & ~pi0237;
  assign n34787 = ~n34619 & ~n34786;
  assign n34788 = ~n34765 & n34786;
  assign n34789 = ~n34787 & ~n34788;
  assign n34790 = ~pi0203 & ~n34789;
  assign n34791 = n34774 & n34786;
  assign n34792 = pi0203 & ~n34791;
  assign po0360 = ~n34790 & ~n34792;
  assign n34794 = n2572 & n6310;
  assign n34795 = n2521 & n34794;
  assign n34796 = ~pi0332 & ~n34795;
  assign n34797 = n6304 & ~n34796;
  assign n34798 = n34590 & ~n34797;
  assign n34799 = pi0055 & n34796;
  assign n34800 = ~pi0468 & pi0602;
  assign n34801 = pi0468 & n6195;
  assign n34802 = ~n34800 & ~n34801;
  assign n34803 = ~pi0299 & ~n34802;
  assign n34804 = ~n6324 & ~n34803;
  assign n34805 = n2521 & ~n34804;
  assign n34806 = ~pi0332 & ~n34805;
  assign n34807 = n15625 & ~n34806;
  assign n34808 = ~pi0299 & ~pi0602;
  assign n34809 = pi0299 & ~pi0907;
  assign n34810 = ~pi0468 & ~n34808;
  assign n34811 = ~n34809 & n34810;
  assign n34812 = ~n34801 & ~n34811;
  assign n34813 = n34597 & ~n34812;
  assign n34814 = ~pi0332 & ~n34813;
  assign n34815 = n7363 & ~n34814;
  assign n34816 = ~n34807 & ~n34815;
  assign n34817 = ~pi0074 & ~n34816;
  assign n34818 = n34596 & ~n34609;
  assign n34819 = ~n34817 & n34818;
  assign n34820 = n2529 & ~n34799;
  assign n34821 = ~n34819 & n34820;
  assign n34822 = n34593 & ~n34821;
  assign n34823 = ~pi0057 & ~n34798;
  assign n34824 = ~n34822 & n34823;
  assign n34825 = ~n34584 & ~n34824;
  assign n34826 = ~n34583 & ~n34825;
  assign n34827 = ~pi0332 & ~n6195;
  assign n34828 = ~pi0907 & ~n34827;
  assign n34829 = n6195 & ~n34635;
  assign n34830 = n34828 & ~n34829;
  assign n34831 = n6195 & ~n34634;
  assign n34832 = ~n6195 & n34641;
  assign n34833 = pi0907 & ~n34831;
  assign n34834 = ~n34832 & n34833;
  assign n34835 = ~n34830 & ~n34834;
  assign n34836 = pi0057 & ~n34835;
  assign n34837 = ~n6304 & n34835;
  assign n34838 = ~n2572 & n34835;
  assign n34839 = n6195 & ~n34662;
  assign n34840 = ~n6195 & n34668;
  assign n34841 = pi0907 & ~n34839;
  assign n34842 = ~n34840 & n34841;
  assign n34843 = pi0332 & ~n16657;
  assign n34844 = pi0680 & ~n34843;
  assign n34845 = ~n34663 & n34844;
  assign n34846 = n34828 & ~n34845;
  assign n34847 = ~n34842 & ~n34846;
  assign n34848 = n2572 & n34847;
  assign n34849 = ~n34838 & ~n34848;
  assign n34850 = n6304 & ~n34849;
  assign n34851 = pi0059 & ~n34837;
  assign n34852 = ~n34850 & n34851;
  assign n34853 = ~n2529 & n34835;
  assign n34854 = pi0055 & n34849;
  assign n34855 = pi0299 & n34847;
  assign n34856 = n6195 & n34682;
  assign n34857 = pi0332 & ~n34856;
  assign n34858 = ~pi0299 & ~n34857;
  assign n34859 = n6326 & n34742;
  assign n34860 = n34858 & ~n34859;
  assign n34861 = ~n34855 & ~n34860;
  assign n34862 = n15625 & ~n34861;
  assign n34863 = n6326 & n34723;
  assign n34864 = n34858 & ~n34863;
  assign n34865 = n6195 & ~n34707;
  assign n34866 = n34828 & ~n34865;
  assign n34867 = n6195 & ~n34706;
  assign n34868 = ~n6195 & n34712;
  assign n34869 = pi0907 & ~n34867;
  assign n34870 = ~n34868 & n34869;
  assign n34871 = pi0299 & ~n34866;
  assign n34872 = ~n34870 & n34871;
  assign n34873 = ~n34864 & ~n34872;
  assign n34874 = n7363 & ~n34873;
  assign n34875 = ~n34862 & ~n34874;
  assign n34876 = ~pi0074 & ~n34875;
  assign n34877 = pi0299 & ~n34835;
  assign n34878 = n34686 & ~n34802;
  assign n34879 = ~n34857 & ~n34878;
  assign n34880 = ~pi0299 & ~n34879;
  assign n34881 = ~n34680 & ~n34880;
  assign n34882 = ~n34877 & n34881;
  assign n34883 = ~pi0055 & ~n34882;
  assign n34884 = ~n34876 & n34883;
  assign n34885 = n2529 & ~n34854;
  assign n34886 = ~n34884 & n34885;
  assign n34887 = ~pi0059 & ~n34853;
  assign n34888 = ~n34886 & n34887;
  assign n34889 = ~n34852 & ~n34888;
  assign n34890 = ~pi0057 & ~n34889;
  assign n34891 = ~n34836 & ~n34890;
  assign n34892 = n34583 & ~n34891;
  assign n34893 = ~n34826 & ~n34892;
  assign n34894 = ~pi0204 & ~n34893;
  assign n34895 = ~n6310 & ~n16479;
  assign n34896 = n6326 & n34682;
  assign n34897 = n16479 & ~n34896;
  assign n34898 = ~n34772 & ~n34895;
  assign n34899 = ~n34897 & n34898;
  assign n34900 = n34583 & n34899;
  assign n34901 = pi0204 & ~n34900;
  assign po0361 = ~n34894 & ~n34901;
  assign n34903 = ~n34778 & ~n34825;
  assign n34904 = n34778 & ~n34891;
  assign n34905 = ~n34903 & ~n34904;
  assign n34906 = ~pi0205 & ~n34905;
  assign n34907 = n34778 & n34899;
  assign n34908 = pi0205 & ~n34907;
  assign po0362 = ~n34906 & ~n34908;
  assign n34910 = pi0233 & ~pi0237;
  assign n34911 = ~n34825 & ~n34910;
  assign n34912 = ~n34891 & n34910;
  assign n34913 = ~n34911 & ~n34912;
  assign n34914 = ~pi0206 & ~n34913;
  assign n34915 = n34899 & n34910;
  assign n34916 = pi0206 & ~n34915;
  assign po0363 = ~n34914 & ~n34916;
  assign n34918 = ~n19146 & n24385;
  assign n34919 = n19151 & n34918;
  assign n34920 = ~n19142 & n34919;
  assign n34921 = pi0207 & ~n34920;
  assign n34922 = n16635 & ~n17059;
  assign n34923 = n2571 & n24388;
  assign n34924 = ~pi0778 & ~n34923;
  assign n34925 = ~pi0625 & ~n17059;
  assign n34926 = pi0625 & ~n34923;
  assign n34927 = ~n34925 & ~n34926;
  assign n34928 = pi1153 & ~n34927;
  assign n34929 = pi0625 & ~n17059;
  assign n34930 = ~pi0625 & ~n34923;
  assign n34931 = ~n34929 & ~n34930;
  assign n34932 = ~pi1153 & ~n34931;
  assign n34933 = ~n34928 & ~n34932;
  assign n34934 = pi0778 & ~n34933;
  assign n34935 = ~n34924 & ~n34934;
  assign n34936 = ~n17075 & ~n34935;
  assign n34937 = ~n17059 & n17075;
  assign n34938 = ~n34936 & ~n34937;
  assign n34939 = ~n16639 & n34938;
  assign n34940 = n16639 & n17059;
  assign n34941 = ~n34939 & ~n34940;
  assign n34942 = ~n16635 & n34941;
  assign n34943 = ~n34922 & ~n34942;
  assign n34944 = ~n16631 & n34943;
  assign n34945 = n16631 & n17059;
  assign n34946 = ~n34944 & ~n34945;
  assign n34947 = ~n19142 & ~n34946;
  assign n34948 = n17059 & n17856;
  assign n34949 = ~n34947 & ~n34948;
  assign n34950 = ~pi0207 & ~n34949;
  assign n34951 = ~n34921 & ~n34950;
  assign n34952 = pi0710 & ~n34951;
  assign n34953 = ~pi0207 & ~n17059;
  assign n34954 = ~pi0710 & ~n34953;
  assign n34955 = ~n34952 & ~n34954;
  assign n34956 = ~pi0787 & ~n34955;
  assign n34957 = ~pi0647 & n34955;
  assign n34958 = pi0647 & n34953;
  assign n34959 = ~pi1157 & ~n34958;
  assign n34960 = ~n34957 & n34959;
  assign n34961 = ~pi0647 & n34953;
  assign n34962 = pi0647 & n34955;
  assign n34963 = pi1157 & ~n34961;
  assign n34964 = ~n34962 & n34963;
  assign n34965 = ~n34960 & ~n34964;
  assign n34966 = pi0787 & ~n34965;
  assign n34967 = ~n34956 & ~n34966;
  assign n34968 = ~pi0644 & n34967;
  assign n34969 = ~pi0630 & n34964;
  assign n34970 = ~n17059 & n17117;
  assign n34971 = n2571 & n19439;
  assign n34972 = ~n17117 & ~n34971;
  assign n34973 = ~n34970 & ~n34972;
  assign n34974 = ~pi0785 & ~n34973;
  assign n34975 = ~n17059 & ~n17296;
  assign n34976 = ~pi0609 & n34972;
  assign n34977 = ~n34975 & ~n34976;
  assign n34978 = ~pi1155 & ~n34977;
  assign n34979 = ~n17059 & ~n17291;
  assign n34980 = pi0609 & n34972;
  assign n34981 = ~n34979 & ~n34980;
  assign n34982 = pi1155 & ~n34981;
  assign n34983 = ~n34978 & ~n34982;
  assign n34984 = pi0785 & ~n34983;
  assign n34985 = ~n34974 & ~n34984;
  assign n34986 = ~pi0781 & ~n34985;
  assign n34987 = ~pi0618 & n34985;
  assign n34988 = pi0618 & n17059;
  assign n34989 = ~pi1154 & ~n34988;
  assign n34990 = ~n34987 & n34989;
  assign n34991 = ~pi0618 & n17059;
  assign n34992 = pi0618 & n34985;
  assign n34993 = pi1154 & ~n34991;
  assign n34994 = ~n34992 & n34993;
  assign n34995 = ~n34990 & ~n34994;
  assign n34996 = pi0781 & ~n34995;
  assign n34997 = ~n34986 & ~n34996;
  assign n34998 = ~pi0789 & ~n34997;
  assign n34999 = ~pi0619 & n34997;
  assign n35000 = pi0619 & n17059;
  assign n35001 = ~pi1159 & ~n35000;
  assign n35002 = ~n34999 & n35001;
  assign n35003 = ~pi0619 & n17059;
  assign n35004 = pi0619 & n34997;
  assign n35005 = pi1159 & ~n35003;
  assign n35006 = ~n35004 & n35005;
  assign n35007 = ~n35002 & ~n35006;
  assign n35008 = pi0789 & ~n35007;
  assign n35009 = ~n34998 & ~n35008;
  assign n35010 = ~n17969 & n35009;
  assign n35011 = n17059 & n17969;
  assign n35012 = ~n35010 & ~n35011;
  assign n35013 = ~n17779 & ~n35012;
  assign n35014 = n17059 & n17779;
  assign n35015 = ~n35013 & ~n35014;
  assign n35016 = ~pi0207 & ~n35015;
  assign n35017 = n2571 & ~n24447;
  assign n35018 = ~n17117 & n35017;
  assign n35019 = ~n20225 & n35018;
  assign n35020 = ~n20235 & n35019;
  assign n35021 = ~n20231 & n35020;
  assign n35022 = ~n17969 & n35021;
  assign n35023 = ~n17779 & n35022;
  assign n35024 = pi0207 & ~n35023;
  assign n35025 = pi0623 & ~n35024;
  assign n35026 = ~n35016 & n35025;
  assign n35027 = ~pi0623 & n34953;
  assign n35028 = ~n35026 & ~n35027;
  assign n35029 = ~n20559 & n35028;
  assign n35030 = pi0630 & n34960;
  assign n35031 = ~n34969 & ~n35029;
  assign n35032 = ~n35030 & n35031;
  assign n35033 = pi0787 & ~n35032;
  assign n35034 = ~pi0710 & ~n35028;
  assign n35035 = ~pi0628 & ~n17059;
  assign n35036 = pi0628 & n34946;
  assign n35037 = ~n35035 & ~n35036;
  assign n35038 = ~pi0629 & ~n35037;
  assign n35039 = ~n35035 & ~n35038;
  assign n35040 = pi1156 & ~n35039;
  assign n35041 = pi0628 & ~n17059;
  assign n35042 = ~pi1156 & n35041;
  assign n35043 = ~pi0628 & n34946;
  assign n35044 = ~n35041 & ~n35043;
  assign n35045 = n17777 & ~n35044;
  assign n35046 = ~n35042 & ~n35045;
  assign n35047 = ~n35040 & n35046;
  assign n35048 = pi0792 & ~n35047;
  assign n35049 = pi1159 & ~n17059;
  assign n35050 = pi0619 & n34941;
  assign n35051 = pi1154 & ~n17059;
  assign n35052 = pi0618 & ~n34938;
  assign n35053 = pi1155 & ~n17059;
  assign n35054 = pi0609 & ~n34935;
  assign n35055 = n2571 & ~n19477;
  assign n35056 = ~pi0778 & ~n35055;
  assign n35057 = ~pi0625 & ~n35055;
  assign n35058 = ~n34929 & ~n35057;
  assign n35059 = ~pi1153 & ~n35058;
  assign n35060 = ~pi0608 & ~n34928;
  assign n35061 = ~n35059 & n35060;
  assign n35062 = pi0625 & ~n35055;
  assign n35063 = ~n34925 & ~n35062;
  assign n35064 = pi1153 & ~n35063;
  assign n35065 = pi0608 & ~n34932;
  assign n35066 = ~n35064 & n35065;
  assign n35067 = pi0778 & ~n35061;
  assign n35068 = ~n35066 & n35067;
  assign n35069 = ~n35056 & ~n35068;
  assign n35070 = ~pi0609 & ~n35069;
  assign n35071 = ~n35054 & ~n35070;
  assign n35072 = ~pi1155 & ~n35071;
  assign n35073 = ~pi0660 & ~n35053;
  assign n35074 = ~n35072 & n35073;
  assign n35075 = ~pi1155 & ~n17059;
  assign n35076 = ~pi0609 & ~n34935;
  assign n35077 = pi0609 & ~n35069;
  assign n35078 = ~n35076 & ~n35077;
  assign n35079 = pi1155 & ~n35078;
  assign n35080 = pi0660 & ~n35075;
  assign n35081 = ~n35079 & n35080;
  assign n35082 = ~n35074 & ~n35081;
  assign n35083 = pi0785 & ~n35082;
  assign n35084 = ~pi0785 & n35069;
  assign n35085 = ~n35083 & ~n35084;
  assign n35086 = ~pi0618 & n35085;
  assign n35087 = ~n35052 & ~n35086;
  assign n35088 = ~pi1154 & ~n35087;
  assign n35089 = ~pi0627 & ~n35051;
  assign n35090 = ~n35088 & n35089;
  assign n35091 = ~pi1154 & ~n17059;
  assign n35092 = ~pi0618 & ~n34938;
  assign n35093 = pi0618 & n35085;
  assign n35094 = ~n35092 & ~n35093;
  assign n35095 = pi1154 & ~n35094;
  assign n35096 = pi0627 & ~n35091;
  assign n35097 = ~n35095 & n35096;
  assign n35098 = ~n35090 & ~n35097;
  assign n35099 = pi0781 & ~n35098;
  assign n35100 = ~pi0781 & ~n35085;
  assign n35101 = ~n35099 & ~n35100;
  assign n35102 = ~pi0619 & n35101;
  assign n35103 = ~n35050 & ~n35102;
  assign n35104 = ~pi1159 & ~n35103;
  assign n35105 = ~pi0648 & ~n35049;
  assign n35106 = ~n35104 & n35105;
  assign n35107 = ~pi1159 & ~n17059;
  assign n35108 = ~pi0619 & n34941;
  assign n35109 = pi0619 & n35101;
  assign n35110 = ~n35108 & ~n35109;
  assign n35111 = pi1159 & ~n35110;
  assign n35112 = pi0648 & ~n35107;
  assign n35113 = ~n35111 & n35112;
  assign n35114 = ~n35106 & ~n35113;
  assign n35115 = pi0789 & ~n35114;
  assign n35116 = ~pi0789 & ~n35101;
  assign n35117 = ~n35115 & ~n35116;
  assign n35118 = ~pi0788 & ~n35117;
  assign n35119 = pi0641 & ~n17059;
  assign n35120 = pi0626 & n34943;
  assign n35121 = ~pi0626 & ~n35117;
  assign n35122 = ~pi0641 & ~n35120;
  assign n35123 = ~n35121 & n35122;
  assign n35124 = ~pi1158 & ~n35119;
  assign n35125 = ~n35123 & n35124;
  assign n35126 = ~pi0641 & ~n17059;
  assign n35127 = ~pi0626 & n34943;
  assign n35128 = pi0626 & ~n35117;
  assign n35129 = pi0641 & ~n35127;
  assign n35130 = ~n35128 & n35129;
  assign n35131 = pi1158 & ~n35126;
  assign n35132 = ~n35130 & n35131;
  assign n35133 = ~n35125 & ~n35132;
  assign n35134 = pi0788 & ~n35133;
  assign n35135 = ~n20364 & ~n35118;
  assign n35136 = ~n35134 & n35135;
  assign n35137 = ~n35048 & ~n35136;
  assign n35138 = ~pi0207 & ~n35137;
  assign n35139 = pi0609 & ~n34918;
  assign n35140 = ~pi0778 & ~n34080;
  assign n35141 = ~pi0625 & n34080;
  assign n35142 = ~pi1153 & ~n35141;
  assign n35143 = pi0625 & n24385;
  assign n35144 = pi1153 & ~n35143;
  assign n35145 = ~pi0608 & ~n35144;
  assign n35146 = ~n35142 & n35145;
  assign n35147 = pi0625 & n34080;
  assign n35148 = pi1153 & ~n35147;
  assign n35149 = ~pi0625 & n24385;
  assign n35150 = ~pi1153 & ~n35149;
  assign n35151 = pi0608 & ~n35150;
  assign n35152 = ~n35148 & n35151;
  assign n35153 = pi0778 & ~n35146;
  assign n35154 = ~n35152 & n35153;
  assign n35155 = ~n35140 & ~n35154;
  assign n35156 = ~pi0609 & ~n35155;
  assign n35157 = n17073 & ~n35139;
  assign n35158 = ~n35156 & n35157;
  assign n35159 = pi0609 & ~n35155;
  assign n35160 = ~pi0609 & ~n34918;
  assign n35161 = n17072 & ~n35160;
  assign n35162 = ~n35159 & n35161;
  assign n35163 = ~n35158 & ~n35162;
  assign n35164 = pi0785 & ~n35163;
  assign n35165 = ~pi0785 & n35155;
  assign n35166 = ~n35164 & ~n35165;
  assign n35167 = ~pi0781 & n35166;
  assign n35168 = ~pi0618 & n35166;
  assign n35169 = ~n17075 & n34918;
  assign n35170 = pi0618 & ~n35169;
  assign n35171 = n16637 & ~n35170;
  assign n35172 = ~n35168 & n35171;
  assign n35173 = ~pi0618 & ~n35169;
  assign n35174 = pi0618 & n35166;
  assign n35175 = n16636 & ~n35173;
  assign n35176 = ~n35174 & n35175;
  assign n35177 = pi0781 & ~n35172;
  assign n35178 = ~n35176 & n35177;
  assign n35179 = ~n23615 & ~n35167;
  assign n35180 = ~n35178 & n35179;
  assign n35181 = n19150 & n34918;
  assign n35182 = n16634 & n20231;
  assign n35183 = n35181 & n35182;
  assign n35184 = ~n35180 & ~n35183;
  assign n35185 = ~pi0788 & n35184;
  assign n35186 = ~n16635 & n35181;
  assign n35187 = pi0626 & ~n35186;
  assign n35188 = ~pi0641 & ~n35187;
  assign n35189 = ~pi0626 & n35184;
  assign n35190 = ~pi1158 & n35188;
  assign n35191 = ~n35189 & n35190;
  assign n35192 = pi0626 & n35184;
  assign n35193 = ~pi0626 & ~n35186;
  assign n35194 = pi0641 & ~n35193;
  assign n35195 = pi1158 & n35194;
  assign n35196 = ~n35192 & n35195;
  assign n35197 = pi0788 & ~n35191;
  assign n35198 = ~n35196 & n35197;
  assign n35199 = ~n20364 & ~n35185;
  assign n35200 = ~n35198 & n35199;
  assign n35201 = n17779 & n17855;
  assign n35202 = n34919 & n35201;
  assign n35203 = ~n35200 & ~n35202;
  assign n35204 = pi0207 & ~n35203;
  assign n35205 = ~pi0623 & ~n35204;
  assign n35206 = ~n35138 & n35205;
  assign n35207 = ~pi1156 & ~n34919;
  assign n35208 = pi1156 & ~n35022;
  assign n35209 = n20566 & ~n35207;
  assign n35210 = ~n35208 & n35209;
  assign n35211 = pi1156 & ~n34919;
  assign n35212 = ~pi1156 & ~n35022;
  assign n35213 = n20568 & ~n35211;
  assign n35214 = ~n35212 & n35213;
  assign n35215 = ~n35210 & ~n35214;
  assign n35216 = pi0792 & ~n35215;
  assign n35217 = n17868 & n35021;
  assign n35218 = ~pi1159 & ~n35020;
  assign n35219 = pi1159 & ~n35181;
  assign n35220 = ~pi0619 & pi0648;
  assign n35221 = ~n35218 & n35220;
  assign n35222 = ~n35219 & n35221;
  assign n35223 = pi1159 & ~n35020;
  assign n35224 = ~pi1159 & ~n35181;
  assign n35225 = pi0619 & ~pi0648;
  assign n35226 = ~n35223 & n35225;
  assign n35227 = ~n35224 & n35226;
  assign n35228 = pi0789 & ~n35222;
  assign n35229 = ~n35227 & n35228;
  assign n35230 = pi0789 & ~n35229;
  assign n35231 = ~pi1154 & ~n35170;
  assign n35232 = n20233 & n35019;
  assign n35233 = ~pi0627 & ~n35232;
  assign n35234 = ~n35231 & n35233;
  assign n35235 = n20232 & n35019;
  assign n35236 = ~pi0778 & ~n34085;
  assign n35237 = ~pi0625 & n34085;
  assign n35238 = pi0625 & n35017;
  assign n35239 = ~pi1153 & ~n35238;
  assign n35240 = ~n35237 & n35239;
  assign n35241 = n35145 & ~n35240;
  assign n35242 = ~pi0625 & n35017;
  assign n35243 = pi0625 & n34085;
  assign n35244 = pi1153 & ~n35242;
  assign n35245 = ~n35243 & n35244;
  assign n35246 = n35151 & ~n35245;
  assign n35247 = pi0778 & ~n35241;
  assign n35248 = ~n35246 & n35247;
  assign n35249 = ~n35236 & ~n35248;
  assign n35250 = ~pi0785 & ~n35249;
  assign n35251 = n20223 & n35018;
  assign n35252 = ~pi0609 & ~n35249;
  assign n35253 = ~pi1155 & ~n35139;
  assign n35254 = ~n35252 & n35253;
  assign n35255 = ~pi0660 & ~n35251;
  assign n35256 = ~n35254 & n35255;
  assign n35257 = n20222 & n35018;
  assign n35258 = pi0609 & ~n35249;
  assign n35259 = pi1155 & ~n35160;
  assign n35260 = ~n35258 & n35259;
  assign n35261 = pi0660 & ~n35257;
  assign n35262 = ~n35260 & n35261;
  assign n35263 = ~n35256 & ~n35262;
  assign n35264 = pi0785 & ~n35263;
  assign n35265 = ~n35250 & ~n35264;
  assign n35266 = pi0618 & ~n35265;
  assign n35267 = pi1154 & ~n35173;
  assign n35268 = ~n35266 & n35267;
  assign n35269 = pi0627 & ~n35235;
  assign n35270 = ~n35268 & n35269;
  assign n35271 = ~n35234 & ~n35270;
  assign n35272 = pi0781 & ~n35271;
  assign n35273 = ~pi0618 & ~pi0627;
  assign n35274 = pi0781 & ~n35273;
  assign n35275 = ~n35265 & ~n35274;
  assign n35276 = ~n23614 & n35229;
  assign n35277 = ~n35275 & ~n35276;
  assign n35278 = ~n35272 & n35277;
  assign n35279 = ~n35230 & ~n35278;
  assign n35280 = ~pi0626 & n35279;
  assign n35281 = n35188 & ~n35280;
  assign n35282 = ~pi1158 & ~n35217;
  assign n35283 = ~n35281 & n35282;
  assign n35284 = n17869 & n35021;
  assign n35285 = pi0626 & n35279;
  assign n35286 = n35194 & ~n35285;
  assign n35287 = pi1158 & ~n35284;
  assign n35288 = ~n35286 & n35287;
  assign n35289 = ~n35283 & ~n35288;
  assign n35290 = pi0788 & ~n35289;
  assign n35291 = ~pi0788 & n35279;
  assign n35292 = ~n20364 & ~n35291;
  assign n35293 = ~n35290 & n35292;
  assign n35294 = ~n35216 & ~n35293;
  assign n35295 = pi0207 & ~n35294;
  assign n35296 = n2571 & n19488;
  assign n35297 = ~pi0778 & ~n35296;
  assign n35298 = ~pi0625 & n34971;
  assign n35299 = pi0625 & n35296;
  assign n35300 = pi1153 & ~n35299;
  assign n35301 = ~n35298 & n35300;
  assign n35302 = n35065 & ~n35301;
  assign n35303 = ~pi0625 & n35296;
  assign n35304 = pi0625 & n34971;
  assign n35305 = ~pi1153 & ~n35303;
  assign n35306 = ~n35304 & n35305;
  assign n35307 = n35060 & ~n35306;
  assign n35308 = pi0778 & ~n35302;
  assign n35309 = ~n35307 & n35308;
  assign n35310 = ~n35297 & ~n35309;
  assign n35311 = ~pi0609 & ~n35310;
  assign n35312 = ~n35054 & ~n35311;
  assign n35313 = ~pi1155 & ~n35312;
  assign n35314 = ~pi0660 & ~n34982;
  assign n35315 = ~n35313 & n35314;
  assign n35316 = pi0609 & ~n35310;
  assign n35317 = ~n35076 & ~n35316;
  assign n35318 = pi1155 & ~n35317;
  assign n35319 = pi0660 & ~n34978;
  assign n35320 = ~n35318 & n35319;
  assign n35321 = ~n35315 & ~n35320;
  assign n35322 = pi0785 & ~n35321;
  assign n35323 = ~pi0785 & n35310;
  assign n35324 = ~n35322 & ~n35323;
  assign n35325 = ~pi0618 & n35324;
  assign n35326 = ~n35052 & ~n35325;
  assign n35327 = ~pi1154 & ~n35326;
  assign n35328 = ~pi0627 & ~n34994;
  assign n35329 = ~n35327 & n35328;
  assign n35330 = pi0618 & n35324;
  assign n35331 = ~n35092 & ~n35330;
  assign n35332 = pi1154 & ~n35331;
  assign n35333 = pi0627 & ~n34990;
  assign n35334 = ~n35332 & n35333;
  assign n35335 = ~n35329 & ~n35334;
  assign n35336 = pi0781 & ~n35335;
  assign n35337 = ~pi0781 & ~n35324;
  assign n35338 = ~n35336 & ~n35337;
  assign n35339 = ~pi0789 & n35338;
  assign n35340 = ~pi0619 & n35338;
  assign n35341 = ~n35050 & ~n35340;
  assign n35342 = ~pi1159 & ~n35341;
  assign n35343 = ~pi0648 & ~n35006;
  assign n35344 = ~n35342 & n35343;
  assign n35345 = pi0619 & n35338;
  assign n35346 = ~n35108 & ~n35345;
  assign n35347 = pi1159 & ~n35346;
  assign n35348 = pi0648 & ~n35002;
  assign n35349 = ~n35347 & n35348;
  assign n35350 = pi0789 & ~n35344;
  assign n35351 = ~n35349 & n35350;
  assign n35352 = n17970 & ~n35339;
  assign n35353 = ~n35351 & n35352;
  assign n35354 = pi0641 & ~n34943;
  assign n35355 = n17865 & ~n35126;
  assign n35356 = ~n35354 & n35355;
  assign n35357 = ~n16630 & ~n17870;
  assign n35358 = n35009 & n35357;
  assign n35359 = ~pi0641 & ~n34943;
  assign n35360 = n17866 & ~n35119;
  assign n35361 = ~n35359 & n35360;
  assign n35362 = ~n35356 & ~n35361;
  assign n35363 = ~n35358 & n35362;
  assign n35364 = pi0788 & ~n35363;
  assign n35365 = ~n20364 & ~n35364;
  assign n35366 = ~n35353 & n35365;
  assign n35367 = ~n20570 & n35012;
  assign n35368 = pi1156 & n35038;
  assign n35369 = ~n35045 & ~n35367;
  assign n35370 = ~n35368 & n35369;
  assign n35371 = pi0792 & ~n35370;
  assign n35372 = ~n35366 & ~n35371;
  assign n35373 = ~pi0207 & ~n35372;
  assign n35374 = pi0623 & ~n35295;
  assign n35375 = ~n35373 & n35374;
  assign n35376 = pi0710 & ~n35375;
  assign n35377 = ~n35206 & n35376;
  assign n35378 = ~n20206 & ~n35034;
  assign n35379 = ~n35377 & n35378;
  assign n35380 = ~n35033 & ~n35379;
  assign n35381 = pi0644 & n35380;
  assign n35382 = pi0715 & ~n34968;
  assign n35383 = ~n35381 & n35382;
  assign n35384 = n17804 & ~n34953;
  assign n35385 = ~n17804 & n35028;
  assign n35386 = ~n35384 & ~n35385;
  assign n35387 = pi0644 & n35386;
  assign n35388 = ~pi0644 & n34953;
  assign n35389 = ~pi0715 & ~n35388;
  assign n35390 = ~n35387 & n35389;
  assign n35391 = pi1160 & ~n35390;
  assign n35392 = ~n35383 & n35391;
  assign n35393 = pi0644 & n34967;
  assign n35394 = ~pi0644 & n35380;
  assign n35395 = ~pi0715 & ~n35393;
  assign n35396 = ~n35394 & n35395;
  assign n35397 = ~pi0644 & n35386;
  assign n35398 = pi0644 & n34953;
  assign n35399 = pi0715 & ~n35398;
  assign n35400 = ~n35397 & n35399;
  assign n35401 = ~pi1160 & ~n35400;
  assign n35402 = ~n35396 & n35401;
  assign n35403 = ~n35392 & ~n35402;
  assign n35404 = pi0790 & ~n35403;
  assign n35405 = ~pi0790 & n35380;
  assign n35406 = ~n35404 & ~n35405;
  assign n35407 = ~po1038 & ~n35406;
  assign n35408 = ~pi0207 & po1038;
  assign po0364 = n35407 | n35408;
  assign n35410 = pi0208 & ~n34920;
  assign n35411 = ~pi0208 & ~n34949;
  assign n35412 = ~n35410 & ~n35411;
  assign n35413 = pi0638 & ~n35412;
  assign n35414 = ~pi0208 & ~n17059;
  assign n35415 = ~pi0638 & ~n35414;
  assign n35416 = ~n35413 & ~n35415;
  assign n35417 = ~pi0787 & ~n35416;
  assign n35418 = ~pi0647 & n35416;
  assign n35419 = pi0647 & n35414;
  assign n35420 = ~pi1157 & ~n35419;
  assign n35421 = ~n35418 & n35420;
  assign n35422 = ~pi0647 & n35414;
  assign n35423 = pi0647 & n35416;
  assign n35424 = pi1157 & ~n35422;
  assign n35425 = ~n35423 & n35424;
  assign n35426 = ~n35421 & ~n35425;
  assign n35427 = pi0787 & ~n35426;
  assign n35428 = ~n35417 & ~n35427;
  assign n35429 = ~pi0644 & n35428;
  assign n35430 = ~pi0630 & n35425;
  assign n35431 = ~pi0208 & ~n35015;
  assign n35432 = pi0208 & ~n35023;
  assign n35433 = pi0607 & ~n35432;
  assign n35434 = ~n35431 & n35433;
  assign n35435 = ~pi0607 & n35414;
  assign n35436 = ~n35434 & ~n35435;
  assign n35437 = ~n20559 & n35436;
  assign n35438 = pi0630 & n35421;
  assign n35439 = ~n35430 & ~n35437;
  assign n35440 = ~n35438 & n35439;
  assign n35441 = pi0787 & ~n35440;
  assign n35442 = ~pi0638 & ~n35436;
  assign n35443 = ~pi0208 & ~n35137;
  assign n35444 = pi0208 & ~n35203;
  assign n35445 = ~pi0607 & ~n35444;
  assign n35446 = ~n35443 & n35445;
  assign n35447 = pi0208 & ~n35294;
  assign n35448 = ~pi0208 & ~n35372;
  assign n35449 = pi0607 & ~n35447;
  assign n35450 = ~n35448 & n35449;
  assign n35451 = pi0638 & ~n35450;
  assign n35452 = ~n35446 & n35451;
  assign n35453 = ~n20206 & ~n35442;
  assign n35454 = ~n35452 & n35453;
  assign n35455 = ~n35441 & ~n35454;
  assign n35456 = pi0644 & n35455;
  assign n35457 = pi0715 & ~n35429;
  assign n35458 = ~n35456 & n35457;
  assign n35459 = n17804 & ~n35414;
  assign n35460 = ~n17804 & n35436;
  assign n35461 = ~n35459 & ~n35460;
  assign n35462 = pi0644 & n35461;
  assign n35463 = ~pi0644 & n35414;
  assign n35464 = ~pi0715 & ~n35463;
  assign n35465 = ~n35462 & n35464;
  assign n35466 = pi1160 & ~n35465;
  assign n35467 = ~n35458 & n35466;
  assign n35468 = pi0644 & n35428;
  assign n35469 = ~pi0644 & n35455;
  assign n35470 = ~pi0715 & ~n35468;
  assign n35471 = ~n35469 & n35470;
  assign n35472 = ~pi0644 & n35461;
  assign n35473 = pi0644 & n35414;
  assign n35474 = pi0715 & ~n35473;
  assign n35475 = ~n35472 & n35474;
  assign n35476 = ~pi1160 & ~n35475;
  assign n35477 = ~n35471 & n35476;
  assign n35478 = ~n35467 & ~n35477;
  assign n35479 = pi0790 & ~n35478;
  assign n35480 = ~pi0790 & n35455;
  assign n35481 = ~n35479 & ~n35480;
  assign n35482 = ~po1038 & ~n35481;
  assign n35483 = ~pi0208 & po1038;
  assign po0365 = n35482 | n35483;
  assign n35485 = n10197 & n17052;
  assign n35486 = ~pi0639 & n35485;
  assign n35487 = pi0715 & n17059;
  assign n35488 = ~n20206 & ~n35137;
  assign n35489 = ~pi0647 & ~n17059;
  assign n35490 = pi0647 & n34949;
  assign n35491 = ~n35489 & ~n35490;
  assign n35492 = ~pi0630 & ~n35491;
  assign n35493 = ~n35489 & ~n35492;
  assign n35494 = pi1157 & ~n35493;
  assign n35495 = pi0647 & ~n17059;
  assign n35496 = ~pi1157 & n35495;
  assign n35497 = ~pi0647 & n34949;
  assign n35498 = ~n35495 & ~n35497;
  assign n35499 = n17802 & ~n35498;
  assign n35500 = ~n35496 & ~n35499;
  assign n35501 = ~n35494 & n35500;
  assign n35502 = pi0787 & ~n35501;
  assign n35503 = ~n35488 & ~n35502;
  assign n35504 = ~pi0644 & ~n35503;
  assign n35505 = ~n19342 & n34949;
  assign n35506 = ~n17059 & n19342;
  assign n35507 = ~n35505 & ~n35506;
  assign n35508 = pi0644 & ~n35507;
  assign n35509 = ~pi0715 & ~n35508;
  assign n35510 = ~n35504 & n35509;
  assign n35511 = ~pi1160 & ~n35487;
  assign n35512 = ~n35510 & n35511;
  assign n35513 = ~pi0715 & n17059;
  assign n35514 = pi0644 & ~n35503;
  assign n35515 = ~pi0644 & ~n35507;
  assign n35516 = pi0715 & ~n35515;
  assign n35517 = ~n35514 & n35516;
  assign n35518 = pi1160 & ~n35513;
  assign n35519 = ~n35517 & n35518;
  assign n35520 = ~n35512 & ~n35519;
  assign n35521 = pi0790 & ~n35520;
  assign n35522 = ~pi0790 & ~n35503;
  assign n35523 = ~po1038 & ~n35522;
  assign n35524 = ~n35521 & n35523;
  assign n35525 = pi0639 & n35524;
  assign n35526 = ~pi0622 & ~n35486;
  assign n35527 = ~n35525 & n35526;
  assign n35528 = ~n17059 & n17804;
  assign n35529 = ~n17804 & n35015;
  assign n35530 = ~n35528 & ~n35529;
  assign n35531 = ~pi0790 & ~n35530;
  assign n35532 = pi0644 & ~n35530;
  assign n35533 = ~pi0644 & ~n17059;
  assign n35534 = ~n35532 & ~n35533;
  assign n35535 = pi1160 & n35534;
  assign n35536 = ~pi0644 & ~n35530;
  assign n35537 = pi0644 & ~n17059;
  assign n35538 = ~n35536 & ~n35537;
  assign n35539 = ~pi1160 & n35538;
  assign n35540 = pi0790 & ~n35535;
  assign n35541 = ~n35539 & n35540;
  assign n35542 = ~po1038 & ~n35531;
  assign n35543 = ~n35541 & n35542;
  assign n35544 = ~pi0639 & n35543;
  assign n35545 = pi0715 & n35538;
  assign n35546 = ~n20206 & ~n35372;
  assign n35547 = ~n20559 & n35015;
  assign n35548 = pi1157 & n35492;
  assign n35549 = ~n35499 & ~n35547;
  assign n35550 = ~n35548 & n35549;
  assign n35551 = pi0787 & ~n35550;
  assign n35552 = ~n35546 & ~n35551;
  assign n35553 = ~pi0644 & ~n35552;
  assign n35554 = n35509 & ~n35553;
  assign n35555 = ~pi1160 & ~n35545;
  assign n35556 = ~n35554 & n35555;
  assign n35557 = ~pi0715 & n35534;
  assign n35558 = pi0644 & ~n35552;
  assign n35559 = n35516 & ~n35558;
  assign n35560 = pi1160 & ~n35557;
  assign n35561 = ~n35559 & n35560;
  assign n35562 = ~n35556 & ~n35561;
  assign n35563 = pi0790 & ~n35562;
  assign n35564 = ~pi0790 & ~n35552;
  assign n35565 = ~po1038 & ~n35564;
  assign n35566 = ~n35563 & n35565;
  assign n35567 = pi0639 & n35566;
  assign n35568 = pi0622 & ~n35544;
  assign n35569 = ~n35567 & n35568;
  assign n35570 = ~n35527 & ~n35569;
  assign n35571 = ~pi0209 & ~n35570;
  assign n35572 = ~pi0644 & pi1160;
  assign n35573 = pi0644 & ~pi1160;
  assign n35574 = ~n35572 & ~n35573;
  assign n35575 = pi0790 & ~n35574;
  assign n35576 = n23684 & n35022;
  assign n35577 = ~po1038 & ~n35575;
  assign n35578 = n35576 & n35577;
  assign n35579 = pi0622 & n35578;
  assign n35580 = ~pi0639 & ~n35579;
  assign n35581 = ~n20206 & ~n35203;
  assign n35582 = n17804 & n19341;
  assign n35583 = n34920 & n35582;
  assign n35584 = ~n35581 & ~n35583;
  assign n35585 = ~pi0790 & n35584;
  assign n35586 = ~n19342 & n34920;
  assign n35587 = ~pi0644 & ~n35586;
  assign n35588 = pi0715 & ~n35587;
  assign n35589 = pi0644 & n35584;
  assign n35590 = pi1160 & n35588;
  assign n35591 = ~n35589 & n35590;
  assign n35592 = pi0644 & ~n35586;
  assign n35593 = ~pi0715 & ~n35592;
  assign n35594 = ~pi0644 & n35584;
  assign n35595 = ~pi1160 & n35593;
  assign n35596 = ~n35594 & n35595;
  assign n35597 = pi0790 & ~n35591;
  assign n35598 = ~n35596 & n35597;
  assign n35599 = ~po1038 & ~n35585;
  assign n35600 = ~n35598 & n35599;
  assign n35601 = ~pi0622 & ~n35600;
  assign n35602 = ~pi0644 & pi0715;
  assign n35603 = n35576 & n35602;
  assign n35604 = pi0647 & n34920;
  assign n35605 = pi1157 & ~n35604;
  assign n35606 = pi0647 & n35023;
  assign n35607 = ~pi0647 & ~n35294;
  assign n35608 = ~pi1157 & ~n35606;
  assign n35609 = ~n35607 & n35608;
  assign n35610 = ~pi0630 & ~n35605;
  assign n35611 = ~n35609 & n35610;
  assign n35612 = ~pi0647 & n34920;
  assign n35613 = ~pi1157 & ~n35612;
  assign n35614 = ~pi0647 & n35023;
  assign n35615 = pi0647 & ~n35294;
  assign n35616 = pi1157 & ~n35614;
  assign n35617 = ~n35615 & n35616;
  assign n35618 = pi0630 & ~n35613;
  assign n35619 = ~n35617 & n35618;
  assign n35620 = ~n35611 & ~n35619;
  assign n35621 = pi0787 & ~n35620;
  assign n35622 = ~pi0787 & ~n35294;
  assign n35623 = ~n35621 & ~n35622;
  assign n35624 = ~pi0644 & n35623;
  assign n35625 = n35593 & ~n35624;
  assign n35626 = ~pi1160 & ~n35603;
  assign n35627 = ~n35625 & n35626;
  assign n35628 = pi0644 & ~pi0715;
  assign n35629 = n35576 & n35628;
  assign n35630 = pi0644 & n35623;
  assign n35631 = n35588 & ~n35630;
  assign n35632 = pi1160 & ~n35629;
  assign n35633 = ~n35631 & n35632;
  assign n35634 = ~n35627 & ~n35633;
  assign n35635 = pi0790 & ~n35634;
  assign n35636 = ~pi0790 & n35623;
  assign n35637 = ~po1038 & ~n35636;
  assign n35638 = ~n35635 & n35637;
  assign n35639 = pi0622 & pi0639;
  assign n35640 = ~n35638 & n35639;
  assign n35641 = pi0209 & ~n35580;
  assign n35642 = ~n35601 & n35641;
  assign n35643 = ~n35640 & n35642;
  assign po0366 = n35571 | n35643;
  assign n35645 = pi0210 & ~n16641;
  assign n35646 = pi0634 & n20902;
  assign n35647 = pi0633 & pi0947;
  assign n35648 = ~n35646 & ~n35647;
  assign n35649 = n16641 & ~n35648;
  assign n35650 = pi0038 & ~n35645;
  assign n35651 = ~n35649 & n35650;
  assign n35652 = ~n16939 & ~n35648;
  assign n35653 = pi0299 & ~n35652;
  assign n35654 = ~n16940 & n35653;
  assign n35655 = pi0210 & ~n16930;
  assign n35656 = n16930 & ~n35648;
  assign n35657 = ~pi0299 & ~n35655;
  assign n35658 = ~n35656 & n35657;
  assign n35659 = ~pi0039 & ~n35654;
  assign n35660 = ~n35658 & n35659;
  assign n35661 = pi0210 & ~n16653;
  assign n35662 = ~n33589 & ~n35661;
  assign n35663 = n6227 & n35662;
  assign n35664 = pi0947 & ~n35663;
  assign n35665 = pi0210 & n16721;
  assign n35666 = pi0633 & ~n16721;
  assign n35667 = ~n35665 & ~n35666;
  assign n35668 = ~n6227 & n35667;
  assign n35669 = n35664 & ~n35668;
  assign n35670 = pi0634 & n16653;
  assign n35671 = ~n35661 & ~n35670;
  assign n35672 = n6227 & n35671;
  assign n35673 = pi0907 & ~n35672;
  assign n35674 = ~n33430 & ~n35665;
  assign n35675 = ~n6227 & n35674;
  assign n35676 = n35673 & ~n35675;
  assign n35677 = n6227 & n16652;
  assign n35678 = n2926 & n35677;
  assign n35679 = n35665 & ~n35678;
  assign n35680 = ~n35676 & ~n35679;
  assign n35681 = ~pi0947 & ~n35680;
  assign n35682 = ~n6205 & ~n35669;
  assign n35683 = ~n35681 & n35682;
  assign n35684 = ~po1101 & n35662;
  assign n35685 = pi0947 & ~n35684;
  assign n35686 = ~n6197 & ~n35667;
  assign n35687 = po1101 & n35662;
  assign n35688 = ~n6198 & ~n35687;
  assign n35689 = ~n35686 & ~n35688;
  assign n35690 = n35685 & ~n35689;
  assign n35691 = ~n6198 & ~n35671;
  assign n35692 = pi0907 & ~n35691;
  assign n35693 = n6198 & ~n35674;
  assign n35694 = n35692 & ~n35693;
  assign n35695 = ~po1101 & n35661;
  assign n35696 = pi0210 & po1101;
  assign n35697 = ~n16797 & n35696;
  assign n35698 = ~n35695 & ~n35697;
  assign n35699 = ~pi0907 & n35698;
  assign n35700 = ~pi0947 & ~n35694;
  assign n35701 = ~n35699 & n35700;
  assign n35702 = n6205 & ~n35690;
  assign n35703 = ~n35701 & n35702;
  assign n35704 = pi0223 & ~n35683;
  assign n35705 = ~n35703 & n35704;
  assign n35706 = n16653 & ~n35648;
  assign n35707 = ~n35661 & ~n35706;
  assign n35708 = n2603 & n35707;
  assign n35709 = pi0210 & n16681;
  assign n35710 = pi0633 & ~n16681;
  assign n35711 = ~n35709 & ~n35710;
  assign n35712 = ~n6197 & ~n35711;
  assign n35713 = ~n35688 & ~n35712;
  assign n35714 = n35685 & ~n35713;
  assign n35715 = pi0634 & ~n16681;
  assign n35716 = ~n35709 & ~n35715;
  assign n35717 = n6198 & ~n35716;
  assign n35718 = n35692 & ~n35717;
  assign n35719 = ~n16684 & n35696;
  assign n35720 = ~n35695 & ~n35719;
  assign n35721 = ~pi0907 & n35720;
  assign n35722 = ~pi0947 & ~n35718;
  assign n35723 = ~n35721 & n35722;
  assign n35724 = n6205 & ~n35714;
  assign n35725 = ~n35723 & n35724;
  assign n35726 = ~n6227 & n35716;
  assign n35727 = n35673 & ~n35726;
  assign n35728 = pi0210 & ~n17143;
  assign n35729 = ~pi0907 & n35728;
  assign n35730 = ~n35727 & ~n35729;
  assign n35731 = ~pi0947 & ~n35730;
  assign n35732 = ~n6227 & n35711;
  assign n35733 = n35664 & ~n35732;
  assign n35734 = ~n6205 & ~n35733;
  assign n35735 = ~n35731 & n35734;
  assign n35736 = ~n35725 & ~n35735;
  assign n35737 = ~n2603 & ~n35736;
  assign n35738 = ~pi0223 & ~n35708;
  assign n35739 = ~n35737 & n35738;
  assign n35740 = ~pi0299 & ~n35705;
  assign n35741 = ~n35739 & n35740;
  assign n35742 = ~n6241 & ~n35679;
  assign n35743 = n6241 & n35698;
  assign n35744 = ~pi0907 & ~n35742;
  assign n35745 = ~n35743 & n35744;
  assign n35746 = ~n35676 & ~n35745;
  assign n35747 = ~pi0947 & ~n35746;
  assign n35748 = ~n35669 & ~n35747;
  assign n35749 = pi0215 & ~n35748;
  assign n35750 = n3448 & n35707;
  assign n35751 = ~n6241 & ~n35728;
  assign n35752 = n6241 & n35720;
  assign n35753 = ~pi0907 & ~n35752;
  assign n35754 = ~n35751 & n35753;
  assign n35755 = ~n35727 & ~n35754;
  assign n35756 = ~pi0947 & ~n35755;
  assign n35757 = ~n3448 & ~n35733;
  assign n35758 = ~n35756 & n35757;
  assign n35759 = ~pi0215 & ~n35750;
  assign n35760 = ~n35758 & n35759;
  assign n35761 = pi0299 & ~n35749;
  assign n35762 = ~n35760 & n35761;
  assign n35763 = pi0039 & ~n35762;
  assign n35764 = ~n35741 & n35763;
  assign n35765 = ~pi0038 & ~n35660;
  assign n35766 = ~n35764 & n35765;
  assign n35767 = ~n35651 & ~n35766;
  assign n35768 = n10197 & ~n35767;
  assign n35769 = ~pi0210 & ~n10197;
  assign po0367 = ~n35768 & ~n35769;
  assign n35771 = n2571 & ~n21641;
  assign n35772 = ~pi0606 & n35771;
  assign n35773 = n2571 & ~n21637;
  assign n35774 = pi0606 & n35773;
  assign n35775 = pi0643 & ~n35772;
  assign n35776 = ~n35774 & n35775;
  assign n35777 = ~pi0606 & n17059;
  assign n35778 = n2571 & ~n21010;
  assign n35779 = pi0606 & n35778;
  assign n35780 = ~pi0643 & ~n35777;
  assign n35781 = ~n35779 & n35780;
  assign n35782 = ~po1038 & ~n35781;
  assign n35783 = ~n35776 & n35782;
  assign n35784 = pi0211 & ~n35783;
  assign n35785 = n2571 & n21628;
  assign n35786 = ~pi0606 & ~n35785;
  assign n35787 = n2571 & n21625;
  assign n35788 = pi0606 & ~n35787;
  assign n35789 = pi0643 & ~n35786;
  assign n35790 = ~n35788 & n35789;
  assign n35791 = n2571 & n21034;
  assign n35792 = pi0606 & ~pi0643;
  assign n35793 = n35791 & n35792;
  assign n35794 = ~n35790 & ~n35793;
  assign n35795 = ~pi0211 & ~po1038;
  assign n35796 = ~n35794 & n35795;
  assign po0368 = n35784 | n35796;
  assign n35798 = ~pi0607 & n35771;
  assign n35799 = pi0607 & n35773;
  assign n35800 = pi0638 & ~n35798;
  assign n35801 = ~n35799 & n35800;
  assign n35802 = ~pi0607 & n17059;
  assign n35803 = pi0607 & n35778;
  assign n35804 = ~pi0638 & ~n35802;
  assign n35805 = ~n35803 & n35804;
  assign n35806 = ~po1038 & ~n35805;
  assign n35807 = ~n35801 & n35806;
  assign n35808 = ~pi0212 & ~n35807;
  assign n35809 = pi0607 & ~n35787;
  assign n35810 = ~pi0607 & ~n35785;
  assign n35811 = pi0638 & ~n35809;
  assign n35812 = ~n35810 & n35811;
  assign n35813 = pi0607 & ~pi0638;
  assign n35814 = n35791 & n35813;
  assign n35815 = ~n35812 & ~n35814;
  assign n35816 = pi0212 & ~po1038;
  assign n35817 = ~n35815 & n35816;
  assign po0369 = n35808 | n35817;
  assign n35819 = pi0213 & ~po1038;
  assign n35820 = pi0622 & ~n35787;
  assign n35821 = ~pi0622 & ~n35785;
  assign n35822 = pi0639 & ~n35820;
  assign n35823 = ~n35821 & n35822;
  assign n35824 = pi0622 & ~pi0639;
  assign n35825 = n35791 & n35824;
  assign n35826 = ~n35823 & ~n35825;
  assign n35827 = n35819 & ~n35826;
  assign n35828 = ~pi0639 & n35778;
  assign n35829 = pi0639 & n35773;
  assign n35830 = pi0622 & ~n35828;
  assign n35831 = ~n35829 & n35830;
  assign n35832 = ~pi0639 & n17059;
  assign n35833 = pi0639 & n35771;
  assign n35834 = ~pi0622 & ~n35832;
  assign n35835 = ~n35833 & n35834;
  assign n35836 = ~po1038 & ~n35835;
  assign n35837 = ~n35831 & n35836;
  assign n35838 = ~pi0213 & ~n35837;
  assign po0370 = n35827 | n35838;
  assign n35840 = ~pi0623 & n35771;
  assign n35841 = pi0623 & n35773;
  assign n35842 = pi0710 & ~n35840;
  assign n35843 = ~n35841 & n35842;
  assign n35844 = ~pi0623 & n17059;
  assign n35845 = pi0623 & n35778;
  assign n35846 = ~pi0710 & ~n35844;
  assign n35847 = ~n35845 & n35846;
  assign n35848 = ~po1038 & ~n35847;
  assign n35849 = ~n35843 & n35848;
  assign n35850 = ~pi0214 & ~n35849;
  assign n35851 = pi0623 & ~n35787;
  assign n35852 = ~pi0623 & ~n35785;
  assign n35853 = pi0710 & ~n35851;
  assign n35854 = ~n35852 & n35853;
  assign n35855 = pi0623 & ~pi0710;
  assign n35856 = n35791 & n35855;
  assign n35857 = ~n35854 & ~n35856;
  assign n35858 = pi0214 & ~po1038;
  assign n35859 = ~n35857 & n35858;
  assign po0371 = n35850 | n35859;
  assign n35861 = pi0215 & ~n10197;
  assign n35862 = pi0681 & pi0907;
  assign n35863 = ~pi0947 & n35862;
  assign n35864 = pi0642 & pi0947;
  assign n35865 = ~n35863 & ~n35864;
  assign n35866 = n16641 & ~n35865;
  assign n35867 = pi0215 & ~n16641;
  assign n35868 = pi0038 & ~n35866;
  assign n35869 = ~n35867 & n35868;
  assign n35870 = pi0215 & ~n16941;
  assign n35871 = n16941 & ~n35865;
  assign n35872 = pi0299 & ~n35870;
  assign n35873 = ~n35871 & n35872;
  assign n35874 = n16930 & ~n35865;
  assign n35875 = pi0215 & ~n16930;
  assign n35876 = ~pi0299 & ~n35874;
  assign n35877 = ~n35875 & n35876;
  assign n35878 = ~pi0039 & ~n35873;
  assign n35879 = ~n35877 & n35878;
  assign n35880 = ~pi0947 & n21326;
  assign n35881 = n16656 & n16963;
  assign n35882 = ~n6195 & ~n16814;
  assign n35883 = ~pi0642 & ~n35881;
  assign n35884 = ~n35882 & n35883;
  assign n35885 = pi0947 & ~n35884;
  assign n35886 = ~n35863 & ~n35885;
  assign n35887 = ~n35880 & n35886;
  assign n35888 = pi0299 & ~n35887;
  assign n35889 = n2603 & ~n35865;
  assign n35890 = n2603 & ~n16653;
  assign n35891 = n21431 & ~n35862;
  assign n35892 = ~pi0642 & n17143;
  assign n35893 = ~n6205 & ~n35892;
  assign n35894 = ~pi0642 & n16684;
  assign n35895 = n6195 & ~n35894;
  assign n35896 = n16769 & n17167;
  assign n35897 = ~n6191 & n16653;
  assign n35898 = ~pi0642 & n35897;
  assign n35899 = ~n6195 & ~n35898;
  assign n35900 = ~n35896 & n35899;
  assign n35901 = ~n35895 & ~n35900;
  assign n35902 = n6205 & ~n35901;
  assign n35903 = pi0947 & ~n35893;
  assign n35904 = ~n35902 & n35903;
  assign n35905 = ~n2603 & ~n35904;
  assign n35906 = ~n35891 & n35905;
  assign n35907 = ~pi0223 & ~n35889;
  assign n35908 = ~n35890 & n35907;
  assign n35909 = ~n35906 & n35908;
  assign n35910 = ~n6205 & ~n35884;
  assign n35911 = n6195 & ~n16797;
  assign n35912 = ~n6195 & ~n16803;
  assign n35913 = ~pi0642 & ~n35911;
  assign n35914 = ~n35912 & n35913;
  assign n35915 = n6205 & ~n35914;
  assign n35916 = pi0947 & ~n35910;
  assign n35917 = ~n35915 & n35916;
  assign n35918 = ~n21052 & ~n35917;
  assign n35919 = pi0223 & ~n35863;
  assign n35920 = ~n35918 & n35919;
  assign n35921 = ~pi0299 & ~n35920;
  assign n35922 = ~n35909 & n35921;
  assign n35923 = ~n35888 & ~n35922;
  assign n35924 = pi0215 & ~n35923;
  assign n35925 = n16653 & n35889;
  assign n35926 = n16702 & n35862;
  assign n35927 = ~pi0947 & ~n35926;
  assign n35928 = pi0642 & n16657;
  assign n35929 = ~n6195 & n16699;
  assign n35930 = ~n17142 & ~n35929;
  assign n35931 = n35928 & n35930;
  assign n35932 = pi0642 & ~n16657;
  assign n35933 = ~n16699 & n35932;
  assign n35934 = pi0947 & ~n35933;
  assign n35935 = ~n35931 & n35934;
  assign n35936 = ~n35927 & ~n35935;
  assign n35937 = ~n6205 & ~n35936;
  assign n35938 = n16653 & n35932;
  assign n35939 = ~n16974 & n35928;
  assign n35940 = ~n16995 & n35939;
  assign n35941 = ~n35938 & ~n35940;
  assign n35942 = pi0947 & ~n35941;
  assign n35943 = n16776 & n35863;
  assign n35944 = n6205 & ~n35942;
  assign n35945 = ~n35943 & n35944;
  assign n35946 = ~n2603 & ~n35937;
  assign n35947 = ~n35945 & n35946;
  assign n35948 = ~pi0223 & ~n35925;
  assign n35949 = ~n35947 & n35948;
  assign n35950 = n6205 & ~n16803;
  assign n35951 = n35862 & ~n35950;
  assign n35952 = ~pi0947 & ~n35951;
  assign n35953 = pi0947 & ~n16723;
  assign n35954 = ~n16814 & ~n35953;
  assign n35955 = ~n6205 & n35954;
  assign n35956 = ~n16973 & n35939;
  assign n35957 = pi0947 & ~n35938;
  assign n35958 = ~n35956 & n35957;
  assign n35959 = ~n35955 & ~n35958;
  assign n35960 = ~n35952 & n35959;
  assign n35961 = pi0223 & ~n35960;
  assign n35962 = ~n35949 & ~n35961;
  assign n35963 = ~pi0299 & ~n35962;
  assign n35964 = n17026 & ~n35865;
  assign n35965 = ~n3448 & n35936;
  assign n35966 = pi0299 & ~n35964;
  assign n35967 = ~n35965 & n35966;
  assign n35968 = ~pi0215 & ~n35967;
  assign n35969 = ~n35963 & n35968;
  assign n35970 = ~n35924 & ~n35969;
  assign n35971 = pi0039 & ~n35970;
  assign n35972 = ~pi0038 & ~n35879;
  assign n35973 = ~n35971 & n35972;
  assign n35974 = n10197 & ~n35869;
  assign n35975 = ~n35973 & n35974;
  assign po0372 = n35861 | n35975;
  assign n35977 = pi0662 & pi0907;
  assign n35978 = ~pi0947 & n35977;
  assign n35979 = pi0614 & pi0947;
  assign n35980 = ~n35978 & ~n35979;
  assign n35981 = n16641 & ~n35980;
  assign n35982 = pi0216 & ~n16641;
  assign n35983 = pi0038 & ~n35981;
  assign n35984 = ~n35982 & n35983;
  assign n35985 = pi0216 & ~n16941;
  assign n35986 = n16941 & ~n35980;
  assign n35987 = pi0299 & ~n35985;
  assign n35988 = ~n35986 & n35987;
  assign n35989 = n16930 & ~n35980;
  assign n35990 = pi0216 & ~n16930;
  assign n35991 = ~pi0299 & ~n35989;
  assign n35992 = ~n35990 & n35991;
  assign n35993 = ~pi0039 & ~n35988;
  assign n35994 = ~n35992 & n35993;
  assign n35995 = ~n35950 & n35977;
  assign n35996 = ~pi0947 & ~n35995;
  assign n35997 = ~n16973 & n16997;
  assign n35998 = pi0947 & ~n17000;
  assign n35999 = ~n35997 & n35998;
  assign n36000 = ~n35955 & ~n35999;
  assign n36001 = ~n35996 & n36000;
  assign n36002 = pi0223 & ~n36001;
  assign n36003 = n2603 & ~n35980;
  assign n36004 = n16653 & n36003;
  assign n36005 = n35930 & n35979;
  assign n36006 = n16702 & n35978;
  assign n36007 = ~n36005 & ~n36006;
  assign n36008 = ~n6205 & n36007;
  assign n36009 = n16776 & n35978;
  assign n36010 = pi0947 & ~n17001;
  assign n36011 = n6205 & ~n36010;
  assign n36012 = ~n36009 & n36011;
  assign n36013 = ~n2603 & ~n36008;
  assign n36014 = ~n36012 & n36013;
  assign n36015 = ~pi0223 & ~n36004;
  assign n36016 = ~n36014 & n36015;
  assign n36017 = ~pi0216 & ~n36002;
  assign n36018 = ~n36016 & n36017;
  assign n36019 = ~pi0616 & n16799;
  assign n36020 = ~n6195 & ~n16978;
  assign n36021 = ~n36019 & n36020;
  assign n36022 = ~pi0614 & ~n35911;
  assign n36023 = ~n36021 & n36022;
  assign n36024 = n6205 & ~n36023;
  assign n36025 = ~n17452 & ~n33382;
  assign n36026 = ~n33383 & n36025;
  assign n36027 = n17002 & ~n36026;
  assign n36028 = ~pi0614 & ~n16721;
  assign n36029 = n6195 & n36028;
  assign n36030 = ~n36027 & ~n36029;
  assign n36031 = ~n6205 & n36030;
  assign n36032 = pi0947 & ~n36031;
  assign n36033 = ~n36024 & n36032;
  assign n36034 = ~n21052 & ~n36033;
  assign n36035 = pi0223 & ~n35978;
  assign n36036 = ~n36034 & n36035;
  assign n36037 = ~pi0614 & n17143;
  assign n36038 = pi0947 & ~n36037;
  assign n36039 = ~pi0947 & ~n17018;
  assign n36040 = ~n6205 & ~n35978;
  assign n36041 = ~n36038 & n36040;
  assign n36042 = ~n36039 & n36041;
  assign n36043 = pi0947 & ~n17008;
  assign n36044 = ~pi0947 & n17011;
  assign n36045 = ~n35977 & n36044;
  assign n36046 = ~n36043 & ~n36045;
  assign n36047 = n6205 & ~n36046;
  assign n36048 = ~n2603 & ~n36042;
  assign n36049 = ~n36047 & n36048;
  assign n36050 = ~pi0223 & ~n36003;
  assign n36051 = ~n35890 & n36050;
  assign n36052 = ~n36049 & n36051;
  assign n36053 = pi0216 & ~n36036;
  assign n36054 = ~n36052 & n36053;
  assign n36055 = ~pi0299 & ~n36018;
  assign n36056 = ~n36054 & n36055;
  assign n36057 = n5777 & ~n36007;
  assign n36058 = n17026 & ~n35980;
  assign n36059 = ~pi0947 & n20994;
  assign n36060 = ~n35978 & ~n36038;
  assign n36061 = ~n36059 & n36060;
  assign n36062 = pi0216 & ~n36061;
  assign n36063 = ~n36057 & ~n36058;
  assign n36064 = ~n36062 & n36063;
  assign n36065 = ~pi0215 & ~n36064;
  assign n36066 = n16814 & n35977;
  assign n36067 = ~pi0947 & ~n36066;
  assign n36068 = pi0947 & n16723;
  assign n36069 = ~n35999 & ~n36068;
  assign n36070 = ~n36067 & n36069;
  assign n36071 = ~pi0216 & ~n36070;
  assign n36072 = pi0947 & n36030;
  assign n36073 = pi0216 & ~n35978;
  assign n36074 = ~n36072 & n36073;
  assign n36075 = ~n35880 & n36074;
  assign n36076 = pi0215 & ~n36071;
  assign n36077 = ~n36075 & n36076;
  assign n36078 = pi0299 & ~n36077;
  assign n36079 = ~n36065 & n36078;
  assign n36080 = pi0039 & ~n36056;
  assign n36081 = ~n36079 & n36080;
  assign n36082 = ~pi0038 & ~n35994;
  assign n36083 = ~n36081 & n36082;
  assign n36084 = ~n35984 & ~n36083;
  assign n36085 = n10197 & ~n36084;
  assign n36086 = ~pi0216 & ~n10197;
  assign po0373 = ~n36085 & ~n36086;
  assign n36088 = ~pi0695 & n35600;
  assign n36089 = pi0217 & ~n36088;
  assign n36090 = pi0695 & ~n35485;
  assign n36091 = ~pi0695 & ~n35524;
  assign n36092 = ~pi0217 & ~n36090;
  assign n36093 = ~n36091 & n36092;
  assign n36094 = ~pi0612 & ~n36089;
  assign n36095 = ~n36093 & n36094;
  assign n36096 = ~pi0695 & n35638;
  assign n36097 = pi0695 & n35578;
  assign n36098 = pi0217 & ~n36097;
  assign n36099 = ~n36096 & n36098;
  assign n36100 = pi0695 & ~n35543;
  assign n36101 = ~pi0695 & ~n35566;
  assign n36102 = ~pi0217 & ~n36100;
  assign n36103 = ~n36101 & n36102;
  assign n36104 = pi0612 & ~n36099;
  assign n36105 = ~n36103 & n36104;
  assign po0374 = n36095 | n36105;
  assign n36107 = ~n34786 & ~n34825;
  assign n36108 = n34786 & ~n34891;
  assign n36109 = ~n36107 & ~n36108;
  assign n36110 = ~pi0218 & ~n36109;
  assign n36111 = n34786 & n34899;
  assign n36112 = pi0218 & ~n36111;
  assign po0375 = ~n36110 & ~n36112;
  assign n36114 = ~pi0219 & ~po1038;
  assign n36115 = pi0617 & ~n35787;
  assign n36116 = ~pi0617 & ~n35785;
  assign n36117 = pi0637 & ~n36115;
  assign n36118 = ~n36116 & n36117;
  assign n36119 = pi0617 & ~pi0637;
  assign n36120 = n35791 & n36119;
  assign n36121 = ~n36118 & ~n36120;
  assign n36122 = n36114 & ~n36121;
  assign n36123 = ~pi0617 & n35771;
  assign n36124 = pi0617 & n35773;
  assign n36125 = pi0637 & ~n36123;
  assign n36126 = ~n36124 & n36125;
  assign n36127 = ~pi0617 & n17059;
  assign n36128 = pi0617 & n35778;
  assign n36129 = ~pi0637 & ~n36127;
  assign n36130 = ~n36128 & n36129;
  assign n36131 = ~po1038 & ~n36130;
  assign n36132 = ~n36126 & n36131;
  assign n36133 = pi0219 & ~n36132;
  assign po0376 = n36122 | n36133;
  assign n36135 = ~n34619 & ~n34910;
  assign n36136 = ~n34765 & n34910;
  assign n36137 = ~n36135 & ~n36136;
  assign n36138 = ~pi0220 & ~n36137;
  assign n36139 = n34774 & n34910;
  assign n36140 = pi0220 & ~n36139;
  assign po0377 = ~n36138 & ~n36140;
  assign n36142 = pi0661 & pi0907;
  assign n36143 = ~pi0947 & n36142;
  assign n36144 = pi0616 & pi0947;
  assign n36145 = ~n36143 & ~n36144;
  assign n36146 = n16641 & ~n36145;
  assign n36147 = pi0221 & ~n16641;
  assign n36148 = pi0038 & ~n36146;
  assign n36149 = ~n36147 & n36148;
  assign n36150 = pi0221 & ~n16941;
  assign n36151 = n16941 & ~n36145;
  assign n36152 = pi0299 & ~n36150;
  assign n36153 = ~n36151 & n36152;
  assign n36154 = n16930 & ~n36145;
  assign n36155 = pi0221 & ~n16930;
  assign n36156 = ~pi0299 & ~n36154;
  assign n36157 = ~n36155 & n36156;
  assign n36158 = ~pi0039 & ~n36153;
  assign n36159 = ~n36157 & n36158;
  assign n36160 = pi0947 & ~n16980;
  assign n36161 = ~n36143 & ~n36160;
  assign n36162 = n35950 & ~n36160;
  assign n36163 = ~n35955 & ~n36161;
  assign n36164 = ~n36162 & n36163;
  assign n36165 = pi0223 & ~n36164;
  assign n36166 = n16653 & ~n36145;
  assign n36167 = n2603 & n36166;
  assign n36168 = ~pi0223 & ~n36167;
  assign n36169 = n16976 & ~n16995;
  assign n36170 = ~n16979 & ~n36169;
  assign n36171 = pi0947 & ~n36170;
  assign n36172 = n16776 & n36143;
  assign n36173 = n6205 & ~n36171;
  assign n36174 = ~n36172 & n36173;
  assign n36175 = n35930 & n36144;
  assign n36176 = n16702 & n36143;
  assign n36177 = ~n36175 & ~n36176;
  assign n36178 = ~n6205 & n36177;
  assign n36179 = ~n2603 & ~n36178;
  assign n36180 = ~n36174 & n36179;
  assign n36181 = n36168 & ~n36180;
  assign n36182 = ~pi0221 & ~n36165;
  assign n36183 = ~n36181 & n36182;
  assign n36184 = ~n35892 & ~n35931;
  assign n36185 = n16984 & ~n36184;
  assign n36186 = ~n6197 & n16774;
  assign n36187 = ~n16697 & ~n36186;
  assign n36188 = n16981 & ~n36187;
  assign n36189 = pi0947 & ~n36185;
  assign n36190 = ~n36188 & n36189;
  assign n36191 = ~n36039 & ~n36190;
  assign n36192 = ~n6205 & ~n36191;
  assign n36193 = n16774 & n16981;
  assign n36194 = ~n16998 & n17008;
  assign n36195 = n16984 & ~n36194;
  assign n36196 = ~n36193 & ~n36195;
  assign n36197 = pi0947 & ~n36196;
  assign n36198 = n6205 & ~n36044;
  assign n36199 = ~n36197 & n36198;
  assign n36200 = ~n36143 & ~n36192;
  assign n36201 = ~n36199 & n36200;
  assign n36202 = ~n2603 & ~n36201;
  assign n36203 = ~n35890 & n36168;
  assign n36204 = ~n36202 & n36203;
  assign n36205 = ~pi0947 & n16990;
  assign n36206 = pi0947 & ~n16987;
  assign n36207 = n6205 & ~n36206;
  assign n36208 = ~n36205 & n36207;
  assign n36209 = ~pi0947 & ~n16970;
  assign n36210 = ~n16723 & ~n16800;
  assign n36211 = ~n6195 & ~n36210;
  assign n36212 = ~pi0616 & ~n35881;
  assign n36213 = ~n36211 & n36212;
  assign n36214 = pi0947 & ~n36213;
  assign n36215 = ~n36209 & ~n36214;
  assign n36216 = ~n6205 & ~n36215;
  assign n36217 = pi0223 & ~n36143;
  assign n36218 = ~n36208 & n36217;
  assign n36219 = ~n36216 & n36218;
  assign n36220 = pi0221 & ~n36219;
  assign n36221 = ~n36204 & n36220;
  assign n36222 = ~pi0299 & ~n36183;
  assign n36223 = ~n36221 & n36222;
  assign n36224 = ~n20994 & ~n36142;
  assign n36225 = ~pi0947 & ~n36224;
  assign n36226 = pi0221 & ~n36190;
  assign n36227 = ~n36225 & n36226;
  assign n36228 = pi0216 & ~n36177;
  assign n36229 = ~pi0216 & n36166;
  assign n36230 = ~pi0221 & ~n36229;
  assign n36231 = ~n36228 & n36230;
  assign n36232 = ~pi0215 & ~n36231;
  assign n36233 = ~n36227 & n36232;
  assign n36234 = pi0221 & ~n36143;
  assign n36235 = ~n36214 & n36234;
  assign n36236 = ~n35880 & n36235;
  assign n36237 = ~n35954 & ~n36161;
  assign n36238 = ~pi0221 & ~n36237;
  assign n36239 = pi0215 & ~n36238;
  assign n36240 = ~n36236 & n36239;
  assign n36241 = pi0299 & ~n36240;
  assign n36242 = ~n36233 & n36241;
  assign n36243 = pi0039 & ~n36223;
  assign n36244 = ~n36242 & n36243;
  assign n36245 = ~pi0038 & ~n36159;
  assign n36246 = ~n36244 & n36245;
  assign n36247 = ~n36149 & ~n36246;
  assign n36248 = n10197 & ~n36247;
  assign n36249 = ~pi0221 & ~n10197;
  assign po0378 = ~n36248 & ~n36249;
  assign n36251 = ~pi0223 & ~n17020;
  assign n36252 = ~n16993 & ~n36251;
  assign n36253 = ~pi0299 & ~n36252;
  assign n36254 = pi0039 & ~n36253;
  assign n36255 = ~n17045 & n36254;
  assign n36256 = ~pi0038 & ~n18147;
  assign n36257 = ~n36255 & n36256;
  assign n36258 = n18591 & ~n36257;
  assign n36259 = pi0222 & ~n36258;
  assign n36260 = ~n19149 & ~n36259;
  assign n36261 = pi0222 & ~n2571;
  assign n36262 = pi0222 & ~n16641;
  assign n36263 = pi0038 & ~n36262;
  assign n36264 = pi0661 & n16646;
  assign n36265 = n36263 & ~n36264;
  assign n36266 = pi0661 & pi0680;
  assign n36267 = n16918 & ~n36266;
  assign n36268 = ~pi0222 & ~n16918;
  assign n36269 = pi0222 & n16935;
  assign n36270 = ~pi0299 & ~n36269;
  assign n36271 = ~n36267 & n36270;
  assign n36272 = ~n36268 & n36271;
  assign n36273 = pi0222 & n16944;
  assign n36274 = n16923 & ~n36266;
  assign n36275 = ~pi0222 & ~n16923;
  assign n36276 = pi0299 & ~n36273;
  assign n36277 = ~n36274 & n36276;
  assign n36278 = ~n36275 & n36277;
  assign n36279 = ~pi0039 & ~n36272;
  assign n36280 = ~n36278 & n36279;
  assign n36281 = ~pi0661 & ~n17018;
  assign n36282 = pi0680 & n16758;
  assign n36283 = ~n16753 & ~n36282;
  assign n36284 = pi0661 & ~n36283;
  assign n36285 = ~n36281 & ~n36284;
  assign n36286 = ~n6205 & n36285;
  assign n36287 = ~pi0661 & n16994;
  assign n36288 = ~n6193 & ~n16776;
  assign n36289 = ~pi0662 & n16995;
  assign n36290 = ~n36288 & ~n36289;
  assign n36291 = n16656 & ~n36290;
  assign n36292 = pi0661 & ~n16786;
  assign n36293 = ~n36287 & ~n36291;
  assign n36294 = ~n36292 & n36293;
  assign n36295 = n6205 & n36294;
  assign n36296 = pi0222 & ~n36286;
  assign n36297 = ~n36295 & n36296;
  assign n36298 = ~n16690 & n36266;
  assign n36299 = n6205 & n36298;
  assign n36300 = pi0661 & n16703;
  assign n36301 = ~n6205 & n36300;
  assign n36302 = pi0224 & ~n36299;
  assign n36303 = ~n36301 & n36302;
  assign n36304 = pi0661 & n16739;
  assign n36305 = ~pi0224 & ~n36304;
  assign n36306 = ~pi0222 & ~n36305;
  assign n36307 = ~n36303 & n36306;
  assign n36308 = ~pi0223 & ~n36307;
  assign n36309 = ~n36297 & n36308;
  assign n36310 = ~pi0222 & pi0661;
  assign n36311 = n16729 & n36310;
  assign n36312 = ~pi0661 & n16960;
  assign n36313 = n16656 & n16966;
  assign n36314 = pi0661 & ~n16818;
  assign n36315 = ~n36312 & ~n36314;
  assign n36316 = ~n36313 & n36315;
  assign n36317 = ~n6205 & n36316;
  assign n36318 = ~pi0661 & ~n16990;
  assign n36319 = ~n16804 & ~n16809;
  assign n36320 = pi0661 & ~n36319;
  assign n36321 = ~n36318 & ~n36320;
  assign n36322 = n6205 & n36321;
  assign n36323 = pi0222 & ~n36317;
  assign n36324 = ~n36322 & n36323;
  assign n36325 = pi0223 & ~n36311;
  assign n36326 = ~n36324 & n36325;
  assign n36327 = ~n36309 & ~n36326;
  assign n36328 = ~pi0299 & ~n36327;
  assign n36329 = n16744 & n36310;
  assign n36330 = ~n6242 & n36316;
  assign n36331 = n6242 & n36321;
  assign n36332 = pi0222 & ~n36330;
  assign n36333 = ~n36331 & n36332;
  assign n36334 = ~n36329 & ~n36333;
  assign n36335 = pi0215 & ~n36334;
  assign n36336 = pi0222 & ~n16653;
  assign n36337 = n3448 & ~n36336;
  assign n36338 = ~n36304 & n36337;
  assign n36339 = ~n6242 & n36285;
  assign n36340 = n6242 & n36294;
  assign n36341 = pi0222 & ~n36339;
  assign n36342 = ~n36340 & n36341;
  assign n36343 = ~n6242 & ~n36300;
  assign n36344 = n6242 & ~n36298;
  assign n36345 = ~pi0222 & ~n36343;
  assign n36346 = ~n36344 & n36345;
  assign n36347 = ~n3448 & ~n36346;
  assign n36348 = ~n36342 & n36347;
  assign n36349 = ~pi0215 & ~n36338;
  assign n36350 = ~n36348 & n36349;
  assign n36351 = pi0299 & ~n36335;
  assign n36352 = ~n36350 & n36351;
  assign n36353 = ~n36328 & ~n36352;
  assign n36354 = pi0039 & ~n36353;
  assign n36355 = ~n36280 & ~n36354;
  assign n36356 = ~pi0038 & ~n36355;
  assign n36357 = n2571 & ~n36265;
  assign n36358 = ~n36356 & n36357;
  assign n36359 = ~n36261 & ~n36358;
  assign n36360 = ~pi0778 & ~n36359;
  assign n36361 = pi0625 & n36359;
  assign n36362 = ~pi0625 & ~n36259;
  assign n36363 = pi1153 & ~n36362;
  assign n36364 = ~n36361 & n36363;
  assign n36365 = ~pi0625 & n36359;
  assign n36366 = pi0625 & ~n36259;
  assign n36367 = ~pi1153 & ~n36366;
  assign n36368 = ~n36365 & n36367;
  assign n36369 = ~n36364 & ~n36368;
  assign n36370 = pi0778 & ~n36369;
  assign n36371 = ~n36360 & ~n36370;
  assign n36372 = ~n17075 & ~n36371;
  assign n36373 = n17075 & n36259;
  assign n36374 = ~n36372 & ~n36373;
  assign n36375 = ~n16639 & ~n36374;
  assign n36376 = n16639 & n36259;
  assign n36377 = ~n36375 & ~n36376;
  assign n36378 = ~n16635 & n36377;
  assign n36379 = ~n16631 & n36378;
  assign n36380 = ~n36260 & ~n36379;
  assign n36381 = ~n19142 & ~n36380;
  assign n36382 = n17856 & ~n36259;
  assign n36383 = ~n36381 & ~n36382;
  assign n36384 = ~pi0787 & n36383;
  assign n36385 = ~pi0647 & ~n36383;
  assign n36386 = pi0647 & ~n36259;
  assign n36387 = ~pi1157 & ~n36386;
  assign n36388 = ~n36385 & n36387;
  assign n36389 = pi0647 & ~n36383;
  assign n36390 = ~pi0647 & ~n36259;
  assign n36391 = pi1157 & ~n36390;
  assign n36392 = ~n36389 & n36391;
  assign n36393 = ~n36388 & ~n36392;
  assign n36394 = pi0787 & ~n36393;
  assign n36395 = ~n36384 & ~n36394;
  assign n36396 = ~pi0644 & n36395;
  assign n36397 = pi0628 & ~n36259;
  assign n36398 = ~pi0628 & ~n36380;
  assign n36399 = n17777 & ~n36397;
  assign n36400 = ~n36398 & n36399;
  assign n36401 = n17969 & ~n36259;
  assign n36402 = pi0616 & n17280;
  assign n36403 = n36263 & ~n36402;
  assign n36404 = ~pi0616 & n17233;
  assign n36405 = ~pi0222 & ~n17233;
  assign n36406 = pi0222 & n17139;
  assign n36407 = ~pi0039 & ~n36404;
  assign n36408 = ~n36405 & n36407;
  assign n36409 = ~n36406 & n36408;
  assign n36410 = ~n6195 & n17235;
  assign n36411 = ~n17236 & ~n36410;
  assign n36412 = pi0616 & ~n36411;
  assign n36413 = ~pi0222 & n36412;
  assign n36414 = ~n16743 & n36413;
  assign n36415 = pi0616 & ~n17182;
  assign n36416 = n16814 & ~n36415;
  assign n36417 = ~n16656 & ~n36416;
  assign n36418 = ~n6193 & ~n16814;
  assign n36419 = ~n16963 & ~n36415;
  assign n36420 = ~n36418 & n36419;
  assign n36421 = n16656 & ~n36420;
  assign n36422 = ~n36417 & ~n36421;
  assign n36423 = ~n6242 & n36422;
  assign n36424 = pi0616 & ~n17169;
  assign n36425 = ~n16802 & ~n36424;
  assign n36426 = ~n16656 & ~n36425;
  assign n36427 = pi0616 & n17168;
  assign n36428 = n6193 & ~n36427;
  assign n36429 = n16797 & n36428;
  assign n36430 = ~n6193 & n36425;
  assign n36431 = n16656 & ~n36429;
  assign n36432 = ~n36430 & n36431;
  assign n36433 = ~n36426 & ~n36432;
  assign n36434 = n6242 & n36433;
  assign n36435 = pi0222 & ~n36423;
  assign n36436 = ~n36434 & n36435;
  assign n36437 = ~n36414 & ~n36436;
  assign n36438 = pi0215 & ~n36437;
  assign n36439 = n16978 & n17168;
  assign n36440 = n36337 & ~n36439;
  assign n36441 = ~n16775 & ~n36424;
  assign n36442 = ~n16656 & ~n36441;
  assign n36443 = n16684 & n36428;
  assign n36444 = ~n6193 & n36441;
  assign n36445 = n16656 & ~n36443;
  assign n36446 = ~n36444 & n36445;
  assign n36447 = ~n36442 & ~n36446;
  assign n36448 = n6242 & n36447;
  assign n36449 = pi0616 & ~n17154;
  assign n36450 = ~pi0616 & n36187;
  assign n36451 = ~n36449 & ~n36450;
  assign n36452 = ~n16656 & ~n36451;
  assign n36453 = n17147 & ~n36427;
  assign n36454 = ~n17145 & ~n36453;
  assign n36455 = n6193 & ~n36454;
  assign n36456 = ~n6193 & n36451;
  assign n36457 = n16656 & ~n36455;
  assign n36458 = ~n36456 & n36457;
  assign n36459 = ~n36452 & ~n36458;
  assign n36460 = ~n6242 & n36459;
  assign n36461 = pi0222 & ~n36448;
  assign n36462 = ~n36460 & n36461;
  assign n36463 = ~n17247 & ~n36410;
  assign n36464 = pi0616 & ~n36463;
  assign n36465 = n6242 & ~n36464;
  assign n36466 = ~n16699 & n36427;
  assign n36467 = ~n16656 & ~n36466;
  assign n36468 = pi0616 & n6193;
  assign n36469 = n17375 & n36468;
  assign n36470 = ~n6193 & n36466;
  assign n36471 = n16656 & ~n36469;
  assign n36472 = ~n36470 & n36471;
  assign n36473 = ~n36467 & ~n36472;
  assign n36474 = ~n6242 & ~n36473;
  assign n36475 = ~pi0222 & ~n36465;
  assign n36476 = ~n36474 & n36475;
  assign n36477 = ~n3448 & ~n36476;
  assign n36478 = ~n36462 & n36477;
  assign n36479 = ~pi0215 & ~n36440;
  assign n36480 = ~n36478 & n36479;
  assign n36481 = pi0299 & ~n36438;
  assign n36482 = ~n36480 & n36481;
  assign n36483 = n6205 & n36464;
  assign n36484 = ~n6205 & n36473;
  assign n36485 = pi0224 & ~n36483;
  assign n36486 = ~n36484 & n36485;
  assign n36487 = ~pi0224 & ~n36439;
  assign n36488 = ~pi0222 & ~n36487;
  assign n36489 = ~n36486 & n36488;
  assign n36490 = n6205 & n36447;
  assign n36491 = ~n6205 & n36459;
  assign n36492 = pi0222 & ~n36490;
  assign n36493 = ~n36491 & n36492;
  assign n36494 = ~pi0223 & ~n36489;
  assign n36495 = ~n36493 & n36494;
  assign n36496 = ~n16724 & n36413;
  assign n36497 = ~n6205 & n36422;
  assign n36498 = n6205 & n36433;
  assign n36499 = pi0222 & ~n36497;
  assign n36500 = ~n36498 & n36499;
  assign n36501 = pi0223 & ~n36496;
  assign n36502 = ~n36500 & n36501;
  assign n36503 = ~n36495 & ~n36502;
  assign n36504 = ~pi0299 & ~n36503;
  assign n36505 = pi0039 & ~n36482;
  assign n36506 = ~n36504 & n36505;
  assign n36507 = ~pi0038 & ~n36409;
  assign n36508 = ~n36506 & n36507;
  assign n36509 = n2571 & ~n36403;
  assign n36510 = ~n36508 & n36509;
  assign n36511 = ~n36261 & ~n36510;
  assign n36512 = ~n17117 & ~n36511;
  assign n36513 = n17117 & n36259;
  assign n36514 = ~n36512 & ~n36513;
  assign n36515 = ~pi0785 & ~n36514;
  assign n36516 = pi0609 & n36514;
  assign n36517 = ~pi0609 & ~n36259;
  assign n36518 = pi1155 & ~n36517;
  assign n36519 = ~n36516 & n36518;
  assign n36520 = ~pi0609 & n36514;
  assign n36521 = pi0609 & ~n36259;
  assign n36522 = ~pi1155 & ~n36521;
  assign n36523 = ~n36520 & n36522;
  assign n36524 = ~n36519 & ~n36523;
  assign n36525 = pi0785 & ~n36524;
  assign n36526 = ~n36515 & ~n36525;
  assign n36527 = ~pi0781 & ~n36526;
  assign n36528 = pi0618 & n36526;
  assign n36529 = ~pi0618 & ~n36259;
  assign n36530 = pi1154 & ~n36529;
  assign n36531 = ~n36528 & n36530;
  assign n36532 = ~pi0618 & n36526;
  assign n36533 = pi0618 & ~n36259;
  assign n36534 = ~pi1154 & ~n36533;
  assign n36535 = ~n36532 & n36534;
  assign n36536 = ~n36531 & ~n36535;
  assign n36537 = pi0781 & ~n36536;
  assign n36538 = ~n36527 & ~n36537;
  assign n36539 = ~pi0789 & ~n36538;
  assign n36540 = pi0619 & n36538;
  assign n36541 = ~pi0619 & ~n36259;
  assign n36542 = pi1159 & ~n36541;
  assign n36543 = ~n36540 & n36542;
  assign n36544 = ~pi0619 & n36538;
  assign n36545 = pi0619 & ~n36259;
  assign n36546 = ~pi1159 & ~n36545;
  assign n36547 = ~n36544 & n36546;
  assign n36548 = ~n36543 & ~n36547;
  assign n36549 = pi0789 & ~n36548;
  assign n36550 = ~n36539 & ~n36549;
  assign n36551 = ~n17969 & n36550;
  assign n36552 = ~n36401 & ~n36551;
  assign n36553 = ~n20570 & n36552;
  assign n36554 = ~pi0628 & ~n36259;
  assign n36555 = pi0628 & ~n36380;
  assign n36556 = n17776 & ~n36554;
  assign n36557 = ~n36555 & n36556;
  assign n36558 = ~n36400 & ~n36557;
  assign n36559 = ~n36553 & n36558;
  assign n36560 = pi0792 & ~n36559;
  assign n36561 = pi0609 & n36371;
  assign n36562 = n16667 & n17493;
  assign n36563 = ~pi0222 & ~pi0616;
  assign n36564 = ~pi0039 & pi0616;
  assign n36565 = n36266 & n36564;
  assign n36566 = ~n36563 & ~n36565;
  assign n36567 = n36562 & ~n36566;
  assign n36568 = ~n36266 & ~n36427;
  assign n36569 = ~pi0616 & ~n17355;
  assign n36570 = ~n36568 & ~n36569;
  assign n36571 = n16641 & n36570;
  assign n36572 = ~n36262 & ~n36571;
  assign n36573 = ~n36567 & ~n36572;
  assign n36574 = pi0038 & ~n36573;
  assign n36575 = ~pi0661 & pi0681;
  assign n36576 = ~n36425 & n36575;
  assign n36577 = ~pi0680 & n36425;
  assign n36578 = pi0616 & ~n17504;
  assign n36579 = pi0680 & ~n36578;
  assign n36580 = ~n17347 & n36579;
  assign n36581 = pi0661 & ~n36577;
  assign n36582 = ~n36580 & n36581;
  assign n36583 = ~n36432 & ~n36576;
  assign n36584 = ~n36582 & n36583;
  assign n36585 = n6242 & ~n36584;
  assign n36586 = ~n36416 & n36575;
  assign n36587 = ~pi0680 & n36416;
  assign n36588 = ~n17324 & n17493;
  assign n36589 = pi0616 & ~n36588;
  assign n36590 = pi0680 & ~n36589;
  assign n36591 = n17330 & n36590;
  assign n36592 = pi0661 & ~n36591;
  assign n36593 = ~n36587 & n36592;
  assign n36594 = ~n36421 & ~n36586;
  assign n36595 = ~n36593 & n36594;
  assign n36596 = ~n6242 & ~n36595;
  assign n36597 = pi0222 & ~n36585;
  assign n36598 = ~n36596 & n36597;
  assign n36599 = n17444 & n36266;
  assign n36600 = ~n36412 & ~n36599;
  assign n36601 = n6242 & ~n36600;
  assign n36602 = pi0616 & n17237;
  assign n36603 = ~pi0661 & ~n36602;
  assign n36604 = ~n16721 & n36439;
  assign n36605 = n6195 & ~n36604;
  assign n36606 = ~pi0680 & n36602;
  assign n36607 = ~n17237 & ~n17559;
  assign n36608 = pi0616 & n36607;
  assign n36609 = pi0680 & ~n36608;
  assign n36610 = n17458 & n36609;
  assign n36611 = pi0661 & ~n36606;
  assign n36612 = ~n36610 & n36611;
  assign n36613 = ~n36603 & ~n36605;
  assign n36614 = ~n36612 & n36613;
  assign n36615 = ~n6242 & n36614;
  assign n36616 = ~pi0222 & ~n36601;
  assign n36617 = ~n36615 & n36616;
  assign n36618 = pi0215 & ~n36617;
  assign n36619 = ~n36598 & n36618;
  assign n36620 = pi0616 & ~n17548;
  assign n36621 = ~pi0616 & ~n17407;
  assign n36622 = ~n36620 & ~n36621;
  assign n36623 = ~n36568 & n36622;
  assign n36624 = n36337 & ~n36623;
  assign n36625 = ~n36451 & n36575;
  assign n36626 = pi0603 & n16681;
  assign n36627 = n6197 & n16754;
  assign n36628 = ~n16756 & ~n36627;
  assign n36629 = ~pi0603 & n36628;
  assign n36630 = ~n17368 & ~n36626;
  assign n36631 = ~n36629 & n36630;
  assign n36632 = ~pi0642 & n36631;
  assign n36633 = ~n17577 & n36628;
  assign n36634 = pi0642 & ~n36633;
  assign n36635 = n6191 & ~n36632;
  assign n36636 = ~n36634 & n36635;
  assign n36637 = n17452 & n36633;
  assign n36638 = n17493 & ~n36628;
  assign n36639 = pi0616 & ~n36638;
  assign n36640 = pi0680 & ~n36639;
  assign n36641 = ~n36637 & n36640;
  assign n36642 = ~n36636 & n36641;
  assign n36643 = ~pi0680 & n36451;
  assign n36644 = pi0661 & ~n36642;
  assign n36645 = ~n36643 & n36644;
  assign n36646 = ~n36458 & ~n36625;
  assign n36647 = ~n36645 & n36646;
  assign n36648 = ~n6242 & ~n36647;
  assign n36649 = ~n36441 & n36575;
  assign n36650 = ~pi0680 & n36441;
  assign n36651 = ~n17363 & n36579;
  assign n36652 = pi0661 & ~n36650;
  assign n36653 = ~n36651 & n36652;
  assign n36654 = ~n36446 & ~n36649;
  assign n36655 = ~n36653 & n36654;
  assign n36656 = n6242 & ~n36655;
  assign n36657 = pi0222 & ~n36656;
  assign n36658 = ~n36648 & n36657;
  assign n36659 = ~n36466 & n36575;
  assign n36660 = ~pi0680 & n36466;
  assign n36661 = pi0616 & n17578;
  assign n36662 = pi0680 & ~n36661;
  assign n36663 = ~n17433 & n36662;
  assign n36664 = pi0661 & ~n36660;
  assign n36665 = ~n36663 & n36664;
  assign n36666 = ~n36472 & ~n36659;
  assign n36667 = ~n36665 & n36666;
  assign n36668 = ~n6242 & n36667;
  assign n36669 = ~n6193 & n36439;
  assign n36670 = n17246 & n36468;
  assign n36671 = n16656 & ~n36669;
  assign n36672 = ~n36670 & n36671;
  assign n36673 = ~n36439 & n36575;
  assign n36674 = ~pi0680 & n36439;
  assign n36675 = pi0680 & ~n17417;
  assign n36676 = ~n36620 & n36675;
  assign n36677 = pi0661 & ~n36674;
  assign n36678 = ~n36676 & n36677;
  assign n36679 = ~n36672 & ~n36673;
  assign n36680 = ~n36678 & n36679;
  assign n36681 = n6242 & n36680;
  assign n36682 = ~pi0222 & ~n36681;
  assign n36683 = ~n36668 & n36682;
  assign n36684 = ~n36658 & ~n36683;
  assign n36685 = ~n3448 & ~n36684;
  assign n36686 = ~pi0215 & ~n36624;
  assign n36687 = ~n36685 & n36686;
  assign n36688 = pi0299 & ~n36619;
  assign n36689 = ~n36687 & n36688;
  assign n36690 = n36266 & ~n36622;
  assign n36691 = ~n36266 & ~n36439;
  assign n36692 = ~pi0222 & ~n36691;
  assign n36693 = ~n36690 & n36692;
  assign n36694 = ~n3351 & ~n36693;
  assign n36695 = ~n6205 & n36667;
  assign n36696 = n6205 & n36680;
  assign n36697 = pi0224 & ~n36696;
  assign n36698 = ~n36695 & n36697;
  assign n36699 = ~n36694 & ~n36698;
  assign n36700 = n6205 & n36655;
  assign n36701 = ~n6205 & n36647;
  assign n36702 = pi0222 & ~n36700;
  assign n36703 = ~n36701 & n36702;
  assign n36704 = ~n36699 & ~n36703;
  assign n36705 = ~pi0223 & ~n36704;
  assign n36706 = n6205 & ~n36584;
  assign n36707 = ~n6205 & ~n36595;
  assign n36708 = pi0222 & ~n36706;
  assign n36709 = ~n36707 & n36708;
  assign n36710 = n6205 & ~n36600;
  assign n36711 = ~n6205 & n36614;
  assign n36712 = ~pi0222 & ~n36710;
  assign n36713 = ~n36711 & n36712;
  assign n36714 = pi0223 & ~n36713;
  assign n36715 = ~n36709 & n36714;
  assign n36716 = ~pi0299 & ~n36715;
  assign n36717 = ~n36705 & n36716;
  assign n36718 = pi0039 & ~n36717;
  assign n36719 = ~n36689 & n36718;
  assign n36720 = pi0661 & n17618;
  assign n36721 = pi0616 & n17226;
  assign n36722 = ~pi0222 & ~n36721;
  assign n36723 = ~n36720 & n36722;
  assign n36724 = ~pi0616 & n17226;
  assign n36725 = n17617 & ~n36266;
  assign n36726 = ~pi0603 & ~n16935;
  assign n36727 = ~n17367 & ~n17614;
  assign n36728 = ~n36726 & n36727;
  assign n36729 = ~n36724 & ~n36728;
  assign n36730 = ~n36725 & n36729;
  assign n36731 = pi0222 & ~n36730;
  assign n36732 = ~n36723 & ~n36731;
  assign n36733 = ~pi0299 & ~n36732;
  assign n36734 = ~pi0616 & n17231;
  assign n36735 = n17622 & ~n36266;
  assign n36736 = ~pi0603 & ~n16944;
  assign n36737 = ~n17123 & ~n17367;
  assign n36738 = ~n36736 & n36737;
  assign n36739 = ~n36734 & ~n36738;
  assign n36740 = ~n36735 & n36739;
  assign n36741 = pi0222 & ~n36740;
  assign n36742 = pi0661 & n17623;
  assign n36743 = pi0616 & n17231;
  assign n36744 = ~pi0222 & ~n36743;
  assign n36745 = ~n36742 & n36744;
  assign n36746 = ~n36741 & ~n36745;
  assign n36747 = pi0299 & ~n36746;
  assign n36748 = ~pi0039 & ~n36733;
  assign n36749 = ~n36747 & n36748;
  assign n36750 = ~pi0038 & ~n36749;
  assign n36751 = ~n36719 & n36750;
  assign n36752 = n2571 & ~n36574;
  assign n36753 = ~n36751 & n36752;
  assign n36754 = ~n36261 & ~n36753;
  assign n36755 = ~pi0625 & n36754;
  assign n36756 = pi0625 & n36511;
  assign n36757 = ~pi1153 & ~n36756;
  assign n36758 = ~n36755 & n36757;
  assign n36759 = ~pi0608 & ~n36364;
  assign n36760 = ~n36758 & n36759;
  assign n36761 = ~pi0625 & n36511;
  assign n36762 = pi0625 & n36754;
  assign n36763 = pi1153 & ~n36761;
  assign n36764 = ~n36762 & n36763;
  assign n36765 = pi0608 & ~n36368;
  assign n36766 = ~n36764 & n36765;
  assign n36767 = ~n36760 & ~n36766;
  assign n36768 = pi0778 & ~n36767;
  assign n36769 = ~pi0778 & n36754;
  assign n36770 = ~n36768 & ~n36769;
  assign n36771 = ~pi0609 & ~n36770;
  assign n36772 = ~pi1155 & ~n36561;
  assign n36773 = ~n36771 & n36772;
  assign n36774 = ~pi0660 & ~n36519;
  assign n36775 = ~n36773 & n36774;
  assign n36776 = ~pi0609 & n36371;
  assign n36777 = pi0609 & ~n36770;
  assign n36778 = pi1155 & ~n36776;
  assign n36779 = ~n36777 & n36778;
  assign n36780 = pi0660 & ~n36523;
  assign n36781 = ~n36779 & n36780;
  assign n36782 = ~n36775 & ~n36781;
  assign n36783 = pi0785 & ~n36782;
  assign n36784 = ~pi0785 & ~n36770;
  assign n36785 = ~n36783 & ~n36784;
  assign n36786 = ~pi0618 & ~n36785;
  assign n36787 = pi0618 & n36374;
  assign n36788 = ~pi1154 & ~n36787;
  assign n36789 = ~n36786 & n36788;
  assign n36790 = ~pi0627 & ~n36531;
  assign n36791 = ~n36789 & n36790;
  assign n36792 = ~pi0618 & n36374;
  assign n36793 = pi0618 & ~n36785;
  assign n36794 = pi1154 & ~n36792;
  assign n36795 = ~n36793 & n36794;
  assign n36796 = pi0627 & ~n36535;
  assign n36797 = ~n36795 & n36796;
  assign n36798 = ~n36791 & ~n36797;
  assign n36799 = pi0781 & ~n36798;
  assign n36800 = ~pi0781 & ~n36785;
  assign n36801 = ~n36799 & ~n36800;
  assign n36802 = ~pi0789 & n36801;
  assign n36803 = ~pi0626 & n36550;
  assign n36804 = pi0626 & ~n36259;
  assign n36805 = n16629 & ~n36804;
  assign n36806 = ~n36803 & n36805;
  assign n36807 = n16635 & ~n36259;
  assign n36808 = n17871 & ~n36807;
  assign n36809 = ~n36378 & n36808;
  assign n36810 = pi0626 & n36550;
  assign n36811 = ~pi0626 & ~n36259;
  assign n36812 = n16628 & ~n36811;
  assign n36813 = ~n36810 & n36812;
  assign n36814 = ~n36806 & ~n36809;
  assign n36815 = ~n36813 & n36814;
  assign n36816 = pi0788 & ~n36815;
  assign n36817 = ~pi0619 & ~n36801;
  assign n36818 = pi0619 & n36377;
  assign n36819 = ~pi1159 & ~n36818;
  assign n36820 = ~n36817 & n36819;
  assign n36821 = ~pi0648 & ~n36543;
  assign n36822 = ~n36820 & n36821;
  assign n36823 = pi0619 & ~n36801;
  assign n36824 = ~pi0619 & n36377;
  assign n36825 = pi1159 & ~n36824;
  assign n36826 = ~n36823 & n36825;
  assign n36827 = pi0648 & ~n36547;
  assign n36828 = ~n36826 & n36827;
  assign n36829 = pi0789 & ~n36822;
  assign n36830 = ~n36828 & n36829;
  assign n36831 = ~n36802 & ~n36816;
  assign n36832 = ~n36830 & n36831;
  assign n36833 = ~n17970 & n36815;
  assign n36834 = ~n20364 & ~n36833;
  assign n36835 = ~n36832 & n36834;
  assign n36836 = ~n36560 & ~n36835;
  assign n36837 = ~n20206 & ~n36836;
  assign n36838 = ~pi0630 & n36392;
  assign n36839 = ~n17779 & n36552;
  assign n36840 = n17779 & n36259;
  assign n36841 = ~n36839 & ~n36840;
  assign n36842 = ~n20559 & ~n36841;
  assign n36843 = pi0630 & n36388;
  assign n36844 = ~n36838 & ~n36843;
  assign n36845 = ~n36842 & n36844;
  assign n36846 = pi0787 & ~n36845;
  assign n36847 = ~n36837 & ~n36846;
  assign n36848 = pi0644 & n36847;
  assign n36849 = pi0715 & ~n36396;
  assign n36850 = ~n36848 & n36849;
  assign n36851 = n17804 & ~n36259;
  assign n36852 = ~n17804 & n36841;
  assign n36853 = ~n36851 & ~n36852;
  assign n36854 = pi0644 & ~n36853;
  assign n36855 = ~pi0644 & ~n36259;
  assign n36856 = ~pi0715 & ~n36855;
  assign n36857 = ~n36854 & n36856;
  assign n36858 = pi1160 & ~n36857;
  assign n36859 = ~n36850 & n36858;
  assign n36860 = pi0644 & n36395;
  assign n36861 = ~pi0644 & n36847;
  assign n36862 = ~pi0715 & ~n36860;
  assign n36863 = ~n36861 & n36862;
  assign n36864 = ~pi0644 & ~n36853;
  assign n36865 = pi0644 & ~n36259;
  assign n36866 = pi0715 & ~n36865;
  assign n36867 = ~n36864 & n36866;
  assign n36868 = ~pi1160 & ~n36867;
  assign n36869 = ~n36863 & n36868;
  assign n36870 = ~n36859 & ~n36869;
  assign n36871 = pi0790 & ~n36870;
  assign n36872 = ~pi0790 & n36847;
  assign n36873 = ~n36871 & ~n36872;
  assign n36874 = ~po1038 & ~n36873;
  assign n36875 = ~pi0222 & po1038;
  assign po0379 = ~n36874 & ~n36875;
  assign n36877 = ~pi0299 & ~n16992;
  assign n36878 = pi0039 & ~n36877;
  assign n36879 = ~n17045 & n36878;
  assign n36880 = n14873 & ~n18147;
  assign n36881 = ~n36879 & n36880;
  assign n36882 = n18591 & ~n36881;
  assign n36883 = pi0223 & ~n36882;
  assign n36884 = ~n19149 & ~n36883;
  assign n36885 = n17075 & ~n36883;
  assign n36886 = pi0223 & ~n2571;
  assign n36887 = pi0680 & pi0681;
  assign n36888 = n16918 & ~n36887;
  assign n36889 = ~pi0223 & ~n16918;
  assign n36890 = pi0223 & n16935;
  assign n36891 = ~pi0299 & ~n36890;
  assign n36892 = ~n36888 & n36891;
  assign n36893 = ~n36889 & n36892;
  assign n36894 = pi0223 & n16944;
  assign n36895 = n16923 & ~n36887;
  assign n36896 = ~pi0223 & ~n16923;
  assign n36897 = pi0299 & ~n36894;
  assign n36898 = ~n36895 & n36897;
  assign n36899 = ~n36896 & n36898;
  assign n36900 = ~pi0039 & ~n36893;
  assign n36901 = ~n36899 & n36900;
  assign n36902 = pi0681 & n16739;
  assign n36903 = n2603 & ~n36902;
  assign n36904 = ~n16690 & n36887;
  assign n36905 = n6205 & n36904;
  assign n36906 = pi0681 & n16703;
  assign n36907 = ~n6205 & n36906;
  assign n36908 = ~n2603 & ~n36905;
  assign n36909 = ~n36907 & n36908;
  assign n36910 = ~n36903 & ~n36909;
  assign n36911 = ~pi0223 & ~n36910;
  assign n36912 = pi0681 & ~n36319;
  assign n36913 = ~n16989 & ~n36912;
  assign n36914 = n6205 & ~n36913;
  assign n36915 = pi0681 & ~n16818;
  assign n36916 = ~n16969 & ~n36915;
  assign n36917 = ~n6205 & ~n36916;
  assign n36918 = pi0223 & ~n36914;
  assign n36919 = ~n36917 & n36918;
  assign n36920 = ~pi0299 & ~n36919;
  assign n36921 = ~n36911 & n36920;
  assign n36922 = ~pi0223 & pi0681;
  assign n36923 = n16744 & n36922;
  assign n36924 = n6242 & n36913;
  assign n36925 = ~n6242 & n36916;
  assign n36926 = pi0223 & ~n36924;
  assign n36927 = ~n36925 & n36926;
  assign n36928 = pi0215 & ~n36923;
  assign n36929 = ~n36927 & n36928;
  assign n36930 = pi0223 & ~n16653;
  assign n36931 = n3448 & ~n36930;
  assign n36932 = ~n36902 & n36931;
  assign n36933 = pi0681 & ~n36283;
  assign n36934 = ~n6242 & ~n17017;
  assign n36935 = ~n36933 & n36934;
  assign n36936 = pi0681 & ~n16786;
  assign n36937 = n6242 & ~n17010;
  assign n36938 = ~n36936 & n36937;
  assign n36939 = pi0223 & ~n36935;
  assign n36940 = ~n36938 & n36939;
  assign n36941 = ~n6242 & ~n36906;
  assign n36942 = n6242 & ~n36904;
  assign n36943 = ~pi0223 & ~n36941;
  assign n36944 = ~n36942 & n36943;
  assign n36945 = ~n3448 & ~n36944;
  assign n36946 = ~n36940 & n36945;
  assign n36947 = ~n36932 & ~n36946;
  assign n36948 = ~pi0215 & ~n36947;
  assign n36949 = pi0299 & ~n36929;
  assign n36950 = ~n36948 & n36949;
  assign n36951 = pi0039 & ~n36921;
  assign n36952 = ~n36950 & n36951;
  assign n36953 = ~n36901 & ~n36952;
  assign n36954 = ~pi0038 & ~n36953;
  assign n36955 = pi0681 & n16646;
  assign n36956 = pi0223 & ~n16641;
  assign n36957 = pi0038 & ~n36955;
  assign n36958 = ~n36956 & n36957;
  assign n36959 = n2571 & ~n36958;
  assign n36960 = ~n36954 & n36959;
  assign n36961 = ~n36886 & ~n36960;
  assign n36962 = ~pi0778 & ~n36961;
  assign n36963 = pi0625 & n36961;
  assign n36964 = ~pi0625 & ~n36883;
  assign n36965 = pi1153 & ~n36964;
  assign n36966 = ~n36963 & n36965;
  assign n36967 = ~pi0625 & n36961;
  assign n36968 = pi0625 & ~n36883;
  assign n36969 = ~pi1153 & ~n36968;
  assign n36970 = ~n36967 & n36969;
  assign n36971 = ~n36966 & ~n36970;
  assign n36972 = pi0778 & ~n36971;
  assign n36973 = ~n36962 & ~n36972;
  assign n36974 = ~n17075 & n36973;
  assign n36975 = ~n36885 & ~n36974;
  assign n36976 = ~n16639 & n36975;
  assign n36977 = n16639 & n36883;
  assign n36978 = ~n36976 & ~n36977;
  assign n36979 = ~n16635 & n36978;
  assign n36980 = ~n16631 & n36979;
  assign n36981 = ~n36884 & ~n36980;
  assign n36982 = ~n19142 & ~n36981;
  assign n36983 = n17856 & ~n36883;
  assign n36984 = ~n36982 & ~n36983;
  assign n36985 = ~pi0787 & n36984;
  assign n36986 = ~pi0647 & ~n36984;
  assign n36987 = pi0647 & ~n36883;
  assign n36988 = ~pi1157 & ~n36987;
  assign n36989 = ~n36986 & n36988;
  assign n36990 = pi0647 & ~n36984;
  assign n36991 = ~pi0647 & ~n36883;
  assign n36992 = pi1157 & ~n36991;
  assign n36993 = ~n36990 & n36992;
  assign n36994 = ~n36989 & ~n36993;
  assign n36995 = pi0787 & ~n36994;
  assign n36996 = ~n36985 & ~n36995;
  assign n36997 = ~pi0644 & n36996;
  assign n36998 = ~pi0630 & n36993;
  assign n36999 = n17969 & ~n36883;
  assign n37000 = n17117 & ~n36883;
  assign n37001 = pi0039 & pi0223;
  assign n37002 = pi0038 & ~n37001;
  assign n37003 = pi0642 & n17168;
  assign n37004 = n16667 & ~n37003;
  assign n37005 = ~pi0223 & ~n16667;
  assign n37006 = ~pi0039 & ~n37005;
  assign n37007 = ~n37004 & n37006;
  assign n37008 = n37002 & ~n37007;
  assign n37009 = ~pi0223 & pi0642;
  assign n37010 = n17226 & n37009;
  assign n37011 = ~pi0299 & ~n37010;
  assign n37012 = ~pi0642 & n17226;
  assign n37013 = pi0223 & ~n37012;
  assign n37014 = n17137 & n37013;
  assign n37015 = n37011 & ~n37014;
  assign n37016 = n17231 & n37009;
  assign n37017 = pi0299 & ~n37016;
  assign n37018 = n6190 & n17230;
  assign n37019 = pi0223 & ~n17124;
  assign n37020 = ~n37018 & n37019;
  assign n37021 = n37017 & ~n37020;
  assign n37022 = ~pi0039 & ~n37021;
  assign n37023 = ~n37015 & n37022;
  assign n37024 = n35897 & ~n37003;
  assign n37025 = pi0642 & ~n17169;
  assign n37026 = n36425 & ~n37025;
  assign n37027 = ~n37024 & ~n37026;
  assign n37028 = pi0681 & n37027;
  assign n37029 = n6194 & n37004;
  assign n37030 = n16797 & n37029;
  assign n37031 = ~n6194 & ~n37027;
  assign n37032 = ~pi0681 & ~n37030;
  assign n37033 = ~n37031 & n37032;
  assign n37034 = ~n37028 & ~n37033;
  assign n37035 = n6205 & n37034;
  assign n37036 = ~pi0642 & ~n16814;
  assign n37037 = pi0642 & ~n17183;
  assign n37038 = ~n37036 & ~n37037;
  assign n37039 = ~n6194 & n37038;
  assign n37040 = pi0642 & ~n17182;
  assign n37041 = n6194 & ~n37040;
  assign n37042 = ~n16721 & n37041;
  assign n37043 = ~pi0681 & ~n37042;
  assign n37044 = ~n37039 & n37043;
  assign n37045 = pi0681 & ~n37038;
  assign n37046 = ~n37044 & ~n37045;
  assign n37047 = ~n6205 & n37046;
  assign n37048 = pi0223 & ~n37047;
  assign n37049 = ~n37035 & n37048;
  assign n37050 = pi0642 & n17235;
  assign n37051 = n2603 & ~n37050;
  assign n37052 = ~n6194 & n37050;
  assign n37053 = ~pi0681 & ~n37052;
  assign n37054 = pi0642 & n6194;
  assign n37055 = n17246 & n37054;
  assign n37056 = n37053 & ~n37055;
  assign n37057 = pi0681 & ~n37050;
  assign n37058 = ~n37056 & ~n37057;
  assign n37059 = n6205 & n37058;
  assign n37060 = ~n16699 & n37003;
  assign n37061 = pi0681 & ~n37060;
  assign n37062 = n17375 & n37054;
  assign n37063 = ~n6194 & n37060;
  assign n37064 = ~pi0681 & ~n37062;
  assign n37065 = ~n37063 & n37064;
  assign n37066 = ~n37061 & ~n37065;
  assign n37067 = ~n6205 & n37066;
  assign n37068 = ~n2603 & ~n37059;
  assign n37069 = ~n37067 & n37068;
  assign n37070 = ~pi0223 & ~n37051;
  assign n37071 = ~n37069 & n37070;
  assign n37072 = ~pi0299 & ~n37049;
  assign n37073 = ~n37071 & n37072;
  assign n37074 = n17236 & n37054;
  assign n37075 = n37053 & ~n37074;
  assign n37076 = n16723 & n37043;
  assign n37077 = ~n37075 & ~n37076;
  assign n37078 = pi0642 & n17237;
  assign n37079 = pi0681 & ~n37078;
  assign n37080 = n37077 & ~n37079;
  assign n37081 = pi0947 & ~n37080;
  assign n37082 = n6242 & ~n37075;
  assign n37083 = n37050 & n37082;
  assign n37084 = ~n20923 & n37080;
  assign n37085 = ~pi0947 & ~n37083;
  assign n37086 = ~n37084 & n37085;
  assign n37087 = ~pi0223 & ~n37081;
  assign n37088 = ~n37086 & n37087;
  assign n37089 = ~n6242 & n37046;
  assign n37090 = n6242 & n37034;
  assign n37091 = pi0223 & ~n37089;
  assign n37092 = ~n37090 & n37091;
  assign n37093 = ~n37088 & ~n37092;
  assign n37094 = pi0215 & ~n37093;
  assign n37095 = n36931 & ~n37050;
  assign n37096 = pi0947 & ~n37066;
  assign n37097 = n20923 & n37058;
  assign n37098 = ~n20923 & n37066;
  assign n37099 = ~pi0947 & ~n37097;
  assign n37100 = ~n37098 & n37099;
  assign n37101 = ~pi0223 & ~n37096;
  assign n37102 = ~n37100 & n37101;
  assign n37103 = pi0642 & ~n17154;
  assign n37104 = ~pi0642 & ~n16702;
  assign n37105 = ~n37103 & ~n37104;
  assign n37106 = pi0681 & ~n37105;
  assign n37107 = ~n6194 & n37105;
  assign n37108 = n17014 & ~n37003;
  assign n37109 = ~pi0681 & ~n37108;
  assign n37110 = ~n37107 & n37109;
  assign n37111 = ~n6242 & ~n37110;
  assign n37112 = ~n37106 & n37111;
  assign n37113 = n6191 & ~n37025;
  assign n37114 = ~n16770 & n37113;
  assign n37115 = ~n37024 & ~n37114;
  assign n37116 = pi0681 & n37115;
  assign n37117 = ~n6194 & ~n37115;
  assign n37118 = ~n17164 & ~n35894;
  assign n37119 = n6194 & ~n37118;
  assign n37120 = ~pi0681 & ~n37119;
  assign n37121 = ~n37117 & n37120;
  assign n37122 = n6242 & ~n37121;
  assign n37123 = ~n37116 & n37122;
  assign n37124 = pi0223 & ~n37112;
  assign n37125 = ~n37123 & n37124;
  assign n37126 = ~n3448 & ~n37102;
  assign n37127 = ~n37125 & n37126;
  assign n37128 = ~pi0215 & ~n37095;
  assign n37129 = ~n37127 & n37128;
  assign n37130 = pi0299 & ~n37094;
  assign n37131 = ~n37129 & n37130;
  assign n37132 = pi0039 & ~n37073;
  assign n37133 = ~n37131 & n37132;
  assign n37134 = ~pi0038 & ~n37023;
  assign n37135 = ~n37133 & n37134;
  assign n37136 = n2571 & ~n37008;
  assign n37137 = ~n37135 & n37136;
  assign n37138 = ~n36886 & ~n37137;
  assign n37139 = ~n17117 & n37138;
  assign n37140 = ~n37000 & ~n37139;
  assign n37141 = ~pi0785 & n37140;
  assign n37142 = pi0609 & ~n37140;
  assign n37143 = ~pi0609 & ~n36883;
  assign n37144 = pi1155 & ~n37143;
  assign n37145 = ~n37142 & n37144;
  assign n37146 = ~pi0609 & ~n37140;
  assign n37147 = pi0609 & ~n36883;
  assign n37148 = ~pi1155 & ~n37147;
  assign n37149 = ~n37146 & n37148;
  assign n37150 = ~n37145 & ~n37149;
  assign n37151 = pi0785 & ~n37150;
  assign n37152 = ~n37141 & ~n37151;
  assign n37153 = ~pi0781 & ~n37152;
  assign n37154 = pi0618 & n37152;
  assign n37155 = ~pi0618 & ~n36883;
  assign n37156 = pi1154 & ~n37155;
  assign n37157 = ~n37154 & n37156;
  assign n37158 = ~pi0618 & n37152;
  assign n37159 = pi0618 & ~n36883;
  assign n37160 = ~pi1154 & ~n37159;
  assign n37161 = ~n37158 & n37160;
  assign n37162 = ~n37157 & ~n37161;
  assign n37163 = pi0781 & ~n37162;
  assign n37164 = ~n37153 & ~n37163;
  assign n37165 = ~pi0789 & ~n37164;
  assign n37166 = pi0619 & n37164;
  assign n37167 = ~pi0619 & ~n36883;
  assign n37168 = pi1159 & ~n37167;
  assign n37169 = ~n37166 & n37168;
  assign n37170 = ~pi0619 & n37164;
  assign n37171 = pi0619 & ~n36883;
  assign n37172 = ~pi1159 & ~n37171;
  assign n37173 = ~n37170 & n37172;
  assign n37174 = ~n37169 & ~n37173;
  assign n37175 = pi0789 & ~n37174;
  assign n37176 = ~n37165 & ~n37175;
  assign n37177 = ~n17969 & n37176;
  assign n37178 = ~n36999 & ~n37177;
  assign n37179 = ~n17779 & n37178;
  assign n37180 = n17779 & n36883;
  assign n37181 = ~n37179 & ~n37180;
  assign n37182 = ~n20559 & ~n37181;
  assign n37183 = pi0630 & n36989;
  assign n37184 = ~n36998 & ~n37183;
  assign n37185 = ~n37182 & n37184;
  assign n37186 = pi0787 & ~n37185;
  assign n37187 = pi0628 & ~n36883;
  assign n37188 = ~pi0628 & ~n36981;
  assign n37189 = n17777 & ~n37187;
  assign n37190 = ~n37188 & n37189;
  assign n37191 = ~n20570 & n37178;
  assign n37192 = ~pi0628 & ~n36883;
  assign n37193 = pi0628 & ~n36981;
  assign n37194 = n17776 & ~n37192;
  assign n37195 = ~n37193 & n37194;
  assign n37196 = ~n37190 & ~n37195;
  assign n37197 = ~n37191 & n37196;
  assign n37198 = pi0792 & ~n37197;
  assign n37199 = n16635 & ~n36883;
  assign n37200 = ~n36979 & ~n37199;
  assign n37201 = n17871 & ~n37200;
  assign n37202 = ~pi0626 & n36883;
  assign n37203 = pi0626 & ~n37176;
  assign n37204 = n16628 & ~n37202;
  assign n37205 = ~n37203 & n37204;
  assign n37206 = pi0626 & n36883;
  assign n37207 = ~pi0626 & ~n37176;
  assign n37208 = n16629 & ~n37206;
  assign n37209 = ~n37207 & n37208;
  assign n37210 = ~n37201 & ~n37205;
  assign n37211 = ~n37209 & n37210;
  assign n37212 = pi0788 & ~n37211;
  assign n37213 = pi0609 & n36973;
  assign n37214 = ~n36887 & n37003;
  assign n37215 = ~pi0642 & ~n17336;
  assign n37216 = n36887 & ~n37215;
  assign n37217 = ~n36562 & n37216;
  assign n37218 = ~n37214 & ~n37217;
  assign n37219 = ~n36887 & n37004;
  assign n37220 = pi0642 & n17493;
  assign n37221 = ~n37215 & ~n37220;
  assign n37222 = n16667 & ~n37221;
  assign n37223 = n36887 & n37222;
  assign n37224 = pi0223 & ~n37219;
  assign n37225 = ~n37223 & n37224;
  assign n37226 = n37218 & ~n37225;
  assign n37227 = n37006 & ~n37226;
  assign n37228 = n37002 & ~n37227;
  assign n37229 = n17618 & n36922;
  assign n37230 = n17617 & ~n36887;
  assign n37231 = ~n36728 & n37013;
  assign n37232 = ~n37230 & n37231;
  assign n37233 = n37011 & ~n37229;
  assign n37234 = ~n37232 & n37233;
  assign n37235 = n17623 & n36922;
  assign n37236 = n17622 & ~n36887;
  assign n37237 = pi0223 & ~n37018;
  assign n37238 = ~n36738 & n37237;
  assign n37239 = ~n37236 & n37238;
  assign n37240 = n37017 & ~n37235;
  assign n37241 = ~n37239 & n37240;
  assign n37242 = ~pi0039 & ~n37234;
  assign n37243 = ~n37241 & n37242;
  assign n37244 = ~n36887 & ~n37028;
  assign n37245 = ~n16650 & n37222;
  assign n37246 = ~n6191 & ~n37245;
  assign n37247 = pi0680 & ~n37246;
  assign n37248 = pi0642 & ~n17504;
  assign n37249 = ~pi0614 & n17343;
  assign n37250 = ~n37248 & ~n37249;
  assign n37251 = ~pi0616 & ~n37250;
  assign n37252 = n37247 & ~n37251;
  assign n37253 = ~n37244 & ~n37252;
  assign n37254 = ~n37033 & ~n37253;
  assign n37255 = n6242 & ~n37254;
  assign n37256 = ~pi0680 & n37038;
  assign n37257 = pi0642 & ~n36588;
  assign n37258 = ~n6191 & n17325;
  assign n37259 = pi0680 & ~n17329;
  assign n37260 = ~n37257 & n37259;
  assign n37261 = ~n37258 & n37260;
  assign n37262 = pi0681 & ~n37261;
  assign n37263 = ~n37256 & n37262;
  assign n37264 = ~n37044 & ~n37263;
  assign n37265 = ~n6242 & ~n37264;
  assign n37266 = pi0223 & ~n37265;
  assign n37267 = ~n37255 & n37266;
  assign n37268 = ~pi0680 & ~n37050;
  assign n37269 = ~n17336 & ~n37248;
  assign n37270 = n35897 & ~n37269;
  assign n37271 = pi0680 & ~n37270;
  assign n37272 = pi0642 & ~n17548;
  assign n37273 = n6191 & ~n37272;
  assign n37274 = ~n17455 & n37273;
  assign n37275 = n37271 & ~n37274;
  assign n37276 = ~n37268 & ~n37275;
  assign n37277 = pi0681 & ~n37276;
  assign n37278 = n37082 & ~n37277;
  assign n37279 = ~n36887 & ~n37079;
  assign n37280 = ~pi0642 & ~n6191;
  assign n37281 = ~n17450 & n37280;
  assign n37282 = n17454 & n17559;
  assign n37283 = n17167 & ~n37282;
  assign n37284 = pi0642 & n36607;
  assign n37285 = pi0680 & ~n37281;
  assign n37286 = ~n37284 & n37285;
  assign n37287 = ~n37283 & n37286;
  assign n37288 = ~n37279 & ~n37287;
  assign n37289 = ~n6242 & n37077;
  assign n37290 = ~n37288 & n37289;
  assign n37291 = ~pi0223 & ~n37278;
  assign n37292 = ~n37290 & n37291;
  assign n37293 = pi0215 & ~n37292;
  assign n37294 = ~n37267 & n37293;
  assign n37295 = ~n36887 & ~n37116;
  assign n37296 = ~n17359 & ~n37248;
  assign n37297 = n6191 & ~n37296;
  assign n37298 = n37247 & ~n37297;
  assign n37299 = ~n37295 & ~n37298;
  assign n37300 = n37122 & ~n37299;
  assign n37301 = ~n36887 & ~n37106;
  assign n37302 = pi0642 & ~n36638;
  assign n37303 = n17167 & ~n36631;
  assign n37304 = n36633 & n37280;
  assign n37305 = pi0680 & ~n37302;
  assign n37306 = ~n37303 & n37305;
  assign n37307 = ~n37304 & n37306;
  assign n37308 = ~n37301 & ~n37307;
  assign n37309 = n37111 & ~n37308;
  assign n37310 = pi0223 & ~n37309;
  assign n37311 = ~n37300 & n37310;
  assign n37312 = ~pi0642 & ~n17414;
  assign n37313 = n37273 & ~n37312;
  assign n37314 = n37271 & ~n37313;
  assign n37315 = ~n37268 & ~n37314;
  assign n37316 = pi0681 & ~n37315;
  assign n37317 = ~n37056 & ~n37316;
  assign n37318 = n6242 & ~n37317;
  assign n37319 = ~n36887 & ~n37061;
  assign n37320 = pi0642 & n17578;
  assign n37321 = ~n17422 & n37280;
  assign n37322 = pi0680 & ~n37320;
  assign n37323 = ~n17430 & n37322;
  assign n37324 = ~n37321 & n37323;
  assign n37325 = ~n37319 & ~n37324;
  assign n37326 = ~n37065 & ~n37325;
  assign n37327 = ~n6242 & ~n37326;
  assign n37328 = ~pi0223 & ~n37318;
  assign n37329 = ~n37327 & n37328;
  assign n37330 = ~n3448 & ~n37311;
  assign n37331 = ~n37329 & n37330;
  assign n37332 = n16653 & ~n37218;
  assign n37333 = ~pi0223 & n37332;
  assign n37334 = n36931 & ~n37225;
  assign n37335 = ~n37333 & n37334;
  assign n37336 = ~pi0215 & ~n37335;
  assign n37337 = ~n37331 & n37336;
  assign n37338 = pi0299 & ~n37294;
  assign n37339 = ~n37337 & n37338;
  assign n37340 = n6205 & n37254;
  assign n37341 = ~n6205 & n37264;
  assign n37342 = pi0223 & ~n37341;
  assign n37343 = ~n37340 & n37342;
  assign n37344 = n2603 & ~n37332;
  assign n37345 = ~n6205 & n37326;
  assign n37346 = n6205 & n37317;
  assign n37347 = ~n2603 & ~n37345;
  assign n37348 = ~n37346 & n37347;
  assign n37349 = ~pi0223 & ~n37344;
  assign n37350 = ~n37348 & n37349;
  assign n37351 = ~pi0299 & ~n37343;
  assign n37352 = ~n37350 & n37351;
  assign n37353 = pi0039 & ~n37352;
  assign n37354 = ~n37339 & n37353;
  assign n37355 = ~pi0038 & ~n37243;
  assign n37356 = ~n37354 & n37355;
  assign n37357 = n2571 & ~n37228;
  assign n37358 = ~n37356 & n37357;
  assign n37359 = ~n36886 & ~n37358;
  assign n37360 = ~pi0625 & n37359;
  assign n37361 = pi0625 & n37138;
  assign n37362 = ~pi1153 & ~n37361;
  assign n37363 = ~n37360 & n37362;
  assign n37364 = ~pi0608 & ~n37363;
  assign n37365 = ~n36966 & n37364;
  assign n37366 = ~pi0625 & n37138;
  assign n37367 = pi0625 & n37359;
  assign n37368 = pi1153 & ~n37366;
  assign n37369 = ~n37367 & n37368;
  assign n37370 = pi0608 & ~n37369;
  assign n37371 = ~n36970 & n37370;
  assign n37372 = ~n37365 & ~n37371;
  assign n37373 = pi0778 & ~n37372;
  assign n37374 = ~pi0778 & n37359;
  assign n37375 = ~n37373 & ~n37374;
  assign n37376 = ~pi0609 & ~n37375;
  assign n37377 = ~pi1155 & ~n37213;
  assign n37378 = ~n37376 & n37377;
  assign n37379 = ~pi0660 & ~n37145;
  assign n37380 = ~n37378 & n37379;
  assign n37381 = ~pi0609 & n36973;
  assign n37382 = pi0609 & ~n37375;
  assign n37383 = pi1155 & ~n37381;
  assign n37384 = ~n37382 & n37383;
  assign n37385 = pi0660 & ~n37149;
  assign n37386 = ~n37384 & n37385;
  assign n37387 = ~n37380 & ~n37386;
  assign n37388 = pi0785 & ~n37387;
  assign n37389 = ~pi0785 & ~n37375;
  assign n37390 = ~n37388 & ~n37389;
  assign n37391 = ~pi0618 & ~n37390;
  assign n37392 = pi0618 & ~n36975;
  assign n37393 = ~pi1154 & ~n37392;
  assign n37394 = ~n37391 & n37393;
  assign n37395 = ~pi0627 & ~n37157;
  assign n37396 = ~n37394 & n37395;
  assign n37397 = pi0618 & ~n37390;
  assign n37398 = ~pi0618 & ~n36975;
  assign n37399 = pi1154 & ~n37398;
  assign n37400 = ~n37397 & n37399;
  assign n37401 = pi0627 & ~n37161;
  assign n37402 = ~n37400 & n37401;
  assign n37403 = ~n37396 & ~n37402;
  assign n37404 = pi0781 & ~n37403;
  assign n37405 = ~pi0781 & ~n37390;
  assign n37406 = ~n37404 & ~n37405;
  assign n37407 = ~pi0789 & n37406;
  assign n37408 = ~pi0619 & ~n37406;
  assign n37409 = pi0619 & n36978;
  assign n37410 = ~pi1159 & ~n37409;
  assign n37411 = ~n37408 & n37410;
  assign n37412 = ~pi0648 & ~n37169;
  assign n37413 = ~n37411 & n37412;
  assign n37414 = ~pi0619 & n36978;
  assign n37415 = pi0619 & ~n37406;
  assign n37416 = pi1159 & ~n37414;
  assign n37417 = ~n37415 & n37416;
  assign n37418 = pi0648 & ~n37173;
  assign n37419 = ~n37417 & n37418;
  assign n37420 = pi0789 & ~n37413;
  assign n37421 = ~n37419 & n37420;
  assign n37422 = n17970 & ~n37407;
  assign n37423 = ~n37421 & n37422;
  assign n37424 = ~n37212 & ~n37423;
  assign n37425 = ~n37198 & ~n37424;
  assign n37426 = n20364 & n37197;
  assign n37427 = ~n20206 & ~n37426;
  assign n37428 = ~n37425 & n37427;
  assign n37429 = ~n37186 & ~n37428;
  assign n37430 = pi0644 & n37429;
  assign n37431 = pi0715 & ~n36997;
  assign n37432 = ~n37430 & n37431;
  assign n37433 = n17804 & ~n36883;
  assign n37434 = ~n17804 & n37181;
  assign n37435 = ~n37433 & ~n37434;
  assign n37436 = pi0644 & ~n37435;
  assign n37437 = ~pi0644 & ~n36883;
  assign n37438 = ~pi0715 & ~n37437;
  assign n37439 = ~n37436 & n37438;
  assign n37440 = pi1160 & ~n37439;
  assign n37441 = ~n37432 & n37440;
  assign n37442 = pi0644 & n36996;
  assign n37443 = ~pi0644 & n37429;
  assign n37444 = ~pi0715 & ~n37442;
  assign n37445 = ~n37443 & n37444;
  assign n37446 = ~pi0644 & ~n37435;
  assign n37447 = pi0644 & ~n36883;
  assign n37448 = pi0715 & ~n37447;
  assign n37449 = ~n37446 & n37448;
  assign n37450 = ~pi1160 & ~n37449;
  assign n37451 = ~n37445 & n37450;
  assign n37452 = ~n37441 & ~n37451;
  assign n37453 = pi0790 & ~n37452;
  assign n37454 = ~pi0790 & n37429;
  assign n37455 = ~n37453 & ~n37454;
  assign n37456 = ~po1038 & ~n37455;
  assign n37457 = ~pi0223 & po1038;
  assign po0380 = ~n37456 & ~n37457;
  assign n37459 = pi0224 & ~n36258;
  assign n37460 = ~n19149 & ~n37459;
  assign n37461 = pi0224 & ~n2571;
  assign n37462 = pi0224 & ~n16641;
  assign n37463 = pi0038 & ~n37462;
  assign n37464 = pi0662 & n16646;
  assign n37465 = n37463 & ~n37464;
  assign n37466 = pi0662 & pi0680;
  assign n37467 = n16918 & ~n37466;
  assign n37468 = ~pi0224 & ~n16918;
  assign n37469 = pi0224 & n16935;
  assign n37470 = ~pi0299 & ~n37469;
  assign n37471 = ~n37467 & n37470;
  assign n37472 = ~n37468 & n37471;
  assign n37473 = pi0224 & n16944;
  assign n37474 = n16923 & ~n37466;
  assign n37475 = ~pi0224 & ~n16923;
  assign n37476 = pi0299 & ~n37473;
  assign n37477 = ~n37474 & n37476;
  assign n37478 = ~n37475 & n37477;
  assign n37479 = ~pi0039 & ~n37472;
  assign n37480 = ~n37478 & n37479;
  assign n37481 = pi0662 & n16655;
  assign n37482 = ~n6193 & ~n36283;
  assign n37483 = n17018 & ~n37482;
  assign n37484 = ~n6205 & n37483;
  assign n37485 = pi0662 & ~n16786;
  assign n37486 = ~pi0662 & ~n17011;
  assign n37487 = ~n37485 & ~n37486;
  assign n37488 = n6205 & n37487;
  assign n37489 = pi0224 & ~n37484;
  assign n37490 = ~n37488 & n37489;
  assign n37491 = pi0662 & n16703;
  assign n37492 = ~n6205 & ~n37491;
  assign n37493 = ~n16690 & n37466;
  assign n37494 = n6205 & ~n37493;
  assign n37495 = n5810 & ~n37492;
  assign n37496 = ~n37494 & n37495;
  assign n37497 = ~pi0223 & ~n37481;
  assign n37498 = ~n37496 & n37497;
  assign n37499 = ~n37490 & n37498;
  assign n37500 = ~pi0224 & pi0662;
  assign n37501 = n16729 & n37500;
  assign n37502 = ~pi0662 & ~n16990;
  assign n37503 = pi0662 & ~n36319;
  assign n37504 = ~n37502 & ~n37503;
  assign n37505 = n6205 & n37504;
  assign n37506 = ~pi0662 & ~n16970;
  assign n37507 = pi0662 & ~n16818;
  assign n37508 = ~n37506 & ~n37507;
  assign n37509 = ~n6205 & n37508;
  assign n37510 = pi0224 & ~n37505;
  assign n37511 = ~n37509 & n37510;
  assign n37512 = pi0223 & ~n37501;
  assign n37513 = ~n37511 & n37512;
  assign n37514 = ~pi0299 & ~n37513;
  assign n37515 = ~n37499 & n37514;
  assign n37516 = pi0224 & ~n16653;
  assign n37517 = n3448 & ~n37516;
  assign n37518 = n16658 & n37466;
  assign n37519 = n37517 & ~n37518;
  assign n37520 = ~n6242 & n37483;
  assign n37521 = n6242 & n37487;
  assign n37522 = pi0224 & ~n37520;
  assign n37523 = ~n37521 & n37522;
  assign n37524 = ~n6242 & ~n37491;
  assign n37525 = n6242 & ~n37493;
  assign n37526 = ~pi0224 & ~n37524;
  assign n37527 = ~n37525 & n37526;
  assign n37528 = ~n3448 & ~n37527;
  assign n37529 = ~n37523 & n37528;
  assign n37530 = ~n37519 & ~n37529;
  assign n37531 = ~pi0215 & ~n37530;
  assign n37532 = n16744 & n37500;
  assign n37533 = n6242 & n37504;
  assign n37534 = ~n6242 & n37508;
  assign n37535 = pi0224 & ~n37533;
  assign n37536 = ~n37534 & n37535;
  assign n37537 = pi0215 & ~n37532;
  assign n37538 = ~n37536 & n37537;
  assign n37539 = pi0299 & ~n37538;
  assign n37540 = ~n37531 & n37539;
  assign n37541 = pi0039 & ~n37515;
  assign n37542 = ~n37540 & n37541;
  assign n37543 = ~n37480 & ~n37542;
  assign n37544 = ~pi0038 & ~n37543;
  assign n37545 = n2571 & ~n37465;
  assign n37546 = ~n37544 & n37545;
  assign n37547 = ~n37461 & ~n37546;
  assign n37548 = ~pi0778 & ~n37547;
  assign n37549 = pi0625 & n37547;
  assign n37550 = ~pi0625 & ~n37459;
  assign n37551 = pi1153 & ~n37550;
  assign n37552 = ~n37549 & n37551;
  assign n37553 = ~pi0625 & n37547;
  assign n37554 = pi0625 & ~n37459;
  assign n37555 = ~pi1153 & ~n37554;
  assign n37556 = ~n37553 & n37555;
  assign n37557 = ~n37552 & ~n37556;
  assign n37558 = pi0778 & ~n37557;
  assign n37559 = ~n37548 & ~n37558;
  assign n37560 = ~n17075 & ~n37559;
  assign n37561 = n17075 & n37459;
  assign n37562 = ~n37560 & ~n37561;
  assign n37563 = ~n16639 & ~n37562;
  assign n37564 = n16639 & n37459;
  assign n37565 = ~n37563 & ~n37564;
  assign n37566 = ~n16635 & n37565;
  assign n37567 = ~n16631 & n37566;
  assign n37568 = ~n37460 & ~n37567;
  assign n37569 = ~n19142 & ~n37568;
  assign n37570 = n17856 & ~n37459;
  assign n37571 = ~n37569 & ~n37570;
  assign n37572 = ~pi0787 & n37571;
  assign n37573 = ~pi0647 & ~n37571;
  assign n37574 = pi0647 & ~n37459;
  assign n37575 = ~pi1157 & ~n37574;
  assign n37576 = ~n37573 & n37575;
  assign n37577 = pi0647 & ~n37571;
  assign n37578 = ~pi0647 & ~n37459;
  assign n37579 = pi1157 & ~n37578;
  assign n37580 = ~n37577 & n37579;
  assign n37581 = ~n37576 & ~n37580;
  assign n37582 = pi0787 & ~n37581;
  assign n37583 = ~n37572 & ~n37582;
  assign n37584 = ~pi0644 & n37583;
  assign n37585 = pi0628 & ~n37459;
  assign n37586 = ~pi0628 & ~n37568;
  assign n37587 = n17777 & ~n37585;
  assign n37588 = ~n37586 & n37587;
  assign n37589 = n17969 & ~n37459;
  assign n37590 = pi0614 & n17280;
  assign n37591 = n37463 & ~n37590;
  assign n37592 = pi0614 & n17226;
  assign n37593 = ~pi0224 & n37592;
  assign n37594 = ~pi0614 & n17226;
  assign n37595 = pi0224 & ~n37594;
  assign n37596 = n17137 & n37595;
  assign n37597 = ~pi0299 & ~n37593;
  assign n37598 = ~n37596 & n37597;
  assign n37599 = pi0614 & n17231;
  assign n37600 = pi0224 & n17122;
  assign n37601 = n37599 & ~n37600;
  assign n37602 = pi0224 & ~n16941;
  assign n37603 = ~n37601 & ~n37602;
  assign n37604 = pi0299 & n37603;
  assign n37605 = ~pi0039 & ~n37598;
  assign n37606 = ~n37604 & n37605;
  assign n37607 = pi0614 & ~n36411;
  assign n37608 = ~pi0224 & n37607;
  assign n37609 = ~n16743 & n37608;
  assign n37610 = pi0614 & ~n17183;
  assign n37611 = ~n36026 & ~n37610;
  assign n37612 = ~pi0680 & ~n37611;
  assign n37613 = pi0680 & ~n17187;
  assign n37614 = ~n36028 & n37613;
  assign n37615 = ~n37612 & ~n37614;
  assign n37616 = n16657 & ~n37615;
  assign n37617 = ~n16657 & ~n37611;
  assign n37618 = ~n37616 & ~n37617;
  assign n37619 = ~n6242 & n37618;
  assign n37620 = pi0614 & n17168;
  assign n37621 = n16653 & ~n37620;
  assign n37622 = ~n6192 & ~n37621;
  assign n37623 = ~n16802 & ~n37622;
  assign n37624 = ~n16657 & ~n37623;
  assign n37625 = ~pi0680 & ~n37623;
  assign n37626 = pi0680 & n37620;
  assign n37627 = ~n16973 & ~n37626;
  assign n37628 = ~n37625 & n37627;
  assign n37629 = n16657 & ~n37628;
  assign n37630 = ~n37624 & ~n37629;
  assign n37631 = n6242 & n37630;
  assign n37632 = pi0224 & ~n37619;
  assign n37633 = ~n37631 & n37632;
  assign n37634 = ~n37609 & ~n37633;
  assign n37635 = pi0215 & ~n37634;
  assign n37636 = n16999 & n17168;
  assign n37637 = n37517 & ~n37636;
  assign n37638 = pi0614 & ~n17154;
  assign n37639 = ~pi0614 & pi0616;
  assign n37640 = n16699 & n37639;
  assign n37641 = ~n6197 & n16772;
  assign n37642 = n6191 & ~n16697;
  assign n37643 = ~n37641 & n37642;
  assign n37644 = ~n37638 & ~n37640;
  assign n37645 = ~n37643 & n37644;
  assign n37646 = ~n16657 & ~n37645;
  assign n37647 = ~pi0680 & ~n37645;
  assign n37648 = pi0614 & n17375;
  assign n37649 = pi0680 & ~n37648;
  assign n37650 = n16681 & n37649;
  assign n37651 = ~n37626 & ~n37650;
  assign n37652 = ~n37647 & n37651;
  assign n37653 = n16657 & ~n37652;
  assign n37654 = ~n37646 & ~n37653;
  assign n37655 = ~n6242 & n37654;
  assign n37656 = ~n16775 & ~n37622;
  assign n37657 = ~n16657 & ~n37656;
  assign n37658 = ~pi0680 & ~n37656;
  assign n37659 = ~n16995 & ~n37626;
  assign n37660 = ~n37658 & n37659;
  assign n37661 = n16657 & ~n37660;
  assign n37662 = ~n37657 & ~n37661;
  assign n37663 = n6242 & n37662;
  assign n37664 = pi0224 & ~n37655;
  assign n37665 = ~n37663 & n37664;
  assign n37666 = ~n16699 & n37620;
  assign n37667 = ~pi0680 & ~n37666;
  assign n37668 = ~n37649 & ~n37667;
  assign n37669 = n16657 & ~n37668;
  assign n37670 = ~n16657 & ~n37666;
  assign n37671 = ~n37669 & ~n37670;
  assign n37672 = ~n6242 & ~n37671;
  assign n37673 = pi0614 & ~n36463;
  assign n37674 = n6242 & ~n37673;
  assign n37675 = ~pi0224 & ~n37674;
  assign n37676 = ~n37672 & n37675;
  assign n37677 = ~n3448 & ~n37676;
  assign n37678 = ~n37665 & n37677;
  assign n37679 = ~pi0215 & ~n37637;
  assign n37680 = ~n37678 & n37679;
  assign n37681 = pi0299 & ~n37635;
  assign n37682 = ~n37680 & n37681;
  assign n37683 = ~n16724 & n37608;
  assign n37684 = ~n6205 & n37618;
  assign n37685 = n6205 & n37630;
  assign n37686 = pi0224 & ~n37684;
  assign n37687 = ~n37685 & n37686;
  assign n37688 = pi0223 & ~n37683;
  assign n37689 = ~n37687 & n37688;
  assign n37690 = pi0614 & n17268;
  assign n37691 = n6205 & ~n37673;
  assign n37692 = ~n6205 & ~n37671;
  assign n37693 = n5810 & ~n37691;
  assign n37694 = ~n37692 & n37693;
  assign n37695 = ~n6205 & n37654;
  assign n37696 = n6205 & n37662;
  assign n37697 = pi0224 & ~n37695;
  assign n37698 = ~n37696 & n37697;
  assign n37699 = ~pi0223 & ~n37690;
  assign n37700 = ~n37694 & n37699;
  assign n37701 = ~n37698 & n37700;
  assign n37702 = ~n37689 & ~n37701;
  assign n37703 = ~pi0299 & ~n37702;
  assign n37704 = pi0039 & ~n37682;
  assign n37705 = ~n37703 & n37704;
  assign n37706 = ~pi0038 & ~n37606;
  assign n37707 = ~n37705 & n37706;
  assign n37708 = n2571 & ~n37591;
  assign n37709 = ~n37707 & n37708;
  assign n37710 = ~n37461 & ~n37709;
  assign n37711 = ~n17117 & ~n37710;
  assign n37712 = n17117 & n37459;
  assign n37713 = ~n37711 & ~n37712;
  assign n37714 = ~pi0785 & ~n37713;
  assign n37715 = pi0609 & n37713;
  assign n37716 = ~pi0609 & ~n37459;
  assign n37717 = pi1155 & ~n37716;
  assign n37718 = ~n37715 & n37717;
  assign n37719 = ~pi0609 & n37713;
  assign n37720 = pi0609 & ~n37459;
  assign n37721 = ~pi1155 & ~n37720;
  assign n37722 = ~n37719 & n37721;
  assign n37723 = ~n37718 & ~n37722;
  assign n37724 = pi0785 & ~n37723;
  assign n37725 = ~n37714 & ~n37724;
  assign n37726 = ~pi0781 & ~n37725;
  assign n37727 = pi0618 & n37725;
  assign n37728 = ~pi0618 & ~n37459;
  assign n37729 = pi1154 & ~n37728;
  assign n37730 = ~n37727 & n37729;
  assign n37731 = ~pi0618 & n37725;
  assign n37732 = pi0618 & ~n37459;
  assign n37733 = ~pi1154 & ~n37732;
  assign n37734 = ~n37731 & n37733;
  assign n37735 = ~n37730 & ~n37734;
  assign n37736 = pi0781 & ~n37735;
  assign n37737 = ~n37726 & ~n37736;
  assign n37738 = ~pi0789 & ~n37737;
  assign n37739 = pi0619 & n37737;
  assign n37740 = ~pi0619 & ~n37459;
  assign n37741 = pi1159 & ~n37740;
  assign n37742 = ~n37739 & n37741;
  assign n37743 = ~pi0619 & n37737;
  assign n37744 = pi0619 & ~n37459;
  assign n37745 = ~pi1159 & ~n37744;
  assign n37746 = ~n37743 & n37745;
  assign n37747 = ~n37742 & ~n37746;
  assign n37748 = pi0789 & ~n37747;
  assign n37749 = ~n37738 & ~n37748;
  assign n37750 = ~n17969 & n37749;
  assign n37751 = ~n37589 & ~n37750;
  assign n37752 = ~n20570 & n37751;
  assign n37753 = ~pi0628 & ~n37459;
  assign n37754 = pi0628 & ~n37568;
  assign n37755 = n17776 & ~n37753;
  assign n37756 = ~n37754 & n37755;
  assign n37757 = ~n37588 & ~n37756;
  assign n37758 = ~n37752 & n37757;
  assign n37759 = pi0792 & ~n37758;
  assign n37760 = pi0609 & n37559;
  assign n37761 = pi0662 & n17355;
  assign n37762 = n16641 & n37761;
  assign n37763 = n37591 & ~n37762;
  assign n37764 = n17617 & n37466;
  assign n37765 = ~n37592 & ~n37764;
  assign n37766 = ~pi0224 & ~n37765;
  assign n37767 = n17617 & ~n37466;
  assign n37768 = ~n36728 & n37595;
  assign n37769 = ~n37767 & n37768;
  assign n37770 = ~n37766 & ~n37769;
  assign n37771 = ~pi0299 & ~n37770;
  assign n37772 = ~n37466 & n37603;
  assign n37773 = ~pi0614 & n17231;
  assign n37774 = ~n36738 & ~n37773;
  assign n37775 = pi0224 & ~n37774;
  assign n37776 = ~pi0224 & ~n17622;
  assign n37777 = ~n37599 & n37776;
  assign n37778 = ~n37775 & ~n37777;
  assign n37779 = n37466 & ~n37778;
  assign n37780 = pi0299 & ~n37772;
  assign n37781 = ~n37779 & n37780;
  assign n37782 = ~n37771 & ~n37781;
  assign n37783 = ~pi0039 & ~n37782;
  assign n37784 = n17407 & n37466;
  assign n37785 = ~n37636 & ~n37784;
  assign n37786 = ~pi0224 & ~n37785;
  assign n37787 = ~pi0222 & n37786;
  assign n37788 = ~n17407 & n37639;
  assign n37789 = ~n36620 & ~n37788;
  assign n37790 = pi0680 & ~n37789;
  assign n37791 = ~n36675 & ~n37636;
  assign n37792 = ~n37790 & ~n37791;
  assign n37793 = pi0662 & ~n37792;
  assign n37794 = ~pi0662 & ~n37673;
  assign n37795 = ~n37793 & ~n37794;
  assign n37796 = n6205 & ~n37795;
  assign n37797 = ~pi0662 & ~n16656;
  assign n37798 = ~n37666 & n37797;
  assign n37799 = ~pi0614 & n17434;
  assign n37800 = pi0614 & ~n17578;
  assign n37801 = pi0680 & ~n37800;
  assign n37802 = ~n37799 & n37801;
  assign n37803 = ~n37667 & ~n37802;
  assign n37804 = pi0662 & ~n37803;
  assign n37805 = ~n37669 & ~n37798;
  assign n37806 = ~n37804 & n37805;
  assign n37807 = ~n6205 & ~n37806;
  assign n37808 = n5810 & ~n37796;
  assign n37809 = ~n37807 & n37808;
  assign n37810 = ~n37656 & n37797;
  assign n37811 = ~pi0614 & ~n24055;
  assign n37812 = pi0614 & ~n36562;
  assign n37813 = ~n37811 & ~n37812;
  assign n37814 = ~n16650 & n37813;
  assign n37815 = pi0616 & ~n37814;
  assign n37816 = pi0614 & ~n17504;
  assign n37817 = ~n17361 & ~n37816;
  assign n37818 = ~pi0616 & ~n37817;
  assign n37819 = ~n37815 & ~n37818;
  assign n37820 = pi0680 & ~n37819;
  assign n37821 = ~n37658 & ~n37820;
  assign n37822 = pi0662 & ~n37821;
  assign n37823 = ~n37661 & ~n37810;
  assign n37824 = ~n37822 & n37823;
  assign n37825 = n6205 & n37824;
  assign n37826 = ~n37645 & n37797;
  assign n37827 = pi0614 & ~n36638;
  assign n37828 = n36633 & n37639;
  assign n37829 = ~n37827 & ~n37828;
  assign n37830 = ~n36636 & n37829;
  assign n37831 = pi0680 & ~n37830;
  assign n37832 = ~n37647 & ~n37831;
  assign n37833 = pi0662 & ~n37832;
  assign n37834 = ~n37653 & ~n37826;
  assign n37835 = ~n37833 & n37834;
  assign n37836 = ~n6205 & n37835;
  assign n37837 = pi0224 & ~n37836;
  assign n37838 = ~n37825 & n37837;
  assign n37839 = ~pi0223 & ~n37787;
  assign n37840 = ~n37809 & n37839;
  assign n37841 = ~n37838 & n37840;
  assign n37842 = pi0680 & ~n17445;
  assign n37843 = ~n37636 & ~n37842;
  assign n37844 = ~n37790 & ~n37843;
  assign n37845 = pi0662 & ~n37844;
  assign n37846 = ~pi0662 & ~n37607;
  assign n37847 = ~n37845 & ~n37846;
  assign n37848 = ~pi0224 & ~n37847;
  assign n37849 = ~n37623 & n37797;
  assign n37850 = ~n17345 & ~n37816;
  assign n37851 = ~pi0616 & ~n37850;
  assign n37852 = ~n37815 & ~n37851;
  assign n37853 = pi0680 & ~n37852;
  assign n37854 = ~n37625 & ~n37853;
  assign n37855 = pi0662 & ~n37854;
  assign n37856 = ~n37629 & ~n37849;
  assign n37857 = ~n37855 & n37856;
  assign n37858 = pi0224 & n37857;
  assign n37859 = n6205 & ~n37848;
  assign n37860 = ~n37858 & n37859;
  assign n37861 = ~n37611 & n37797;
  assign n37862 = pi0614 & ~n36588;
  assign n37863 = n17330 & ~n37862;
  assign n37864 = pi0680 & ~n37863;
  assign n37865 = ~n37612 & ~n37864;
  assign n37866 = pi0662 & ~n37865;
  assign n37867 = ~n37616 & ~n37861;
  assign n37868 = ~n37866 & n37867;
  assign n37869 = pi0224 & n37868;
  assign n37870 = ~n16723 & n37607;
  assign n37871 = ~pi0662 & ~n37870;
  assign n37872 = pi0614 & ~pi0680;
  assign n37873 = n17237 & n37872;
  assign n37874 = pi0614 & n36607;
  assign n37875 = ~pi0614 & n17451;
  assign n37876 = pi0680 & ~n37874;
  assign n37877 = ~n37875 & n37876;
  assign n37878 = ~n17457 & n37877;
  assign n37879 = pi0662 & ~n37873;
  assign n37880 = ~n37878 & n37879;
  assign n37881 = ~n37871 & ~n37880;
  assign n37882 = ~pi0224 & ~n37881;
  assign n37883 = ~n6205 & ~n37882;
  assign n37884 = ~n37869 & n37883;
  assign n37885 = pi0223 & ~n37884;
  assign n37886 = ~n37860 & n37885;
  assign n37887 = ~n37841 & ~n37886;
  assign n37888 = ~pi0299 & ~n37887;
  assign n37889 = ~n6242 & ~n37868;
  assign n37890 = n6242 & ~n37857;
  assign n37891 = pi0224 & ~n37889;
  assign n37892 = ~n37890 & n37891;
  assign n37893 = n6242 & n37847;
  assign n37894 = ~n6242 & n37881;
  assign n37895 = ~pi0224 & ~n37894;
  assign n37896 = ~n37893 & n37895;
  assign n37897 = pi0215 & ~n37896;
  assign n37898 = ~n37892 & n37897;
  assign n37899 = n37466 & n37813;
  assign n37900 = ~n37466 & ~n37620;
  assign n37901 = n16667 & n37900;
  assign n37902 = pi0224 & ~n37901;
  assign n37903 = ~n37899 & n37902;
  assign n37904 = n37517 & ~n37903;
  assign n37905 = ~n37786 & n37904;
  assign n37906 = ~pi0224 & ~n37795;
  assign n37907 = pi0224 & n37824;
  assign n37908 = n6242 & ~n37906;
  assign n37909 = ~n37907 & n37908;
  assign n37910 = ~pi0224 & ~n37806;
  assign n37911 = pi0224 & n37835;
  assign n37912 = ~n6242 & ~n37910;
  assign n37913 = ~n37911 & n37912;
  assign n37914 = ~n3448 & ~n37909;
  assign n37915 = ~n37913 & n37914;
  assign n37916 = ~pi0215 & ~n37905;
  assign n37917 = ~n37915 & n37916;
  assign n37918 = pi0299 & ~n37898;
  assign n37919 = ~n37917 & n37918;
  assign n37920 = pi0039 & ~n37888;
  assign n37921 = ~n37919 & n37920;
  assign n37922 = ~pi0038 & ~n37783;
  assign n37923 = ~n37921 & n37922;
  assign n37924 = n2571 & ~n37763;
  assign n37925 = ~n37923 & n37924;
  assign n37926 = ~n37461 & ~n37925;
  assign n37927 = ~pi0625 & n37926;
  assign n37928 = pi0625 & n37710;
  assign n37929 = ~pi1153 & ~n37928;
  assign n37930 = ~n37927 & n37929;
  assign n37931 = ~pi0608 & ~n37552;
  assign n37932 = ~n37930 & n37931;
  assign n37933 = ~pi0625 & n37710;
  assign n37934 = pi0625 & n37926;
  assign n37935 = pi1153 & ~n37933;
  assign n37936 = ~n37934 & n37935;
  assign n37937 = pi0608 & ~n37556;
  assign n37938 = ~n37936 & n37937;
  assign n37939 = ~n37932 & ~n37938;
  assign n37940 = pi0778 & ~n37939;
  assign n37941 = ~pi0778 & n37926;
  assign n37942 = ~n37940 & ~n37941;
  assign n37943 = ~pi0609 & ~n37942;
  assign n37944 = ~pi1155 & ~n37760;
  assign n37945 = ~n37943 & n37944;
  assign n37946 = ~pi0660 & ~n37718;
  assign n37947 = ~n37945 & n37946;
  assign n37948 = ~pi0609 & n37559;
  assign n37949 = pi0609 & ~n37942;
  assign n37950 = pi1155 & ~n37948;
  assign n37951 = ~n37949 & n37950;
  assign n37952 = pi0660 & ~n37722;
  assign n37953 = ~n37951 & n37952;
  assign n37954 = ~n37947 & ~n37953;
  assign n37955 = pi0785 & ~n37954;
  assign n37956 = ~pi0785 & ~n37942;
  assign n37957 = ~n37955 & ~n37956;
  assign n37958 = ~pi0618 & ~n37957;
  assign n37959 = pi0618 & n37562;
  assign n37960 = ~pi1154 & ~n37959;
  assign n37961 = ~n37958 & n37960;
  assign n37962 = ~pi0627 & ~n37730;
  assign n37963 = ~n37961 & n37962;
  assign n37964 = ~pi0618 & n37562;
  assign n37965 = pi0618 & ~n37957;
  assign n37966 = pi1154 & ~n37964;
  assign n37967 = ~n37965 & n37966;
  assign n37968 = pi0627 & ~n37734;
  assign n37969 = ~n37967 & n37968;
  assign n37970 = ~n37963 & ~n37969;
  assign n37971 = pi0781 & ~n37970;
  assign n37972 = ~pi0781 & ~n37957;
  assign n37973 = ~n37971 & ~n37972;
  assign n37974 = ~pi0789 & n37973;
  assign n37975 = ~pi0619 & ~n37973;
  assign n37976 = pi0619 & n37565;
  assign n37977 = ~pi1159 & ~n37976;
  assign n37978 = ~n37975 & n37977;
  assign n37979 = ~pi0648 & ~n37742;
  assign n37980 = ~n37978 & n37979;
  assign n37981 = pi0619 & ~n37973;
  assign n37982 = ~pi0619 & n37565;
  assign n37983 = pi1159 & ~n37982;
  assign n37984 = ~n37981 & n37983;
  assign n37985 = pi0648 & ~n37746;
  assign n37986 = ~n37984 & n37985;
  assign n37987 = pi0789 & ~n37980;
  assign n37988 = ~n37986 & n37987;
  assign n37989 = n17970 & ~n37974;
  assign n37990 = ~n37988 & n37989;
  assign n37991 = n16635 & ~n37459;
  assign n37992 = ~n37566 & ~n37991;
  assign n37993 = n17871 & ~n37992;
  assign n37994 = ~pi0626 & n37459;
  assign n37995 = pi0626 & ~n37749;
  assign n37996 = n16628 & ~n37994;
  assign n37997 = ~n37995 & n37996;
  assign n37998 = pi0626 & n37459;
  assign n37999 = ~pi0626 & ~n37749;
  assign n38000 = n16629 & ~n37998;
  assign n38001 = ~n37999 & n38000;
  assign n38002 = ~n37993 & ~n37997;
  assign n38003 = ~n38001 & n38002;
  assign n38004 = pi0788 & ~n38003;
  assign n38005 = ~n20364 & ~n38004;
  assign n38006 = ~n37990 & n38005;
  assign n38007 = ~n37759 & ~n38006;
  assign n38008 = ~n20206 & ~n38007;
  assign n38009 = ~pi0630 & n37580;
  assign n38010 = ~n17779 & n37751;
  assign n38011 = n17779 & n37459;
  assign n38012 = ~n38010 & ~n38011;
  assign n38013 = ~n20559 & ~n38012;
  assign n38014 = pi0630 & n37576;
  assign n38015 = ~n38009 & ~n38014;
  assign n38016 = ~n38013 & n38015;
  assign n38017 = pi0787 & ~n38016;
  assign n38018 = ~n38008 & ~n38017;
  assign n38019 = pi0644 & n38018;
  assign n38020 = pi0715 & ~n37584;
  assign n38021 = ~n38019 & n38020;
  assign n38022 = n17804 & ~n37459;
  assign n38023 = ~n17804 & n38012;
  assign n38024 = ~n38022 & ~n38023;
  assign n38025 = pi0644 & ~n38024;
  assign n38026 = ~pi0644 & ~n37459;
  assign n38027 = ~pi0715 & ~n38026;
  assign n38028 = ~n38025 & n38027;
  assign n38029 = pi1160 & ~n38028;
  assign n38030 = ~n38021 & n38029;
  assign n38031 = pi0644 & n37583;
  assign n38032 = ~pi0644 & n38018;
  assign n38033 = ~pi0715 & ~n38031;
  assign n38034 = ~n38032 & n38033;
  assign n38035 = ~pi0644 & ~n38024;
  assign n38036 = pi0644 & ~n37459;
  assign n38037 = pi0715 & ~n38036;
  assign n38038 = ~n38035 & n38037;
  assign n38039 = ~pi1160 & ~n38038;
  assign n38040 = ~n38034 & n38039;
  assign n38041 = ~n38030 & ~n38040;
  assign n38042 = pi0790 & ~n38041;
  assign n38043 = ~pi0790 & n38018;
  assign n38044 = ~n38042 & ~n38043;
  assign n38045 = ~po1038 & ~n38044;
  assign n38046 = ~pi0224 & po1038;
  assign po0381 = ~n38045 & ~n38046;
  assign n38048 = n2547 & n2625;
  assign n38049 = n3330 & n38048;
  assign n38050 = ~pi0062 & n38049;
  assign n38051 = ~n3328 & ~n38050;
  assign n38052 = pi0062 & n38049;
  assign n38053 = n2534 & n38048;
  assign n38054 = pi0054 & ~n38053;
  assign n38055 = pi0092 & n2533;
  assign n38056 = n38048 & n38055;
  assign n38057 = ~n6169 & n6263;
  assign n38058 = ~pi0137 & ~n38057;
  assign n38059 = n7301 & ~n38058;
  assign n38060 = pi0075 & ~n38059;
  assign n38061 = pi0087 & n38048;
  assign n38062 = n6286 & ~n38058;
  assign n38063 = pi0038 & ~pi0137;
  assign n38064 = pi0039 & n2547;
  assign n38065 = ~n2741 & ~n2979;
  assign n38066 = pi0137 & ~n38065;
  assign n38067 = ~n2740 & ~n38066;
  assign n38068 = ~pi0332 & ~n38067;
  assign n38069 = n2517 & n11417;
  assign n38070 = n2738 & ~n38069;
  assign n38071 = ~pi0137 & n2713;
  assign n38072 = ~n38070 & n38071;
  assign n38073 = n3168 & ~n11417;
  assign n38074 = ~n2903 & n38073;
  assign n38075 = n2746 & ~n38074;
  assign n38076 = n2744 & ~n38075;
  assign n38077 = ~n2712 & ~n38076;
  assign n38078 = ~pi0095 & ~n38077;
  assign n38079 = n3088 & ~n38078;
  assign n38080 = pi0332 & ~n38072;
  assign n38081 = ~n38079 & n38080;
  assign n38082 = ~n38068 & ~n38081;
  assign n38083 = pi0210 & ~n38082;
  assign n38084 = n2922 & ~n38070;
  assign n38085 = pi1093 & ~n38084;
  assign n38086 = n2922 & n2933;
  assign n38087 = n2517 & ~n7455;
  assign n38088 = ~n2960 & n38087;
  assign n38089 = ~pi0032 & ~n38088;
  assign n38090 = n38086 & ~n38089;
  assign n38091 = ~pi1093 & ~n38090;
  assign n38092 = ~n2933 & n38084;
  assign n38093 = n11416 & n38087;
  assign n38094 = n38086 & n38093;
  assign n38095 = ~n38092 & ~n38094;
  assign n38096 = n38091 & n38095;
  assign n38097 = ~n38085 & ~n38096;
  assign n38098 = n11549 & ~n38097;
  assign n38099 = ~n2921 & ~n38076;
  assign n38100 = ~pi0095 & ~n38099;
  assign n38101 = ~n2741 & ~n38100;
  assign n38102 = pi0137 & ~n38101;
  assign n38103 = ~n2933 & n3023;
  assign n38104 = n38091 & ~n38103;
  assign n38105 = ~n2997 & n38087;
  assign n38106 = ~pi0032 & ~n38105;
  assign n38107 = n38086 & ~n38106;
  assign n38108 = pi1093 & ~n38103;
  assign n38109 = ~n38107 & n38108;
  assign n38110 = ~n38104 & ~n38109;
  assign n38111 = n11517 & ~n38110;
  assign n38112 = n38095 & n38111;
  assign n38113 = ~n38098 & ~n38112;
  assign n38114 = ~n38102 & n38113;
  assign n38115 = pi0332 & ~n38114;
  assign n38116 = ~n2741 & ~n2986;
  assign n38117 = pi0137 & ~n38116;
  assign n38118 = pi1093 & ~n3023;
  assign n38119 = ~n38104 & ~n38118;
  assign n38120 = n11549 & ~n38119;
  assign n38121 = ~n38111 & ~n38120;
  assign n38122 = ~n38117 & n38121;
  assign n38123 = ~pi0332 & ~n38122;
  assign n38124 = ~n38115 & ~n38123;
  assign n38125 = ~n2640 & n38124;
  assign n38126 = ~pi0137 & ~n38084;
  assign n38127 = ~n38102 & ~n38126;
  assign n38128 = pi0332 & ~n38127;
  assign n38129 = ~n3024 & ~n38117;
  assign n38130 = ~pi0332 & ~n38129;
  assign n38131 = ~n38128 & ~n38130;
  assign n38132 = n2640 & n38131;
  assign n38133 = ~pi0210 & ~n38125;
  assign n38134 = ~n38132 & n38133;
  assign n38135 = pi0299 & ~n38083;
  assign n38136 = ~n38134 & n38135;
  assign n38137 = pi0198 & ~n38082;
  assign n38138 = n6260 & n38131;
  assign n38139 = ~n6260 & n38124;
  assign n38140 = ~pi0198 & ~n38138;
  assign n38141 = ~n38139 & n38140;
  assign n38142 = ~pi0299 & ~n38137;
  assign n38143 = ~n38141 & n38142;
  assign n38144 = ~n38136 & ~n38143;
  assign n38145 = ~pi0039 & ~n38144;
  assign n38146 = ~pi0038 & ~n38064;
  assign n38147 = ~n38145 & n38146;
  assign n38148 = n6137 & ~n38063;
  assign n38149 = ~n38147 & n38148;
  assign n38150 = ~n38062 & ~n38149;
  assign n38151 = ~pi0087 & ~n38150;
  assign n38152 = ~pi0075 & ~n38061;
  assign n38153 = ~n38151 & n38152;
  assign n38154 = ~pi0092 & ~n38060;
  assign n38155 = ~n38153 & n38154;
  assign n38156 = ~pi0054 & ~n38056;
  assign n38157 = ~n38155 & n38156;
  assign n38158 = ~pi0074 & ~n38054;
  assign n38159 = ~n38157 & n38158;
  assign n38160 = pi0074 & n6128;
  assign n38161 = n38048 & n38160;
  assign n38162 = ~pi0055 & ~n38161;
  assign n38163 = ~n38159 & n38162;
  assign n38164 = n7348 & ~n38163;
  assign n38165 = pi0056 & n2536;
  assign n38166 = n38048 & n38165;
  assign n38167 = ~n38164 & ~n38166;
  assign n38168 = ~pi0062 & ~n38167;
  assign n38169 = n3328 & ~n38052;
  assign n38170 = ~n38168 & n38169;
  assign n38171 = ~n6120 & ~n38051;
  assign po0382 = ~n38170 & n38171;
  assign n38173 = pi0228 & pi0231;
  assign n38174 = ~n7360 & ~n38173;
  assign n38175 = pi0056 & ~n38174;
  assign n38176 = pi0055 & ~n38173;
  assign n38177 = ~n7364 & ~n38173;
  assign n38178 = pi0074 & ~n38177;
  assign n38179 = pi0054 & ~n38173;
  assign n38180 = ~n13971 & ~n38173;
  assign n38181 = pi0075 & ~n38180;
  assign n38182 = pi0087 & ~n38173;
  assign n38183 = ~n7356 & n38182;
  assign n38184 = ~n13975 & ~n38173;
  assign n38185 = pi0100 & ~n38184;
  assign n38186 = ~n2730 & ~n3123;
  assign n38187 = ~pi0070 & ~n38186;
  assign n38188 = ~pi0051 & ~n38187;
  assign n38189 = n2748 & ~n38188;
  assign n38190 = n3168 & ~n38189;
  assign n38191 = n2746 & ~n38190;
  assign n38192 = n2744 & ~n38191;
  assign n38193 = ~n6176 & ~n38192;
  assign n38194 = ~pi0095 & ~n38193;
  assign n38195 = n2742 & ~n38194;
  assign n38196 = ~pi0039 & ~n38195;
  assign n38197 = ~pi0038 & ~n3402;
  assign n38198 = ~n38196 & n38197;
  assign n38199 = ~pi0228 & n38198;
  assign n38200 = ~n38173 & ~n38199;
  assign n38201 = ~pi0100 & ~n38200;
  assign n38202 = ~pi0087 & ~n38185;
  assign n38203 = ~n38201 & n38202;
  assign n38204 = ~pi0075 & ~n38183;
  assign n38205 = ~n38203 & n38204;
  assign n38206 = ~pi0092 & ~n38181;
  assign n38207 = ~n38205 & n38206;
  assign n38208 = pi0092 & ~n38173;
  assign n38209 = ~n7369 & n38208;
  assign n38210 = ~n38207 & ~n38209;
  assign n38211 = ~pi0054 & ~n38210;
  assign n38212 = ~pi0074 & ~n38179;
  assign n38213 = ~n38211 & n38212;
  assign n38214 = ~pi0055 & ~n38178;
  assign n38215 = ~n38213 & n38214;
  assign n38216 = ~pi0056 & ~n38176;
  assign n38217 = ~n38215 & n38216;
  assign n38218 = ~pi0062 & ~n38175;
  assign n38219 = ~n38217 & n38218;
  assign n38220 = pi0062 & ~n38173;
  assign n38221 = ~n7357 & n38220;
  assign n38222 = ~n38219 & ~n38221;
  assign n38223 = n3328 & ~n38222;
  assign n38224 = ~n3328 & ~n38173;
  assign po0383 = ~n38223 & ~n38224;
  assign n38226 = n13080 & ~n13116;
  assign n38227 = n6480 & n38226;
  assign n38228 = ~n6395 & ~n38227;
  assign n38229 = pi1093 & ~n38228;
  assign n38230 = n2708 & n6420;
  assign n38231 = ~pi0091 & ~n2761;
  assign n38232 = n38230 & ~n38231;
  assign n38233 = ~pi0072 & ~n38232;
  assign n38234 = n11022 & n38230;
  assign n38235 = ~n7417 & n38234;
  assign n38236 = ~n8903 & n38233;
  assign n38237 = ~n38235 & n38236;
  assign n38238 = n6480 & ~n38237;
  assign n38239 = ~n38229 & ~n38238;
  assign n38240 = n38233 & ~n38234;
  assign n38241 = n6480 & ~n38240;
  assign n38242 = n10074 & ~n38241;
  assign n38243 = ~n2932 & n11022;
  assign n38244 = n2754 & n11031;
  assign n38245 = n11029 & n38244;
  assign n38246 = n38231 & ~n38243;
  assign n38247 = ~n38245 & n38246;
  assign n38248 = n38230 & ~n38247;
  assign n38249 = ~pi0072 & ~n38248;
  assign n38250 = n6480 & ~n38249;
  assign n38251 = pi0829 & ~n6215;
  assign n38252 = ~n38250 & n38251;
  assign n38253 = ~n38239 & ~n38242;
  assign n38254 = ~n38252 & n38253;
  assign n38255 = ~pi0039 & ~n38254;
  assign po0384 = ~n11471 | n38255;
  assign n38257 = ~pi0039 & pi0228;
  assign n38258 = ~n11420 & ~n11425;
  assign n38259 = pi0039 & ~n38258;
  assign n38260 = n6391 & n38259;
  assign n38261 = ~n2930 & ~n8904;
  assign n38262 = ~pi0032 & n10235;
  assign n38263 = ~n38261 & n38262;
  assign n38264 = n2967 & n38263;
  assign n38265 = ~n11487 & n38264;
  assign n38266 = ~n38260 & ~n38265;
  assign n38267 = n10200 & ~n38266;
  assign po0385 = n38257 | n38267;
  assign n38269 = ~n6136 & n10197;
  assign n38270 = pi0120 & n6218;
  assign n38271 = n16652 & ~n38270;
  assign n38272 = ~n35677 & ~n38271;
  assign n38273 = ~n6205 & ~n38272;
  assign n38274 = ~n6198 & n16652;
  assign n38275 = ~n38271 & ~n38274;
  assign n38276 = n6205 & ~n38275;
  assign n38277 = pi0223 & ~n38273;
  assign n38278 = ~n38276 & n38277;
  assign n38279 = n2603 & n16652;
  assign n38280 = ~n6213 & n7517;
  assign n38281 = n16661 & n38280;
  assign n38282 = n16649 & ~n38280;
  assign n38283 = pi1091 & ~n38281;
  assign n38284 = ~n38282 & n38283;
  assign n38285 = n6383 & n16661;
  assign n38286 = ~n6383 & n16649;
  assign n38287 = ~pi1091 & ~n38285;
  assign n38288 = ~n38286 & n38287;
  assign n38289 = ~n38284 & ~n38288;
  assign n38290 = ~pi0120 & ~n38289;
  assign n38291 = ~n16651 & ~n38290;
  assign n38292 = ~n6227 & n38291;
  assign n38293 = ~n35677 & ~n38292;
  assign n38294 = ~n6205 & n38293;
  assign n38295 = n6198 & n38291;
  assign n38296 = ~n38274 & ~n38295;
  assign n38297 = n6205 & n38296;
  assign n38298 = ~n2603 & ~n38294;
  assign n38299 = ~n38297 & n38298;
  assign n38300 = ~pi0223 & ~n38279;
  assign n38301 = ~n38299 & n38300;
  assign n38302 = ~pi0299 & ~n38278;
  assign n38303 = ~n38301 & n38302;
  assign n38304 = ~n6242 & ~n38272;
  assign n38305 = n6242 & ~n38275;
  assign n38306 = pi0215 & ~n38304;
  assign n38307 = ~n38305 & n38306;
  assign n38308 = ~n6242 & n38293;
  assign n38309 = n6242 & n38296;
  assign n38310 = ~n3448 & ~n38308;
  assign n38311 = ~n38309 & n38310;
  assign n38312 = ~pi0215 & ~n16825;
  assign n38313 = ~n38311 & n38312;
  assign n38314 = pi0299 & ~n38307;
  assign n38315 = ~n38313 & n38314;
  assign n38316 = ~n38303 & ~n38315;
  assign n38317 = pi0039 & ~n38316;
  assign n38318 = n6170 & n16854;
  assign n38319 = ~n16856 & n38318;
  assign n38320 = ~pi0040 & ~n38319;
  assign n38321 = n10289 & ~n38320;
  assign n38322 = pi0252 & ~n38321;
  assign n38323 = n6277 & ~n16853;
  assign n38324 = ~n38322 & n38323;
  assign n38325 = ~n6277 & n16866;
  assign n38326 = ~pi1093 & ~n38324;
  assign n38327 = ~n38325 & n38326;
  assign n38328 = ~n6169 & ~n6387;
  assign n38329 = ~n7417 & n16866;
  assign n38330 = ~n16883 & ~n38329;
  assign n38331 = n38328 & ~n38330;
  assign n38332 = pi0829 & pi1091;
  assign n38333 = n16907 & n38332;
  assign n38334 = ~pi0824 & ~n38333;
  assign n38335 = pi0824 & ~n16902;
  assign n38336 = ~n6387 & ~n38334;
  assign n38337 = ~n38335 & n38336;
  assign n38338 = ~n16866 & ~n38337;
  assign n38339 = n38332 & n38334;
  assign n38340 = ~n38335 & ~n38339;
  assign n38341 = n2932 & ~n6387;
  assign n38342 = ~n38340 & n38341;
  assign n38343 = ~n38328 & ~n38338;
  assign n38344 = ~n38342 & n38343;
  assign n38345 = pi1093 & ~n38331;
  assign n38346 = ~n38344 & n38345;
  assign n38347 = ~pi0039 & ~n38327;
  assign n38348 = ~n38346 & n38347;
  assign n38349 = ~pi0038 & ~n38317;
  assign n38350 = ~n38348 & n38349;
  assign po0387 = n38269 & ~n38350;
  assign n38352 = ~pi0081 & ~n2865;
  assign n38353 = n6443 & ~n38352;
  assign n38354 = n2462 & ~n38353;
  assign n38355 = n2873 & ~n38354;
  assign n38356 = n2785 & ~n38355;
  assign n38357 = n2877 & ~n38356;
  assign n38358 = n2719 & ~n38357;
  assign n38359 = ~n2722 & ~n38358;
  assign n38360 = ~pi0086 & ~n38359;
  assign n38361 = n2783 & ~n38360;
  assign n38362 = n2781 & ~n38361;
  assign n38363 = ~n2776 & ~n38362;
  assign n38364 = ~pi0108 & ~n38363;
  assign n38365 = n2775 & ~n38364;
  assign n38366 = n2889 & ~n38365;
  assign n38367 = ~n2766 & ~n38366;
  assign n38368 = n2765 & ~n38367;
  assign n38369 = n2764 & ~n38368;
  assign n38370 = n2757 & ~n38369;
  assign n38371 = n3108 & ~n38370;
  assign n38372 = n2504 & ~n38371;
  assign n38373 = n15635 & ~n38372;
  assign n38374 = ~pi0070 & ~n38373;
  assign n38375 = ~n3099 & ~n38374;
  assign n38376 = ~pi0051 & ~n38375;
  assign n38377 = n2748 & ~n38376;
  assign n38378 = n3168 & ~n38377;
  assign n38379 = n2746 & ~n38378;
  assign n38380 = ~pi1082 & n2743;
  assign n38381 = ~pi0032 & ~n38380;
  assign n38382 = ~n38379 & n38381;
  assign n38383 = ~n3412 & ~n38382;
  assign n38384 = ~pi0095 & ~n38383;
  assign n38385 = ~n2741 & ~n38384;
  assign n38386 = ~pi0039 & ~n38385;
  assign n38387 = ~n7307 & ~n7309;
  assign po0950 = ~n2932 | ~n6217;
  assign n38389 = n6381 & ~po0950;
  assign n38390 = ~n38387 & n38389;
  assign n38391 = n6185 & n11369;
  assign n38392 = ~n38390 & n38391;
  assign n38393 = ~n3402 & ~n38392;
  assign n38394 = ~n38386 & n38393;
  assign n38395 = ~pi0038 & ~n38394;
  assign n38396 = n6137 & ~n38395;
  assign n38397 = ~pi0087 & ~n6286;
  assign n38398 = ~n38396 & n38397;
  assign n38399 = ~n6132 & ~n38398;
  assign n38400 = n2569 & ~n38399;
  assign n38401 = n7306 & ~n38400;
  assign n38402 = ~pi0054 & ~n38401;
  assign n38403 = ~n7341 & ~n38402;
  assign n38404 = n8879 & ~n38403;
  assign n38405 = n15712 & ~n38404;
  assign n38406 = ~pi0056 & ~n38405;
  assign n38407 = ~n6127 & ~n38406;
  assign n38408 = ~pi0062 & ~n38407;
  assign n38409 = ~n6299 & ~n38408;
  assign n38410 = n3328 & ~n38409;
  assign po0389 = n6123 & ~n38410;
  assign n38412 = ~pi0230 & ~pi0233;
  assign n38413 = ~pi0212 & ~pi0214;
  assign n38414 = ~pi0211 & ~n38413;
  assign n38415 = pi0219 & ~n38414;
  assign n38416 = po1038 & ~n38415;
  assign n38417 = pi1142 & ~n10486;
  assign n38418 = pi0211 & pi1143;
  assign n38419 = ~pi0211 & pi1144;
  assign n38420 = ~n38418 & ~n38419;
  assign n38421 = ~pi0212 & pi0214;
  assign n38422 = pi0212 & ~pi0214;
  assign n38423 = ~n38421 & ~n38422;
  assign n38424 = ~n38420 & ~n38423;
  assign n38425 = ~pi0211 & pi1143;
  assign n38426 = n10843 & n38425;
  assign n38427 = ~n38424 & ~n38426;
  assign n38428 = ~pi0219 & ~n38427;
  assign n38429 = ~n38417 & ~n38428;
  assign n38430 = n38416 & ~n38429;
  assign n38431 = pi0299 & ~n38420;
  assign n38432 = pi0199 & pi1142;
  assign n38433 = ~pi0200 & ~n38432;
  assign n38434 = ~pi0199 & pi1144;
  assign n38435 = n38433 & ~n38434;
  assign n38436 = ~pi0199 & pi1143;
  assign n38437 = pi0200 & ~n38436;
  assign n38438 = ~n38435 & ~n38437;
  assign n38439 = ~pi0299 & ~n38438;
  assign n38440 = ~pi0207 & ~n38439;
  assign n38441 = pi0207 & ~pi0299;
  assign n38442 = n38433 & ~n38436;
  assign n38443 = ~pi0199 & pi1142;
  assign n38444 = pi0200 & ~n38443;
  assign n38445 = n38441 & ~n38444;
  assign n38446 = ~n38442 & n38445;
  assign n38447 = ~n38440 & ~n38446;
  assign n38448 = pi0208 & ~n38447;
  assign n38449 = pi0207 & ~pi0208;
  assign n38450 = n38438 & n38449;
  assign n38451 = ~n38448 & ~n38450;
  assign n38452 = ~pi0299 & ~n38451;
  assign n38453 = ~pi0214 & ~n38452;
  assign n38454 = ~n38431 & n38453;
  assign n38455 = pi0211 & pi1142;
  assign n38456 = ~n38425 & ~n38455;
  assign n38457 = pi0299 & ~n38456;
  assign n38458 = pi0214 & ~n38457;
  assign n38459 = ~n38452 & n38458;
  assign n38460 = pi0212 & ~n38459;
  assign n38461 = ~n38454 & n38460;
  assign n38462 = ~n38431 & ~n38452;
  assign n38463 = ~pi0212 & ~n38453;
  assign n38464 = ~n38462 & n38463;
  assign n38465 = ~pi0219 & ~n38461;
  assign n38466 = ~n38464 & n38465;
  assign n38467 = ~n38414 & n38452;
  assign n38468 = ~pi0299 & n38451;
  assign n38469 = pi0299 & ~pi1142;
  assign n38470 = n38414 & ~n38469;
  assign n38471 = ~n38468 & n38470;
  assign n38472 = pi0219 & ~n38467;
  assign n38473 = ~n38471 & n38472;
  assign n38474 = ~po1038 & ~n38473;
  assign n38475 = ~n38466 & n38474;
  assign n38476 = ~n38430 & ~n38475;
  assign n38477 = pi0213 & n38476;
  assign n38478 = ~pi0211 & pi1157;
  assign n38479 = pi0211 & pi1156;
  assign n38480 = ~n38478 & ~n38479;
  assign n38481 = pi0214 & ~n38480;
  assign n38482 = ~pi0212 & ~n38481;
  assign n38483 = ~pi0211 & pi1156;
  assign n38484 = pi0211 & pi1155;
  assign n38485 = ~n38483 & ~n38484;
  assign n38486 = ~pi0214 & ~n38485;
  assign n38487 = ~pi0211 & pi1155;
  assign n38488 = pi0211 & pi1154;
  assign n38489 = ~n38487 & ~n38488;
  assign n38490 = pi0214 & ~n38489;
  assign n38491 = ~n38486 & ~n38490;
  assign n38492 = pi0212 & n38491;
  assign n38493 = ~n38482 & ~n38492;
  assign n38494 = ~pi0219 & ~n38493;
  assign n38495 = ~pi0211 & pi1154;
  assign n38496 = ~pi0214 & ~n38495;
  assign n38497 = ~pi0211 & pi1153;
  assign n38498 = n10843 & ~n38497;
  assign n38499 = ~pi0211 & pi0214;
  assign n38500 = pi1155 & n38499;
  assign n38501 = ~pi0212 & ~n38500;
  assign n38502 = ~n38496 & ~n38498;
  assign n38503 = ~n38501 & n38502;
  assign n38504 = pi0219 & ~n38503;
  assign n38505 = po1038 & ~n38504;
  assign n38506 = ~n38494 & n38505;
  assign n38507 = ~pi0213 & ~n38506;
  assign n38508 = ~pi0219 & pi0299;
  assign n38509 = n38493 & n38508;
  assign n38510 = pi0299 & pi1155;
  assign n38511 = n38421 & n38510;
  assign n38512 = pi0299 & pi1153;
  assign n38513 = pi0214 & ~n38512;
  assign n38514 = pi0299 & pi1154;
  assign n38515 = ~pi0214 & ~n38514;
  assign n38516 = pi0212 & ~n38513;
  assign n38517 = ~n38515 & n38516;
  assign n38518 = ~n38511 & ~n38517;
  assign n38519 = ~pi0211 & pi0219;
  assign n38520 = ~n38518 & n38519;
  assign n38521 = ~n38509 & ~n38520;
  assign n38522 = ~n38452 & n38521;
  assign n38523 = ~po1038 & ~n38522;
  assign n38524 = n38507 & ~n38523;
  assign n38525 = pi0209 & ~n38524;
  assign n38526 = ~n38477 & n38525;
  assign n38527 = ~pi0211 & n10843;
  assign n38528 = pi0299 & ~pi1143;
  assign n38529 = ~pi0200 & pi1155;
  assign n38530 = pi0199 & n38529;
  assign n38531 = ~pi0299 & n38530;
  assign n38532 = ~pi1156 & ~n38531;
  assign n38533 = ~pi0299 & ~n11444;
  assign n38534 = pi1156 & ~n38530;
  assign n38535 = n38533 & n38534;
  assign n38536 = ~n38532 & ~n38535;
  assign n38537 = pi0207 & n38536;
  assign n38538 = ~pi0299 & ~n38537;
  assign n38539 = ~pi0208 & ~n38538;
  assign n38540 = ~pi1157 & n38539;
  assign n38541 = ~n38528 & n38540;
  assign n38542 = ~pi0208 & pi1157;
  assign n38543 = pi0299 & pi1143;
  assign n38544 = ~pi1155 & ~n10810;
  assign n38545 = pi0200 & ~pi0299;
  assign n38546 = pi1155 & ~n38545;
  assign n38547 = ~n38544 & ~n38546;
  assign n38548 = pi0199 & ~pi1155;
  assign n38549 = pi0199 & pi0200;
  assign n38550 = ~pi0299 & ~n38549;
  assign n38551 = pi1156 & ~n38548;
  assign n38552 = n38550 & n38551;
  assign n38553 = n38547 & ~n38552;
  assign n38554 = pi0207 & ~n38528;
  assign n38555 = ~n38553 & n38554;
  assign n38556 = ~n38543 & ~n38555;
  assign n38557 = n38542 & ~n38556;
  assign n38558 = pi1153 & ~n38550;
  assign n38559 = pi1154 & ~n38558;
  assign n38560 = n11384 & n38529;
  assign n38561 = ~n10809 & ~n38549;
  assign n38562 = ~pi1153 & ~n11384;
  assign n38563 = pi1154 & n38561;
  assign n38564 = ~n38562 & n38563;
  assign n38565 = ~n38560 & ~n38564;
  assign n38566 = n38559 & ~n38565;
  assign n38567 = ~pi0199 & ~pi1155;
  assign n38568 = ~pi0200 & ~pi0299;
  assign n38569 = pi0199 & ~pi1153;
  assign n38570 = n38568 & ~n38569;
  assign n38571 = ~pi1154 & ~n38567;
  assign n38572 = n38570 & n38571;
  assign n38573 = ~n38566 & ~n38572;
  assign n38574 = pi0207 & n38573;
  assign n38575 = ~n38543 & n38574;
  assign n38576 = ~pi0199 & pi1155;
  assign n38577 = n38545 & n38576;
  assign n38578 = ~pi1154 & ~n38577;
  assign n38579 = ~n38543 & n38578;
  assign n38580 = ~pi1155 & n38543;
  assign n38581 = ~pi0299 & ~n38561;
  assign n38582 = pi1155 & ~n38581;
  assign n38583 = ~n38528 & n38582;
  assign n38584 = ~pi0200 & ~pi1155;
  assign n38585 = n11373 & n38584;
  assign n38586 = pi1154 & ~n38585;
  assign n38587 = ~n38580 & n38586;
  assign n38588 = ~n38583 & n38587;
  assign n38589 = ~pi1156 & ~n38579;
  assign n38590 = ~n38588 & n38589;
  assign n38591 = pi0200 & ~n38576;
  assign n38592 = ~pi0299 & ~n38591;
  assign n38593 = pi1154 & ~n38592;
  assign n38594 = ~n38543 & n38593;
  assign n38595 = pi1155 & ~n11373;
  assign n38596 = ~n38544 & ~n38595;
  assign n38597 = ~n38528 & ~n38596;
  assign n38598 = ~pi1154 & ~n38597;
  assign n38599 = pi1156 & ~n38594;
  assign n38600 = ~n38598 & n38599;
  assign n38601 = ~n38590 & ~n38600;
  assign n38602 = ~pi0207 & n38601;
  assign n38603 = pi0208 & ~n38575;
  assign n38604 = ~n38602 & n38603;
  assign n38605 = ~n38541 & ~n38557;
  assign n38606 = ~n38604 & n38605;
  assign n38607 = n38527 & n38606;
  assign n38608 = ~n10843 & ~n38413;
  assign n38609 = pi0211 & ~n38606;
  assign n38610 = pi0299 & ~pi1144;
  assign n38611 = n38540 & ~n38610;
  assign n38612 = pi0299 & pi1144;
  assign n38613 = pi0207 & ~n38610;
  assign n38614 = ~n38553 & n38613;
  assign n38615 = ~n38612 & ~n38614;
  assign n38616 = n38542 & ~n38615;
  assign n38617 = n38574 & ~n38612;
  assign n38618 = n38578 & ~n38612;
  assign n38619 = ~pi1155 & n38612;
  assign n38620 = n38582 & ~n38610;
  assign n38621 = n38586 & ~n38619;
  assign n38622 = ~n38620 & n38621;
  assign n38623 = ~pi1156 & ~n38618;
  assign n38624 = ~n38622 & n38623;
  assign n38625 = n38593 & ~n38612;
  assign n38626 = ~n38596 & ~n38610;
  assign n38627 = ~pi1154 & ~n38626;
  assign n38628 = pi1156 & ~n38625;
  assign n38629 = ~n38627 & n38628;
  assign n38630 = ~n38624 & ~n38629;
  assign n38631 = ~pi0207 & n38630;
  assign n38632 = pi0208 & ~n38617;
  assign n38633 = ~n38631 & n38632;
  assign n38634 = ~n38611 & ~n38616;
  assign n38635 = ~n38633 & n38634;
  assign n38636 = ~pi0211 & ~n38635;
  assign n38637 = n38608 & ~n38609;
  assign n38638 = ~n38636 & n38637;
  assign n38639 = ~n38607 & ~n38638;
  assign n38640 = ~pi0219 & ~n38639;
  assign n38641 = ~pi0299 & n38561;
  assign n38642 = ~n38584 & n38641;
  assign n38643 = ~n38532 & n38642;
  assign n38644 = pi0207 & n38643;
  assign n38645 = ~pi0208 & ~n38644;
  assign n38646 = n10810 & ~n38591;
  assign n38647 = ~n38578 & n38646;
  assign n38648 = pi0200 & ~pi1155;
  assign n38649 = n11384 & ~n38648;
  assign n38650 = pi1156 & n38649;
  assign n38651 = ~n38647 & ~n38650;
  assign n38652 = ~pi0207 & n38651;
  assign n38653 = ~n38574 & ~n38652;
  assign n38654 = pi0208 & ~n38653;
  assign n38655 = ~n38645 & ~n38654;
  assign n38656 = ~pi1157 & ~n38655;
  assign n38657 = ~pi1156 & ~n38548;
  assign n38658 = n38568 & n38657;
  assign n38659 = ~n38552 & ~n38658;
  assign n38660 = pi0207 & ~n38659;
  assign n38661 = ~pi0208 & ~n38660;
  assign n38662 = ~n38654 & ~n38661;
  assign n38663 = pi1157 & ~n38662;
  assign n38664 = ~n38656 & ~n38663;
  assign n38665 = ~pi0219 & ~n38413;
  assign n38666 = ~n38414 & ~n38665;
  assign n38667 = ~n38664 & n38666;
  assign n38668 = ~pi1157 & ~n38539;
  assign n38669 = ~pi1156 & ~n38547;
  assign n38670 = n11373 & ~n38529;
  assign n38671 = pi1156 & ~n38670;
  assign n38672 = ~n38669 & ~n38671;
  assign n38673 = pi0207 & n38672;
  assign n38674 = ~pi0207 & ~pi0299;
  assign n38675 = ~pi0208 & ~n38674;
  assign n38676 = ~n38673 & n38675;
  assign n38677 = pi1157 & ~n38676;
  assign n38678 = ~n38469 & ~n38668;
  assign n38679 = ~n38677 & n38678;
  assign n38680 = pi0299 & pi1142;
  assign n38681 = pi1153 & n38585;
  assign n38682 = pi1153 & ~n38545;
  assign n38683 = ~pi1153 & ~n10810;
  assign n38684 = ~n38682 & ~n38683;
  assign n38685 = pi1155 & ~n38684;
  assign n38686 = ~n38681 & ~n38685;
  assign n38687 = ~pi1154 & ~n38686;
  assign n38688 = ~n38569 & n38641;
  assign n38689 = ~n38595 & ~n38688;
  assign n38690 = pi1154 & ~n38689;
  assign n38691 = ~n38687 & ~n38690;
  assign n38692 = ~pi0299 & ~n38691;
  assign n38693 = pi0207 & ~n38680;
  assign n38694 = ~n38692 & n38693;
  assign n38695 = ~n38577 & ~n38680;
  assign n38696 = ~pi1154 & ~pi1156;
  assign n38697 = ~n38695 & n38696;
  assign n38698 = pi1156 & ~n38596;
  assign n38699 = pi0199 & ~pi0200;
  assign n38700 = ~pi0299 & ~n38699;
  assign n38701 = ~pi1155 & ~n38700;
  assign n38702 = ~n38582 & ~n38701;
  assign n38703 = pi1154 & ~n38702;
  assign n38704 = ~n38698 & ~n38703;
  assign n38705 = ~n38469 & ~n38704;
  assign n38706 = ~pi0207 & ~n38697;
  assign n38707 = ~n38705 & n38706;
  assign n38708 = pi0208 & ~n38707;
  assign n38709 = ~n38694 & n38708;
  assign n38710 = ~n10486 & ~n38666;
  assign n38711 = ~n38679 & n38710;
  assign n38712 = ~n38709 & n38711;
  assign n38713 = ~po1038 & ~n38712;
  assign n38714 = ~n38667 & n38713;
  assign n38715 = ~n38640 & n38714;
  assign n38716 = pi0213 & ~n38430;
  assign n38717 = ~n38715 & n38716;
  assign n38718 = pi0211 & ~n38664;
  assign n38719 = ~pi0214 & ~n38664;
  assign n38720 = ~pi0212 & ~n38719;
  assign n38721 = ~pi0207 & ~n38510;
  assign n38722 = ~pi0208 & ~n38721;
  assign n38723 = ~n11384 & ~n38546;
  assign n38724 = pi1156 & ~n38723;
  assign n38725 = ~pi1156 & ~n38545;
  assign n38726 = ~n38701 & n38725;
  assign n38727 = ~n38724 & ~n38726;
  assign n38728 = pi0207 & n38727;
  assign n38729 = pi1157 & n38722;
  assign n38730 = ~n38728 & n38729;
  assign n38731 = ~pi1155 & ~n11384;
  assign n38732 = ~pi0299 & n38532;
  assign n38733 = ~n38581 & ~n38731;
  assign n38734 = ~n38732 & n38733;
  assign n38735 = n38722 & n38734;
  assign n38736 = pi0207 & n38691;
  assign n38737 = n38651 & n38721;
  assign n38738 = pi0208 & ~n38737;
  assign n38739 = ~n38736 & n38738;
  assign n38740 = ~n38730 & ~n38735;
  assign n38741 = ~n38739 & n38740;
  assign n38742 = n38499 & n38741;
  assign n38743 = n38720 & ~n38742;
  assign n38744 = ~pi0211 & ~pi0214;
  assign n38745 = pi0299 & ~pi1154;
  assign n38746 = pi1157 & ~n38745;
  assign n38747 = n38676 & n38746;
  assign n38748 = n38651 & ~n38703;
  assign n38749 = ~pi0207 & ~n38748;
  assign n38750 = ~pi0299 & n38689;
  assign n38751 = pi1154 & ~n38750;
  assign n38752 = ~n38572 & ~n38751;
  assign n38753 = pi0207 & ~n38752;
  assign n38754 = ~n38749 & ~n38753;
  assign n38755 = pi0208 & ~n38754;
  assign n38756 = ~n38514 & ~n38644;
  assign n38757 = ~pi0208 & ~n38756;
  assign n38758 = ~pi1157 & n38757;
  assign n38759 = ~n38747 & ~n38758;
  assign n38760 = ~n38755 & n38759;
  assign n38761 = n38744 & n38760;
  assign n38762 = pi1153 & ~n38700;
  assign n38763 = n38565 & ~n38762;
  assign n38764 = pi0207 & ~n38763;
  assign n38765 = pi0299 & ~pi1155;
  assign n38766 = pi1155 & ~n38533;
  assign n38767 = ~n38765 & ~n38766;
  assign n38768 = n38704 & n38767;
  assign n38769 = pi0299 & ~pi1153;
  assign n38770 = ~pi0207 & ~n38769;
  assign n38771 = ~n38768 & n38770;
  assign n38772 = ~n38764 & ~n38771;
  assign n38773 = pi0208 & ~n38772;
  assign n38774 = ~n38668 & ~n38769;
  assign n38775 = ~n38677 & n38774;
  assign n38776 = n38499 & ~n38773;
  assign n38777 = ~n38775 & n38776;
  assign n38778 = pi0212 & ~n38761;
  assign n38779 = ~n38777 & n38778;
  assign n38780 = ~n38743 & ~n38779;
  assign n38781 = ~n38718 & ~n38780;
  assign n38782 = pi0219 & ~n38781;
  assign n38783 = ~n10484 & ~n38744;
  assign n38784 = ~n38741 & n38783;
  assign n38785 = n10484 & ~n38760;
  assign n38786 = ~n38532 & n38539;
  assign n38787 = pi0299 & pi1156;
  assign n38788 = ~n38660 & ~n38787;
  assign n38789 = n38542 & ~n38788;
  assign n38790 = pi0207 & ~n38573;
  assign n38791 = ~n38647 & ~n38698;
  assign n38792 = ~pi0207 & ~n38791;
  assign n38793 = pi0207 & n38787;
  assign n38794 = ~n38792 & ~n38793;
  assign n38795 = ~n38790 & n38794;
  assign n38796 = pi0208 & ~n38795;
  assign n38797 = ~n38786 & ~n38789;
  assign n38798 = ~n38796 & n38797;
  assign n38799 = n38744 & ~n38798;
  assign n38800 = ~n38784 & ~n38799;
  assign n38801 = ~n38785 & n38800;
  assign n38802 = pi0212 & ~n38801;
  assign n38803 = pi0211 & ~n38798;
  assign n38804 = ~pi0207 & n38768;
  assign n38805 = n38441 & n38763;
  assign n38806 = pi0208 & ~n38805;
  assign n38807 = ~n38804 & n38806;
  assign n38808 = n38677 & ~n38807;
  assign n38809 = ~pi0211 & ~n38808;
  assign n38810 = ~n38656 & n38809;
  assign n38811 = pi0214 & ~n38803;
  assign n38812 = ~n38810 & n38811;
  assign n38813 = n38720 & ~n38812;
  assign n38814 = ~pi0219 & ~n38802;
  assign n38815 = ~n38813 & n38814;
  assign n38816 = ~po1038 & ~n38815;
  assign n38817 = ~n38782 & n38816;
  assign n38818 = n38507 & ~n38817;
  assign n38819 = ~pi0209 & ~n38717;
  assign n38820 = ~n38818 & n38819;
  assign n38821 = ~n38526 & ~n38820;
  assign n38822 = pi0230 & ~n38821;
  assign po0390 = n38412 | n38822;
  assign n38824 = ~n10487 & n38651;
  assign n38825 = ~pi0207 & ~pi0208;
  assign n38826 = ~n10487 & ~n38825;
  assign n38827 = ~pi0199 & n38584;
  assign n38828 = ~pi1154 & ~n38560;
  assign n38829 = n38550 & ~n38827;
  assign n38830 = ~n38828 & n38829;
  assign n38831 = pi0207 & n38830;
  assign n38832 = ~n38826 & ~n38831;
  assign n38833 = ~n38824 & ~n38832;
  assign n38834 = ~n38414 & n38833;
  assign n38835 = pi0219 & ~n38834;
  assign n38836 = ~pi0207 & n38514;
  assign n38837 = pi0207 & ~n38748;
  assign n38838 = ~n38836 & ~n38837;
  assign n38839 = ~pi0208 & ~n38838;
  assign n38840 = ~pi1155 & n10809;
  assign n38841 = ~n38549 & ~n38840;
  assign n38842 = ~pi0299 & ~n38841;
  assign n38843 = ~n38828 & ~n38842;
  assign n38844 = pi0207 & n38843;
  assign n38845 = ~n38749 & ~n38844;
  assign n38846 = pi0208 & ~n38845;
  assign n38847 = ~n38839 & ~n38846;
  assign n38848 = ~pi0211 & ~n38847;
  assign n38849 = ~n38413 & n38848;
  assign n38850 = n38835 & ~n38849;
  assign n38851 = ~pi0214 & ~n38833;
  assign n38852 = ~pi0212 & ~n38851;
  assign n38853 = pi0207 & ~n38791;
  assign n38854 = ~n38787 & ~n38853;
  assign n38855 = ~pi0208 & ~n38854;
  assign n38856 = n38794 & ~n38831;
  assign n38857 = pi0208 & ~n38856;
  assign n38858 = ~n38855 & ~n38857;
  assign n38859 = ~pi0211 & ~n38858;
  assign n38860 = ~n38510 & n38651;
  assign n38861 = n38722 & ~n38860;
  assign n38862 = pi0207 & ~n38510;
  assign n38863 = ~n38830 & n38862;
  assign n38864 = pi0208 & ~n38863;
  assign n38865 = ~n38737 & n38864;
  assign n38866 = ~n38861 & ~n38865;
  assign n38867 = pi0211 & ~n38866;
  assign n38868 = ~n38859 & ~n38867;
  assign n38869 = pi0214 & n38868;
  assign n38870 = n38852 & ~n38869;
  assign n38871 = pi0211 & ~n38847;
  assign n38872 = ~pi0211 & ~n38866;
  assign n38873 = pi0214 & ~n38872;
  assign n38874 = ~n38871 & n38873;
  assign n38875 = ~pi0214 & n38868;
  assign n38876 = pi0212 & ~n38874;
  assign n38877 = ~n38875 & n38876;
  assign n38878 = ~pi0219 & ~n38870;
  assign n38879 = ~n38877 & n38878;
  assign n38880 = n35819 & ~n38850;
  assign n38881 = ~n38879 & n38880;
  assign n38882 = pi0211 & pi1153;
  assign n38883 = ~n38495 & ~n38882;
  assign n38884 = ~n10843 & n38883;
  assign n38885 = n38665 & ~n38884;
  assign n38886 = ~n38498 & n38885;
  assign n38887 = po1038 & n38886;
  assign n38888 = ~pi1152 & ~n38887;
  assign n38889 = pi0207 & n38767;
  assign n38890 = n38704 & n38889;
  assign n38891 = n38675 & ~n38890;
  assign n38892 = n38441 & ~n38843;
  assign n38893 = pi0208 & ~n38892;
  assign n38894 = ~n38804 & n38893;
  assign n38895 = ~n38891 & ~n38894;
  assign n38896 = ~n38769 & ~n38895;
  assign n38897 = pi0211 & n38896;
  assign n38898 = ~n38848 & ~n38897;
  assign n38899 = pi0214 & n38898;
  assign n38900 = n38852 & ~n38899;
  assign n38901 = ~pi0219 & ~n38900;
  assign n38902 = ~pi0214 & ~n38898;
  assign n38903 = ~pi0211 & ~n38896;
  assign n38904 = pi0214 & ~n38903;
  assign n38905 = pi0211 & ~n38833;
  assign n38906 = n38904 & ~n38905;
  assign n38907 = ~n38902 & ~n38906;
  assign n38908 = pi0212 & ~n38907;
  assign n38909 = n38901 & ~n38908;
  assign n38910 = pi0219 & ~n38833;
  assign n38911 = ~po1038 & ~n38910;
  assign n38912 = ~n38909 & n38911;
  assign n38913 = n38888 & ~n38912;
  assign n38914 = pi1153 & ~n38744;
  assign n38915 = ~n38496 & ~n38499;
  assign n38916 = ~n38914 & ~n38915;
  assign n38917 = pi0212 & ~n38916;
  assign n38918 = n38421 & ~n38883;
  assign n38919 = ~pi0219 & ~n38918;
  assign n38920 = ~n38917 & n38919;
  assign n38921 = n38416 & ~n38920;
  assign n38922 = pi1152 & ~n38921;
  assign n38923 = ~n38895 & n38904;
  assign n38924 = ~n38902 & ~n38923;
  assign n38925 = pi0212 & ~n38924;
  assign n38926 = n38901 & ~n38925;
  assign n38927 = n38414 & ~n38895;
  assign n38928 = n38835 & ~n38927;
  assign n38929 = ~po1038 & ~n38928;
  assign n38930 = ~n38926 & n38929;
  assign n38931 = n38922 & ~n38930;
  assign n38932 = ~pi0213 & ~n38913;
  assign n38933 = ~n38931 & n38932;
  assign n38934 = pi0209 & ~n38881;
  assign n38935 = ~n38933 & n38934;
  assign n38936 = ~pi0199 & pi1153;
  assign n38937 = pi0200 & n38936;
  assign n38938 = ~pi0299 & n38937;
  assign n38939 = ~pi1154 & ~n38938;
  assign n38940 = pi1154 & n38545;
  assign n38941 = ~n38936 & n38940;
  assign n38942 = ~n38939 & ~n38941;
  assign n38943 = n38700 & ~n38942;
  assign n38944 = n38675 & ~n38943;
  assign n38945 = ~pi0200 & ~pi1153;
  assign n38946 = ~pi0199 & ~n38945;
  assign n38947 = ~pi0299 & ~n38946;
  assign n38948 = ~n38699 & n38947;
  assign n38949 = pi0207 & n38948;
  assign n38950 = ~pi0207 & n38943;
  assign n38951 = pi0208 & ~n38949;
  assign n38952 = ~n38950 & n38951;
  assign n38953 = ~n38944 & ~n38952;
  assign n38954 = ~pi0211 & n38953;
  assign n38955 = ~pi0299 & n10809;
  assign n38956 = ~pi1153 & ~n38955;
  assign n38957 = n38559 & ~n38956;
  assign n38958 = ~pi0199 & ~pi1153;
  assign n38959 = n38641 & ~n38958;
  assign n38960 = ~n38957 & ~n38959;
  assign n38961 = ~n10487 & n38960;
  assign n38962 = ~pi1153 & n10809;
  assign n38963 = n38550 & ~n38962;
  assign n38964 = n10487 & ~n38963;
  assign n38965 = ~n38825 & ~n38964;
  assign n38966 = ~n38961 & n38965;
  assign n38967 = pi0211 & ~n38966;
  assign n38968 = ~n38954 & ~n38967;
  assign n38969 = ~n38413 & n38968;
  assign n38970 = pi0219 & ~n38413;
  assign n38971 = pi0219 & ~n38966;
  assign n38972 = ~n38970 & ~n38971;
  assign n38973 = ~n38969 & ~n38972;
  assign n38974 = ~po1038 & ~n38973;
  assign n38975 = ~pi0207 & n38512;
  assign n38976 = ~pi1153 & ~n38568;
  assign n38977 = ~n38581 & ~n38976;
  assign n38978 = pi1154 & ~n11373;
  assign n38979 = ~n38976 & n38978;
  assign n38980 = ~n38977 & ~n38979;
  assign n38981 = pi0207 & ~n38980;
  assign n38982 = ~n38975 & ~n38981;
  assign n38983 = ~pi0208 & ~n38982;
  assign n38984 = ~pi0207 & ~n38980;
  assign n38985 = ~pi0299 & n38549;
  assign n38986 = pi0207 & ~n38985;
  assign n38987 = ~n38683 & n38986;
  assign n38988 = ~n38984 & ~n38987;
  assign n38989 = pi0208 & ~n38988;
  assign n38990 = ~n38983 & ~n38989;
  assign n38991 = ~pi0211 & ~n38990;
  assign n38992 = pi0211 & ~n38953;
  assign n38993 = pi0214 & ~n38991;
  assign n38994 = ~n38992 & n38993;
  assign n38995 = pi0207 & ~n38960;
  assign n38996 = ~n38514 & ~n38995;
  assign n38997 = ~pi0208 & ~n38996;
  assign n38998 = pi0207 & ~n38948;
  assign n38999 = ~n38745 & n38998;
  assign n39000 = pi1154 & ~n10810;
  assign n39001 = ~n38957 & ~n39000;
  assign n39002 = ~n38959 & n39001;
  assign n39003 = ~pi0207 & ~n39002;
  assign n39004 = ~n38999 & ~n39003;
  assign n39005 = pi0208 & ~n39004;
  assign n39006 = ~n38997 & ~n39005;
  assign n39007 = ~pi0211 & ~n39006;
  assign n39008 = pi0211 & ~n38990;
  assign n39009 = ~n39007 & ~n39008;
  assign n39010 = ~pi0214 & n39009;
  assign n39011 = pi0212 & ~n38994;
  assign n39012 = ~n39010 & n39011;
  assign n39013 = ~pi0214 & ~n38966;
  assign n39014 = ~pi0212 & ~n39013;
  assign n39015 = pi0214 & n39009;
  assign n39016 = n39014 & ~n39015;
  assign n39017 = ~pi0219 & ~n39012;
  assign n39018 = ~n39016 & n39017;
  assign n39019 = n38974 & ~n39018;
  assign n39020 = n38922 & ~n39019;
  assign n39021 = pi0200 & ~pi1153;
  assign n39022 = n11384 & ~n39021;
  assign n39023 = pi1154 & ~n39022;
  assign n39024 = ~n38939 & ~n39023;
  assign n39025 = n38826 & n39024;
  assign n39026 = pi0208 & n38441;
  assign n39027 = pi1153 & ~n10810;
  assign n39028 = n39026 & n39027;
  assign n39029 = ~n39025 & ~n39028;
  assign n39030 = pi0219 & n39029;
  assign n39031 = ~po1038 & ~n39030;
  assign n39032 = pi1153 & ~pi1154;
  assign n39033 = ~n38533 & n39032;
  assign n39034 = ~n38979 & ~n39033;
  assign n39035 = pi0207 & ~n39034;
  assign n39036 = ~n38975 & ~n39035;
  assign n39037 = ~pi0208 & ~n39036;
  assign n39038 = ~pi0207 & ~n39034;
  assign n39039 = pi0207 & ~n10810;
  assign n39040 = pi1153 & n39039;
  assign n39041 = ~n39038 & ~n39040;
  assign n39042 = pi0208 & ~n39041;
  assign n39043 = ~n39037 & ~n39042;
  assign n39044 = n38527 & n39043;
  assign n39045 = pi1153 & ~n11373;
  assign n39046 = ~n38683 & ~n39045;
  assign n39047 = pi1154 & ~n39046;
  assign n39048 = ~n38938 & ~n39047;
  assign n39049 = pi0207 & ~n39048;
  assign n39050 = ~n38836 & ~n39049;
  assign n39051 = ~pi0208 & ~n39050;
  assign n39052 = ~pi0299 & ~pi1153;
  assign n39053 = ~n10810 & ~n39052;
  assign n39054 = ~n38745 & n39053;
  assign n39055 = pi0207 & ~n39054;
  assign n39056 = ~pi0207 & n39048;
  assign n39057 = pi0208 & ~n39055;
  assign n39058 = ~n39056 & n39057;
  assign n39059 = ~n39051 & ~n39058;
  assign n39060 = ~pi0211 & n39059;
  assign n39061 = pi0211 & n39043;
  assign n39062 = ~n39060 & ~n39061;
  assign n39063 = n38608 & ~n39062;
  assign n39064 = ~n39044 & ~n39063;
  assign n39065 = ~pi0219 & ~n39064;
  assign n39066 = ~n38499 & ~n38608;
  assign n39067 = n39029 & n39066;
  assign n39068 = n39031 & ~n39067;
  assign n39069 = ~n39065 & n39068;
  assign n39070 = n38888 & ~n39069;
  assign n39071 = ~n39020 & ~n39070;
  assign n39072 = ~pi0213 & n39071;
  assign n39073 = ~pi1152 & ~po1038;
  assign n39074 = n38413 & ~n39029;
  assign n39075 = ~pi0299 & ~n38937;
  assign n39076 = ~pi1154 & ~n39075;
  assign n39077 = ~n38765 & n39076;
  assign n39078 = ~n38731 & n39047;
  assign n39079 = ~n39077 & ~n39078;
  assign n39080 = pi0207 & n39079;
  assign n39081 = n38722 & ~n39080;
  assign n39082 = ~pi0207 & n39079;
  assign n39083 = ~n38765 & n39053;
  assign n39084 = pi0207 & ~n39083;
  assign n39085 = pi0208 & ~n39084;
  assign n39086 = ~n39082 & n39085;
  assign n39087 = ~n39081 & ~n39086;
  assign n39088 = ~pi0211 & n39087;
  assign n39089 = pi0211 & n39059;
  assign n39090 = n10843 & ~n39088;
  assign n39091 = ~n39089 & n39090;
  assign n39092 = ~pi0211 & ~n38787;
  assign n39093 = n39029 & n39092;
  assign n39094 = pi0211 & n39087;
  assign n39095 = ~n38423 & ~n39093;
  assign n39096 = ~n39094 & n39095;
  assign n39097 = ~n39091 & ~n39096;
  assign n39098 = ~pi0219 & ~n39097;
  assign n39099 = pi0211 & n39029;
  assign n39100 = n38970 & ~n39099;
  assign n39101 = ~n39060 & n39100;
  assign n39102 = ~n39074 & ~n39101;
  assign n39103 = ~n39098 & n39102;
  assign n39104 = n39073 & ~n39103;
  assign n39105 = ~n38414 & n38966;
  assign n39106 = ~n38413 & n39007;
  assign n39107 = ~n39105 & ~n39106;
  assign n39108 = pi0219 & ~n39107;
  assign n39109 = ~pi0212 & n39013;
  assign n39110 = pi0211 & ~n39006;
  assign n39111 = ~pi0199 & ~pi1154;
  assign n39112 = ~pi0200 & n39111;
  assign n39113 = n38674 & n39112;
  assign n39114 = n38722 & ~n38943;
  assign n39115 = ~n38952 & ~n39114;
  assign n39116 = ~n38765 & ~n39113;
  assign n39117 = ~n39115 & n39116;
  assign n39118 = ~pi0211 & n39117;
  assign n39119 = n10843 & ~n39118;
  assign n39120 = ~n39110 & n39119;
  assign n39121 = ~pi0208 & ~n38787;
  assign n39122 = ~n38995 & n39121;
  assign n39123 = pi0299 & ~pi1156;
  assign n39124 = n38998 & ~n39123;
  assign n39125 = ~n38787 & n38960;
  assign n39126 = ~pi0207 & ~n39125;
  assign n39127 = pi0208 & ~n39124;
  assign n39128 = ~n39126 & n39127;
  assign n39129 = ~pi0211 & ~n39122;
  assign n39130 = ~n39128 & n39129;
  assign n39131 = pi0211 & n39117;
  assign n39132 = ~n38423 & ~n39130;
  assign n39133 = ~n39131 & n39132;
  assign n39134 = ~pi0219 & ~n39109;
  assign n39135 = ~n39133 & n39134;
  assign n39136 = ~n39120 & n39135;
  assign n39137 = ~n39108 & ~n39136;
  assign n39138 = pi1152 & ~po1038;
  assign n39139 = ~n39137 & n39138;
  assign n39140 = ~n39104 & ~n39139;
  assign n39141 = pi0213 & ~n39140;
  assign n39142 = ~pi0209 & ~n39141;
  assign n39143 = ~n39072 & n39142;
  assign n39144 = ~n38935 & ~n39143;
  assign n39145 = pi0219 & ~n38495;
  assign n39146 = pi0212 & ~n38491;
  assign n39147 = pi0214 & ~n38485;
  assign n39148 = ~pi0212 & n39147;
  assign n39149 = ~pi0219 & ~n39148;
  assign n39150 = ~n39146 & n39149;
  assign n39151 = pi0213 & ~n39145;
  assign n39152 = n38416 & n39151;
  assign n39153 = ~n39150 & n39152;
  assign n39154 = ~n39144 & ~n39153;
  assign n39155 = pi0230 & ~n39154;
  assign n39156 = ~pi0230 & pi0234;
  assign po0391 = n39155 | n39156;
  assign n39158 = pi0219 & ~n38487;
  assign n39159 = pi0219 & ~n38608;
  assign n39160 = ~pi0212 & n38481;
  assign n39161 = ~pi0214 & ~n38480;
  assign n39162 = ~n39147 & ~n39161;
  assign n39163 = pi0212 & ~n39162;
  assign n39164 = ~pi0219 & ~n39163;
  assign n39165 = ~n39160 & n39164;
  assign n39166 = ~n39158 & ~n39159;
  assign n39167 = po1038 & n39166;
  assign n39168 = ~n39165 & n39167;
  assign n39169 = pi0208 & pi1157;
  assign n39170 = ~n38650 & ~n38766;
  assign n39171 = pi0207 & ~n39170;
  assign n39172 = ~pi0207 & ~n38727;
  assign n39173 = ~n39171 & ~n39172;
  assign n39174 = n39169 & ~n39173;
  assign n39175 = ~pi0207 & n38734;
  assign n39176 = ~n39171 & ~n39175;
  assign n39177 = pi0208 & ~n39176;
  assign n39178 = ~n38735 & ~n39177;
  assign n39179 = ~pi1157 & ~n39178;
  assign n39180 = ~n38730 & ~n39174;
  assign n39181 = ~n39179 & n39180;
  assign n39182 = pi0211 & ~n39181;
  assign n39183 = ~pi1156 & n38577;
  assign n39184 = ~n38698 & ~n39183;
  assign n39185 = pi0207 & ~n39184;
  assign n39186 = ~n38658 & ~n38671;
  assign n39187 = ~pi0207 & ~n39186;
  assign n39188 = ~n39185 & ~n39187;
  assign n39189 = n39169 & ~n39188;
  assign n39190 = ~pi0207 & n38536;
  assign n39191 = ~n39185 & ~n39190;
  assign n39192 = pi0208 & ~n39191;
  assign n39193 = ~n38786 & ~n39192;
  assign n39194 = ~pi1157 & ~n39193;
  assign n39195 = ~n38789 & ~n39189;
  assign n39196 = ~n39194 & n39195;
  assign n39197 = ~pi0211 & ~n39196;
  assign n39198 = n10843 & ~n39182;
  assign n39199 = ~n39197 & n39198;
  assign n39200 = n10487 & ~n38650;
  assign n39201 = ~n39183 & n39200;
  assign n39202 = ~pi0207 & ~n38643;
  assign n39203 = ~n39201 & ~n39202;
  assign n39204 = ~n38645 & n39203;
  assign n39205 = ~pi1157 & ~n39204;
  assign n39206 = ~pi0207 & n38659;
  assign n39207 = ~n39201 & ~n39206;
  assign n39208 = ~n38661 & n39207;
  assign n39209 = pi1157 & ~n39208;
  assign n39210 = ~n39205 & ~n39209;
  assign n39211 = n38413 & ~n39210;
  assign n39212 = pi0211 & ~n39196;
  assign n39213 = ~pi0207 & n38672;
  assign n39214 = pi0208 & ~n39213;
  assign n39215 = ~n38698 & n38889;
  assign n39216 = n39214 & ~n39215;
  assign n39217 = ~n38676 & ~n39216;
  assign n39218 = pi1157 & n39217;
  assign n39219 = ~pi0211 & ~n39205;
  assign n39220 = ~n39218 & n39219;
  assign n39221 = n38608 & ~n39220;
  assign n39222 = ~n39212 & n39221;
  assign n39223 = ~n39211 & ~n39222;
  assign n39224 = ~n39199 & n39223;
  assign n39225 = ~pi0219 & ~n39224;
  assign n39226 = ~pi0211 & n39181;
  assign n39227 = pi0211 & ~n39210;
  assign n39228 = ~n38423 & ~n39227;
  assign n39229 = ~n39226 & n39228;
  assign n39230 = n38423 & n39210;
  assign n39231 = pi0219 & ~n39230;
  assign n39232 = ~n39229 & n39231;
  assign n39233 = pi0209 & ~n39232;
  assign n39234 = ~n39225 & n39233;
  assign n39235 = ~n38691 & n38722;
  assign n39236 = ~pi0207 & n38691;
  assign n39237 = pi0208 & ~n39080;
  assign n39238 = ~n39236 & n39237;
  assign n39239 = ~n39235 & ~n39238;
  assign n39240 = pi0211 & ~n39239;
  assign n39241 = n10487 & ~n39024;
  assign n39242 = ~n38573 & ~n38825;
  assign n39243 = ~n10487 & ~n39242;
  assign n39244 = ~n39241 & ~n39243;
  assign n39245 = ~n38787 & ~n39244;
  assign n39246 = ~pi0211 & ~n39245;
  assign n39247 = n10843 & ~n39240;
  assign n39248 = ~n39246 & n39247;
  assign n39249 = n38413 & ~n39244;
  assign n39250 = n38675 & ~n38805;
  assign n39251 = n38674 & n38763;
  assign n39252 = ~n39047 & ~n39076;
  assign n39253 = pi0207 & n39252;
  assign n39254 = pi0208 & ~n39251;
  assign n39255 = ~n39253 & n39254;
  assign n39256 = ~n39250 & ~n39255;
  assign n39257 = pi1157 & ~n39256;
  assign n39258 = ~pi1157 & n39244;
  assign n39259 = ~pi0211 & ~n39257;
  assign n39260 = ~n39258 & n39259;
  assign n39261 = pi0211 & n39245;
  assign n39262 = ~n39260 & ~n39261;
  assign n39263 = n38608 & ~n39262;
  assign n39264 = ~n39248 & ~n39249;
  assign n39265 = ~n39263 & n39264;
  assign n39266 = ~pi0219 & ~n39265;
  assign n39267 = ~pi0211 & n39239;
  assign n39268 = pi0211 & ~n39244;
  assign n39269 = ~n38423 & ~n39268;
  assign n39270 = ~n39267 & n39269;
  assign n39271 = n38423 & n39244;
  assign n39272 = pi0219 & ~n39271;
  assign n39273 = ~n39270 & n39272;
  assign n39274 = ~pi0209 & ~n39273;
  assign n39275 = ~n39266 & n39274;
  assign n39276 = ~n39234 & ~n39275;
  assign n39277 = ~po1038 & ~n39276;
  assign n39278 = pi0213 & ~n39168;
  assign n39279 = ~n39277 & n39278;
  assign n39280 = pi0219 & ~n38497;
  assign n39281 = po1038 & ~n39280;
  assign n39282 = ~n38489 & n38608;
  assign n39283 = n10843 & ~n38883;
  assign n39284 = ~pi0219 & ~n39282;
  assign n39285 = ~n39283 & n39284;
  assign n39286 = ~n39159 & n39281;
  assign n39287 = ~n39285 & n39286;
  assign n39288 = pi1157 & ~n39217;
  assign n39289 = pi0299 & ~pi1157;
  assign n39290 = ~n39194 & ~n39289;
  assign n39291 = ~n39288 & n39290;
  assign n39292 = ~n38769 & ~n39291;
  assign n39293 = ~pi0211 & ~n39292;
  assign n39294 = n39228 & ~n39293;
  assign n39295 = n39231 & ~n39294;
  assign n39296 = ~n38578 & ~n38767;
  assign n39297 = ~n38650 & ~n39296;
  assign n39298 = pi0207 & ~n39297;
  assign n39299 = pi1154 & ~n38535;
  assign n39300 = ~n38642 & ~n39299;
  assign n39301 = ~pi0207 & ~n38732;
  assign n39302 = ~n39300 & n39301;
  assign n39303 = ~n39298 & ~n39302;
  assign n39304 = pi0208 & ~n39303;
  assign n39305 = ~n38757 & ~n39304;
  assign n39306 = ~pi1157 & ~n39305;
  assign n39307 = n38746 & ~n39217;
  assign n39308 = ~n39306 & ~n39307;
  assign n39309 = ~pi0211 & ~n39308;
  assign n39310 = pi0211 & n39292;
  assign n39311 = n10843 & ~n39309;
  assign n39312 = ~n39310 & n39311;
  assign n39313 = pi0211 & n39308;
  assign n39314 = ~n39226 & ~n39313;
  assign n39315 = n38608 & ~n39314;
  assign n39316 = ~n39211 & ~n39315;
  assign n39317 = ~n39312 & n39316;
  assign n39318 = ~pi0219 & ~n39317;
  assign n39319 = ~n39295 & ~n39318;
  assign n39320 = pi0209 & ~n39319;
  assign n39321 = ~n38764 & ~n38975;
  assign n39322 = ~pi0208 & ~n39321;
  assign n39323 = ~pi0207 & ~n38763;
  assign n39324 = ~n39035 & ~n39323;
  assign n39325 = pi0208 & ~n39324;
  assign n39326 = ~n39322 & ~n39325;
  assign n39327 = ~pi0211 & n39326;
  assign n39328 = n39269 & ~n39327;
  assign n39329 = n39272 & ~n39328;
  assign n39330 = ~n38753 & ~n38836;
  assign n39331 = ~pi0208 & ~n39330;
  assign n39332 = ~pi0207 & ~n38752;
  assign n39333 = ~n39049 & ~n39332;
  assign n39334 = pi0208 & ~n39333;
  assign n39335 = ~n39331 & ~n39334;
  assign n39336 = pi0211 & n39335;
  assign n39337 = ~n39267 & ~n39336;
  assign n39338 = ~n38423 & ~n39337;
  assign n39339 = ~pi0211 & ~n39335;
  assign n39340 = pi0211 & ~n39326;
  assign n39341 = n10843 & ~n39340;
  assign n39342 = ~n39339 & n39341;
  assign n39343 = ~n39249 & ~n39342;
  assign n39344 = ~n39338 & n39343;
  assign n39345 = ~pi0219 & ~n39344;
  assign n39346 = ~n39329 & ~n39345;
  assign n39347 = ~pi0209 & ~n39346;
  assign n39348 = ~po1038 & ~n39347;
  assign n39349 = ~n39320 & n39348;
  assign n39350 = ~pi0213 & ~n39287;
  assign n39351 = ~n39349 & n39350;
  assign n39352 = ~n39279 & ~n39351;
  assign n39353 = pi0230 & ~n39352;
  assign n39354 = ~pi0230 & ~pi0235;
  assign po0392 = ~n39353 & ~n39354;
  assign n39356 = ~pi0100 & n38198;
  assign n39357 = n38397 & ~n39356;
  assign n39358 = ~n6132 & ~n39357;
  assign n39359 = ~pi0075 & ~n39358;
  assign n39360 = ~n7302 & ~n39359;
  assign n39361 = ~pi0092 & ~n39360;
  assign n39362 = n13654 & ~n39361;
  assign n39363 = ~pi0074 & ~n39362;
  assign n39364 = n6131 & ~n39363;
  assign n39365 = ~pi0056 & ~n39364;
  assign n39366 = ~n6127 & ~n39365;
  assign n39367 = ~pi0062 & ~n39366;
  assign po0393 = n13662 & ~n39367;
  assign n39369 = pi0211 & pi1157;
  assign n39370 = ~pi0211 & pi1158;
  assign n39371 = ~n39369 & ~n39370;
  assign n39372 = n38421 & ~n39371;
  assign n39373 = n39164 & ~n39372;
  assign n39374 = ~pi0219 & po1038;
  assign n39375 = n38421 & n38483;
  assign n39376 = po1038 & n39375;
  assign n39377 = ~n39374 & ~n39376;
  assign n39378 = pi0214 & n38495;
  assign n39379 = pi1155 & n38744;
  assign n39380 = ~n39378 & ~n39379;
  assign n39381 = pi0212 & ~n39380;
  assign n39382 = po1038 & n39381;
  assign n39383 = n39377 & ~n39382;
  assign n39384 = ~n39373 & ~n39383;
  assign n39385 = ~pi0213 & ~n39384;
  assign n39386 = n38508 & ~n39373;
  assign n39387 = pi0199 & pi1143;
  assign n39388 = ~pi0200 & ~n39387;
  assign n39389 = ~n38434 & n39388;
  assign n39390 = ~n38437 & n39026;
  assign n39391 = ~n39389 & n39390;
  assign n39392 = pi0200 & ~n38434;
  assign n39393 = ~pi0199 & pi1145;
  assign n39394 = n39388 & ~n39393;
  assign n39395 = n38826 & ~n39392;
  assign n39396 = ~n39394 & n39395;
  assign n39397 = ~n39391 & ~n39396;
  assign n39398 = ~pi0299 & ~n39397;
  assign n39399 = n38421 & n38787;
  assign n39400 = pi0214 & ~n38514;
  assign n39401 = ~pi0214 & ~n38510;
  assign n39402 = pi0212 & ~n39400;
  assign n39403 = ~n39401 & n39402;
  assign n39404 = ~n39399 & ~n39403;
  assign n39405 = n38519 & ~n39404;
  assign n39406 = ~n39398 & ~n39405;
  assign n39407 = ~n39386 & n39406;
  assign n39408 = ~po1038 & ~n39407;
  assign n39409 = n39385 & ~n39408;
  assign n39410 = pi0219 & ~n38425;
  assign n39411 = n10843 & n38420;
  assign n39412 = ~pi0211 & pi1145;
  assign n39413 = pi0211 & pi1144;
  assign n39414 = ~n39412 & ~n39413;
  assign n39415 = ~n10843 & n39414;
  assign n39416 = ~n38413 & ~n39411;
  assign n39417 = ~n39415 & n39416;
  assign n39418 = ~pi0219 & ~n39417;
  assign n39419 = n38416 & ~n39410;
  assign n39420 = ~n39418 & n39419;
  assign n39421 = n38508 & n39417;
  assign n39422 = pi0299 & n38970;
  assign n39423 = n38425 & n39422;
  assign n39424 = ~n39398 & ~n39423;
  assign n39425 = ~n39421 & n39424;
  assign n39426 = ~po1038 & ~n39425;
  assign n39427 = ~n39420 & ~n39426;
  assign n39428 = pi0213 & n39427;
  assign n39429 = pi0209 & ~n39409;
  assign n39430 = ~n39428 & n39429;
  assign n39431 = n38449 & n38568;
  assign n39432 = pi1158 & n38955;
  assign n39433 = ~pi0199 & ~pi1158;
  assign n39434 = pi1156 & ~n39433;
  assign n39435 = ~n39432 & ~n39434;
  assign n39436 = n39431 & ~n39435;
  assign n39437 = pi0207 & n38651;
  assign n39438 = pi0208 & ~n39202;
  assign n39439 = ~n39437 & n39438;
  assign n39440 = ~n39436 & ~n39439;
  assign n39441 = ~pi1157 & ~n39440;
  assign n39442 = pi1156 & n38699;
  assign n39443 = ~pi0200 & ~pi1158;
  assign n39444 = ~pi0199 & ~n39443;
  assign n39445 = ~n39442 & ~n39444;
  assign n39446 = n38441 & ~n39445;
  assign n39447 = ~pi0208 & n39446;
  assign n39448 = pi0208 & ~n39206;
  assign n39449 = ~n39437 & n39448;
  assign n39450 = ~n39447 & ~n39449;
  assign n39451 = pi1157 & ~n39450;
  assign n39452 = ~n39441 & ~n39451;
  assign n39453 = ~n38414 & n39452;
  assign n39454 = ~pi0200 & pi0207;
  assign n39455 = ~n39435 & n39454;
  assign n39456 = ~pi1157 & ~n39455;
  assign n39457 = pi1156 & ~n38985;
  assign n39458 = ~pi1158 & ~n38641;
  assign n39459 = n39457 & ~n39458;
  assign n39460 = ~n39444 & ~n39459;
  assign n39461 = n38441 & ~n39460;
  assign n39462 = ~pi0208 & ~n39456;
  assign n39463 = n39461 & n39462;
  assign n39464 = ~pi0208 & ~n39463;
  assign n39465 = ~n38543 & n39464;
  assign n39466 = ~pi0299 & ~n38536;
  assign n39467 = ~pi0200 & pi1157;
  assign n39468 = ~pi0199 & n39467;
  assign n39469 = n39466 & ~n39468;
  assign n39470 = ~pi0207 & ~n38528;
  assign n39471 = ~n39469 & n39470;
  assign n39472 = pi0207 & ~n38601;
  assign n39473 = pi0208 & ~n39471;
  assign n39474 = ~n39472 & n39473;
  assign n39475 = ~n39465 & ~n39474;
  assign n39476 = n38414 & ~n39475;
  assign n39477 = ~n39453 & ~n39476;
  assign n39478 = pi0219 & ~n39477;
  assign n39479 = ~pi0214 & n39452;
  assign n39480 = ~pi0212 & ~n39479;
  assign n39481 = pi0299 & ~pi1145;
  assign n39482 = ~pi0207 & ~n39481;
  assign n39483 = ~n39469 & n39482;
  assign n39484 = pi0299 & pi1145;
  assign n39485 = n38578 & ~n39484;
  assign n39486 = ~n38702 & ~n39481;
  assign n39487 = pi1154 & ~n39486;
  assign n39488 = ~pi1156 & ~n39485;
  assign n39489 = ~n39487 & n39488;
  assign n39490 = n38593 & ~n39484;
  assign n39491 = ~n38596 & ~n39481;
  assign n39492 = ~pi1154 & ~n39491;
  assign n39493 = pi1156 & ~n39490;
  assign n39494 = ~n39492 & n39493;
  assign n39495 = ~n39489 & ~n39494;
  assign n39496 = pi0207 & ~n39495;
  assign n39497 = pi0208 & ~n39483;
  assign n39498 = ~n39496 & n39497;
  assign n39499 = n38641 & ~n38725;
  assign n39500 = pi1157 & ~n39432;
  assign n39501 = ~n39499 & n39500;
  assign n39502 = pi0207 & ~n39501;
  assign n39503 = ~pi0299 & n39442;
  assign n39504 = ~pi1157 & ~n39432;
  assign n39505 = ~n39503 & n39504;
  assign n39506 = n39502 & ~n39505;
  assign n39507 = ~pi0208 & ~n39484;
  assign n39508 = ~n39506 & n39507;
  assign n39509 = ~n39498 & ~n39508;
  assign n39510 = ~pi0211 & ~n39509;
  assign n39511 = ~n38612 & n39464;
  assign n39512 = ~pi0207 & ~n38610;
  assign n39513 = ~n39469 & n39512;
  assign n39514 = pi0207 & ~n38630;
  assign n39515 = pi0208 & ~n39513;
  assign n39516 = ~n39514 & n39515;
  assign n39517 = ~n39511 & ~n39516;
  assign n39518 = pi0211 & ~n39517;
  assign n39519 = ~n39510 & ~n39518;
  assign n39520 = pi0214 & ~n39519;
  assign n39521 = n39480 & ~n39520;
  assign n39522 = ~pi0211 & n39517;
  assign n39523 = pi0211 & n39475;
  assign n39524 = pi0214 & ~n39522;
  assign n39525 = ~n39523 & n39524;
  assign n39526 = ~pi0214 & ~n39519;
  assign n39527 = pi0212 & ~n39525;
  assign n39528 = ~n39526 & n39527;
  assign n39529 = ~pi0219 & ~n39521;
  assign n39530 = ~n39528 & n39529;
  assign n39531 = ~po1038 & ~n39478;
  assign n39532 = ~n39530 & n39531;
  assign n39533 = pi0213 & ~n39420;
  assign n39534 = ~n39532 & n39533;
  assign n39535 = ~n38853 & ~n39187;
  assign n39536 = n39169 & ~n39535;
  assign n39537 = ~n38787 & ~n39446;
  assign n39538 = n38542 & ~n39537;
  assign n39539 = n39121 & ~n39455;
  assign n39540 = pi0208 & ~n39190;
  assign n39541 = ~n38853 & n39540;
  assign n39542 = ~pi1157 & ~n39539;
  assign n39543 = ~n39541 & n39542;
  assign n39544 = ~n39536 & ~n39538;
  assign n39545 = ~n39543 & n39544;
  assign n39546 = n38421 & n39545;
  assign n39547 = pi0207 & ~n38860;
  assign n39548 = ~n39172 & ~n39547;
  assign n39549 = n39169 & ~n39548;
  assign n39550 = ~n38510 & ~n39461;
  assign n39551 = n38542 & ~n39550;
  assign n39552 = ~n39175 & ~n39547;
  assign n39553 = pi0208 & ~n39552;
  assign n39554 = ~pi0208 & n38510;
  assign n39555 = ~n39436 & ~n39554;
  assign n39556 = ~n39553 & n39555;
  assign n39557 = ~pi1157 & ~n39556;
  assign n39558 = ~n39549 & ~n39551;
  assign n39559 = ~n39557 & n39558;
  assign n39560 = ~pi0214 & ~n39559;
  assign n39561 = ~pi0207 & ~n38672;
  assign n39562 = ~n38745 & n39561;
  assign n39563 = pi1157 & ~n39562;
  assign n39564 = ~pi1157 & ~n39436;
  assign n39565 = ~n39302 & n39564;
  assign n39566 = ~n39563 & ~n39565;
  assign n39567 = pi0208 & ~n38837;
  assign n39568 = ~n39566 & n39567;
  assign n39569 = n39461 & ~n39564;
  assign n39570 = ~pi0208 & ~n38514;
  assign n39571 = ~n39569 & n39570;
  assign n39572 = pi0214 & ~n39571;
  assign n39573 = ~n39568 & n39572;
  assign n39574 = pi0212 & ~n39573;
  assign n39575 = ~n39560 & n39574;
  assign n39576 = ~n39546 & ~n39575;
  assign n39577 = ~pi0211 & ~n39576;
  assign n39578 = ~n39453 & ~n39577;
  assign n39579 = pi0219 & ~n39578;
  assign n39580 = ~pi0299 & n39445;
  assign n39581 = n38675 & ~n39580;
  assign n39582 = ~n38890 & n39214;
  assign n39583 = ~n39581 & ~n39582;
  assign n39584 = pi1157 & ~n39583;
  assign n39585 = ~n39441 & ~n39584;
  assign n39586 = pi0211 & n39585;
  assign n39587 = n38441 & n39442;
  assign n39588 = ~pi0299 & ~n39039;
  assign n39589 = pi1158 & ~n39588;
  assign n39590 = ~pi0208 & ~n39587;
  assign n39591 = ~n39589 & n39590;
  assign n39592 = ~pi1158 & n38651;
  assign n39593 = pi1158 & n38768;
  assign n39594 = pi0207 & ~n39592;
  assign n39595 = ~n39593 & n39594;
  assign n39596 = pi0299 & ~pi1158;
  assign n39597 = ~pi0207 & ~n39596;
  assign n39598 = ~n39466 & n39597;
  assign n39599 = pi0208 & ~n39598;
  assign n39600 = ~n39595 & n39599;
  assign n39601 = ~pi1157 & ~n39591;
  assign n39602 = ~n39600 & n39601;
  assign n39603 = n39561 & ~n39596;
  assign n39604 = ~n39595 & ~n39603;
  assign n39605 = n39169 & ~n39604;
  assign n39606 = ~n39502 & ~n39589;
  assign n39607 = n38542 & ~n39606;
  assign n39608 = ~pi0211 & ~n39607;
  assign n39609 = ~n39602 & n39608;
  assign n39610 = ~n39605 & n39609;
  assign n39611 = ~n39586 & ~n39610;
  assign n39612 = pi0214 & ~n39611;
  assign n39613 = n39480 & ~n39612;
  assign n39614 = n38783 & ~n39545;
  assign n39615 = n10484 & ~n39559;
  assign n39616 = n38744 & ~n39585;
  assign n39617 = ~n39614 & ~n39615;
  assign n39618 = ~n39616 & n39617;
  assign n39619 = pi0212 & ~n39618;
  assign n39620 = ~pi0219 & ~n39619;
  assign n39621 = ~n39613 & n39620;
  assign n39622 = ~po1038 & ~n39579;
  assign n39623 = ~n39621 & n39622;
  assign n39624 = n39385 & ~n39623;
  assign n39625 = ~pi0209 & ~n39534;
  assign n39626 = ~n39624 & n39625;
  assign n39627 = ~n39430 & ~n39626;
  assign n39628 = pi0230 & ~n39627;
  assign n39629 = ~pi0230 & ~pi0237;
  assign po0394 = n39628 | n39629;
  assign n39631 = ~pi0211 & ~pi1153;
  assign n39632 = pi0219 & n39631;
  assign n39633 = n38416 & ~n39632;
  assign n39634 = ~n39285 & n39633;
  assign n39635 = ~pi1151 & ~po1038;
  assign n39636 = n10809 & n38826;
  assign n39637 = ~pi0299 & ~n39636;
  assign n39638 = ~n13061 & ~n39637;
  assign n39639 = n38826 & n38955;
  assign n39640 = ~pi0214 & ~n39639;
  assign n39641 = ~pi0212 & n39640;
  assign n39642 = n39638 & ~n39641;
  assign n39643 = pi1153 & n39642;
  assign n39644 = ~n38665 & ~n39643;
  assign n39645 = n38882 & ~n39637;
  assign n39646 = pi1153 & n39639;
  assign n39647 = ~n38514 & ~n39646;
  assign n39648 = ~pi0211 & ~n39647;
  assign n39649 = n10843 & ~n39645;
  assign n39650 = ~n39648 & n39649;
  assign n39651 = pi0299 & ~n38489;
  assign n39652 = ~n38423 & ~n39651;
  assign n39653 = ~n39646 & n39652;
  assign n39654 = ~n39650 & ~n39653;
  assign n39655 = ~pi0219 & ~n39654;
  assign n39656 = n39635 & ~n39644;
  assign n39657 = ~n39655 & n39656;
  assign n39658 = ~n10487 & n38568;
  assign n39659 = ~n38825 & n39658;
  assign n39660 = n38561 & n39026;
  assign n39661 = ~n39659 & ~n39660;
  assign n39662 = ~n38962 & ~n39661;
  assign n39663 = ~pi0214 & ~n39662;
  assign n39664 = ~pi0212 & ~n39663;
  assign n39665 = n38568 & ~n38958;
  assign n39666 = ~pi1153 & ~n38700;
  assign n39667 = ~n38682 & ~n39666;
  assign n39668 = pi1155 & ~n39667;
  assign n39669 = ~n39665 & ~n39668;
  assign n39670 = n38441 & ~n38561;
  assign n39671 = pi0208 & ~n39670;
  assign n39672 = ~n38722 & ~n39671;
  assign n39673 = ~n39669 & ~n39672;
  assign n39674 = ~n39660 & ~n39673;
  assign n39675 = ~pi0299 & ~n39674;
  assign n39676 = pi0214 & ~n39651;
  assign n39677 = ~n39675 & n39676;
  assign n39678 = n39664 & ~n39677;
  assign n39679 = ~n38514 & n38783;
  assign n39680 = ~n39662 & n39679;
  assign n39681 = n38744 & n39674;
  assign n39682 = ~pi0299 & ~n39454;
  assign n39683 = ~pi0208 & ~n39682;
  assign n39684 = pi0200 & n38674;
  assign n39685 = n39671 & ~n39684;
  assign n39686 = ~n39683 & ~n39685;
  assign n39687 = ~n38683 & ~n39686;
  assign n39688 = n10484 & ~n39687;
  assign n39689 = pi0212 & ~n39680;
  assign n39690 = ~n39688 & n39689;
  assign n39691 = ~n39681 & n39690;
  assign n39692 = ~pi0219 & ~n39691;
  assign n39693 = ~n39678 & n39692;
  assign n39694 = pi1151 & ~po1038;
  assign n39695 = ~pi0211 & ~n39686;
  assign n39696 = pi0211 & ~n39661;
  assign n39697 = ~n39695 & ~n39696;
  assign n39698 = ~n38683 & ~n39697;
  assign n39699 = n38413 & ~n39662;
  assign n39700 = n39698 & ~n39699;
  assign n39701 = pi0219 & ~n39700;
  assign n39702 = n39694 & ~n39701;
  assign n39703 = ~n39693 & n39702;
  assign n39704 = ~pi1152 & ~n39657;
  assign n39705 = ~n39703 & n39704;
  assign n39706 = ~n11445 & ~n39045;
  assign n39707 = pi0207 & ~n39706;
  assign n39708 = ~n38975 & ~n39707;
  assign n39709 = ~pi0208 & ~n39708;
  assign n39710 = pi0200 & pi0207;
  assign n39711 = ~pi0199 & ~n39710;
  assign n39712 = ~pi0299 & ~n39711;
  assign n39713 = pi0208 & ~n39712;
  assign n39714 = ~pi0207 & n10809;
  assign n39715 = ~pi0299 & ~n39714;
  assign n39716 = ~pi1153 & ~n39715;
  assign n39717 = n39713 & ~n39716;
  assign n39718 = ~n39709 & ~n39717;
  assign n39719 = pi0211 & ~n39718;
  assign n39720 = ~pi0207 & ~n38947;
  assign n39721 = ~n39039 & ~n39720;
  assign n39722 = pi0208 & ~n39721;
  assign n39723 = n38675 & ~n38947;
  assign n39724 = ~n39722 & ~n39723;
  assign n39725 = ~pi0211 & ~n38745;
  assign n39726 = ~n39724 & n39725;
  assign n39727 = ~n39719 & ~n39726;
  assign n39728 = n10843 & ~n39727;
  assign n39729 = pi0299 & n38489;
  assign n39730 = ~n38423 & ~n39724;
  assign n39731 = ~n39729 & n39730;
  assign n39732 = ~n39728 & ~n39731;
  assign n39733 = ~pi0219 & ~n39732;
  assign n39734 = ~n10487 & n38945;
  assign n39735 = ~n38826 & ~n39454;
  assign n39736 = n11384 & ~n39735;
  assign n39737 = ~n39734 & n39736;
  assign n39738 = ~pi0211 & n38512;
  assign n39739 = ~n38413 & n39738;
  assign n39740 = ~n39737 & ~n39739;
  assign n39741 = ~n38665 & ~n39740;
  assign n39742 = ~n39733 & ~n39741;
  assign n39743 = n39635 & ~n39742;
  assign n39744 = n38441 & n38561;
  assign n39745 = pi0208 & n38550;
  assign n39746 = ~n39714 & n39745;
  assign n39747 = ~n39744 & ~n39746;
  assign n39748 = ~pi0214 & n39747;
  assign n39749 = ~n39646 & n39748;
  assign n39750 = ~pi0212 & ~n39749;
  assign n39751 = ~pi0214 & n39750;
  assign n39752 = n38948 & ~n38986;
  assign n39753 = pi0208 & ~n39752;
  assign n39754 = n38675 & ~n38949;
  assign n39755 = ~n39753 & ~n39754;
  assign n39756 = ~pi0211 & ~n39755;
  assign n39757 = ~n38765 & n39756;
  assign n39758 = pi0211 & ~n39755;
  assign n39759 = ~n38745 & n39758;
  assign n39760 = ~n39757 & ~n39759;
  assign n39761 = ~n38423 & ~n39760;
  assign n39762 = ~n39645 & n39747;
  assign n39763 = ~n39726 & n39762;
  assign n39764 = n10843 & ~n39763;
  assign n39765 = ~pi0219 & ~n39751;
  assign n39766 = ~n39764 & n39765;
  assign n39767 = ~n39761 & n39766;
  assign n39768 = pi0219 & n39747;
  assign n39769 = ~n39643 & n39768;
  assign n39770 = n39694 & ~n39769;
  assign n39771 = ~n39767 & n39770;
  assign n39772 = pi1152 & ~n39771;
  assign n39773 = ~n39743 & n39772;
  assign n39774 = ~n39705 & ~n39773;
  assign n39775 = ~pi0209 & ~n39774;
  assign n39776 = n38641 & n39032;
  assign n39777 = n10487 & ~n39776;
  assign n39778 = ~n38957 & n39777;
  assign n39779 = ~n39243 & ~n39778;
  assign n39780 = ~pi0214 & ~n39779;
  assign n39781 = ~pi0212 & n39780;
  assign n39782 = pi0211 & n39779;
  assign n39783 = pi1153 & ~n38581;
  assign n39784 = ~n38957 & ~n39783;
  assign n39785 = pi0207 & ~n39784;
  assign n39786 = ~n39323 & ~n39785;
  assign n39787 = pi0208 & ~n39786;
  assign n39788 = ~n39322 & ~n39787;
  assign n39789 = ~pi0211 & ~n39788;
  assign n39790 = ~n39782 & ~n39789;
  assign n39791 = n38970 & n39790;
  assign n39792 = ~n38550 & n39084;
  assign n39793 = ~pi1154 & ~n39052;
  assign n39794 = ~n38581 & n39793;
  assign n39795 = pi0207 & ~n39794;
  assign n39796 = n39001 & n39795;
  assign n39797 = pi0208 & ~n39796;
  assign n39798 = ~n39792 & n39797;
  assign n39799 = ~n39236 & n39798;
  assign n39800 = ~n39235 & ~n39799;
  assign n39801 = ~pi0211 & ~n39800;
  assign n39802 = n39001 & ~n39776;
  assign n39803 = pi0207 & ~n39802;
  assign n39804 = ~n39332 & ~n39803;
  assign n39805 = pi0208 & ~n39804;
  assign n39806 = ~n39331 & ~n39805;
  assign n39807 = pi0211 & ~n39806;
  assign n39808 = n38421 & ~n39801;
  assign n39809 = ~n39807 & n39808;
  assign n39810 = n10484 & ~n39788;
  assign n39811 = n38744 & ~n39800;
  assign n39812 = n38783 & ~n39806;
  assign n39813 = pi0212 & ~n39810;
  assign n39814 = ~n39811 & n39813;
  assign n39815 = ~n39812 & n39814;
  assign n39816 = ~n39809 & ~n39815;
  assign n39817 = ~pi0219 & ~n39816;
  assign n39818 = ~po1038 & ~n39781;
  assign n39819 = ~n39791 & n39818;
  assign n39820 = ~n39817 & n39819;
  assign n39821 = pi0209 & ~n39820;
  assign n39822 = ~n39775 & ~n39821;
  assign n39823 = ~n39634 & ~n39822;
  assign n39824 = pi0213 & ~n39823;
  assign n39825 = ~pi0211 & n38608;
  assign n39826 = pi1153 & n39825;
  assign n39827 = n39374 & n39826;
  assign n39828 = ~pi1151 & ~n39827;
  assign n39829 = pi0219 & ~n39639;
  assign n39830 = ~po1038 & ~n39829;
  assign n39831 = ~n13061 & ~n39646;
  assign n39832 = pi0212 & ~n39640;
  assign n39833 = ~n39831 & n39832;
  assign n39834 = ~pi0219 & ~n39833;
  assign n39835 = n39640 & n39643;
  assign n39836 = n38421 & n39738;
  assign n39837 = ~n39639 & ~n39836;
  assign n39838 = n39834 & n39837;
  assign n39839 = ~n39835 & n39838;
  assign n39840 = n39643 & n39830;
  assign n39841 = ~n39839 & n39840;
  assign n39842 = n39828 & ~n39841;
  assign n39843 = n10486 & ~n39826;
  assign n39844 = n38416 & ~n39843;
  assign n39845 = pi1151 & ~n39844;
  assign n39846 = ~pi0214 & n39698;
  assign n39847 = ~n39662 & n39831;
  assign n39848 = pi0214 & ~n39847;
  assign n39849 = pi0212 & ~n39848;
  assign n39850 = ~n39846 & n39849;
  assign n39851 = ~pi0212 & ~n39700;
  assign n39852 = ~n39850 & ~n39851;
  assign n39853 = ~pi0219 & ~n39852;
  assign n39854 = ~pi0211 & pi0299;
  assign n39855 = ~n39646 & ~n39854;
  assign n39856 = ~n39662 & n39855;
  assign n39857 = ~n39699 & ~n39856;
  assign n39858 = pi0219 & ~n39857;
  assign n39859 = ~po1038 & ~n39858;
  assign n39860 = ~n39853 & n39859;
  assign n39861 = n39845 & ~n39860;
  assign n39862 = ~pi1152 & ~n39842;
  assign n39863 = ~n39861 & n39862;
  assign n39864 = ~n10485 & n38665;
  assign n39865 = po1038 & n39864;
  assign n39866 = ~n10843 & ~n39631;
  assign n39867 = ~n38527 & ~n39866;
  assign n39868 = n39865 & ~n39867;
  assign n39869 = ~n10486 & n38416;
  assign n39870 = pi1151 & ~n39869;
  assign n39871 = ~n39868 & n39870;
  assign n39872 = ~n39646 & n39747;
  assign n39873 = ~n39756 & n39872;
  assign n39874 = pi0214 & n39873;
  assign n39875 = ~n39749 & ~n39874;
  assign n39876 = ~pi0212 & ~n39875;
  assign n39877 = ~n39873 & ~n39876;
  assign n39878 = pi0219 & ~n39877;
  assign n39879 = ~po1038 & ~n39878;
  assign n39880 = pi1153 & ~n39637;
  assign n39881 = ~n39758 & ~n39880;
  assign n39882 = pi0214 & n39747;
  assign n39883 = n39881 & n39882;
  assign n39884 = n39750 & ~n39883;
  assign n39885 = pi0214 & n39755;
  assign n39886 = n39748 & n39881;
  assign n39887 = pi0212 & ~n39885;
  assign n39888 = ~n39886 & n39887;
  assign n39889 = ~pi0219 & ~n39884;
  assign n39890 = ~n39888 & n39889;
  assign n39891 = n39879 & ~n39890;
  assign n39892 = n39871 & ~n39891;
  assign n39893 = ~pi1151 & ~n39868;
  assign n39894 = pi0219 & ~n39737;
  assign n39895 = ~po1038 & ~n39894;
  assign n39896 = ~pi0211 & n39718;
  assign n39897 = n39730 & ~n39896;
  assign n39898 = ~n38608 & n39737;
  assign n39899 = pi0299 & n38527;
  assign n39900 = ~pi0219 & ~n39899;
  assign n39901 = ~n39898 & n39900;
  assign n39902 = ~n39897 & n39901;
  assign n39903 = n39895 & ~n39902;
  assign n39904 = n39893 & ~n39903;
  assign n39905 = pi1152 & ~n39904;
  assign n39906 = ~n39892 & n39905;
  assign n39907 = ~n39863 & ~n39906;
  assign n39908 = ~pi0209 & n39907;
  assign n39909 = ~pi0219 & n38608;
  assign n39910 = ~n39779 & ~n39909;
  assign n39911 = n39790 & n39909;
  assign n39912 = ~po1038 & ~n39910;
  assign n39913 = ~n39911 & n39912;
  assign n39914 = n39828 & ~n39913;
  assign n39915 = ~n39251 & n39797;
  assign n39916 = ~n39250 & ~n39915;
  assign n39917 = ~pi0211 & ~n39916;
  assign n39918 = ~n39782 & ~n39917;
  assign n39919 = ~n38413 & n39918;
  assign n39920 = ~n39781 & ~n39919;
  assign n39921 = pi0219 & ~n39920;
  assign n39922 = ~po1038 & ~n39921;
  assign n39923 = pi0214 & n39790;
  assign n39924 = ~n39780 & ~n39923;
  assign n39925 = ~pi0212 & ~n39924;
  assign n39926 = ~pi0214 & ~n39790;
  assign n39927 = pi0211 & ~n39916;
  assign n39928 = ~pi0211 & n39779;
  assign n39929 = ~n39927 & ~n39928;
  assign n39930 = pi0214 & ~n39929;
  assign n39931 = pi0212 & ~n39926;
  assign n39932 = ~n39930 & n39931;
  assign n39933 = ~n39925 & ~n39932;
  assign n39934 = ~pi0219 & ~n39933;
  assign n39935 = n39922 & ~n39934;
  assign n39936 = n39845 & ~n39935;
  assign n39937 = ~pi1152 & ~n39914;
  assign n39938 = ~n39936 & n39937;
  assign n39939 = ~n39789 & ~n39927;
  assign n39940 = ~pi0214 & ~n39939;
  assign n39941 = pi0214 & ~n39918;
  assign n39942 = ~n39940 & ~n39941;
  assign n39943 = pi0212 & ~n39942;
  assign n39944 = pi0214 & n39939;
  assign n39945 = ~pi0212 & ~n39780;
  assign n39946 = ~n39944 & n39945;
  assign n39947 = ~pi0219 & ~n39946;
  assign n39948 = ~n39943 & n39947;
  assign n39949 = pi0219 & ~n39779;
  assign n39950 = ~po1038 & ~n39949;
  assign n39951 = ~n39948 & n39950;
  assign n39952 = n39893 & ~n39951;
  assign n39953 = pi0214 & ~n39916;
  assign n39954 = ~n39940 & ~n39953;
  assign n39955 = pi0212 & ~n39954;
  assign n39956 = n39947 & ~n39955;
  assign n39957 = n39922 & ~n39956;
  assign n39958 = n39871 & ~n39957;
  assign n39959 = pi1152 & ~n39952;
  assign n39960 = ~n39958 & n39959;
  assign n39961 = pi0209 & ~n39938;
  assign n39962 = ~n39960 & n39961;
  assign n39963 = ~pi0213 & ~n39908;
  assign n39964 = ~n39962 & n39963;
  assign n39965 = ~n39824 & ~n39964;
  assign n39966 = pi0230 & ~n39965;
  assign n39967 = ~pi0230 & pi0238;
  assign po0395 = n39966 | n39967;
  assign n39969 = n38449 & ~n38651;
  assign n39970 = pi0212 & ~n39969;
  assign n39971 = ~po1038 & ~n39970;
  assign n39972 = ~pi0214 & n39969;
  assign n39973 = ~pi0212 & ~n39972;
  assign n39974 = ~pi0219 & n39973;
  assign n39975 = pi0299 & pi1158;
  assign n39976 = ~n38449 & n39975;
  assign n39977 = ~pi0208 & n39595;
  assign n39978 = ~n39976 & ~n39977;
  assign n39979 = ~pi0211 & ~n39978;
  assign n39980 = ~pi1157 & ~n39969;
  assign n39981 = pi0208 & pi0299;
  assign n39982 = pi1157 & ~n39981;
  assign n39983 = ~n38891 & n39982;
  assign n39984 = pi0211 & ~n39980;
  assign n39985 = ~n39983 & n39984;
  assign n39986 = ~n39979 & ~n39985;
  assign n39987 = pi0214 & ~n39986;
  assign n39988 = n39974 & ~n39987;
  assign n39989 = pi0219 & n39973;
  assign n39990 = pi0211 & ~n39969;
  assign n39991 = pi0214 & ~n39990;
  assign n39992 = ~n38855 & n39092;
  assign n39993 = n39991 & ~n39992;
  assign n39994 = n39989 & ~n39993;
  assign n39995 = ~pi0209 & n39971;
  assign n39996 = ~n39994 & n39995;
  assign n39997 = ~n39988 & n39996;
  assign n39998 = ~pi0219 & ~n39372;
  assign n39999 = ~n39377 & ~n39998;
  assign n40000 = n39447 & ~n39564;
  assign n40001 = ~pi0214 & n40000;
  assign n40002 = ~pi0212 & ~n40001;
  assign n40003 = ~pi0219 & n40002;
  assign n40004 = ~n39581 & n39982;
  assign n40005 = ~n39564 & ~n40004;
  assign n40006 = pi0211 & ~n40005;
  assign n40007 = pi0208 & ~n39975;
  assign n40008 = ~n38542 & ~n40007;
  assign n40009 = ~n39591 & n40008;
  assign n40010 = n39608 & ~n40009;
  assign n40011 = pi0214 & ~n40006;
  assign n40012 = ~n40010 & n40011;
  assign n40013 = n40003 & ~n40012;
  assign n40014 = pi0212 & ~n40000;
  assign n40015 = ~po1038 & ~n40014;
  assign n40016 = pi0219 & n40002;
  assign n40017 = pi0211 & ~n40000;
  assign n40018 = n39092 & ~n40000;
  assign n40019 = pi0214 & ~n40018;
  assign n40020 = ~n40017 & n40019;
  assign n40021 = n40016 & ~n40020;
  assign n40022 = pi0209 & n40015;
  assign n40023 = ~n40021 & n40022;
  assign n40024 = ~n40013 & n40023;
  assign n40025 = pi0213 & ~n39999;
  assign n40026 = ~n40024 & n40025;
  assign n40027 = ~n39997 & n40026;
  assign n40028 = po1038 & ~n39145;
  assign n40029 = n38421 & ~n39149;
  assign n40030 = n40028 & n40029;
  assign n40031 = pi0211 & ~n38510;
  assign n40032 = ~n39463 & n40031;
  assign n40033 = n40019 & ~n40032;
  assign n40034 = n40003 & ~n40033;
  assign n40035 = ~pi0211 & ~n38514;
  assign n40036 = ~n39463 & n40035;
  assign n40037 = pi0214 & ~n40017;
  assign n40038 = ~n40036 & n40037;
  assign n40039 = n40016 & ~n40038;
  assign n40040 = n40015 & ~n40034;
  assign n40041 = ~n40039 & n40040;
  assign n40042 = pi0209 & ~n40041;
  assign n40043 = ~n38514 & ~n38839;
  assign n40044 = n39991 & ~n40043;
  assign n40045 = n39989 & ~n40044;
  assign n40046 = ~n38861 & n40031;
  assign n40047 = pi0214 & ~n40046;
  assign n40048 = ~n39992 & n40047;
  assign n40049 = n39974 & ~n40048;
  assign n40050 = n39971 & ~n40049;
  assign n40051 = ~n40045 & n40050;
  assign n40052 = ~pi0209 & ~n40051;
  assign n40053 = ~n40042 & ~n40052;
  assign n40054 = ~pi0213 & ~n40030;
  assign n40055 = ~n40053 & n40054;
  assign n40056 = ~n40027 & ~n40055;
  assign n40057 = pi0230 & ~n40056;
  assign n40058 = ~pi0230 & ~pi0239;
  assign po0396 = ~n40057 & ~n40058;
  assign n40060 = ~po1038 & n39736;
  assign n40061 = ~n39830 & ~n40060;
  assign n40062 = ~pi0214 & ~n39736;
  assign n40063 = ~pi0212 & ~n40062;
  assign n40064 = n11384 & n38449;
  assign n40065 = ~pi0299 & ~n40064;
  assign n40066 = ~n39713 & n40065;
  assign n40067 = pi0214 & n40066;
  assign n40068 = n40063 & ~n40067;
  assign n40069 = ~pi0219 & ~n40068;
  assign n40070 = pi0211 & n39736;
  assign n40071 = ~pi0211 & ~n40066;
  assign n40072 = pi0214 & ~n40070;
  assign n40073 = ~n40071 & n40072;
  assign n40074 = pi0212 & ~n40073;
  assign n40075 = ~n40066 & n40074;
  assign n40076 = n40069 & ~n40075;
  assign n40077 = ~n40061 & ~n40076;
  assign n40078 = ~n39865 & ~n40077;
  assign n40079 = ~pi1147 & n40078;
  assign n40080 = ~pi0211 & po1038;
  assign n40081 = ~n39374 & ~n40080;
  assign n40082 = ~n38413 & ~n40081;
  assign n40083 = pi0299 & ~n38413;
  assign n40084 = ~po1038 & ~n38415;
  assign n40085 = n40083 & n40084;
  assign n40086 = n38550 & ~n38825;
  assign n40087 = ~po1038 & n40086;
  assign n40088 = ~n40085 & ~n40087;
  assign n40089 = ~n40082 & n40088;
  assign n40090 = pi1147 & n40089;
  assign n40091 = pi1149 & ~n40090;
  assign n40092 = ~n40079 & n40091;
  assign n40093 = pi0211 & n38421;
  assign n40094 = pi0212 & n38783;
  assign n40095 = ~n40093 & ~n40094;
  assign n40096 = n39374 & ~n40095;
  assign n40097 = ~n38826 & ~n39039;
  assign n40098 = ~n10487 & n38533;
  assign n40099 = ~n40097 & ~n40098;
  assign n40100 = n39715 & n40099;
  assign n40101 = pi0299 & n10484;
  assign n40102 = ~n40100 & ~n40101;
  assign n40103 = ~pi0212 & ~n40102;
  assign n40104 = ~pi0219 & ~n40103;
  assign n40105 = ~pi0299 & ~n40099;
  assign n40106 = pi0214 & ~n40105;
  assign n40107 = ~pi0214 & n40100;
  assign n40108 = ~pi0212 & ~n40107;
  assign n40109 = ~n40106 & n40108;
  assign n40110 = ~pi0211 & ~n40105;
  assign n40111 = ~n40100 & ~n40110;
  assign n40112 = pi0214 & ~n40111;
  assign n40113 = pi0212 & ~n40112;
  assign n40114 = ~pi0214 & ~n40105;
  assign n40115 = n40113 & ~n40114;
  assign n40116 = ~n40109 & ~n40115;
  assign n40117 = ~n13061 & ~n40100;
  assign n40118 = ~n40106 & n40117;
  assign n40119 = pi0212 & ~n40118;
  assign n40120 = n40116 & n40119;
  assign n40121 = n40104 & ~n40120;
  assign n40122 = pi0219 & ~n40100;
  assign n40123 = ~po1038 & ~n40122;
  assign n40124 = ~n40121 & n40123;
  assign n40125 = ~n40096 & ~n40124;
  assign n40126 = ~pi1147 & n40125;
  assign n40127 = ~po1038 & ~n39747;
  assign n40128 = pi0212 & ~n38744;
  assign n40129 = ~pi0219 & ~n40093;
  assign n40130 = ~n40128 & n40129;
  assign n40131 = n38416 & ~n40130;
  assign n40132 = n40085 & ~n40130;
  assign n40133 = ~n40127 & ~n40131;
  assign n40134 = ~n40132 & n40133;
  assign n40135 = pi1147 & n40134;
  assign n40136 = ~pi1149 & ~n40135;
  assign n40137 = ~n40126 & n40136;
  assign n40138 = ~n40092 & ~n40137;
  assign n40139 = pi1148 & ~n40138;
  assign n40140 = n16479 & n39636;
  assign n40141 = ~pi0219 & ~n16479;
  assign n40142 = n39825 & n40141;
  assign n40143 = ~n40140 & ~n40142;
  assign n40144 = ~pi1147 & n40143;
  assign n40145 = n10486 & ~n39825;
  assign n40146 = n38416 & ~n40145;
  assign n40147 = ~pi0211 & ~n39661;
  assign n40148 = pi0211 & ~n39686;
  assign n40149 = pi0214 & ~n40148;
  assign n40150 = ~n40147 & n40149;
  assign n40151 = n10843 & ~n40150;
  assign n40152 = ~pi0214 & n39661;
  assign n40153 = ~pi0212 & ~n40152;
  assign n40154 = pi0214 & n39697;
  assign n40155 = n40153 & ~n40154;
  assign n40156 = ~pi0219 & ~n40155;
  assign n40157 = pi0212 & ~n40150;
  assign n40158 = ~n39697 & n40157;
  assign n40159 = n40156 & ~n40158;
  assign n40160 = ~n40151 & n40159;
  assign n40161 = pi0212 & ~n39697;
  assign n40162 = pi0219 & ~n40161;
  assign n40163 = ~n40155 & n40162;
  assign n40164 = ~po1038 & ~n40163;
  assign n40165 = ~n40160 & n40164;
  assign n40166 = ~n40146 & ~n40165;
  assign n40167 = pi1147 & n40166;
  assign n40168 = pi1149 & ~n40144;
  assign n40169 = ~n40167 & n40168;
  assign n40170 = ~pi0212 & ~n40101;
  assign n40171 = n39747 & n40170;
  assign n40172 = n39747 & ~n39854;
  assign n40173 = ~n39748 & ~n40172;
  assign n40174 = ~pi0214 & n13061;
  assign n40175 = pi0212 & ~n40174;
  assign n40176 = ~n40173 & n40175;
  assign n40177 = ~n40171 & ~n40176;
  assign n40178 = ~pi0219 & ~n40177;
  assign n40179 = n38700 & ~n39710;
  assign n40180 = pi0208 & ~n40179;
  assign n40181 = ~pi0199 & ~n40180;
  assign n40182 = ~n39747 & ~n40181;
  assign n40183 = ~pi0299 & ~n40182;
  assign n40184 = ~pi0219 & n40183;
  assign n40185 = ~n40178 & ~n40184;
  assign n40186 = ~pi0211 & ~n40185;
  assign n40187 = ~n13061 & n39882;
  assign n40188 = ~pi0214 & n40172;
  assign n40189 = pi0212 & ~n40188;
  assign n40190 = ~n40187 & n40189;
  assign n40191 = ~pi0212 & n40173;
  assign n40192 = ~pi0219 & ~n40191;
  assign n40193 = ~n40190 & n40192;
  assign n40194 = pi0219 & ~n39854;
  assign n40195 = n40084 & ~n40194;
  assign n40196 = ~n40127 & ~n40195;
  assign n40197 = ~n40193 & ~n40196;
  assign n40198 = ~n40183 & n40197;
  assign n40199 = ~n40186 & n40198;
  assign n40200 = ~n39869 & ~n40199;
  assign n40201 = pi1147 & ~pi1149;
  assign n40202 = ~n40200 & n40201;
  assign n40203 = ~n40169 & ~n40202;
  assign n40204 = ~pi1148 & ~n40203;
  assign n40205 = ~n40139 & ~n40204;
  assign n40206 = pi0213 & ~n40205;
  assign n40207 = n10846 & n38665;
  assign n40208 = po1038 & n40207;
  assign n40209 = ~pi0211 & pi1146;
  assign n40210 = pi0211 & pi1145;
  assign n40211 = ~n40209 & ~n40210;
  assign n40212 = pi0214 & ~n40211;
  assign n40213 = pi0211 & pi1146;
  assign n40214 = ~pi0214 & n40213;
  assign n40215 = ~n40212 & ~n40214;
  assign n40216 = pi0212 & ~n40215;
  assign n40217 = n38421 & n40213;
  assign n40218 = ~n40216 & ~n40217;
  assign n40219 = ~n38970 & n40218;
  assign n40220 = po1038 & n39412;
  assign n40221 = ~n39374 & ~n40220;
  assign n40222 = ~n40219 & ~n40221;
  assign n40223 = pi1147 & ~n40208;
  assign n40224 = ~n40222 & n40223;
  assign n40225 = ~pi0211 & n39484;
  assign n40226 = pi0219 & ~n40225;
  assign n40227 = n40084 & ~n40226;
  assign n40228 = ~n40127 & ~n40227;
  assign n40229 = n38413 & ~n39747;
  assign n40230 = ~pi0219 & ~n40229;
  assign n40231 = pi0299 & ~n40211;
  assign n40232 = n39747 & ~n40231;
  assign n40233 = n10843 & ~n40232;
  assign n40234 = pi0299 & pi1146;
  assign n40235 = pi0211 & n40234;
  assign n40236 = ~n39854 & ~n40235;
  assign n40237 = n39747 & n40236;
  assign n40238 = n38608 & ~n40237;
  assign n40239 = n40230 & ~n40233;
  assign n40240 = ~n40238 & n40239;
  assign n40241 = ~n40228 & ~n40240;
  assign n40242 = n40224 & ~n40241;
  assign n40243 = ~po1038 & n40100;
  assign n40244 = ~pi1147 & ~n40222;
  assign n40245 = pi0219 & n40227;
  assign n40246 = pi0299 & ~n40218;
  assign n40247 = n36114 & n40246;
  assign n40248 = ~n40245 & ~n40247;
  assign n40249 = n40244 & n40248;
  assign n40250 = ~n40243 & n40249;
  assign n40251 = pi1148 & ~n40242;
  assign n40252 = ~n40250 & n40251;
  assign n40253 = n39412 & n39422;
  assign n40254 = ~n38665 & n40182;
  assign n40255 = ~pi1146 & n13061;
  assign n40256 = n38608 & ~n40255;
  assign n40257 = ~n40233 & ~n40256;
  assign n40258 = ~pi0219 & ~n40183;
  assign n40259 = ~n40257 & n40258;
  assign n40260 = ~n40253 & ~n40254;
  assign n40261 = ~n40259 & n40260;
  assign n40262 = ~po1038 & ~n40261;
  assign n40263 = n40224 & ~n40262;
  assign n40264 = ~pi1148 & ~n40249;
  assign n40265 = ~n40263 & n40264;
  assign n40266 = ~n40252 & ~n40265;
  assign n40267 = ~pi1149 & ~n40266;
  assign n40268 = pi0219 & n39661;
  assign n40269 = ~po1038 & ~n40268;
  assign n40270 = ~n40227 & ~n40269;
  assign n40271 = ~pi0299 & n39685;
  assign n40272 = ~n39431 & ~n40271;
  assign n40273 = ~n40234 & n40272;
  assign n40274 = pi0211 & ~n40273;
  assign n40275 = ~n39695 & ~n40274;
  assign n40276 = pi0214 & n40275;
  assign n40277 = n40153 & ~n40276;
  assign n40278 = pi0214 & ~n40231;
  assign n40279 = n40272 & n40278;
  assign n40280 = ~pi0214 & n40275;
  assign n40281 = pi0212 & ~n40279;
  assign n40282 = ~n40280 & n40281;
  assign n40283 = ~pi0219 & ~n40277;
  assign n40284 = ~n40282 & n40283;
  assign n40285 = ~n40270 & ~n40284;
  assign n40286 = n40224 & ~n40285;
  assign n40287 = ~n40140 & n40249;
  assign n40288 = ~pi1148 & ~n40287;
  assign n40289 = ~n40286 & n40288;
  assign n40290 = pi0219 & ~n40086;
  assign n40291 = ~po1038 & ~n40290;
  assign n40292 = pi0211 & ~n40086;
  assign n40293 = pi0214 & pi0299;
  assign n40294 = ~n40086 & ~n40293;
  assign n40295 = ~pi0212 & ~n40294;
  assign n40296 = ~n40292 & n40295;
  assign n40297 = ~pi0299 & ~n40086;
  assign n40298 = pi0212 & ~n40297;
  assign n40299 = pi0299 & n40128;
  assign n40300 = n40298 & ~n40299;
  assign n40301 = ~pi0219 & ~n40296;
  assign n40302 = ~n40300 & n40301;
  assign n40303 = n40291 & ~n40302;
  assign n40304 = n40224 & n40248;
  assign n40305 = ~n40303 & n40304;
  assign n40306 = ~n38414 & n39736;
  assign n40307 = ~n38413 & n40071;
  assign n40308 = pi0219 & ~n40306;
  assign n40309 = ~n40307 & n40308;
  assign n40310 = ~po1038 & ~n40309;
  assign n40311 = n11384 & n40310;
  assign n40312 = ~n40227 & ~n40311;
  assign n40313 = ~n39736 & ~n40235;
  assign n40314 = n40063 & ~n40313;
  assign n40315 = pi0212 & ~n40066;
  assign n40316 = ~n39736 & n40215;
  assign n40317 = n40315 & ~n40316;
  assign n40318 = ~pi0219 & ~n40314;
  assign n40319 = ~n40317 & n40318;
  assign n40320 = ~n40312 & ~n40319;
  assign n40321 = n40244 & ~n40320;
  assign n40322 = pi1148 & ~n40305;
  assign n40323 = ~n40321 & n40322;
  assign n40324 = ~n40289 & ~n40323;
  assign n40325 = pi1149 & ~n40324;
  assign n40326 = ~n40267 & ~n40325;
  assign n40327 = ~pi0213 & ~n40326;
  assign n40328 = pi0209 & ~n40327;
  assign n40329 = ~n40206 & n40328;
  assign n40330 = pi0200 & ~n39393;
  assign n40331 = pi0199 & pi1145;
  assign n40332 = ~pi0200 & ~n40331;
  assign n40333 = ~pi0199 & pi1146;
  assign n40334 = n40332 & ~n40333;
  assign n40335 = n38441 & ~n40330;
  assign n40336 = ~n40334 & n40335;
  assign n40337 = ~n38826 & ~n40336;
  assign n40338 = pi0200 & ~n40333;
  assign n40339 = ~pi0299 & ~n40338;
  assign n40340 = ~n40332 & n40339;
  assign n40341 = ~n10487 & ~n40340;
  assign n40342 = ~n40337 & ~n40341;
  assign n40343 = n38413 & n40342;
  assign n40344 = pi0219 & ~n40343;
  assign n40345 = ~n38413 & n40342;
  assign n40346 = ~n38414 & ~n40345;
  assign n40347 = n38699 & ~n40331;
  assign n40348 = n40339 & ~n40347;
  assign n40349 = ~pi0207 & n40348;
  assign n40350 = n40332 & n40349;
  assign n40351 = ~n40234 & ~n40336;
  assign n40352 = ~n40349 & n40351;
  assign n40353 = pi0208 & ~n40352;
  assign n40354 = ~n40350 & n40353;
  assign n40355 = n38449 & n40340;
  assign n40356 = ~n40354 & ~n40355;
  assign n40357 = ~pi0299 & ~n40356;
  assign n40358 = ~pi0211 & ~n39484;
  assign n40359 = ~n40357 & n40358;
  assign n40360 = ~n40346 & ~n40359;
  assign n40361 = n40344 & ~n40360;
  assign n40362 = ~n40235 & ~n40342;
  assign n40363 = ~pi0214 & ~n40342;
  assign n40364 = ~pi0212 & ~n40363;
  assign n40365 = ~n40362 & n40364;
  assign n40366 = ~pi0219 & ~n40365;
  assign n40367 = n40278 & ~n40357;
  assign n40368 = ~pi0214 & n40362;
  assign n40369 = pi0212 & ~n40368;
  assign n40370 = ~n40367 & n40369;
  assign n40371 = n40366 & ~n40370;
  assign n40372 = ~po1038 & ~n40361;
  assign n40373 = ~n40371 & n40372;
  assign n40374 = n40244 & ~n40373;
  assign n40375 = ~n10487 & ~n40348;
  assign n40376 = ~n40337 & ~n40375;
  assign n40377 = ~n38414 & n40376;
  assign n40378 = pi0219 & ~n40377;
  assign n40379 = n38449 & n40348;
  assign n40380 = ~n40353 & ~n40379;
  assign n40381 = ~pi0299 & n40380;
  assign n40382 = ~pi0211 & ~n40381;
  assign n40383 = ~n39481 & n40382;
  assign n40384 = ~n38413 & n40383;
  assign n40385 = n40378 & ~n40384;
  assign n40386 = ~n40376 & ~n40382;
  assign n40387 = ~pi0214 & ~n40376;
  assign n40388 = ~pi0212 & ~n40387;
  assign n40389 = ~n40386 & n40388;
  assign n40390 = pi0211 & ~n40381;
  assign n40391 = ~n39481 & n40390;
  assign n40392 = n40278 & n40380;
  assign n40393 = n10484 & ~n40381;
  assign n40394 = ~n40392 & ~n40393;
  assign n40395 = ~n40391 & ~n40394;
  assign n40396 = ~pi0214 & n40236;
  assign n40397 = n40380 & n40396;
  assign n40398 = pi0212 & ~n40397;
  assign n40399 = ~n40395 & n40398;
  assign n40400 = n40366 & ~n40389;
  assign n40401 = ~n40399 & n40400;
  assign n40402 = ~po1038 & ~n40385;
  assign n40403 = ~n40401 & n40402;
  assign n40404 = n40224 & ~n40403;
  assign n40405 = ~n40374 & ~n40404;
  assign n40406 = ~pi0213 & n40405;
  assign n40407 = pi1147 & ~n40131;
  assign n40408 = ~n38413 & n40382;
  assign n40409 = n40378 & ~n40408;
  assign n40410 = ~po1038 & ~n40409;
  assign n40411 = ~pi0299 & n40356;
  assign n40412 = pi0214 & ~n40411;
  assign n40413 = ~n40390 & ~n40412;
  assign n40414 = pi0212 & ~n40413;
  assign n40415 = ~pi0219 & ~n40376;
  assign n40416 = ~n40393 & n40415;
  assign n40417 = ~n40414 & n40416;
  assign n40418 = n40410 & ~n40417;
  assign n40419 = n40407 & ~n40418;
  assign n40420 = ~n40343 & n40417;
  assign n40421 = pi0219 & ~n40342;
  assign n40422 = pi0214 & n40386;
  assign n40423 = ~n40411 & ~n40422;
  assign n40424 = pi0212 & ~n40423;
  assign n40425 = ~pi0214 & n40342;
  assign n40426 = ~pi0212 & ~n40425;
  assign n40427 = ~n40412 & n40426;
  assign n40428 = ~n40424 & ~n40427;
  assign n40429 = ~pi0219 & ~n40428;
  assign n40430 = ~po1038 & ~n40421;
  assign n40431 = ~n40429 & n40430;
  assign n40432 = ~n40420 & n40431;
  assign n40433 = ~pi1147 & ~n40096;
  assign n40434 = ~n40432 & n40433;
  assign n40435 = ~pi1149 & ~n40419;
  assign n40436 = ~n40434 & n40435;
  assign n40437 = ~n40083 & n40415;
  assign n40438 = n40410 & ~n40437;
  assign n40439 = pi1147 & ~n40082;
  assign n40440 = ~n40438 & n40439;
  assign n40441 = ~pi1147 & ~n39865;
  assign n40442 = ~n40431 & n40441;
  assign n40443 = pi1149 & ~n40440;
  assign n40444 = ~n40442 & n40443;
  assign n40445 = pi1148 & ~n40444;
  assign n40446 = ~n40436 & n40445;
  assign n40447 = ~pi1147 & ~po1038;
  assign n40448 = n40342 & n40447;
  assign n40449 = pi0214 & ~n40376;
  assign n40450 = ~n40390 & n40449;
  assign n40451 = ~n40382 & n40387;
  assign n40452 = pi0212 & ~n40450;
  assign n40453 = ~n40451 & n40452;
  assign n40454 = ~pi0219 & ~n40389;
  assign n40455 = ~n40453 & n40454;
  assign n40456 = n40418 & ~n40455;
  assign n40457 = ~n39869 & ~n40456;
  assign n40458 = pi1147 & ~n40457;
  assign n40459 = ~n40448 & ~n40458;
  assign n40460 = ~pi1149 & ~n40459;
  assign n40461 = n40410 & ~n40455;
  assign n40462 = ~n40146 & ~n40461;
  assign n40463 = pi1147 & ~n40462;
  assign n40464 = ~pi1147 & n40207;
  assign n40465 = ~n40448 & ~n40464;
  assign n40466 = n16479 & n40207;
  assign n40467 = n40356 & n40466;
  assign n40468 = ~n40465 & ~n40467;
  assign n40469 = ~n40463 & ~n40468;
  assign n40470 = pi1149 & ~n40469;
  assign n40471 = ~pi1148 & ~n40470;
  assign n40472 = ~n40460 & n40471;
  assign n40473 = pi0213 & ~n40446;
  assign n40474 = ~n40472 & n40473;
  assign n40475 = ~pi0209 & ~n40406;
  assign n40476 = ~n40474 & n40475;
  assign n40477 = ~n40329 & ~n40476;
  assign n40478 = pi0230 & ~n40477;
  assign n40479 = ~pi0230 & ~pi0240;
  assign po0397 = ~n40478 & ~n40479;
  assign n40481 = pi0213 & ~n39907;
  assign n40482 = n39635 & n39646;
  assign n40483 = n38508 & n39825;
  assign n40484 = ~n39662 & ~n40483;
  assign n40485 = po1038 & ~n40207;
  assign n40486 = pi1151 & ~n40485;
  assign n40487 = ~n40484 & n40486;
  assign n40488 = ~n40482 & ~n40487;
  assign n40489 = ~pi1152 & ~n40488;
  assign n40490 = ~n39755 & n40207;
  assign n40491 = n39872 & ~n40490;
  assign n40492 = pi1152 & ~n40491;
  assign n40493 = ~po1038 & ~n40492;
  assign n40494 = n40486 & ~n40493;
  assign n40495 = pi1152 & n39635;
  assign n40496 = n39737 & n40495;
  assign n40497 = ~n40489 & ~n40496;
  assign n40498 = ~n40494 & n40497;
  assign n40499 = ~pi1150 & ~n40498;
  assign n40500 = pi1151 & ~n39865;
  assign n40501 = pi0219 & ~n39646;
  assign n40502 = ~po1038 & ~n40501;
  assign n40503 = ~n40127 & ~n40502;
  assign n40504 = n39750 & ~n39885;
  assign n40505 = ~pi0219 & ~n40504;
  assign n40506 = ~pi0214 & n39755;
  assign n40507 = pi0212 & ~n40506;
  assign n40508 = ~n39874 & n40507;
  assign n40509 = n40505 & ~n40508;
  assign n40510 = pi1152 & ~n40509;
  assign n40511 = ~pi0299 & ~n39687;
  assign n40512 = ~pi0214 & n39686;
  assign n40513 = pi0212 & ~n40512;
  assign n40514 = ~n40154 & n40513;
  assign n40515 = ~n39664 & ~n40514;
  assign n40516 = ~n40511 & ~n40515;
  assign n40517 = ~pi0219 & ~n40516;
  assign n40518 = ~pi1152 & ~n40268;
  assign n40519 = ~n40517 & n40518;
  assign n40520 = ~n40510 & ~n40519;
  assign n40521 = ~n40503 & ~n40520;
  assign n40522 = n40500 & ~n40521;
  assign n40523 = ~pi1151 & ~n40096;
  assign n40524 = ~pi0212 & ~n39637;
  assign n40525 = ~n39640 & n40524;
  assign n40526 = ~n39854 & n40525;
  assign n40527 = ~pi0219 & ~n40526;
  assign n40528 = pi0214 & ~n39638;
  assign n40529 = ~pi0211 & n39640;
  assign n40530 = pi0212 & ~n39637;
  assign n40531 = ~n40529 & n40530;
  assign n40532 = ~n40528 & n40531;
  assign n40533 = n40527 & ~n40532;
  assign n40534 = ~n39646 & n39834;
  assign n40535 = ~pi0299 & n40534;
  assign n40536 = ~n40533 & ~n40535;
  assign n40537 = n40502 & n40536;
  assign n40538 = ~pi1152 & ~n40537;
  assign n40539 = ~n39737 & ~n40536;
  assign n40540 = n39895 & ~n40539;
  assign n40541 = pi1152 & ~n40540;
  assign n40542 = ~n40538 & ~n40541;
  assign n40543 = n40523 & ~n40542;
  assign n40544 = pi1150 & ~n40543;
  assign n40545 = ~n40522 & n40544;
  assign n40546 = ~n40499 & ~n40545;
  assign n40547 = ~pi1149 & ~n40546;
  assign n40548 = pi1151 & ~n40146;
  assign n40549 = ~pi0214 & ~n39856;
  assign n40550 = n39849 & ~n40549;
  assign n40551 = ~pi0212 & ~n39857;
  assign n40552 = ~n40550 & ~n40551;
  assign n40553 = ~pi0219 & ~n40552;
  assign n40554 = ~pi1152 & n39859;
  assign n40555 = ~n40553 & n40554;
  assign n40556 = ~n38783 & ~n39755;
  assign n40557 = pi0212 & n39872;
  assign n40558 = ~n40556 & n40557;
  assign n40559 = ~n39876 & ~n40558;
  assign n40560 = ~pi0219 & ~n40559;
  assign n40561 = pi1152 & ~n40560;
  assign n40562 = n39879 & n40561;
  assign n40563 = n40548 & ~n40555;
  assign n40564 = ~n40562 & n40563;
  assign n40565 = ~pi1151 & ~n39869;
  assign n40566 = ~n40195 & ~n40502;
  assign n40567 = ~n40534 & ~n40566;
  assign n40568 = ~pi1152 & n40567;
  assign n40569 = ~n39895 & n40566;
  assign n40570 = ~n39737 & n39834;
  assign n40571 = pi1152 & ~n40569;
  assign n40572 = ~n40570 & n40571;
  assign n40573 = n40565 & ~n40568;
  assign n40574 = ~n40572 & n40573;
  assign n40575 = ~pi1150 & ~n40574;
  assign n40576 = ~n40564 & n40575;
  assign n40577 = ~pi1151 & ~n40131;
  assign n40578 = n10843 & n39724;
  assign n40579 = ~n39641 & ~n39831;
  assign n40580 = ~n10843 & ~n39737;
  assign n40581 = ~n40579 & n40580;
  assign n40582 = ~n40578 & ~n40581;
  assign n40583 = ~pi0219 & ~n40582;
  assign n40584 = ~n40569 & ~n40583;
  assign n40585 = pi1152 & ~n40584;
  assign n40586 = n40538 & ~n40567;
  assign n40587 = ~n40585 & ~n40586;
  assign n40588 = n40577 & ~n40587;
  assign n40589 = pi0212 & ~n39755;
  assign n40590 = n40505 & ~n40589;
  assign n40591 = pi1152 & ~n40590;
  assign n40592 = n39879 & n40591;
  assign n40593 = pi1151 & ~n40082;
  assign n40594 = ~n39699 & ~n40511;
  assign n40595 = ~pi0219 & ~n40594;
  assign n40596 = n40554 & ~n40595;
  assign n40597 = n40593 & ~n40596;
  assign n40598 = ~n40592 & n40597;
  assign n40599 = pi1150 & ~n40588;
  assign n40600 = ~n40598 & n40599;
  assign n40601 = ~n40576 & ~n40600;
  assign n40602 = pi1149 & ~n40601;
  assign n40603 = ~n40547 & ~n40602;
  assign n40604 = ~pi0213 & ~n40603;
  assign n40605 = pi0209 & ~n40481;
  assign n40606 = ~n40604 & n40605;
  assign n40607 = ~pi1150 & pi1151;
  assign n40608 = ~n40143 & n40607;
  assign n40609 = ~n40124 & n40523;
  assign n40610 = ~n40077 & n40500;
  assign n40611 = pi1150 & ~n40610;
  assign n40612 = ~n40609 & n40611;
  assign n40613 = ~pi1149 & ~n40608;
  assign n40614 = ~n40612 & n40613;
  assign n40615 = n40088 & n40593;
  assign n40616 = ~pi1151 & n40134;
  assign n40617 = pi1150 & ~n40615;
  assign n40618 = ~n40616 & n40617;
  assign n40619 = ~n40199 & n40565;
  assign n40620 = ~n40165 & n40548;
  assign n40621 = ~pi1150 & ~n40619;
  assign n40622 = ~n40620 & n40621;
  assign n40623 = pi1149 & ~n40618;
  assign n40624 = ~n40622 & n40623;
  assign n40625 = ~n40614 & ~n40624;
  assign n40626 = ~pi0213 & n40625;
  assign n40627 = ~n40153 & ~n40157;
  assign n40628 = ~n38769 & n39695;
  assign n40629 = ~n39696 & ~n40628;
  assign n40630 = ~n40151 & n40629;
  assign n40631 = ~n40627 & ~n40630;
  assign n40632 = ~pi0219 & ~n40631;
  assign n40633 = n40164 & ~n40632;
  assign n40634 = n39845 & ~n40633;
  assign n40635 = pi0299 & n39631;
  assign n40636 = ~n40182 & ~n40483;
  assign n40637 = ~po1038 & ~n40636;
  assign n40638 = ~n40635 & n40637;
  assign n40639 = n39828 & ~n40638;
  assign n40640 = ~pi1152 & ~n40639;
  assign n40641 = ~n40634 & n40640;
  assign n40642 = ~n40150 & ~n40152;
  assign n40643 = ~pi0219 & ~n40299;
  assign n40644 = ~n39700 & n40643;
  assign n40645 = ~n40642 & n40644;
  assign n40646 = n40164 & ~n40645;
  assign n40647 = n39871 & ~n40646;
  assign n40648 = ~n40083 & ~n40182;
  assign n40649 = ~n38641 & n39867;
  assign n40650 = ~n40648 & ~n40649;
  assign n40651 = ~pi0219 & ~n40650;
  assign n40652 = pi0219 & ~n40182;
  assign n40653 = ~po1038 & ~n40652;
  assign n40654 = ~n40651 & n40653;
  assign n40655 = n39893 & ~n40654;
  assign n40656 = pi1152 & ~n40655;
  assign n40657 = ~n40647 & n40656;
  assign n40658 = ~pi1150 & ~n40657;
  assign n40659 = ~n40641 & n40658;
  assign n40660 = ~pi0219 & ~n40086;
  assign n40661 = ~n40299 & n40660;
  assign n40662 = ~pi1153 & n40661;
  assign n40663 = pi0299 & n10485;
  assign n40664 = ~pi0219 & ~n40663;
  assign n40665 = n40195 & ~n40664;
  assign n40666 = ~n40303 & ~n40665;
  assign n40667 = ~n40662 & ~n40666;
  assign n40668 = n39845 & ~n40667;
  assign n40669 = pi1153 & n40483;
  assign n40670 = n39828 & ~n40669;
  assign n40671 = ~pi1152 & ~n40670;
  assign n40672 = ~pi1151 & ~n40127;
  assign n40673 = ~pi1152 & ~n40672;
  assign n40674 = ~n40671 & ~n40673;
  assign n40675 = ~n40668 & ~n40674;
  assign n40676 = ~pi0211 & n40661;
  assign n40677 = ~n40088 & ~n40676;
  assign n40678 = n39871 & ~n40677;
  assign n40679 = ~n40667 & n40678;
  assign n40680 = ~po1038 & ~n39768;
  assign n40681 = n10843 & ~n40172;
  assign n40682 = ~pi0299 & n39747;
  assign n40683 = ~n38423 & ~n40635;
  assign n40684 = ~n40682 & n40683;
  assign n40685 = n40230 & ~n40681;
  assign n40686 = ~n40684 & n40685;
  assign n40687 = n40680 & ~n40686;
  assign n40688 = n39893 & ~n40687;
  assign n40689 = pi1152 & ~n40688;
  assign n40690 = ~n40679 & n40689;
  assign n40691 = pi1150 & ~n40675;
  assign n40692 = ~n40690 & n40691;
  assign n40693 = pi1149 & ~n40692;
  assign n40694 = ~n40659 & n40693;
  assign n40695 = pi0219 & ~n39642;
  assign n40696 = ~po1038 & ~n40695;
  assign n40697 = ~n39839 & n40696;
  assign n40698 = n39845 & ~n40697;
  assign n40699 = n40671 & ~n40698;
  assign n40700 = pi0299 & n39864;
  assign n40701 = ~n39867 & n40700;
  assign n40702 = n39893 & ~n40701;
  assign n40703 = n40527 & ~n40531;
  assign n40704 = n40696 & ~n40703;
  assign n40705 = n39871 & ~n40697;
  assign n40706 = ~n40704 & n40705;
  assign n40707 = pi1152 & ~n40702;
  assign n40708 = ~n40706 & n40707;
  assign n40709 = ~pi1150 & ~n40699;
  assign n40710 = ~n40708 & n40709;
  assign n40711 = ~n39909 & n40100;
  assign n40712 = ~n38769 & ~n40105;
  assign n40713 = ~pi0211 & ~n40712;
  assign n40714 = n39909 & ~n40111;
  assign n40715 = ~n40713 & n40714;
  assign n40716 = ~n40711 & ~n40715;
  assign n40717 = ~po1038 & ~n40716;
  assign n40718 = n39828 & ~n40717;
  assign n40719 = pi0211 & ~n40066;
  assign n40720 = ~n11373 & n38675;
  assign n40721 = ~n39713 & ~n40720;
  assign n40722 = ~pi0211 & ~n38769;
  assign n40723 = ~n40721 & n40722;
  assign n40724 = ~n40719 & ~n40723;
  assign n40725 = ~n39736 & ~n40719;
  assign n40726 = pi0214 & n40725;
  assign n40727 = n40062 & ~n40071;
  assign n40728 = pi0212 & ~n40727;
  assign n40729 = ~n40726 & n40728;
  assign n40730 = ~n40724 & n40729;
  assign n40731 = ~n40070 & ~n40723;
  assign n40732 = n40063 & ~n40731;
  assign n40733 = ~pi0219 & ~n40732;
  assign n40734 = ~n40730 & n40733;
  assign n40735 = n40310 & ~n40734;
  assign n40736 = n39845 & ~n40735;
  assign n40737 = ~pi1152 & ~n40718;
  assign n40738 = ~n40736 & n40737;
  assign n40739 = pi0214 & n40724;
  assign n40740 = n40063 & ~n40739;
  assign n40741 = ~pi0214 & n40724;
  assign n40742 = n40315 & ~n40741;
  assign n40743 = ~pi0219 & ~n40740;
  assign n40744 = ~n40742 & n40743;
  assign n40745 = n40310 & ~n40744;
  assign n40746 = n39871 & ~n40745;
  assign n40747 = ~n40105 & ~n40635;
  assign n40748 = pi0214 & n40747;
  assign n40749 = n40108 & ~n40748;
  assign n40750 = ~pi0214 & n40747;
  assign n40751 = n40113 & ~n40750;
  assign n40752 = ~n40749 & ~n40751;
  assign n40753 = ~pi0219 & ~n40752;
  assign n40754 = n40123 & ~n40753;
  assign n40755 = n39893 & ~n40754;
  assign n40756 = pi1152 & ~n40746;
  assign n40757 = ~n40755 & n40756;
  assign n40758 = pi1150 & ~n40738;
  assign n40759 = ~n40757 & n40758;
  assign n40760 = ~pi1149 & ~n40710;
  assign n40761 = ~n40759 & n40760;
  assign n40762 = ~n40694 & ~n40761;
  assign n40763 = pi0213 & ~n40762;
  assign n40764 = ~pi0209 & ~n40626;
  assign n40765 = ~n40763 & n40764;
  assign n40766 = ~n40606 & ~n40765;
  assign n40767 = pi0230 & ~n40766;
  assign n40768 = ~pi0230 & ~pi0241;
  assign po0398 = ~n40767 & ~n40768;
  assign n40770 = ~pi0230 & ~pi0242;
  assign n40771 = pi0219 & ~n38419;
  assign n40772 = pi0214 & ~n39414;
  assign n40773 = ~pi0214 & ~n40211;
  assign n40774 = ~n40772 & ~n40773;
  assign n40775 = pi0212 & ~n40774;
  assign n40776 = ~pi0212 & n40212;
  assign n40777 = ~pi0219 & ~n40776;
  assign n40778 = ~n40775 & n40777;
  assign n40779 = n38416 & ~n40771;
  assign n40780 = ~n40778 & n40779;
  assign n40781 = pi0199 & pi1144;
  assign n40782 = ~pi0200 & ~n40781;
  assign n40783 = ~n40333 & n40782;
  assign n40784 = ~pi0299 & ~n40330;
  assign n40785 = ~n40783 & n40784;
  assign n40786 = n38826 & n40785;
  assign n40787 = ~pi0207 & ~n40785;
  assign n40788 = ~pi0299 & ~n39392;
  assign n40789 = ~n39393 & n40782;
  assign n40790 = n40788 & ~n40789;
  assign n40791 = pi0207 & ~n40790;
  assign n40792 = pi0208 & ~n40787;
  assign n40793 = ~n40791 & n40792;
  assign n40794 = ~n40786 & ~n40793;
  assign n40795 = ~pi0214 & n40794;
  assign n40796 = ~pi0212 & ~n40795;
  assign n40797 = n38449 & n40785;
  assign n40798 = ~n40234 & ~n40797;
  assign n40799 = ~n40793 & n40798;
  assign n40800 = ~pi0211 & ~n40799;
  assign n40801 = ~n39484 & ~n40797;
  assign n40802 = ~n40793 & n40801;
  assign n40803 = pi0211 & ~n40802;
  assign n40804 = ~n40800 & ~n40803;
  assign n40805 = pi0214 & n40804;
  assign n40806 = n40796 & ~n40805;
  assign n40807 = ~pi0211 & ~n40802;
  assign n40808 = ~n38612 & ~n40797;
  assign n40809 = ~n40793 & n40808;
  assign n40810 = pi0211 & ~n40809;
  assign n40811 = pi0214 & ~n40807;
  assign n40812 = ~n40810 & n40811;
  assign n40813 = ~pi0214 & n40804;
  assign n40814 = pi0212 & ~n40812;
  assign n40815 = ~n40813 & n40814;
  assign n40816 = ~pi0219 & ~n40806;
  assign n40817 = ~n40815 & n40816;
  assign n40818 = ~n38414 & ~n40794;
  assign n40819 = pi0219 & ~n40818;
  assign n40820 = n38414 & ~n40809;
  assign n40821 = n40819 & ~n40820;
  assign n40822 = ~po1038 & ~n40821;
  assign n40823 = ~n40817 & n40822;
  assign n40824 = ~n40780 & ~n40823;
  assign n40825 = pi0213 & n40824;
  assign n40826 = n38413 & ~n40786;
  assign n40827 = pi0211 & ~n40786;
  assign n40828 = n38414 & ~n38680;
  assign n40829 = ~n40797 & n40828;
  assign n40830 = ~n40827 & ~n40829;
  assign n40831 = pi0219 & ~n40830;
  assign n40832 = n10843 & ~n38457;
  assign n40833 = ~n38431 & n38608;
  assign n40834 = ~n40832 & ~n40833;
  assign n40835 = ~pi0219 & ~n40797;
  assign n40836 = ~n40834 & n40835;
  assign n40837 = ~n40826 & ~n40836;
  assign n40838 = ~n40831 & n40837;
  assign n40839 = ~n40793 & ~n40838;
  assign n40840 = ~po1038 & ~n40839;
  assign n40841 = ~pi0213 & ~n38430;
  assign n40842 = ~n40840 & n40841;
  assign n40843 = ~n40825 & ~n40842;
  assign n40844 = pi0209 & ~n40843;
  assign n40845 = ~pi0213 & ~n38476;
  assign n40846 = pi0219 & n38413;
  assign n40847 = ~n40771 & ~n40846;
  assign n40848 = ~n40778 & n40847;
  assign n40849 = pi0299 & ~n40848;
  assign n40850 = ~po1038 & ~n40849;
  assign n40851 = ~n38468 & n40850;
  assign n40852 = ~n40780 & ~n40851;
  assign n40853 = pi0213 & ~n40852;
  assign n40854 = ~pi0209 & ~n40853;
  assign n40855 = ~n40845 & n40854;
  assign n40856 = ~n40844 & ~n40855;
  assign n40857 = pi0230 & ~n40856;
  assign po0399 = ~n40770 & ~n40857;
  assign n40859 = pi0253 & pi0254;
  assign n40860 = pi0267 & n40859;
  assign n40861 = ~pi0263 & n40860;
  assign n40862 = ~pi0083 & ~pi0085;
  assign n40863 = pi0314 & ~n40862;
  assign n40864 = pi0802 & n40863;
  assign n40865 = pi0276 & n40864;
  assign n40866 = ~pi1091 & n40865;
  assign n40867 = pi0271 & n40866;
  assign n40868 = pi0273 & n40867;
  assign n40869 = pi0243 & n40868;
  assign n40870 = ~pi1091 & ~n40865;
  assign n40871 = pi0271 & ~n40870;
  assign n40872 = ~pi1091 & ~n40871;
  assign n40873 = pi0273 & ~n40872;
  assign n40874 = ~pi1091 & ~n40873;
  assign n40875 = ~pi0243 & n40874;
  assign n40876 = pi0243 & ~pi1091;
  assign n40877 = n38478 & ~n40876;
  assign n40878 = ~n40866 & n40877;
  assign n40879 = ~n40869 & ~n40878;
  assign n40880 = ~n40875 & n40879;
  assign n40881 = pi0219 & ~n40880;
  assign n40882 = ~n38479 & ~n38487;
  assign n40883 = pi1091 & n40882;
  assign n40884 = ~pi0081 & n40862;
  assign n40885 = pi0314 & ~n40884;
  assign n40886 = pi0802 & n40885;
  assign n40887 = pi0276 & n40886;
  assign n40888 = ~pi1091 & n40887;
  assign n40889 = pi0271 & n40888;
  assign n40890 = pi0273 & n40889;
  assign n40891 = ~n40873 & ~n40890;
  assign n40892 = n40876 & n40891;
  assign n40893 = ~pi0243 & n40890;
  assign n40894 = ~pi0219 & ~n40883;
  assign n40895 = ~n40893 & n40894;
  assign n40896 = ~n40892 & n40895;
  assign n40897 = ~n40881 & ~n40896;
  assign n40898 = n40861 & ~n40897;
  assign n40899 = ~pi0243 & ~pi1091;
  assign n40900 = ~pi0219 & ~n40882;
  assign n40901 = pi1157 & n38519;
  assign n40902 = ~n40900 & ~n40901;
  assign n40903 = pi1091 & ~n40902;
  assign n40904 = ~n40899 & ~n40903;
  assign n40905 = ~n40861 & ~n40904;
  assign n40906 = po1038 & ~n40905;
  assign n40907 = ~n40898 & n40906;
  assign n40908 = pi0272 & pi0283;
  assign n40909 = pi0275 & n40908;
  assign n40910 = pi0268 & n40909;
  assign n40911 = ~pi0299 & pi1091;
  assign n40912 = n38841 & n40911;
  assign n40913 = ~n40899 & ~n40912;
  assign n40914 = pi1156 & ~n40913;
  assign n40915 = pi1091 & ~n38955;
  assign n40916 = n39457 & n40915;
  assign n40917 = ~n40914 & ~n40916;
  assign n40918 = ~pi0299 & n38699;
  assign n40919 = pi1091 & ~n40918;
  assign n40920 = ~n40876 & ~n40919;
  assign n40921 = ~pi1155 & ~n40899;
  assign n40922 = ~n40876 & ~n40921;
  assign n40923 = n38568 & n40922;
  assign n40924 = ~n40920 & ~n40923;
  assign n40925 = ~pi1156 & ~n40924;
  assign n40926 = n40917 & ~n40925;
  assign n40927 = pi1157 & ~n40926;
  assign n40928 = ~n40915 & n40922;
  assign n40929 = ~pi1156 & ~n40928;
  assign n40930 = pi1155 & ~n40876;
  assign n40931 = pi0199 & pi1091;
  assign n40932 = ~pi0299 & n40931;
  assign n40933 = n40930 & ~n40932;
  assign n40934 = pi1156 & ~n40933;
  assign n40935 = ~pi1155 & ~n40876;
  assign n40936 = ~n11444 & n40911;
  assign n40937 = n40935 & ~n40936;
  assign n40938 = n40934 & ~n40937;
  assign n40939 = ~pi1157 & ~n40929;
  assign n40940 = ~n40938 & n40939;
  assign n40941 = ~n40927 & ~n40940;
  assign n40942 = pi0211 & ~n40941;
  assign n40943 = pi1091 & ~n11445;
  assign n40944 = n40935 & ~n40943;
  assign n40945 = ~n40933 & ~n40944;
  assign n40946 = pi0200 & ~pi1156;
  assign n40947 = n40911 & n40946;
  assign n40948 = ~n40945 & ~n40947;
  assign n40949 = ~pi1157 & ~n40948;
  assign n40950 = n40913 & n40934;
  assign n40951 = pi0200 & pi1091;
  assign n40952 = ~pi0299 & n40951;
  assign n40953 = n40930 & ~n40952;
  assign n40954 = ~pi1155 & n40920;
  assign n40955 = ~pi1156 & ~n40953;
  assign n40956 = ~n40954 & n40955;
  assign n40957 = ~n40950 & ~n40956;
  assign n40958 = pi1157 & ~n40957;
  assign n40959 = ~pi0211 & ~n40949;
  assign n40960 = ~n40958 & n40959;
  assign n40961 = ~n40942 & ~n40960;
  assign n40962 = ~pi0219 & ~n40961;
  assign n40963 = n39369 & ~n40914;
  assign n40964 = ~n40925 & n40963;
  assign n40965 = pi0299 & pi1091;
  assign n40966 = n40948 & ~n40965;
  assign n40967 = ~pi1157 & ~n40966;
  assign n40968 = pi1091 & n38700;
  assign n40969 = n40935 & ~n40968;
  assign n40970 = ~n40953 & ~n40969;
  assign n40971 = ~pi1156 & ~n40970;
  assign n40972 = n38478 & ~n40971;
  assign n40973 = n40917 & n40972;
  assign n40974 = pi0219 & ~n40964;
  assign n40975 = ~n40967 & ~n40973;
  assign n40976 = n40974 & n40975;
  assign n40977 = ~n40962 & ~n40976;
  assign n40978 = ~n40861 & ~n40977;
  assign n40979 = pi0199 & ~n40874;
  assign n40980 = ~pi1091 & n40891;
  assign n40981 = ~pi0199 & ~n40980;
  assign n40982 = ~n40979 & ~n40981;
  assign n40983 = ~pi0200 & ~n40888;
  assign n40984 = ~n40982 & ~n40983;
  assign n40985 = ~pi0299 & ~n40984;
  assign n40986 = pi0299 & n40874;
  assign n40987 = ~n40890 & n40986;
  assign n40988 = ~n40985 & ~n40987;
  assign n40989 = ~pi0243 & ~n40988;
  assign n40990 = ~pi0200 & ~n40874;
  assign n40991 = n40888 & ~n40982;
  assign n40992 = ~pi0299 & ~n40991;
  assign n40993 = ~n40990 & n40992;
  assign n40994 = pi0299 & ~n40868;
  assign n40995 = ~n40993 & ~n40994;
  assign n40996 = pi0243 & n40995;
  assign n40997 = ~n40989 & ~n40996;
  assign n40998 = pi1155 & ~n40997;
  assign n40999 = ~n40981 & n40985;
  assign n41000 = ~n40986 & ~n40999;
  assign n41001 = ~pi0243 & ~n41000;
  assign n41002 = ~n40979 & n40992;
  assign n41003 = n40995 & ~n41002;
  assign n41004 = pi0243 & n41003;
  assign n41005 = ~n41001 & ~n41004;
  assign n41006 = ~n40998 & n41005;
  assign n41007 = ~pi1156 & ~n41006;
  assign n41008 = ~n40990 & n41002;
  assign n41009 = ~n40986 & ~n41008;
  assign n41010 = ~pi0243 & n41009;
  assign n41011 = ~n40979 & n40985;
  assign n41012 = ~n40981 & n40993;
  assign n41013 = ~n40994 & ~n41012;
  assign n41014 = ~n41011 & n41013;
  assign n41015 = pi0243 & ~n41014;
  assign n41016 = ~n41010 & ~n41015;
  assign n41017 = ~pi1155 & ~n41001;
  assign n41018 = pi1155 & ~n40989;
  assign n41019 = pi0243 & n41013;
  assign n41020 = n41018 & ~n41019;
  assign n41021 = ~n41017 & ~n41020;
  assign n41022 = ~n41016 & ~n41021;
  assign n41023 = pi1156 & ~n41022;
  assign n41024 = n39369 & ~n41007;
  assign n41025 = ~n41023 & n41024;
  assign n41026 = ~n40981 & n40992;
  assign n41027 = n40996 & ~n41026;
  assign n41028 = ~n40986 & ~n41011;
  assign n41029 = ~pi0243 & ~n41028;
  assign n41030 = pi1155 & ~n41029;
  assign n41031 = ~n41027 & n41030;
  assign n41032 = ~n40992 & ~n40994;
  assign n41033 = n40899 & ~n41032;
  assign n41034 = ~pi1155 & ~n41033;
  assign n41035 = pi0243 & n41032;
  assign n41036 = n41034 & ~n41035;
  assign n41037 = ~pi1156 & ~n41036;
  assign n41038 = ~n41031 & n41037;
  assign n41039 = ~n40994 & ~n41026;
  assign n41040 = pi1155 & n41039;
  assign n41041 = ~n40985 & n41039;
  assign n41042 = ~n41040 & ~n41041;
  assign n41043 = pi0243 & ~n41042;
  assign n41044 = pi0299 & ~n40890;
  assign n41045 = ~n40993 & ~n41044;
  assign n41046 = ~pi1155 & n41045;
  assign n41047 = ~n40888 & n41046;
  assign n41048 = ~n40986 & ~n41002;
  assign n41049 = ~pi0243 & ~n41048;
  assign n41050 = ~n41047 & n41049;
  assign n41051 = ~n41043 & ~n41050;
  assign n41052 = pi1156 & ~n41051;
  assign n41053 = ~pi1157 & ~n41038;
  assign n41054 = ~n41052 & n41053;
  assign n41055 = ~n40986 & ~n40993;
  assign n41056 = pi0243 & ~n41055;
  assign n41057 = ~n40994 & ~n40999;
  assign n41058 = ~pi0243 & ~n41057;
  assign n41059 = pi0243 & ~n41002;
  assign n41060 = ~pi1155 & ~n41059;
  assign n41061 = ~n41058 & n41060;
  assign n41062 = ~n40985 & ~n40994;
  assign n41063 = ~pi0243 & pi1155;
  assign n41064 = n41062 & n41063;
  assign n41065 = ~pi1156 & ~n41064;
  assign n41066 = ~n41056 & n41065;
  assign n41067 = ~n41061 & n41066;
  assign n41068 = ~n41014 & n41056;
  assign n41069 = pi1155 & ~n41068;
  assign n41070 = n41010 & n41062;
  assign n41071 = n41069 & ~n41070;
  assign n41072 = ~n41008 & ~n41044;
  assign n41073 = ~n40876 & ~n41072;
  assign n41074 = ~n41001 & ~n41073;
  assign n41075 = ~n41016 & n41074;
  assign n41076 = ~pi1155 & ~n41075;
  assign n41077 = ~n41071 & ~n41076;
  assign n41078 = pi1156 & ~n41077;
  assign n41079 = n38478 & ~n41067;
  assign n41080 = ~n41078 & n41079;
  assign n41081 = ~n41025 & ~n41054;
  assign n41082 = ~n41080 & n41081;
  assign n41083 = pi0219 & ~n41082;
  assign n41084 = ~n40992 & ~n41044;
  assign n41085 = ~pi1155 & n41084;
  assign n41086 = ~n41017 & ~n41085;
  assign n41087 = pi0243 & n41045;
  assign n41088 = ~n41002 & n41087;
  assign n41089 = ~n41086 & ~n41088;
  assign n41090 = ~pi1156 & ~n41089;
  assign n41091 = ~n40985 & ~n41044;
  assign n41092 = ~pi0243 & n41091;
  assign n41093 = ~n40987 & ~n40993;
  assign n41094 = pi0243 & ~n41093;
  assign n41095 = ~n41092 & ~n41094;
  assign n41096 = n41090 & n41095;
  assign n41097 = ~n40987 & ~n41012;
  assign n41098 = pi1155 & n41097;
  assign n41099 = ~n41069 & ~n41098;
  assign n41100 = ~n41008 & n41092;
  assign n41101 = ~n41099 & ~n41100;
  assign n41102 = ~n40999 & ~n41008;
  assign n41103 = ~n40987 & n41102;
  assign n41104 = ~pi0243 & ~n41103;
  assign n41105 = ~n41011 & ~n41044;
  assign n41106 = pi0243 & ~n41012;
  assign n41107 = n41105 & n41106;
  assign n41108 = ~n41104 & ~n41107;
  assign n41109 = ~pi1155 & ~n41108;
  assign n41110 = ~n41101 & ~n41109;
  assign n41111 = pi1156 & ~n41110;
  assign n41112 = pi1157 & ~n41096;
  assign n41113 = ~n41111 & n41112;
  assign n41114 = ~pi1155 & n41093;
  assign n41115 = ~n41091 & n41114;
  assign n41116 = ~n40987 & ~n41026;
  assign n41117 = pi0243 & ~n41116;
  assign n41118 = ~n41002 & ~n41044;
  assign n41119 = ~pi0243 & n41118;
  assign n41120 = ~n41117 & ~n41119;
  assign n41121 = pi1156 & ~n41047;
  assign n41122 = n41120 & n41121;
  assign n41123 = ~n41115 & n41122;
  assign n41124 = pi0243 & n41084;
  assign n41125 = ~n41034 & ~n41085;
  assign n41126 = ~n41124 & ~n41125;
  assign n41127 = ~pi1156 & ~n41126;
  assign n41128 = n41095 & n41120;
  assign n41129 = pi1155 & ~n41128;
  assign n41130 = n41127 & ~n41129;
  assign n41131 = ~pi1157 & ~n41123;
  assign n41132 = ~n41130 & n41131;
  assign n41133 = ~pi0211 & ~n41132;
  assign n41134 = ~n41113 & n41133;
  assign n41135 = n41018 & ~n41087;
  assign n41136 = n40930 & n40979;
  assign n41137 = ~n41135 & ~n41136;
  assign n41138 = n41127 & n41137;
  assign n41139 = ~pi1157 & ~n41122;
  assign n41140 = ~n41138 & n41139;
  assign n41141 = n41090 & ~n41135;
  assign n41142 = ~n41073 & n41110;
  assign n41143 = pi1156 & ~n41142;
  assign n41144 = pi1157 & ~n41141;
  assign n41145 = ~n41143 & n41144;
  assign n41146 = pi0211 & ~n41140;
  assign n41147 = ~n41145 & n41146;
  assign n41148 = ~pi0219 & ~n41134;
  assign n41149 = ~n41147 & n41148;
  assign n41150 = n40861 & ~n41083;
  assign n41151 = ~n41149 & n41150;
  assign n41152 = ~po1038 & ~n40978;
  assign n41153 = ~n41151 & n41152;
  assign n41154 = ~n40907 & n40910;
  assign n41155 = ~n41153 & n41154;
  assign n41156 = ~po1038 & n40977;
  assign n41157 = po1038 & n40904;
  assign n41158 = ~n40910 & ~n41157;
  assign n41159 = ~n41156 & n41158;
  assign n41160 = ~pi0230 & ~n41159;
  assign n41161 = ~n41155 & n41160;
  assign n41162 = ~n16479 & ~n40902;
  assign n41163 = pi0199 & ~n39467;
  assign n41164 = ~n38840 & ~n40946;
  assign n41165 = ~n41163 & n41164;
  assign n41166 = n16479 & n41165;
  assign n41167 = pi0230 & ~n41162;
  assign n41168 = ~n41166 & n41167;
  assign po0400 = ~n41161 & ~n41168;
  assign n41170 = ~pi0230 & ~pi0244;
  assign n41171 = pi0213 & ~n40405;
  assign n41172 = ~pi0211 & ~n38543;
  assign n41173 = ~n40357 & n41172;
  assign n41174 = ~n40346 & ~n41173;
  assign n41175 = n40344 & ~n41174;
  assign n41176 = ~n38610 & n40390;
  assign n41177 = ~n40383 & ~n41176;
  assign n41178 = ~n40411 & ~n41177;
  assign n41179 = pi0214 & ~n41178;
  assign n41180 = n40364 & ~n41179;
  assign n41181 = n38420 & n40293;
  assign n41182 = ~pi0214 & n41177;
  assign n41183 = pi0212 & ~n41181;
  assign n41184 = ~n41182 & n41183;
  assign n41185 = ~n40411 & n41184;
  assign n41186 = ~pi0219 & ~n41180;
  assign n41187 = ~n41185 & n41186;
  assign n41188 = n40447 & ~n41175;
  assign n41189 = ~n41187 & n41188;
  assign n41190 = pi0299 & n39410;
  assign n41191 = pi0214 & n41177;
  assign n41192 = n40388 & ~n41191;
  assign n41193 = ~n40381 & n41184;
  assign n41194 = ~pi0219 & ~n41192;
  assign n41195 = ~n41193 & n41194;
  assign n41196 = pi1147 & ~n41190;
  assign n41197 = n40410 & n41196;
  assign n41198 = ~n41195 & n41197;
  assign n41199 = ~pi0213 & ~n39420;
  assign n41200 = ~n41198 & n41199;
  assign n41201 = ~n41189 & n41200;
  assign n41202 = ~n41171 & ~n41201;
  assign n41203 = pi0209 & ~n41202;
  assign n41204 = ~pi0213 & ~n39427;
  assign n41205 = n40244 & ~n40247;
  assign n41206 = ~n40224 & ~n41205;
  assign n41207 = ~n10843 & n40236;
  assign n41208 = n10843 & ~n40231;
  assign n41209 = n40244 & ~n40246;
  assign n41210 = n38665 & ~n41207;
  assign n41211 = ~n41208 & n41210;
  assign n41212 = ~n41209 & n41211;
  assign n41213 = ~n39398 & ~n40253;
  assign n41214 = ~n41212 & n41213;
  assign n41215 = ~po1038 & ~n41214;
  assign n41216 = ~n41206 & ~n41215;
  assign n41217 = pi0213 & ~n41216;
  assign n41218 = ~pi0209 & ~n41204;
  assign n41219 = ~n41217 & n41218;
  assign n41220 = ~n41203 & ~n41219;
  assign n41221 = pi0230 & ~n41220;
  assign po0401 = ~n41170 & ~n41221;
  assign n41223 = ~pi0213 & ~n40824;
  assign n41224 = pi1146 & n39869;
  assign n41225 = ~pi1147 & ~n41224;
  assign n41226 = n39865 & ~n40145;
  assign n41227 = n41225 & ~n41226;
  assign n41228 = ~n38413 & n40800;
  assign n41229 = n40819 & ~n41228;
  assign n41230 = ~po1038 & ~n41229;
  assign n41231 = pi0214 & ~n40235;
  assign n41232 = ~pi0299 & ~n40804;
  assign n41233 = n41231 & ~n41232;
  assign n41234 = pi0212 & ~n41233;
  assign n41235 = ~pi0299 & n40802;
  assign n41236 = ~pi0211 & ~n41235;
  assign n41237 = n40794 & ~n41236;
  assign n41238 = ~pi0214 & n41237;
  assign n41239 = n41234 & ~n41238;
  assign n41240 = n40796 & ~n41237;
  assign n41241 = ~pi0219 & ~n41240;
  assign n41242 = ~n41239 & n41241;
  assign n41243 = n41230 & ~n41242;
  assign n41244 = n41227 & ~n41243;
  assign n41245 = pi1147 & ~n39865;
  assign n41246 = ~n41224 & n41245;
  assign n41247 = pi0211 & ~n40799;
  assign n41248 = ~n41236 & ~n41247;
  assign n41249 = pi0214 & ~n41248;
  assign n41250 = ~pi0214 & ~n41235;
  assign n41251 = ~n41249 & ~n41250;
  assign n41252 = pi0212 & ~n41251;
  assign n41253 = n40796 & ~n41235;
  assign n41254 = ~pi0219 & ~n41253;
  assign n41255 = ~n41252 & n41254;
  assign n41256 = n41230 & ~n41255;
  assign n41257 = n41246 & ~n41256;
  assign n41258 = pi1148 & ~n41244;
  assign n41259 = ~n41257 & n41258;
  assign n41260 = ~n40407 & ~n41246;
  assign n41261 = ~n13061 & n40794;
  assign n41262 = ~pi0214 & ~n41261;
  assign n41263 = ~n41249 & ~n41262;
  assign n41264 = pi0212 & ~n41263;
  assign n41265 = n40796 & ~n41261;
  assign n41266 = ~pi0219 & ~n41265;
  assign n41267 = ~n41264 & n41266;
  assign n41268 = n41230 & ~n41267;
  assign n41269 = ~n41260 & ~n41268;
  assign n41270 = ~n40795 & n41234;
  assign n41271 = ~pi0212 & ~n40794;
  assign n41272 = ~pi0219 & ~n41271;
  assign n41273 = ~n41270 & n41272;
  assign n41274 = n41230 & ~n41273;
  assign n41275 = n41225 & ~n41274;
  assign n41276 = ~pi1148 & ~n41269;
  assign n41277 = ~n41275 & n41276;
  assign n41278 = ~n41259 & ~n41277;
  assign n41279 = pi0213 & ~n41278;
  assign n41280 = ~pi0209 & ~n41223;
  assign n41281 = ~n41279 & n41280;
  assign n41282 = pi0199 & pi1146;
  assign n41283 = n38699 & ~n41282;
  assign n41284 = n38550 & ~n41283;
  assign n41285 = ~n10487 & ~n41284;
  assign n41286 = n40339 & ~n41283;
  assign n41287 = pi0207 & n41286;
  assign n41288 = ~n38826 & ~n41287;
  assign n41289 = ~n41285 & ~n41288;
  assign n41290 = ~n38414 & n41289;
  assign n41291 = pi0219 & ~n41290;
  assign n41292 = n38449 & n41284;
  assign n41293 = pi0208 & n41286;
  assign n41294 = ~pi0200 & ~n41282;
  assign n41295 = n38550 & ~n41294;
  assign n41296 = ~pi0207 & n41295;
  assign n41297 = ~n40234 & ~n41296;
  assign n41298 = ~n41287 & n41297;
  assign n41299 = pi0208 & ~n41298;
  assign n41300 = ~pi0299 & n41299;
  assign n41301 = ~n41292 & ~n41293;
  assign n41302 = ~n41300 & n41301;
  assign n41303 = ~n40234 & n41302;
  assign n41304 = n38414 & ~n41303;
  assign n41305 = n41291 & ~n41304;
  assign n41306 = ~pi0214 & ~n41289;
  assign n41307 = ~pi0212 & ~n41306;
  assign n41308 = ~pi0299 & n41302;
  assign n41309 = n41307 & ~n41308;
  assign n41310 = ~pi0219 & ~n41309;
  assign n41311 = pi0212 & ~n41308;
  assign n41312 = n10484 & n41303;
  assign n41313 = n41311 & ~n41312;
  assign n41314 = n41310 & ~n41313;
  assign n41315 = ~po1038 & ~n41305;
  assign n41316 = ~n41314 & n41315;
  assign n41317 = n41246 & ~n41316;
  assign n41318 = ~pi0208 & n40234;
  assign n41319 = n40339 & ~n41294;
  assign n41320 = pi0207 & n41319;
  assign n41321 = pi1146 & ~n38700;
  assign n41322 = ~n41320 & ~n41321;
  assign n41323 = pi0208 & ~n41322;
  assign n41324 = ~pi0207 & ~n41293;
  assign n41325 = n39658 & ~n41283;
  assign n41326 = ~n41324 & n41325;
  assign n41327 = ~n41318 & ~n41323;
  assign n41328 = ~n41326 & n41327;
  assign n41329 = ~pi0299 & ~n41328;
  assign n41330 = ~pi0214 & ~n41329;
  assign n41331 = ~pi0212 & ~n41330;
  assign n41332 = ~n10487 & ~n39659;
  assign n41333 = n41319 & ~n41332;
  assign n41334 = pi0211 & ~n41333;
  assign n41335 = ~pi0299 & ~n41319;
  assign n41336 = ~n41328 & ~n41335;
  assign n41337 = ~pi0299 & ~n41336;
  assign n41338 = ~pi0211 & n41337;
  assign n41339 = ~n41334 & ~n41338;
  assign n41340 = ~n41329 & ~n41339;
  assign n41341 = n41331 & ~n41340;
  assign n41342 = ~pi0219 & ~n41341;
  assign n41343 = n41231 & ~n41329;
  assign n41344 = ~pi0214 & n41340;
  assign n41345 = pi0212 & ~n41344;
  assign n41346 = ~n41343 & n41345;
  assign n41347 = n41342 & ~n41346;
  assign n41348 = ~n38414 & n41329;
  assign n41349 = pi0219 & ~n41348;
  assign n41350 = n38414 & ~n41328;
  assign n41351 = n41349 & ~n41350;
  assign n41352 = ~po1038 & ~n41351;
  assign n41353 = ~n41347 & n41352;
  assign n41354 = n41227 & ~n41353;
  assign n41355 = pi1148 & ~n41317;
  assign n41356 = ~n41354 & n41355;
  assign n41357 = ~n40663 & ~n41329;
  assign n41358 = ~n41322 & ~n41357;
  assign n41359 = ~pi0219 & ~n41358;
  assign n41360 = pi0219 & ~n41333;
  assign n41361 = ~n38970 & ~n41360;
  assign n41362 = ~n38413 & ~n41334;
  assign n41363 = n41336 & n41362;
  assign n41364 = ~n41361 & ~n41363;
  assign n41365 = ~po1038 & ~n41364;
  assign n41366 = ~n41359 & n41365;
  assign n41367 = n41225 & ~n41366;
  assign n41368 = ~n10487 & ~n41295;
  assign n41369 = ~n41288 & ~n41368;
  assign n41370 = ~n13061 & ~n41369;
  assign n41371 = pi0214 & ~n41370;
  assign n41372 = ~pi0214 & n41369;
  assign n41373 = ~pi0212 & ~n41372;
  assign n41374 = ~n41371 & n41373;
  assign n41375 = ~pi0214 & ~n41370;
  assign n41376 = n38449 & n41295;
  assign n41377 = ~n41318 & ~n41376;
  assign n41378 = ~n41299 & n41377;
  assign n41379 = ~pi0299 & n41378;
  assign n41380 = pi0214 & ~n41379;
  assign n41381 = ~pi0211 & ~n41308;
  assign n41382 = ~n41289 & ~n41381;
  assign n41383 = n41380 & ~n41382;
  assign n41384 = pi0212 & ~n41383;
  assign n41385 = ~n41375 & n41384;
  assign n41386 = ~n41374 & ~n41385;
  assign n41387 = ~pi0219 & ~n41386;
  assign n41388 = ~pi1146 & ~n38783;
  assign n41389 = n40299 & ~n41388;
  assign n41390 = n41387 & ~n41389;
  assign n41391 = ~n38413 & n41369;
  assign n41392 = ~n38414 & ~n41391;
  assign n41393 = ~n41378 & ~n41392;
  assign n41394 = ~pi0212 & n41372;
  assign n41395 = pi0219 & ~n41394;
  assign n41396 = ~n41393 & n41395;
  assign n41397 = ~po1038 & ~n41396;
  assign n41398 = ~n41390 & n41397;
  assign n41399 = ~n41260 & ~n41398;
  assign n41400 = ~pi1148 & ~n41367;
  assign n41401 = ~n41399 & n41400;
  assign n41402 = ~n41356 & ~n41401;
  assign n41403 = pi0213 & ~n41402;
  assign n41404 = pi1147 & ~po1038;
  assign n41405 = ~n38612 & n41302;
  assign n41406 = n38414 & ~n41405;
  assign n41407 = n41291 & ~n41406;
  assign n41408 = ~n40231 & n41302;
  assign n41409 = pi0214 & n41408;
  assign n41410 = n41307 & ~n41409;
  assign n41411 = pi0299 & ~n40774;
  assign n41412 = n41302 & ~n41411;
  assign n41413 = pi0212 & ~n41412;
  assign n41414 = ~pi0219 & ~n41413;
  assign n41415 = ~n41410 & n41414;
  assign n41416 = n41404 & ~n41407;
  assign n41417 = ~n41415 & n41416;
  assign n41418 = ~pi0299 & n41328;
  assign n41419 = n38414 & ~n41418;
  assign n41420 = ~n38610 & n41419;
  assign n41421 = n41349 & ~n41420;
  assign n41422 = ~n40231 & ~n41329;
  assign n41423 = n41331 & ~n41422;
  assign n41424 = ~n41329 & ~n41411;
  assign n41425 = pi0212 & ~n41424;
  assign n41426 = ~pi0219 & ~n41425;
  assign n41427 = ~n41423 & n41426;
  assign n41428 = n40447 & ~n41421;
  assign n41429 = ~n41427 & n41428;
  assign n41430 = pi1148 & ~n40780;
  assign n41431 = ~n41417 & n41430;
  assign n41432 = ~n41429 & n41431;
  assign n41433 = ~n41379 & n41413;
  assign n41434 = n41380 & ~n41408;
  assign n41435 = ~n41372 & ~n41434;
  assign n41436 = ~pi0212 & ~n41435;
  assign n41437 = ~pi0219 & ~n41433;
  assign n41438 = ~n41436 & n41437;
  assign n41439 = ~n41379 & ~n41405;
  assign n41440 = ~pi0211 & ~n41439;
  assign n41441 = ~n41392 & ~n41440;
  assign n41442 = n41395 & ~n41441;
  assign n41443 = n41404 & ~n41438;
  assign n41444 = ~n41442 & n41443;
  assign n41445 = ~n41335 & n41425;
  assign n41446 = ~pi0214 & n41333;
  assign n41447 = pi0214 & ~n41337;
  assign n41448 = ~n41422 & n41447;
  assign n41449 = ~n41446 & ~n41448;
  assign n41450 = ~pi0212 & ~n41449;
  assign n41451 = ~pi0219 & ~n41445;
  assign n41452 = ~n41450 & n41451;
  assign n41453 = ~n38610 & ~n41337;
  assign n41454 = ~pi0211 & ~n41453;
  assign n41455 = n41362 & ~n41454;
  assign n41456 = ~n41361 & ~n41455;
  assign n41457 = n40447 & ~n41456;
  assign n41458 = ~n41452 & n41457;
  assign n41459 = ~pi1148 & ~n40780;
  assign n41460 = ~n41444 & n41459;
  assign n41461 = ~n41458 & n41460;
  assign n41462 = ~pi0213 & ~n41432;
  assign n41463 = ~n41461 & n41462;
  assign n41464 = pi0209 & ~n41463;
  assign n41465 = ~n41403 & n41464;
  assign n41466 = ~n41281 & ~n41465;
  assign n41467 = pi0230 & ~n41466;
  assign n41468 = ~pi0230 & ~pi0245;
  assign po0402 = ~n41467 & ~n41468;
  assign n41470 = ~pi1150 & n40134;
  assign n41471 = pi1150 & n40089;
  assign n41472 = pi1149 & ~n41470;
  assign n41473 = ~n41471 & n41472;
  assign n41474 = ~pi1150 & n40200;
  assign n41475 = pi1150 & n40166;
  assign n41476 = ~pi1149 & ~n41474;
  assign n41477 = ~n41475 & n41476;
  assign n41478 = ~n41473 & ~n41477;
  assign n41479 = pi1148 & ~n41478;
  assign n41480 = ~pi1150 & n40125;
  assign n41481 = pi1150 & n40078;
  assign n41482 = pi1149 & ~n41481;
  assign n41483 = ~n41480 & n41482;
  assign n41484 = ~pi1149 & pi1150;
  assign n41485 = ~n40143 & n41484;
  assign n41486 = ~n41483 & ~n41485;
  assign n41487 = ~pi1148 & ~n41486;
  assign n41488 = ~n41479 & ~n41487;
  assign n41489 = pi0213 & ~n41488;
  assign n41490 = ~n40184 & ~n40193;
  assign n41491 = n41227 & ~n41490;
  assign n41492 = ~n41227 & ~n41246;
  assign n41493 = pi0219 & ~n40234;
  assign n41494 = n40084 & ~n41493;
  assign n41495 = n40127 & ~n40181;
  assign n41496 = ~n41494 & ~n41495;
  assign n41497 = ~n40183 & ~n40255;
  assign n41498 = n38423 & ~n41497;
  assign n41499 = ~n40648 & ~n41498;
  assign n41500 = ~pi0219 & ~n41499;
  assign n41501 = ~n41496 & ~n41500;
  assign n41502 = ~n41492 & ~n41501;
  assign n41503 = ~pi1150 & ~n41491;
  assign n41504 = ~n41502 & n41503;
  assign n41505 = ~n40269 & ~n41494;
  assign n41506 = ~pi0214 & n39697;
  assign n41507 = pi0214 & ~n40147;
  assign n41508 = ~n40274 & n41507;
  assign n41509 = pi0212 & ~n41506;
  assign n41510 = ~n41508 & n41509;
  assign n41511 = n40156 & ~n41510;
  assign n41512 = ~n41505 & ~n41511;
  assign n41513 = n41227 & ~n41512;
  assign n41514 = ~n40276 & n40513;
  assign n41515 = ~pi0212 & ~n39661;
  assign n41516 = ~pi0219 & ~n41515;
  assign n41517 = ~n40525 & n41516;
  assign n41518 = ~n41514 & n41517;
  assign n41519 = ~n41505 & ~n41518;
  assign n41520 = n41246 & ~n41519;
  assign n41521 = pi1150 & ~n41513;
  assign n41522 = ~n41520 & n41521;
  assign n41523 = ~n41504 & ~n41522;
  assign n41524 = pi1148 & ~n41523;
  assign n41525 = pi1150 & n39639;
  assign n41526 = pi0299 & n40093;
  assign n41527 = ~pi0219 & ~n41526;
  assign n41528 = ~n41389 & n41527;
  assign n41529 = ~n41525 & n41528;
  assign n41530 = ~n41260 & n41529;
  assign n41531 = ~pi0219 & ~n40213;
  assign n41532 = ~n40664 & ~n41531;
  assign n41533 = n41494 & n41532;
  assign n41534 = n41225 & ~n41533;
  assign n41535 = ~n41260 & ~n41494;
  assign n41536 = ~n41534 & ~n41535;
  assign n41537 = pi1150 & n40140;
  assign n41538 = ~n41536 & ~n41537;
  assign n41539 = ~pi1148 & ~n41530;
  assign n41540 = ~n41538 & n41539;
  assign n41541 = ~n41524 & ~n41540;
  assign n41542 = ~pi1149 & ~n41541;
  assign n41543 = ~pi1146 & n40122;
  assign n41544 = n40084 & ~n40105;
  assign n41545 = ~n40123 & ~n41544;
  assign n41546 = n40213 & n40293;
  assign n41547 = ~n40100 & ~n41546;
  assign n41548 = n40121 & n41547;
  assign n41549 = ~n41543 & ~n41545;
  assign n41550 = ~n41548 & n41549;
  assign n41551 = ~n41260 & ~n41550;
  assign n41552 = ~n40102 & ~n40524;
  assign n41553 = ~pi0219 & ~n41552;
  assign n41554 = ~n41545 & ~n41553;
  assign n41555 = ~pi1146 & ~n40100;
  assign n41556 = n41554 & ~n41555;
  assign n41557 = n41225 & ~n41556;
  assign n41558 = ~pi1150 & ~n41557;
  assign n41559 = ~n41551 & n41558;
  assign n41560 = ~n40311 & ~n41494;
  assign n41561 = ~n40062 & ~n40725;
  assign n41562 = ~pi0214 & n40725;
  assign n41563 = n40074 & ~n41562;
  assign n41564 = ~pi0219 & ~n41563;
  assign n41565 = ~n41561 & n41564;
  assign n41566 = ~pi0212 & n41561;
  assign n41567 = n41564 & ~n41566;
  assign n41568 = ~pi0299 & n39713;
  assign n41569 = ~n40064 & ~n40234;
  assign n41570 = ~n41568 & n41569;
  assign n41571 = n41567 & n41570;
  assign n41572 = ~n41560 & ~n41565;
  assign n41573 = ~n41571 & n41572;
  assign n41574 = ~n40060 & ~n41573;
  assign n41575 = n40063 & ~n40073;
  assign n41576 = ~pi0219 & ~n41575;
  assign n41577 = ~n40729 & n41576;
  assign n41578 = n40310 & ~n41577;
  assign n41579 = ~n41574 & n41578;
  assign n41580 = n41225 & ~n41579;
  assign n41581 = ~n41260 & ~n41573;
  assign n41582 = pi1150 & ~n41581;
  assign n41583 = ~n41580 & n41582;
  assign n41584 = ~pi1148 & ~n41583;
  assign n41585 = ~n41559 & n41584;
  assign n41586 = ~n40127 & ~n41494;
  assign n41587 = n39747 & n41231;
  assign n41588 = n40189 & ~n41587;
  assign n41589 = ~n40172 & n40190;
  assign n41590 = ~n40177 & ~n41589;
  assign n41591 = ~n41227 & ~n41590;
  assign n41592 = n40192 & ~n41588;
  assign n41593 = ~n41591 & n41592;
  assign n41594 = ~n41586 & ~n41593;
  assign n41595 = ~n41492 & ~n41594;
  assign n41596 = ~pi1150 & ~n41595;
  assign n41597 = ~n40303 & ~n41533;
  assign n41598 = n41227 & n41597;
  assign n41599 = pi0214 & n40292;
  assign n41600 = n40298 & ~n41599;
  assign n41601 = ~pi0219 & ~n40295;
  assign n41602 = ~n41600 & n41601;
  assign n41603 = n40291 & ~n41602;
  assign n41604 = pi1146 & n40085;
  assign n41605 = n41246 & ~n41604;
  assign n41606 = ~n41603 & n41605;
  assign n41607 = pi1150 & ~n41606;
  assign n41608 = ~n41598 & n41607;
  assign n41609 = pi1148 & ~n41608;
  assign n41610 = ~n41596 & n41609;
  assign n41611 = pi1149 & ~n41610;
  assign n41612 = ~n41585 & n41611;
  assign n41613 = ~n41542 & ~n41612;
  assign n41614 = ~pi0213 & ~n41613;
  assign n41615 = pi0209 & ~n41489;
  assign n41616 = ~n41614 & n41615;
  assign n41617 = ~pi0213 & ~n41402;
  assign n41618 = pi0219 & ~n41369;
  assign n41619 = n41404 & ~n41618;
  assign n41620 = ~n41387 & n41619;
  assign n41621 = ~pi0212 & ~n41446;
  assign n41622 = ~n13061 & ~n41333;
  assign n41623 = pi0214 & ~n41622;
  assign n41624 = n41621 & ~n41623;
  assign n41625 = ~pi0214 & ~n41622;
  assign n41626 = pi0214 & n41339;
  assign n41627 = pi0212 & ~n41626;
  assign n41628 = ~n41625 & n41627;
  assign n41629 = ~n41624 & ~n41628;
  assign n41630 = ~pi0219 & ~n41629;
  assign n41631 = n40447 & ~n41360;
  assign n41632 = ~n41630 & n41631;
  assign n41633 = ~pi1150 & ~n40096;
  assign n41634 = ~n41620 & n41633;
  assign n41635 = ~n41632 & n41634;
  assign n41636 = n41373 & ~n41380;
  assign n41637 = ~pi0214 & ~n41379;
  assign n41638 = n41384 & ~n41637;
  assign n41639 = ~n41636 & ~n41638;
  assign n41640 = ~pi0219 & ~n41639;
  assign n41641 = ~n41618 & ~n41640;
  assign n41642 = pi1147 & ~n41641;
  assign n41643 = ~n41447 & n41621;
  assign n41644 = ~pi0214 & ~n41337;
  assign n41645 = n41627 & ~n41644;
  assign n41646 = ~n41643 & ~n41645;
  assign n41647 = ~pi0219 & ~n41646;
  assign n41648 = ~n41360 & ~n41647;
  assign n41649 = ~pi1147 & ~n41648;
  assign n41650 = ~po1038 & ~n41642;
  assign n41651 = ~n41649 & n41650;
  assign n41652 = pi1150 & ~n39865;
  assign n41653 = ~n41651 & n41652;
  assign n41654 = ~n41635 & ~n41653;
  assign n41655 = pi1149 & ~n41654;
  assign n41656 = pi1150 & n40207;
  assign n41657 = n41333 & ~n41656;
  assign n41658 = ~pi1147 & ~n41657;
  assign n41659 = pi1147 & ~n41369;
  assign n41660 = ~po1038 & ~n41658;
  assign n41661 = ~n41659 & n41660;
  assign n41662 = ~pi1147 & n41336;
  assign n41663 = n16479 & ~n41662;
  assign n41664 = n41656 & ~n41663;
  assign n41665 = ~pi1149 & ~n41661;
  assign n41666 = ~n41664 & n41665;
  assign n41667 = ~n41655 & ~n41666;
  assign n41668 = ~pi1148 & ~n41667;
  assign n41669 = ~n38413 & n41381;
  assign n41670 = n41291 & ~n41669;
  assign n41671 = n41404 & ~n41670;
  assign n41672 = pi0214 & ~n13061;
  assign n41673 = n41302 & n41672;
  assign n41674 = pi0212 & ~n41673;
  assign n41675 = ~n41306 & n41674;
  assign n41676 = ~pi0212 & n41289;
  assign n41677 = ~pi0219 & ~n41676;
  assign n41678 = ~n41675 & n41677;
  assign n41679 = n41671 & ~n41678;
  assign n41680 = n41349 & ~n41419;
  assign n41681 = n40447 & ~n41680;
  assign n41682 = ~pi0219 & n41357;
  assign n41683 = n41681 & ~n41682;
  assign n41684 = ~pi1150 & ~n39869;
  assign n41685 = ~n41679 & n41684;
  assign n41686 = ~n41683 & n41685;
  assign n41687 = ~n41329 & n41622;
  assign n41688 = pi0214 & n41687;
  assign n41689 = n41345 & ~n41688;
  assign n41690 = n41342 & ~n41689;
  assign n41691 = n41681 & ~n41690;
  assign n41692 = ~pi0214 & n41382;
  assign n41693 = n41674 & ~n41692;
  assign n41694 = n41307 & ~n41382;
  assign n41695 = ~pi0219 & ~n41694;
  assign n41696 = ~n41693 & n41695;
  assign n41697 = n41671 & ~n41696;
  assign n41698 = pi1150 & ~n40146;
  assign n41699 = ~n41697 & n41698;
  assign n41700 = ~n41691 & n41699;
  assign n41701 = ~pi1149 & ~n41686;
  assign n41702 = ~n41700 & n41701;
  assign n41703 = pi0057 & n38666;
  assign n41704 = ~n6305 & ~n38666;
  assign n41705 = n41310 & ~n41311;
  assign n41706 = ~n41670 & ~n41705;
  assign n41707 = n6305 & n41706;
  assign n41708 = ~pi0057 & pi1147;
  assign n41709 = ~n41704 & n41708;
  assign n41710 = ~n41707 & n41709;
  assign n41711 = n6305 & ~n38665;
  assign n41712 = n41348 & n41711;
  assign n41713 = ~n38666 & ~n41418;
  assign n41714 = ~pi0057 & ~pi1147;
  assign n41715 = ~n41704 & n41714;
  assign n41716 = ~n41713 & n41715;
  assign n41717 = ~n41712 & n41716;
  assign n41718 = ~n41703 & ~n41717;
  assign n41719 = ~n41710 & n41718;
  assign n41720 = pi1150 & ~n41719;
  assign n41721 = n41331 & ~n41688;
  assign n41722 = ~n41447 & n41687;
  assign n41723 = pi0212 & ~n41722;
  assign n41724 = ~pi0219 & ~n41721;
  assign n41725 = ~n41723 & n41724;
  assign n41726 = n41681 & ~n41725;
  assign n41727 = ~n40676 & n41404;
  assign n41728 = n41706 & n41727;
  assign n41729 = ~pi1150 & ~n40131;
  assign n41730 = ~n41728 & n41729;
  assign n41731 = ~n41726 & n41730;
  assign n41732 = pi1149 & ~n41731;
  assign n41733 = ~n41720 & n41732;
  assign n41734 = pi1148 & ~n41733;
  assign n41735 = ~n41702 & n41734;
  assign n41736 = pi0213 & ~n41735;
  assign n41737 = ~n41668 & n41736;
  assign n41738 = ~pi0209 & ~n41617;
  assign n41739 = ~n41737 & n41738;
  assign n41740 = ~n41616 & ~n41739;
  assign n41741 = pi0230 & ~n41740;
  assign n41742 = ~pi0230 & ~pi0246;
  assign po0403 = ~n41741 & ~n41742;
  assign n41744 = pi0213 & n40625;
  assign n41745 = pi1151 & ~n40131;
  assign n41746 = n40310 & ~n41565;
  assign n41747 = n41745 & ~n41746;
  assign n41748 = n40104 & ~n40119;
  assign n41749 = ~n41545 & ~n41748;
  assign n41750 = ~n40131 & ~n41749;
  assign n41751 = ~pi1151 & n41750;
  assign n41752 = pi1147 & ~n41747;
  assign n41753 = ~n41751 & n41752;
  assign n41754 = ~pi1147 & ~n40609;
  assign n41755 = pi1151 & ~n40096;
  assign n41756 = ~n40061 & ~n41567;
  assign n41757 = n41755 & ~n41756;
  assign n41758 = n41754 & ~n41757;
  assign n41759 = ~pi1149 & ~n41753;
  assign n41760 = ~n41758 & n41759;
  assign n41761 = pi1147 & ~n40615;
  assign n41762 = ~n40082 & ~n40085;
  assign n41763 = n40672 & n41762;
  assign n41764 = n41761 & ~n41763;
  assign n41765 = ~pi1151 & ~n39865;
  assign n41766 = n40192 & ~n41589;
  assign n41767 = n40680 & ~n41766;
  assign n41768 = ~n40178 & n40680;
  assign n41769 = ~n41767 & ~n41768;
  assign n41770 = n41765 & n41769;
  assign n41771 = n40500 & ~n41603;
  assign n41772 = ~pi1147 & ~n41771;
  assign n41773 = ~n41770 & n41772;
  assign n41774 = pi1149 & ~n41764;
  assign n41775 = ~n41773 & n41774;
  assign n41776 = pi1150 & ~n41775;
  assign n41777 = ~n41760 & n41776;
  assign n41778 = ~n40095 & n40141;
  assign n41779 = ~pi1151 & ~n41778;
  assign n41780 = ~pi1147 & ~n41779;
  assign n41781 = n39830 & ~n40533;
  assign n41782 = n41755 & ~n41781;
  assign n41783 = n41780 & ~n41782;
  assign n41784 = ~n40704 & n41745;
  assign n41785 = ~n40132 & n40577;
  assign n41786 = pi1147 & ~n41785;
  assign n41787 = ~n41784 & n41786;
  assign n41788 = ~pi1149 & ~n41783;
  assign n41789 = ~n41787 & n41788;
  assign n41790 = pi0212 & ~n39686;
  assign n41791 = n41517 & ~n41790;
  assign n41792 = n40164 & ~n41791;
  assign n41793 = n40593 & ~n41792;
  assign n41794 = pi1147 & ~n41793;
  assign n41795 = n38423 & ~n40173;
  assign n41796 = ~n40183 & n40653;
  assign n41797 = ~n41795 & n41796;
  assign n41798 = ~pi1151 & ~n40082;
  assign n41799 = ~n41797 & n41798;
  assign n41800 = ~n40198 & n41799;
  assign n41801 = n41794 & ~n41800;
  assign n41802 = n41765 & ~n41797;
  assign n41803 = ~n40514 & n41517;
  assign n41804 = n40269 & ~n41803;
  assign n41805 = ~n39865 & ~n41804;
  assign n41806 = pi1151 & n41805;
  assign n41807 = ~pi1147 & ~n41802;
  assign n41808 = ~n41806 & n41807;
  assign n41809 = pi1149 & ~n41808;
  assign n41810 = ~n41801 & n41809;
  assign n41811 = ~pi1150 & ~n41789;
  assign n41812 = ~n41810 & n41811;
  assign n41813 = ~n41777 & ~n41812;
  assign n41814 = pi1148 & ~n41813;
  assign n41815 = ~pi1151 & ~n40243;
  assign n41816 = ~pi1147 & ~n41815;
  assign n41817 = pi1151 & ~n40060;
  assign n41818 = n41816 & ~n41817;
  assign n41819 = ~n41577 & n41746;
  assign n41820 = n39870 & ~n41819;
  assign n41821 = ~n39869 & ~n41554;
  assign n41822 = ~pi1151 & n41821;
  assign n41823 = pi1147 & ~n41822;
  assign n41824 = ~n41820 & n41823;
  assign n41825 = pi1150 & ~n41818;
  assign n41826 = ~n41824 & n41825;
  assign n41827 = ~pi1147 & pi1151;
  assign n41828 = n40140 & n41827;
  assign n41829 = ~n39639 & n40664;
  assign n41830 = n40696 & ~n41829;
  assign n41831 = n39870 & ~n41830;
  assign n41832 = n40565 & ~n40665;
  assign n41833 = pi1147 & ~n41832;
  assign n41834 = ~n41831 & n41833;
  assign n41835 = ~pi1150 & ~n41828;
  assign n41836 = ~n41834 & n41835;
  assign n41837 = ~n41826 & ~n41836;
  assign n41838 = ~pi1149 & ~n41837;
  assign n41839 = ~pi1151 & ~n40208;
  assign n41840 = ~n40637 & n41839;
  assign n41841 = ~n40159 & n40269;
  assign n41842 = ~n40208 & ~n41841;
  assign n41843 = pi1151 & n41842;
  assign n41844 = ~pi1147 & ~n41840;
  assign n41845 = ~n41843 & n41844;
  assign n41846 = pi1147 & ~n40620;
  assign n41847 = ~pi1151 & ~n40146;
  assign n41848 = ~n40198 & n41847;
  assign n41849 = n41846 & ~n41848;
  assign n41850 = ~pi1150 & ~n41845;
  assign n41851 = ~n41849 & n41850;
  assign n41852 = n40548 & n40666;
  assign n41853 = pi1147 & ~n41852;
  assign n41854 = ~n40146 & ~n40197;
  assign n41855 = ~pi1151 & n41854;
  assign n41856 = n41853 & ~n41855;
  assign n41857 = ~n41767 & n41839;
  assign n41858 = pi1151 & ~n40208;
  assign n41859 = ~n40303 & n41858;
  assign n41860 = ~pi1147 & ~n41859;
  assign n41861 = ~n41857 & n41860;
  assign n41862 = pi1150 & ~n41856;
  assign n41863 = ~n41861 & n41862;
  assign n41864 = ~n41851 & ~n41863;
  assign n41865 = pi1149 & ~n41864;
  assign n41866 = ~pi1148 & ~n41838;
  assign n41867 = ~n41865 & n41866;
  assign n41868 = ~n41814 & ~n41867;
  assign n41869 = ~pi0213 & ~n41868;
  assign n41870 = pi0209 & ~n41744;
  assign n41871 = ~n41869 & n41870;
  assign n41872 = ~pi0213 & ~n40205;
  assign n41873 = ~n41767 & n41858;
  assign n41874 = pi1147 & ~n40672;
  assign n41875 = ~n41873 & n41874;
  assign n41876 = ~po1038 & ~n40711;
  assign n41877 = ~n40714 & n41876;
  assign n41878 = ~n40485 & ~n41877;
  assign n41879 = n41816 & n41878;
  assign n41880 = ~pi1150 & ~n41879;
  assign n41881 = ~n41875 & n41880;
  assign n41882 = n40500 & n41769;
  assign n41883 = n40523 & ~n41768;
  assign n41884 = pi1147 & ~n41883;
  assign n41885 = ~n41882 & n41884;
  assign n41886 = n40116 & n40123;
  assign n41887 = n40500 & ~n41886;
  assign n41888 = n41754 & ~n41887;
  assign n41889 = pi1150 & ~n41885;
  assign n41890 = ~n41888 & n41889;
  assign n41891 = ~n41881 & ~n41890;
  assign n41892 = ~pi1149 & ~n41891;
  assign n41893 = n40565 & ~n41819;
  assign n41894 = ~n40146 & ~n41578;
  assign n41895 = pi1151 & n41894;
  assign n41896 = ~pi1147 & ~n41895;
  assign n41897 = ~n41893 & n41896;
  assign n41898 = ~n40087 & n41832;
  assign n41899 = n41853 & ~n41898;
  assign n41900 = ~pi1150 & ~n41899;
  assign n41901 = ~n41897 & n41900;
  assign n41902 = ~n40131 & ~n40677;
  assign n41903 = ~pi1151 & n41902;
  assign n41904 = n41761 & ~n41903;
  assign n41905 = n40577 & ~n41746;
  assign n41906 = n40069 & ~n40315;
  assign n41907 = n40310 & ~n41906;
  assign n41908 = n40593 & ~n41907;
  assign n41909 = ~pi1147 & ~n41908;
  assign n41910 = ~n41905 & n41909;
  assign n41911 = pi1150 & ~n41904;
  assign n41912 = ~n41910 & n41911;
  assign n41913 = ~n41901 & ~n41912;
  assign n41914 = pi1149 & ~n41913;
  assign n41915 = pi1148 & ~n41914;
  assign n41916 = ~n41892 & n41915;
  assign n41917 = ~n16479 & n39864;
  assign n41918 = pi1151 & ~n41917;
  assign n41919 = n41780 & ~n41918;
  assign n41920 = n40500 & ~n41797;
  assign n41921 = n40185 & n40653;
  assign n41922 = ~n40096 & ~n41921;
  assign n41923 = ~pi1151 & n41922;
  assign n41924 = pi1147 & ~n41920;
  assign n41925 = ~n41923 & n41924;
  assign n41926 = pi1150 & ~n41919;
  assign n41927 = ~n41925 & n41926;
  assign n41928 = n40142 & n41827;
  assign n41929 = ~n40208 & ~n40637;
  assign n41930 = ~pi1151 & ~n41495;
  assign n41931 = pi1147 & ~n41930;
  assign n41932 = ~n41929 & n41931;
  assign n41933 = ~pi1150 & ~n41928;
  assign n41934 = ~n41932 & n41933;
  assign n41935 = ~n41927 & ~n41934;
  assign n41936 = ~pi1149 & ~n41935;
  assign n41937 = n39642 & n39830;
  assign n41938 = ~n10843 & n41937;
  assign n41939 = ~n41830 & ~n41938;
  assign n41940 = n40548 & n41939;
  assign n41941 = n40565 & ~n41830;
  assign n41942 = ~pi1147 & ~n41941;
  assign n41943 = ~n41940 & n41942;
  assign n41944 = ~pi0219 & ~n40531;
  assign n41945 = ~n40642 & n41944;
  assign n41946 = n40164 & ~n41945;
  assign n41947 = ~n40160 & n41946;
  assign n41948 = n40565 & ~n41947;
  assign n41949 = n41846 & ~n41948;
  assign n41950 = ~pi1150 & ~n41943;
  assign n41951 = ~n41949 & n41950;
  assign n41952 = n40593 & ~n41937;
  assign n41953 = ~n40704 & n41952;
  assign n41954 = n40577 & ~n40704;
  assign n41955 = ~pi1147 & ~n41953;
  assign n41956 = ~n41954 & n41955;
  assign n41957 = ~n40131 & ~n41946;
  assign n41958 = ~pi1151 & n41957;
  assign n41959 = n41794 & ~n41958;
  assign n41960 = pi1150 & ~n41956;
  assign n41961 = ~n41959 & n41960;
  assign n41962 = ~n41951 & ~n41961;
  assign n41963 = pi1149 & ~n41962;
  assign n41964 = ~pi1148 & ~n41936;
  assign n41965 = ~n41963 & n41964;
  assign n41966 = ~n41916 & ~n41965;
  assign n41967 = pi0213 & ~n41966;
  assign n41968 = ~pi0209 & ~n41872;
  assign n41969 = ~n41967 & n41968;
  assign n41970 = ~n41871 & ~n41969;
  assign n41971 = pi0230 & ~n41970;
  assign n41972 = ~pi0230 & ~pi0247;
  assign po0404 = ~n41971 & ~n41972;
  assign n41974 = ~pi1151 & ~n40142;
  assign n41975 = ~n40140 & n41974;
  assign n41976 = pi1152 & ~n41975;
  assign n41977 = ~n40610 & n41976;
  assign n41978 = pi1151 & ~pi1152;
  assign n41979 = ~n40125 & n41978;
  assign n41980 = ~pi1150 & ~n41977;
  assign n41981 = ~n41979 & n41980;
  assign n41982 = pi1151 & n40134;
  assign n41983 = ~pi1152 & ~n41982;
  assign n41984 = ~n40619 & n41983;
  assign n41985 = pi1152 & ~n40615;
  assign n41986 = ~n40165 & n41847;
  assign n41987 = n41985 & ~n41986;
  assign n41988 = pi1150 & ~n41984;
  assign n41989 = ~n41987 & n41988;
  assign n41990 = ~n41981 & ~n41989;
  assign n41991 = pi0213 & n41990;
  assign n41992 = pi1152 & ~n41954;
  assign n41993 = ~n41747 & n41992;
  assign n41994 = pi1151 & n41750;
  assign n41995 = ~pi1152 & ~n41785;
  assign n41996 = ~n41994 & n41995;
  assign n41997 = ~pi1150 & ~n41993;
  assign n41998 = ~n41996 & n41997;
  assign n41999 = ~n41792 & n41798;
  assign n42000 = n41985 & ~n41999;
  assign n42001 = pi1151 & ~n40127;
  assign n42002 = n41762 & n42001;
  assign n42003 = ~pi1152 & ~n42002;
  assign n42004 = ~n41800 & n42003;
  assign n42005 = pi1150 & ~n42004;
  assign n42006 = ~n42000 & n42005;
  assign n42007 = pi1148 & ~n41998;
  assign n42008 = ~n42006 & n42007;
  assign n42009 = ~n40124 & n41755;
  assign n42010 = ~pi1152 & ~n42009;
  assign n42011 = ~n41779 & n42010;
  assign n42012 = n40523 & ~n41781;
  assign n42013 = pi1152 & ~n42012;
  assign n42014 = ~n41757 & n42013;
  assign n42015 = ~pi1150 & ~n42014;
  assign n42016 = ~n42011 & n42015;
  assign n42017 = ~pi1151 & n41805;
  assign n42018 = pi1152 & ~n41771;
  assign n42019 = ~n42017 & n42018;
  assign n42020 = ~pi1152 & ~n41802;
  assign n42021 = ~n41882 & n42020;
  assign n42022 = pi1150 & ~n42019;
  assign n42023 = ~n42021 & n42022;
  assign n42024 = ~pi1148 & ~n42023;
  assign n42025 = ~n42016 & n42024;
  assign n42026 = ~n42008 & ~n42025;
  assign n42027 = pi1149 & ~n42026;
  assign n42028 = ~pi1152 & ~n41840;
  assign n42029 = ~n41873 & n42028;
  assign n42030 = ~pi1151 & n41842;
  assign n42031 = pi1152 & ~n41859;
  assign n42032 = ~n42030 & n42031;
  assign n42033 = pi1150 & ~n42029;
  assign n42034 = ~n42032 & n42033;
  assign n42035 = n40243 & n41978;
  assign n42036 = ~pi1151 & ~n40140;
  assign n42037 = pi1152 & ~n41817;
  assign n42038 = ~n42036 & n42037;
  assign n42039 = ~pi1150 & ~n42035;
  assign n42040 = ~n42038 & n42039;
  assign n42041 = ~n42034 & ~n42040;
  assign n42042 = ~pi1148 & ~n42041;
  assign n42043 = pi1152 & ~n41986;
  assign n42044 = ~n41852 & n42043;
  assign n42045 = pi1151 & n41854;
  assign n42046 = ~pi1152 & ~n41848;
  assign n42047 = ~n42045 & n42046;
  assign n42048 = ~n42044 & ~n42047;
  assign n42049 = pi1150 & ~n42048;
  assign n42050 = pi1151 & n41821;
  assign n42051 = ~n41832 & ~n42050;
  assign n42052 = ~pi1152 & ~n42051;
  assign n42053 = ~n41820 & ~n41941;
  assign n42054 = pi1152 & ~n42053;
  assign n42055 = ~pi1150 & ~n42052;
  assign n42056 = ~n42054 & n42055;
  assign n42057 = pi1148 & ~n42056;
  assign n42058 = ~n42049 & n42057;
  assign n42059 = ~pi1149 & ~n42042;
  assign n42060 = ~n42058 & n42059;
  assign n42061 = ~n42027 & ~n42060;
  assign n42062 = ~pi0213 & ~n42061;
  assign n42063 = pi0209 & ~n41991;
  assign n42064 = ~n42062 & n42063;
  assign n42065 = ~pi0213 & ~n41488;
  assign n42066 = n41778 & n41978;
  assign n42067 = pi1152 & ~n41918;
  assign n42068 = ~n41974 & n42067;
  assign n42069 = ~pi1150 & ~n42066;
  assign n42070 = ~n42068 & n42069;
  assign n42071 = ~pi1152 & ~n41941;
  assign n42072 = ~n41784 & n42071;
  assign n42073 = n41847 & n41939;
  assign n42074 = pi1152 & ~n41953;
  assign n42075 = ~n42073 & n42074;
  assign n42076 = pi1150 & ~n42072;
  assign n42077 = ~n42075 & n42076;
  assign n42078 = ~pi1149 & ~n42070;
  assign n42079 = ~n42077 & n42078;
  assign n42080 = ~pi1151 & n41894;
  assign n42081 = pi1152 & ~n41908;
  assign n42082 = ~n42080 & n42081;
  assign n42083 = ~pi1152 & ~n41747;
  assign n42084 = ~n41893 & n42083;
  assign n42085 = pi1150 & ~n42082;
  assign n42086 = ~n42084 & n42085;
  assign n42087 = ~n41815 & n42010;
  assign n42088 = ~pi1151 & ~n41878;
  assign n42089 = pi1152 & ~n42088;
  assign n42090 = ~n41887 & n42089;
  assign n42091 = ~pi1150 & ~n42090;
  assign n42092 = ~n42087 & n42091;
  assign n42093 = pi1149 & ~n42086;
  assign n42094 = ~n42092 & n42093;
  assign n42095 = ~pi1148 & ~n42079;
  assign n42096 = ~n42094 & n42095;
  assign n42097 = n41755 & ~n41768;
  assign n42098 = n40673 & ~n42097;
  assign n42099 = pi1152 & ~n41857;
  assign n42100 = ~n41882 & n42099;
  assign n42101 = ~pi1150 & ~n42098;
  assign n42102 = ~n42100 & n42101;
  assign n42103 = pi1151 & n41902;
  assign n42104 = ~pi1152 & ~n41898;
  assign n42105 = ~n42103 & n42104;
  assign n42106 = n40666 & n41847;
  assign n42107 = n41985 & ~n42106;
  assign n42108 = pi1150 & ~n42105;
  assign n42109 = ~n42107 & n42108;
  assign n42110 = pi1149 & ~n42109;
  assign n42111 = ~n42102 & n42110;
  assign n42112 = pi1151 & n41922;
  assign n42113 = ~pi1152 & ~n41930;
  assign n42114 = ~n42112 & n42113;
  assign n42115 = pi1152 & ~n41840;
  assign n42116 = ~n41920 & n42115;
  assign n42117 = ~pi1150 & ~n42116;
  assign n42118 = ~n42114 & n42117;
  assign n42119 = ~n41793 & n42043;
  assign n42120 = pi1151 & n41957;
  assign n42121 = ~pi1152 & ~n41948;
  assign n42122 = ~n42120 & n42121;
  assign n42123 = pi1150 & ~n42119;
  assign n42124 = ~n42122 & n42123;
  assign n42125 = ~pi1149 & ~n42118;
  assign n42126 = ~n42124 & n42125;
  assign n42127 = pi1148 & ~n42111;
  assign n42128 = ~n42126 & n42127;
  assign n42129 = pi0213 & ~n42096;
  assign n42130 = ~n42128 & n42129;
  assign n42131 = ~pi0209 & ~n42065;
  assign n42132 = ~n42130 & n42131;
  assign n42133 = ~n42064 & ~n42132;
  assign n42134 = pi0230 & ~n42133;
  assign n42135 = ~pi0230 & ~pi0248;
  assign po0405 = ~n42134 & ~n42135;
  assign n42137 = ~pi0213 & n41990;
  assign n42138 = pi0057 & ~n38886;
  assign n42139 = ~n6305 & n38886;
  assign n42140 = ~n39738 & n39882;
  assign n42141 = pi0299 & n38883;
  assign n42142 = ~n40682 & ~n42141;
  assign n42143 = ~pi0214 & ~n42142;
  assign n42144 = pi0212 & ~n42140;
  assign n42145 = ~n42143 & n42144;
  assign n42146 = pi0214 & ~n42142;
  assign n42147 = ~pi0212 & ~n39748;
  assign n42148 = ~n42146 & n42147;
  assign n42149 = ~pi0219 & ~n42145;
  assign n42150 = ~n42148 & n42149;
  assign n42151 = n6305 & ~n39768;
  assign n42152 = ~n42150 & n42151;
  assign n42153 = ~pi0057 & pi1151;
  assign n42154 = ~n42139 & n42153;
  assign n42155 = ~n42152 & n42154;
  assign n42156 = ~n40183 & ~n42141;
  assign n42157 = ~n39748 & n42156;
  assign n42158 = ~pi0212 & ~n42157;
  assign n42159 = ~pi0214 & n42156;
  assign n42160 = ~n39854 & ~n40182;
  assign n42161 = pi0214 & ~n40635;
  assign n42162 = ~n42160 & n42161;
  assign n42163 = pi0212 & ~n42162;
  assign n42164 = ~n42159 & n42163;
  assign n42165 = ~n42158 & ~n42164;
  assign n42166 = ~pi0219 & ~n42165;
  assign n42167 = n6305 & ~n40652;
  assign n42168 = ~n42166 & n42167;
  assign n42169 = ~pi0057 & ~pi1151;
  assign n42170 = ~n42139 & n42169;
  assign n42171 = ~n42168 & n42170;
  assign n42172 = ~n42138 & ~n42155;
  assign n42173 = ~n42171 & n42172;
  assign n42174 = ~pi1152 & ~n42173;
  assign n42175 = pi0299 & ~n38883;
  assign n42176 = ~n10843 & n42175;
  assign n42177 = ~n38917 & ~n42176;
  assign n42178 = n40083 & ~n42177;
  assign n42179 = n40660 & ~n42178;
  assign n42180 = ~n40195 & ~n40291;
  assign n42181 = pi1151 & ~n42180;
  assign n42182 = ~n42179 & n42181;
  assign n42183 = n40525 & ~n42141;
  assign n42184 = ~n39686 & ~n42141;
  assign n42185 = ~pi0214 & ~n42184;
  assign n42186 = n40149 & ~n40628;
  assign n42187 = pi0212 & ~n42185;
  assign n42188 = ~n42186 & n42187;
  assign n42189 = n41516 & ~n42183;
  assign n42190 = ~n42188 & n42189;
  assign n42191 = ~pi1151 & ~n42190;
  assign n42192 = n40164 & n42191;
  assign n42193 = n38922 & ~n42182;
  assign n42194 = ~n42192 & n42193;
  assign n42195 = pi1150 & ~n42194;
  assign n42196 = ~n42174 & n42195;
  assign n42197 = ~pi0212 & n39736;
  assign n42198 = n40062 & ~n42175;
  assign n42199 = pi0212 & ~n42198;
  assign n42200 = ~n40739 & n42199;
  assign n42201 = ~pi0219 & ~n42197;
  assign n42202 = ~n42183 & n42201;
  assign n42203 = ~n42200 & n42202;
  assign n42204 = n39694 & ~n40309;
  assign n42205 = ~n42203 & n42204;
  assign n42206 = ~pi1151 & n41830;
  assign n42207 = ~n39738 & ~n42176;
  assign n42208 = n38885 & n39635;
  assign n42209 = ~n42207 & n42208;
  assign n42210 = n38922 & ~n42209;
  assign n42211 = ~n42206 & n42210;
  assign n42212 = ~n42205 & n42211;
  assign n42213 = n10843 & n40713;
  assign n42214 = n39066 & ~n40100;
  assign n42215 = ~n38745 & n40110;
  assign n42216 = pi0211 & n40712;
  assign n42217 = n38608 & ~n42215;
  assign n42218 = ~n42216 & n42217;
  assign n42219 = ~n42213 & ~n42214;
  assign n42220 = ~n42218 & n42219;
  assign n42221 = ~pi0219 & ~n42220;
  assign n42222 = pi1151 & n40123;
  assign n42223 = ~n42221 & n42222;
  assign n42224 = n38888 & ~n42209;
  assign n42225 = ~n42223 & n42224;
  assign n42226 = ~pi1150 & ~n42212;
  assign n42227 = ~n42225 & n42226;
  assign n42228 = ~n42196 & ~n42227;
  assign n42229 = pi0213 & ~n42228;
  assign n42230 = ~pi0209 & ~n42229;
  assign n42231 = ~n42137 & n42230;
  assign n42232 = pi0213 & n39071;
  assign n42233 = ~n10484 & ~n39029;
  assign n42234 = n38675 & ~n39253;
  assign n42235 = pi0207 & ~n38769;
  assign n42236 = ~n39027 & n42235;
  assign n42237 = ~pi0207 & n39252;
  assign n42238 = pi0208 & ~n42236;
  assign n42239 = ~n42237 & n42238;
  assign n42240 = ~n42234 & ~n42239;
  assign n42241 = pi0211 & ~n42240;
  assign n42242 = pi0214 & n42241;
  assign n42243 = ~n42233 & ~n42242;
  assign n42244 = ~pi0212 & ~n42243;
  assign n42245 = ~pi0219 & ~n42244;
  assign n42246 = ~pi0211 & n42240;
  assign n42247 = ~n39099 & ~n42246;
  assign n42248 = pi0214 & ~n42247;
  assign n42249 = ~pi0211 & ~n39029;
  assign n42250 = ~pi0214 & ~n42249;
  assign n42251 = ~n42241 & n42250;
  assign n42252 = pi0212 & ~n42251;
  assign n42253 = ~n42248 & n42252;
  assign n42254 = n42245 & ~n42253;
  assign n42255 = n39031 & ~n42254;
  assign n42256 = n41755 & ~n42255;
  assign n42257 = ~n39029 & n39073;
  assign n42258 = ~n41978 & ~n42257;
  assign n42259 = ~n42256 & ~n42258;
  assign n42260 = ~n38966 & ~n39909;
  assign n42261 = ~n38968 & n39909;
  assign n42262 = ~po1038 & ~n42260;
  assign n42263 = ~n42261 & n42262;
  assign n42264 = n41839 & ~n42263;
  assign n42265 = pi0214 & n38953;
  assign n42266 = n39014 & ~n42265;
  assign n42267 = ~pi0219 & ~n42266;
  assign n42268 = pi0214 & ~n38968;
  assign n42269 = ~pi0214 & n38953;
  assign n42270 = pi0212 & ~n42269;
  assign n42271 = ~n42268 & n42270;
  assign n42272 = n42267 & ~n42271;
  assign n42273 = ~po1038 & ~n38971;
  assign n42274 = ~n42272 & n42273;
  assign n42275 = n40500 & ~n42274;
  assign n42276 = pi1152 & ~n42264;
  assign n42277 = ~n42275 & n42276;
  assign n42278 = ~n42259 & ~n42277;
  assign n42279 = ~pi1150 & ~n42278;
  assign n42280 = ~n38413 & n42247;
  assign n42281 = pi0219 & ~n39074;
  assign n42282 = ~n42280 & n42281;
  assign n42283 = ~po1038 & ~n42282;
  assign n42284 = pi0212 & ~n42243;
  assign n42285 = ~pi0212 & ~n39029;
  assign n42286 = ~pi0219 & ~n42285;
  assign n42287 = ~n42284 & n42286;
  assign n42288 = n42283 & ~n42287;
  assign n42289 = n40565 & ~n42288;
  assign n42290 = pi0214 & n42240;
  assign n42291 = n42252 & ~n42290;
  assign n42292 = n42245 & ~n42291;
  assign n42293 = n42283 & ~n42292;
  assign n42294 = n41745 & ~n42293;
  assign n42295 = ~pi1152 & ~n42289;
  assign n42296 = ~n42294 & n42295;
  assign n42297 = pi0212 & ~n38953;
  assign n42298 = n42267 & ~n42297;
  assign n42299 = n38974 & ~n42298;
  assign n42300 = n40593 & ~n42299;
  assign n42301 = ~n39013 & ~n42268;
  assign n42302 = ~pi0212 & ~n42301;
  assign n42303 = ~pi0211 & n38966;
  assign n42304 = ~n38992 & ~n42303;
  assign n42305 = pi0214 & ~n42304;
  assign n42306 = ~pi0214 & n38968;
  assign n42307 = pi0212 & ~n42305;
  assign n42308 = ~n42306 & n42307;
  assign n42309 = ~n42302 & ~n42308;
  assign n42310 = ~pi0219 & ~n42309;
  assign n42311 = n38974 & ~n42310;
  assign n42312 = n41847 & ~n42311;
  assign n42313 = pi1152 & ~n42300;
  assign n42314 = ~n42312 & n42313;
  assign n42315 = ~n42296 & ~n42314;
  assign n42316 = pi1150 & ~n42315;
  assign n42317 = ~n42279 & ~n42316;
  assign n42318 = ~pi0213 & ~n42317;
  assign n42319 = pi0209 & ~n42232;
  assign n42320 = ~n42318 & n42319;
  assign n42321 = ~n42231 & ~n42320;
  assign n42322 = pi0230 & ~n42321;
  assign n42323 = ~pi0230 & ~pi0249;
  assign po0406 = ~n42322 & ~n42323;
  assign n42325 = n2531 & n11513;
  assign n42326 = ~n6286 & ~n42325;
  assign n42327 = ~pi0075 & ~n42326;
  assign n42328 = n7333 & n8966;
  assign n42329 = ~n42327 & ~n42328;
  assign n42330 = ~pi0087 & ~pi0250;
  assign n42331 = n8881 & n42330;
  assign po0407 = ~n42329 & n42331;
  assign n42333 = pi0897 & n10809;
  assign n42334 = ~pi0476 & n11444;
  assign n42335 = ~n42333 & ~n42334;
  assign n42336 = ~pi0200 & pi1053;
  assign n42337 = pi0200 & pi1039;
  assign n42338 = ~pi0199 & ~n42336;
  assign n42339 = ~n42337 & n42338;
  assign n42340 = ~n42335 & ~n42339;
  assign n42341 = pi0251 & n42335;
  assign po0408 = n42340 | n42341;
  assign n42343 = ~n10983 & n11552;
  assign n42344 = ~n6198 & n11552;
  assign n42345 = ~pi0979 & ~pi0984;
  assign n42346 = pi1001 & n42345;
  assign n42347 = n6186 & n42346;
  assign n42348 = ~n6213 & n42347;
  assign n42349 = n6380 & n42348;
  assign n42350 = ~pi0252 & ~n42349;
  assign n42351 = pi1092 & ~pi1093;
  assign n42352 = ~n42350 & n42351;
  assign n42353 = n6392 & ~n42352;
  assign n42354 = n6391 & n42352;
  assign n42355 = ~n42353 & ~n42354;
  assign n42356 = n6198 & n42355;
  assign n42357 = ~n42344 & ~n42356;
  assign n42358 = n6242 & ~n42357;
  assign n42359 = ~n6227 & n42355;
  assign n42360 = n6227 & n11552;
  assign n42361 = ~n42359 & ~n42360;
  assign n42362 = ~n6242 & ~n42361;
  assign n42363 = pi0299 & ~n42358;
  assign n42364 = ~n42362 & n42363;
  assign n42365 = n6205 & ~n42357;
  assign n42366 = ~n6205 & ~n42361;
  assign n42367 = ~pi0299 & ~n42365;
  assign n42368 = ~n42366 & n42367;
  assign n42369 = n10983 & ~n42364;
  assign n42370 = ~n42368 & n42369;
  assign n42371 = ~n7643 & ~n42343;
  assign n42372 = ~n42370 & n42371;
  assign n42373 = pi0057 & n11551;
  assign n42374 = n10982 & n42347;
  assign n42375 = n21130 & n42374;
  assign n42376 = n6217 & n42375;
  assign n42377 = ~n38387 & n42376;
  assign n42378 = n6380 & n42377;
  assign n42379 = ~pi0252 & ~n42378;
  assign n42380 = ~pi0057 & pi1092;
  assign n42381 = ~n42379 & n42380;
  assign n42382 = n7643 & ~n42373;
  assign n42383 = ~n42381 & n42382;
  assign po0409 = ~n42372 & ~n42383;
  assign n42385 = ~n13061 & ~n38508;
  assign n42386 = ~n38700 & n42385;
  assign n42387 = ~po1038 & n42386;
  assign n42388 = pi0219 & n40080;
  assign n42389 = ~n42387 & ~n42388;
  assign n42390 = pi1153 & ~n42389;
  assign n42391 = ~pi1151 & ~n42390;
  assign n42392 = n10844 & n38684;
  assign n42393 = pi0211 & ~n38570;
  assign n42394 = ~n42392 & ~n42393;
  assign n42395 = ~n38545 & ~n38562;
  assign n42396 = n38519 & ~n42395;
  assign n42397 = ~po1038 & ~n42396;
  assign n42398 = n42394 & n42397;
  assign n42399 = ~n11446 & n39281;
  assign n42400 = pi1151 & ~n42399;
  assign n42401 = ~n42398 & n42400;
  assign n42402 = ~n42391 & ~n42401;
  assign n42403 = ~pi1152 & ~n42402;
  assign n42404 = n38519 & n39783;
  assign n42405 = ~pi1151 & ~n11447;
  assign n42406 = ~n38688 & n42405;
  assign n42407 = ~n42404 & n42406;
  assign n42408 = ~n11384 & ~n38508;
  assign n42409 = ~n38568 & ~n39854;
  assign n42410 = pi1153 & ~n42409;
  assign n42411 = pi1151 & n42408;
  assign n42412 = ~n42410 & n42411;
  assign n42413 = ~po1038 & ~n42412;
  assign n42414 = ~n42407 & n42413;
  assign n42415 = ~pi1151 & n10844;
  assign n42416 = ~n39280 & ~n42415;
  assign n42417 = po1038 & n42416;
  assign n42418 = pi1152 & ~n42417;
  assign n42419 = ~n42414 & n42418;
  assign n42420 = ~n42403 & ~n42419;
  assign n42421 = pi0230 & ~n42420;
  assign n42422 = ~pi0253 & ~pi1091;
  assign n42423 = po1038 & ~n42422;
  assign n42424 = pi0211 & pi1091;
  assign n42425 = pi1091 & ~pi1153;
  assign n42426 = pi0219 & n42425;
  assign n42427 = ~n42424 & ~n42426;
  assign n42428 = n42423 & n42427;
  assign n42429 = pi1091 & ~n42394;
  assign n42430 = ~pi1153 & ~n40915;
  assign n42431 = pi1153 & ~n40952;
  assign n42432 = n38519 & ~n42431;
  assign n42433 = ~n42430 & n42432;
  assign n42434 = ~n42429 & ~n42433;
  assign n42435 = pi0253 & ~n42434;
  assign n42436 = ~n13064 & ~n42410;
  assign n42437 = pi1091 & ~n42436;
  assign n42438 = ~pi0253 & ~n42437;
  assign n42439 = ~po1038 & ~n42438;
  assign n42440 = ~n42435 & n42439;
  assign n42441 = pi1151 & ~n42428;
  assign n42442 = ~n42440 & n42441;
  assign n42443 = pi0253 & ~pi1091;
  assign n42444 = pi0219 & pi1091;
  assign n42445 = ~n38497 & n42444;
  assign n42446 = n42423 & ~n42445;
  assign n42447 = pi0219 & n42446;
  assign n42448 = pi1091 & pi1153;
  assign n42449 = n42387 & n42448;
  assign n42450 = ~pi1151 & ~n42443;
  assign n42451 = ~n42449 & n42450;
  assign n42452 = ~n42447 & n42451;
  assign n42453 = ~n42442 & ~n42452;
  assign n42454 = ~pi1152 & ~n42453;
  assign n42455 = ~pi0211 & pi1091;
  assign n42456 = ~pi0219 & n42455;
  assign n42457 = n42446 & ~n42456;
  assign n42458 = n11446 & n40911;
  assign n42459 = ~n38688 & n42458;
  assign n42460 = ~pi1153 & ~n40943;
  assign n42461 = ~n38561 & n40911;
  assign n42462 = pi1153 & ~n42461;
  assign n42463 = n38519 & ~n42462;
  assign n42464 = ~n42460 & n42463;
  assign n42465 = pi0253 & ~n42459;
  assign n42466 = ~n42464 & n42465;
  assign n42467 = pi1091 & n39783;
  assign n42468 = pi1091 & n38545;
  assign n42469 = n38958 & n42468;
  assign n42470 = n38519 & ~n42469;
  assign n42471 = ~n42467 & n42470;
  assign n42472 = pi1091 & n38688;
  assign n42473 = pi0211 & ~n40965;
  assign n42474 = ~n42472 & n42473;
  assign n42475 = ~pi0253 & ~n42471;
  assign n42476 = ~n42474 & n42475;
  assign n42477 = ~n42466 & ~n42476;
  assign n42478 = ~n11446 & ~n38519;
  assign n42479 = ~n42443 & n42478;
  assign n42480 = ~n42472 & n42479;
  assign n42481 = n39635 & ~n42480;
  assign n42482 = ~n42477 & n42481;
  assign n42483 = n42409 & ~n42443;
  assign n42484 = ~n42425 & ~n42483;
  assign n42485 = n42408 & ~n42484;
  assign n42486 = ~po1038 & ~n42422;
  assign n42487 = ~n42485 & n42486;
  assign n42488 = ~n42446 & ~n42487;
  assign n42489 = pi1151 & ~n42488;
  assign n42490 = pi1152 & ~n42457;
  assign n42491 = ~n42489 & n42490;
  assign n42492 = ~n42482 & n42491;
  assign n42493 = ~n40910 & ~n42492;
  assign n42494 = ~n42454 & n42493;
  assign n42495 = n40988 & n41072;
  assign n42496 = pi1153 & ~n42495;
  assign n42497 = ~pi1153 & ~n41118;
  assign n42498 = ~pi0219 & ~n42497;
  assign n42499 = ~n42496 & n42498;
  assign n42500 = ~pi1153 & ~n41048;
  assign n42501 = ~n40987 & ~n41011;
  assign n42502 = ~pi0211 & n41044;
  assign n42503 = n42501 & ~n42502;
  assign n42504 = n41000 & ~n41008;
  assign n42505 = n42503 & n42504;
  assign n42506 = pi1153 & ~n42505;
  assign n42507 = pi0219 & ~n42500;
  assign n42508 = ~n42506 & n42507;
  assign n42509 = pi0253 & ~n42499;
  assign n42510 = ~n42508 & n42509;
  assign n42511 = ~n40993 & n41048;
  assign n42512 = ~pi0211 & n42511;
  assign n42513 = ~n41013 & ~n42512;
  assign n42514 = pi1153 & ~n42513;
  assign n42515 = ~n41039 & ~n42514;
  assign n42516 = pi0219 & n42515;
  assign n42517 = ~pi1153 & n41116;
  assign n42518 = pi1153 & n41097;
  assign n42519 = ~pi0219 & ~n42517;
  assign n42520 = ~n42518 & n42519;
  assign n42521 = ~pi0253 & ~n42520;
  assign n42522 = ~n42516 & n42521;
  assign n42523 = ~n42510 & ~n42522;
  assign n42524 = ~po1038 & ~n42523;
  assign n42525 = ~pi0219 & ~n40980;
  assign n42526 = ~pi0211 & ~n40890;
  assign n42527 = n42525 & ~n42526;
  assign n42528 = ~pi0219 & ~n42527;
  assign n42529 = po1038 & n42528;
  assign n42530 = ~n40874 & n42529;
  assign n42531 = ~n40868 & ~n42445;
  assign n42532 = ~n42525 & n42531;
  assign n42533 = pi0253 & ~n42532;
  assign n42534 = ~pi0219 & ~n40890;
  assign n42535 = pi0211 & n40868;
  assign n42536 = ~pi0211 & ~n40874;
  assign n42537 = pi0219 & ~n42535;
  assign n42538 = ~n42536 & n42537;
  assign n42539 = ~n42445 & ~n42534;
  assign n42540 = ~n42538 & n42539;
  assign n42541 = ~pi0253 & ~n42540;
  assign n42542 = po1038 & ~n42533;
  assign n42543 = ~n42541 & n42542;
  assign n42544 = pi1151 & ~n42530;
  assign n42545 = ~n42543 & n42544;
  assign n42546 = ~n42524 & n42545;
  assign n42547 = ~n41072 & ~n42512;
  assign n42548 = n42525 & ~n42547;
  assign n42549 = ~n40987 & ~n40999;
  assign n42550 = ~pi1153 & ~n42549;
  assign n42551 = ~n41102 & ~n42550;
  assign n42552 = n42548 & ~n42551;
  assign n42553 = pi0219 & n41009;
  assign n42554 = ~n41057 & n42506;
  assign n42555 = n42553 & ~n42554;
  assign n42556 = ~n42552 & ~n42555;
  assign n42557 = pi0253 & ~n42556;
  assign n42558 = ~n41012 & n42503;
  assign n42559 = ~n42550 & n42558;
  assign n42560 = ~pi0219 & ~n42559;
  assign n42561 = pi0219 & n41011;
  assign n42562 = ~n42560 & ~n42561;
  assign n42563 = ~n42516 & n42562;
  assign n42564 = ~pi0253 & ~n42563;
  assign n42565 = ~po1038 & ~n42557;
  assign n42566 = ~n42564 & n42565;
  assign n42567 = ~pi1151 & ~n42566;
  assign n42568 = ~n42546 & ~n42567;
  assign n42569 = n42534 & ~n42536;
  assign n42570 = n42525 & ~n42569;
  assign n42571 = pi0219 & ~n40874;
  assign n42572 = po1038 & ~n42571;
  assign n42573 = ~n42570 & n42572;
  assign n42574 = ~n40874 & n42573;
  assign n42575 = ~n42543 & ~n42574;
  assign n42576 = ~n42568 & n42575;
  assign n42577 = pi1152 & ~n42576;
  assign n42578 = pi0219 & ~n42515;
  assign n42579 = ~n42520 & n42548;
  assign n42580 = ~n42578 & ~n42579;
  assign n42581 = ~n40993 & ~n42580;
  assign n42582 = ~pi0253 & ~n42581;
  assign n42583 = pi1153 & ~n40988;
  assign n42584 = n42503 & n42525;
  assign n42585 = ~n42583 & n42584;
  assign n42586 = ~pi1153 & ~n41028;
  assign n42587 = ~n41062 & ~n42505;
  assign n42588 = pi1153 & n42587;
  assign n42589 = pi0219 & ~n42586;
  assign n42590 = ~n42588 & n42589;
  assign n42591 = ~n42585 & ~n42590;
  assign n42592 = pi0253 & ~n42591;
  assign n42593 = ~po1038 & ~n42592;
  assign n42594 = ~n42582 & n42593;
  assign n42595 = n42545 & ~n42594;
  assign n42596 = ~pi1091 & ~n41039;
  assign n42597 = ~pi1153 & ~n42596;
  assign n42598 = ~n41057 & ~n42505;
  assign n42599 = ~pi0219 & n42549;
  assign n42600 = ~n42597 & ~n42599;
  assign n42601 = n42598 & n42600;
  assign n42602 = pi0253 & ~n42601;
  assign n42603 = ~n41002 & n42578;
  assign n42604 = ~pi1153 & ~n41084;
  assign n42605 = ~n40993 & ~n42604;
  assign n42606 = ~pi0219 & n41118;
  assign n42607 = n42605 & n42606;
  assign n42608 = ~pi0253 & ~n42607;
  assign n42609 = ~n42603 & n42608;
  assign n42610 = ~po1038 & ~n42602;
  assign n42611 = ~n42609 & n42610;
  assign n42612 = ~pi1151 & ~n42543;
  assign n42613 = ~n42611 & n42612;
  assign n42614 = ~pi1152 & ~n42613;
  assign n42615 = ~n42595 & n42614;
  assign n42616 = ~n42577 & ~n42615;
  assign n42617 = n40910 & ~n42616;
  assign n42618 = ~pi0230 & ~n42494;
  assign n42619 = ~n42617 & n42618;
  assign po0410 = ~n42421 & ~n42619;
  assign n42621 = ~pi0219 & ~n38882;
  assign n42622 = ~n39145 & ~n42621;
  assign n42623 = po1038 & n42622;
  assign n42624 = pi1154 & n38977;
  assign n42625 = ~n39033 & ~n42624;
  assign n42626 = n11446 & ~n42625;
  assign n42627 = pi0299 & n38519;
  assign n42628 = ~n11446 & n38959;
  assign n42629 = ~n42627 & ~n42628;
  assign n42630 = ~n38939 & ~n42629;
  assign n42631 = ~n42626 & ~n42630;
  assign n42632 = ~po1038 & ~n42631;
  assign n42633 = ~pi1152 & ~n42623;
  assign n42634 = ~n42632 & n42633;
  assign n42635 = n11446 & ~n38882;
  assign n42636 = n40028 & ~n42635;
  assign n42637 = ~pi0200 & pi1154;
  assign n42638 = n11373 & ~n42637;
  assign n42639 = n38976 & ~n39854;
  assign n42640 = ~n42638 & ~n42639;
  assign n42641 = ~pi0219 & ~n42640;
  assign n42642 = ~n38558 & ~n38976;
  assign n42643 = n38488 & ~n42642;
  assign n42644 = ~pi1154 & ~n39022;
  assign n42645 = ~n38941 & ~n42644;
  assign n42646 = ~n42643 & n42645;
  assign n42647 = pi0219 & ~n42646;
  assign n42648 = ~po1038 & ~n42641;
  assign n42649 = ~n42647 & n42648;
  assign n42650 = pi1152 & ~n42636;
  assign n42651 = ~n42649 & n42650;
  assign n42652 = ~n42634 & ~n42651;
  assign n42653 = pi0230 & ~n42652;
  assign n42654 = ~pi0254 & ~pi1091;
  assign n42655 = pi1091 & ~n42622;
  assign n42656 = po1038 & ~n42654;
  assign n42657 = ~n42655 & n42656;
  assign n42658 = po1038 & n42456;
  assign n42659 = ~n42657 & ~n42658;
  assign n42660 = pi1153 & ~n40932;
  assign n42661 = ~pi1154 & ~n42660;
  assign n42662 = ~pi0211 & n38683;
  assign n42663 = ~n42430 & n42661;
  assign n42664 = ~n42662 & n42663;
  assign n42665 = pi1091 & n38488;
  assign n42666 = ~n38568 & n42665;
  assign n42667 = ~n39045 & n42666;
  assign n42668 = ~n42664 & ~n42667;
  assign n42669 = ~pi0219 & ~n42668;
  assign n42670 = pi1154 & n42455;
  assign n42671 = ~n42444 & ~n42670;
  assign n42672 = ~n42646 & ~n42671;
  assign n42673 = ~n42669 & ~n42672;
  assign n42674 = pi0254 & ~n42673;
  assign n42675 = pi1154 & ~n42409;
  assign n42676 = pi0219 & ~n39022;
  assign n42677 = ~n42675 & n42676;
  assign n42678 = ~n42641 & ~n42677;
  assign n42679 = ~pi0254 & ~n42678;
  assign n42680 = ~n42654 & ~n42679;
  assign n42681 = ~n42674 & n42680;
  assign n42682 = ~po1038 & n42681;
  assign n42683 = pi1152 & n42659;
  assign n42684 = ~n42682 & n42683;
  assign n42685 = n40918 & n42425;
  assign n42686 = ~n42467 & ~n42685;
  assign n42687 = pi0211 & ~n42661;
  assign n42688 = ~n42686 & n42687;
  assign n42689 = n11445 & n42448;
  assign n42690 = ~pi1154 & ~n42689;
  assign n42691 = pi1091 & n38959;
  assign n42692 = pi1154 & ~n42691;
  assign n42693 = ~pi0211 & ~n42690;
  assign n42694 = ~n42692 & n42693;
  assign n42695 = ~n42688 & ~n42694;
  assign n42696 = ~pi0219 & ~n42695;
  assign n42697 = pi0211 & n42692;
  assign n42698 = pi1091 & n39666;
  assign n42699 = n38495 & ~n42698;
  assign n42700 = ~n42467 & n42699;
  assign n42701 = pi0219 & ~n42690;
  assign n42702 = ~n42700 & n42701;
  assign n42703 = ~n42697 & n42702;
  assign n42704 = ~n42696 & ~n42703;
  assign n42705 = ~pi0254 & ~n42704;
  assign n42706 = ~pi1153 & ~n40919;
  assign n42707 = ~n42462 & ~n42706;
  assign n42708 = pi1091 & ~pi1154;
  assign n42709 = n38533 & n42708;
  assign n42710 = ~n42707 & ~n42709;
  assign n42711 = n11446 & ~n42710;
  assign n42712 = pi1091 & ~n11446;
  assign n42713 = ~n38938 & n42712;
  assign n42714 = ~pi1154 & ~n42713;
  assign n42715 = n40968 & n42463;
  assign n42716 = pi1091 & ~n38641;
  assign n42717 = ~n42707 & ~n42716;
  assign n42718 = n42478 & ~n42717;
  assign n42719 = pi1154 & ~n42715;
  assign n42720 = ~n42718 & n42719;
  assign n42721 = ~n42714 & ~n42720;
  assign n42722 = pi0254 & ~n42711;
  assign n42723 = ~n42721 & n42722;
  assign n42724 = ~n42705 & ~n42723;
  assign n42725 = ~po1038 & ~n42724;
  assign n42726 = ~pi1152 & ~n42657;
  assign n42727 = ~n42725 & n42726;
  assign n42728 = ~n40910 & ~n42684;
  assign n42729 = ~n42727 & n42728;
  assign n42730 = pi1091 & n39145;
  assign n42731 = ~pi0211 & ~n40866;
  assign n42732 = n42571 & ~n42731;
  assign n42733 = ~pi0219 & n40890;
  assign n42734 = ~n42732 & ~n42733;
  assign n42735 = n11446 & n42425;
  assign n42736 = pi0254 & ~n42735;
  assign n42737 = ~n42730 & n42736;
  assign n42738 = n42734 & n42737;
  assign n42739 = ~n42448 & n42569;
  assign n42740 = ~pi0254 & ~n42730;
  assign n42741 = ~n42538 & n42740;
  assign n42742 = ~n42739 & n42741;
  assign n42743 = pi0253 & ~n42738;
  assign n42744 = ~n42742 & n42743;
  assign n42745 = pi0253 & po1038;
  assign n42746 = n42659 & ~n42745;
  assign n42747 = ~n42744 & ~n42746;
  assign n42748 = ~pi0253 & ~n42681;
  assign n42749 = pi1154 & ~n40985;
  assign n42750 = n42503 & n42749;
  assign n42751 = ~n42496 & n42750;
  assign n42752 = ~pi1153 & n42559;
  assign n42753 = ~n41118 & ~n42752;
  assign n42754 = ~pi1154 & ~n42753;
  assign n42755 = pi0254 & ~n42751;
  assign n42756 = ~n42754 & n42755;
  assign n42757 = pi0211 & n41044;
  assign n42758 = ~n40993 & ~n42757;
  assign n42759 = ~pi1153 & ~n42758;
  assign n42760 = ~n41012 & n41028;
  assign n42761 = pi1154 & n42760;
  assign n42762 = ~n41116 & ~n42761;
  assign n42763 = ~pi0254 & ~n42759;
  assign n42764 = ~n42762 & n42763;
  assign n42765 = ~n42756 & ~n42764;
  assign n42766 = ~pi0219 & ~n42765;
  assign n42767 = pi1154 & ~n42506;
  assign n42768 = ~n42587 & n42767;
  assign n42769 = pi1153 & ~n41048;
  assign n42770 = ~pi1154 & ~n42586;
  assign n42771 = ~n42769 & n42770;
  assign n42772 = pi0254 & ~n42771;
  assign n42773 = ~n42768 & n42772;
  assign n42774 = ~n42500 & n42760;
  assign n42775 = n38495 & ~n42774;
  assign n42776 = ~n40990 & n42775;
  assign n42777 = ~pi1153 & ~n41032;
  assign n42778 = n41041 & ~n42777;
  assign n42779 = ~pi1154 & ~n42778;
  assign n42780 = ~n40993 & n41039;
  assign n42781 = n42779 & ~n42780;
  assign n42782 = pi1153 & n41013;
  assign n42783 = n38488 & ~n40995;
  assign n42784 = ~n42782 & n42783;
  assign n42785 = ~pi0254 & ~n42784;
  assign n42786 = ~n42776 & n42785;
  assign n42787 = ~n42781 & n42786;
  assign n42788 = ~n42773 & ~n42787;
  assign n42789 = pi0219 & ~n42788;
  assign n42790 = pi0253 & ~n42789;
  assign n42791 = ~n42766 & n42790;
  assign n42792 = ~po1038 & ~n42748;
  assign n42793 = ~n42791 & n42792;
  assign n42794 = pi1152 & ~n42747;
  assign n42795 = ~n42793 & n42794;
  assign n42796 = ~n42657 & ~n42745;
  assign n42797 = ~n42570 & n42738;
  assign n42798 = ~n42528 & n42742;
  assign n42799 = pi0253 & ~n42797;
  assign n42800 = ~n42798 & n42799;
  assign n42801 = ~n42796 & ~n42800;
  assign n42802 = ~pi0253 & n42724;
  assign n42803 = n38495 & ~n41057;
  assign n42804 = ~pi1153 & n41000;
  assign n42805 = ~pi1154 & ~n41003;
  assign n42806 = ~pi1154 & ~n42805;
  assign n42807 = ~n42504 & ~n42804;
  assign n42808 = ~n42806 & n42807;
  assign n42809 = pi0219 & ~n42803;
  assign n42810 = ~n42808 & n42809;
  assign n42811 = pi1154 & n40999;
  assign n42812 = n42547 & ~n42804;
  assign n42813 = ~pi0219 & ~n42811;
  assign n42814 = ~n42812 & n42813;
  assign n42815 = ~n42810 & ~n42814;
  assign n42816 = pi0254 & ~n42815;
  assign n42817 = n41014 & ~n42500;
  assign n42818 = n38488 & ~n42817;
  assign n42819 = pi0219 & ~n42775;
  assign n42820 = ~n42779 & n42819;
  assign n42821 = ~n42818 & n42820;
  assign n42822 = pi1154 & n41011;
  assign n42823 = ~n41044 & ~n42822;
  assign n42824 = ~pi0211 & ~n42823;
  assign n42825 = ~n40985 & n41116;
  assign n42826 = ~n42604 & n42825;
  assign n42827 = ~pi1154 & ~n42826;
  assign n42828 = ~n40993 & n41118;
  assign n42829 = pi1154 & ~n42828;
  assign n42830 = ~n42826 & n42829;
  assign n42831 = ~pi0219 & ~n42824;
  assign n42832 = ~n42827 & n42831;
  assign n42833 = ~n42830 & n42832;
  assign n42834 = ~pi0254 & ~n42833;
  assign n42835 = ~n42821 & n42834;
  assign n42836 = ~n42816 & ~n42835;
  assign n42837 = pi0253 & ~n42836;
  assign n42838 = ~po1038 & ~n42802;
  assign n42839 = ~n42837 & n42838;
  assign n42840 = ~pi1152 & ~n42801;
  assign n42841 = ~n42839 & n42840;
  assign n42842 = n40910 & ~n42841;
  assign n42843 = ~n42795 & n42842;
  assign n42844 = ~pi0230 & ~n42729;
  assign n42845 = ~n42843 & n42844;
  assign po0411 = ~n42653 & ~n42845;
  assign n42847 = ~pi0200 & pi1049;
  assign n42848 = pi0200 & pi1036;
  assign n42849 = ~n42847 & ~n42848;
  assign n42850 = ~n42335 & n42849;
  assign n42851 = ~pi0255 & n42335;
  assign po0412 = ~n42850 & ~n42851;
  assign n42853 = ~pi0200 & pi1048;
  assign n42854 = pi0200 & pi1070;
  assign n42855 = ~n42853 & ~n42854;
  assign n42856 = ~n42335 & n42855;
  assign n42857 = ~pi0256 & n42335;
  assign po0413 = ~n42856 & ~n42857;
  assign n42859 = ~pi0200 & pi1084;
  assign n42860 = pi0200 & pi1065;
  assign n42861 = ~n42859 & ~n42860;
  assign n42862 = ~n42335 & n42861;
  assign n42863 = ~pi0257 & n42335;
  assign po0414 = ~n42862 & ~n42863;
  assign n42865 = ~pi0200 & pi1072;
  assign n42866 = pi0200 & pi1062;
  assign n42867 = ~n42865 & ~n42866;
  assign n42868 = ~n42335 & n42867;
  assign n42869 = ~pi0258 & n42335;
  assign po0415 = ~n42868 & ~n42869;
  assign n42871 = ~pi0200 & pi1059;
  assign n42872 = pi0200 & pi1069;
  assign n42873 = ~n42871 & ~n42872;
  assign n42874 = ~n42335 & n42873;
  assign n42875 = ~pi0259 & n42335;
  assign po0416 = ~n42874 & ~n42875;
  assign n42877 = ~pi0200 & pi1044;
  assign n42878 = pi0200 & pi1067;
  assign n42879 = ~pi0199 & ~n42877;
  assign n42880 = ~n42878 & n42879;
  assign n42881 = ~n42335 & ~n42880;
  assign n42882 = pi0260 & n42335;
  assign po0417 = n42881 | n42882;
  assign n42884 = ~pi0200 & pi1037;
  assign n42885 = pi0200 & pi1040;
  assign n42886 = ~pi0199 & ~n42884;
  assign n42887 = ~n42885 & n42886;
  assign n42888 = ~n42335 & ~n42887;
  assign n42889 = pi0261 & n42335;
  assign po0418 = n42888 | n42889;
  assign n42891 = pi1093 & pi1142;
  assign n42892 = ~pi0262 & ~pi1093;
  assign n42893 = ~n42891 & ~n42892;
  assign n42894 = ~pi0228 & ~n42893;
  assign n42895 = ~pi0123 & ~pi1142;
  assign n42896 = pi0123 & pi0262;
  assign n42897 = pi0228 & ~n42895;
  assign n42898 = ~n42896 & n42897;
  assign n42899 = ~n42894 & ~n42898;
  assign n42900 = ~pi0228 & ~pi1093;
  assign n42901 = pi0123 & pi0228;
  assign n42902 = ~n42900 & ~n42901;
  assign n42903 = ~pi0262 & ~n42902;
  assign n42904 = ~n40700 & ~n42903;
  assign n42905 = pi0199 & n42902;
  assign n42906 = n38441 & ~n42905;
  assign n42907 = n42904 & ~n42906;
  assign n42908 = ~n42899 & ~n42907;
  assign n42909 = ~pi0207 & n42903;
  assign n42910 = ~pi0208 & ~n42909;
  assign n42911 = ~n40700 & ~n42910;
  assign n42912 = ~n42908 & ~n42911;
  assign n42913 = ~n39711 & n42902;
  assign n42914 = ~pi0299 & ~n42913;
  assign n42915 = ~n42899 & n42914;
  assign n42916 = pi0299 & ~n42904;
  assign n42917 = pi0208 & ~n42915;
  assign n42918 = ~n42916 & n42917;
  assign n42919 = ~po1038 & ~n42918;
  assign n42920 = ~n42912 & n42919;
  assign n42921 = ~n39864 & n42902;
  assign n42922 = po1038 & ~n42899;
  assign n42923 = ~n42921 & n42922;
  assign po0419 = n42920 | n42923;
  assign n42925 = ~n40915 & ~n42708;
  assign n42926 = ~pi1156 & ~n38577;
  assign n42927 = ~n42925 & n42926;
  assign n42928 = pi1155 & ~n38985;
  assign n42929 = n40952 & ~n42928;
  assign n42930 = ~pi1154 & n42716;
  assign n42931 = ~n42929 & ~n42930;
  assign n42932 = ~n40965 & n42931;
  assign n42933 = n38479 & ~n42932;
  assign n42934 = ~pi1154 & ~n38702;
  assign n42935 = n38545 & ~n38576;
  assign n42936 = pi1154 & ~n42935;
  assign n42937 = pi1091 & n38483;
  assign n42938 = ~n42936 & n42937;
  assign n42939 = ~n42934 & n42938;
  assign n42940 = pi0219 & ~n42927;
  assign n42941 = ~n42939 & n42940;
  assign n42942 = ~n42933 & n42941;
  assign n42943 = ~pi0211 & ~n42931;
  assign n42944 = n38568 & ~n39111;
  assign n42945 = n42424 & ~n42944;
  assign n42946 = ~n38766 & n42945;
  assign n42947 = ~n42943 & ~n42946;
  assign n42948 = pi1156 & ~n42947;
  assign n42949 = ~n38766 & ~n42925;
  assign n42950 = pi0211 & n42949;
  assign n42951 = ~n38577 & ~n39000;
  assign n42952 = n42455 & n42951;
  assign n42953 = ~n42950 & ~n42952;
  assign n42954 = ~pi1156 & ~n42953;
  assign n42955 = ~pi0219 & ~n42954;
  assign n42956 = ~n42948 & n42955;
  assign n42957 = ~n42942 & ~n42956;
  assign n42958 = ~pi0263 & ~n42957;
  assign n42959 = ~pi1154 & n38646;
  assign n42960 = pi1154 & ~n38591;
  assign n42961 = pi1156 & ~n42960;
  assign n42962 = ~pi0299 & ~n42961;
  assign n42963 = ~n39854 & ~n42959;
  assign n42964 = ~n42962 & n42963;
  assign n42965 = pi1156 & ~n42964;
  assign n42966 = ~n42951 & n42962;
  assign n42967 = pi0219 & ~n42966;
  assign n42968 = ~n42965 & n42967;
  assign n42969 = ~n38648 & n39499;
  assign n42970 = ~n39000 & ~n42969;
  assign n42971 = ~pi0211 & ~n42970;
  assign n42972 = ~pi1156 & n42949;
  assign n42973 = ~n38568 & ~n38595;
  assign n42974 = pi1154 & ~n42973;
  assign n42975 = ~n38544 & n42934;
  assign n42976 = pi1156 & ~n42974;
  assign n42977 = ~n42975 & n42976;
  assign n42978 = pi0211 & ~n42972;
  assign n42979 = ~n42977 & n42978;
  assign n42980 = ~pi0219 & ~n42971;
  assign n42981 = ~n42979 & n42980;
  assign n42982 = pi0263 & pi1091;
  assign n42983 = ~n42968 & n42982;
  assign n42984 = ~n42981 & n42983;
  assign n42985 = ~n42958 & ~n42984;
  assign n42986 = ~po1038 & n42985;
  assign n42987 = pi0219 & ~n38483;
  assign n42988 = ~pi0219 & ~n38484;
  assign n42989 = ~n38495 & n42988;
  assign n42990 = ~n42987 & ~n42989;
  assign n42991 = pi1091 & ~n42990;
  assign n42992 = pi0263 & ~pi1091;
  assign n42993 = ~n42991 & ~n42992;
  assign n42994 = po1038 & ~n42993;
  assign n42995 = ~n40910 & ~n42994;
  assign n42996 = ~n42986 & n42995;
  assign n42997 = pi1091 & n42987;
  assign n42998 = pi0211 & n40874;
  assign n42999 = ~pi0211 & ~n42708;
  assign n43000 = ~n38484 & ~n42999;
  assign n43001 = ~n42998 & n43000;
  assign n43002 = ~n40890 & ~n43001;
  assign n43003 = ~pi0219 & ~n43002;
  assign n43004 = ~pi0263 & ~n42732;
  assign n43005 = ~n43003 & n43004;
  assign n43006 = ~n38484 & ~n42670;
  assign n43007 = ~n42998 & ~n43006;
  assign n43008 = n42534 & ~n43007;
  assign n43009 = pi0263 & ~n42538;
  assign n43010 = ~n43008 & n43009;
  assign n43011 = ~n43005 & ~n43010;
  assign n43012 = n40860 & ~n42997;
  assign n43013 = ~n43011 & n43012;
  assign n43014 = ~n40860 & n42993;
  assign n43015 = po1038 & ~n43014;
  assign n43016 = ~n43013 & n43015;
  assign n43017 = ~n40860 & ~n42985;
  assign n43018 = pi1155 & ~n41118;
  assign n43019 = pi1154 & ~n43018;
  assign n43020 = n41105 & n43019;
  assign n43021 = ~pi1155 & n42596;
  assign n43022 = pi1155 & ~n41009;
  assign n43023 = ~pi1154 & ~n43022;
  assign n43024 = ~n43021 & n43023;
  assign n43025 = ~n41116 & n43021;
  assign n43026 = pi1155 & ~n41072;
  assign n43027 = ~pi1154 & ~n43026;
  assign n43028 = ~n43025 & n43027;
  assign n43029 = ~pi1156 & ~n43028;
  assign n43030 = ~n43020 & ~n43024;
  assign n43031 = n43029 & n43030;
  assign n43032 = ~pi1155 & n41000;
  assign n43033 = ~n41044 & n41102;
  assign n43034 = ~n43032 & ~n43033;
  assign n43035 = ~pi1154 & ~n43034;
  assign n43036 = pi1156 & ~n43035;
  assign n43037 = n41000 & n43023;
  assign n43038 = ~n40983 & n43020;
  assign n43039 = ~n43037 & ~n43038;
  assign n43040 = n43036 & n43039;
  assign n43041 = ~pi0211 & ~n43031;
  assign n43042 = ~n43040 & n43041;
  assign n43043 = n40988 & n43019;
  assign n43044 = n43036 & ~n43043;
  assign n43045 = n42501 & n43019;
  assign n43046 = n43029 & ~n43045;
  assign n43047 = pi0211 & ~n43044;
  assign n43048 = ~n43046 & n43047;
  assign n43049 = ~pi0219 & ~n43042;
  assign n43050 = ~n43048 & n43049;
  assign n43051 = pi1155 & n41008;
  assign n43052 = pi1154 & n41028;
  assign n43053 = ~n43051 & n43052;
  assign n43054 = ~n40985 & n43053;
  assign n43055 = ~n43037 & ~n43054;
  assign n43056 = n38479 & ~n43055;
  assign n43057 = ~n43024 & ~n43053;
  assign n43058 = ~pi1156 & ~n43057;
  assign n43059 = ~pi1154 & n41039;
  assign n43060 = ~n41062 & ~n43059;
  assign n43061 = n38483 & ~n43051;
  assign n43062 = ~n43060 & n43061;
  assign n43063 = pi0219 & ~n43062;
  assign n43064 = ~n43056 & n43063;
  assign n43065 = ~n43058 & n43064;
  assign n43066 = ~pi0263 & ~n43065;
  assign n43067 = ~n43050 & n43066;
  assign n43068 = ~n41040 & ~n41055;
  assign n43069 = pi1154 & ~n43068;
  assign n43070 = pi1155 & ~n42760;
  assign n43071 = ~pi1155 & ~n42511;
  assign n43072 = ~pi1154 & ~n43070;
  assign n43073 = ~n43071 & n43072;
  assign n43074 = n38483 & ~n43069;
  assign n43075 = ~n43073 & n43074;
  assign n43076 = ~n41014 & ~n42822;
  assign n43077 = ~n43068 & ~n43076;
  assign n43078 = n38479 & ~n43077;
  assign n43079 = ~n41026 & n43077;
  assign n43080 = ~pi1156 & ~n43079;
  assign n43081 = pi0219 & ~n43075;
  assign n43082 = ~n43078 & n43081;
  assign n43083 = ~n43080 & n43082;
  assign n43084 = pi1154 & ~n41098;
  assign n43085 = ~n41046 & n43084;
  assign n43086 = ~pi1154 & ~n41085;
  assign n43087 = pi1155 & n42825;
  assign n43088 = n43086 & ~n43087;
  assign n43089 = ~n41114 & n43084;
  assign n43090 = ~pi1156 & ~n42811;
  assign n43091 = ~n43089 & n43090;
  assign n43092 = ~pi1156 & ~n43091;
  assign n43093 = ~n43088 & ~n43092;
  assign n43094 = pi1156 & n42828;
  assign n43095 = ~n43093 & ~n43094;
  assign n43096 = ~n43085 & ~n43095;
  assign n43097 = pi0211 & ~n43096;
  assign n43098 = ~n41026 & n41091;
  assign n43099 = pi1155 & n43098;
  assign n43100 = n43086 & ~n43099;
  assign n43101 = ~n42828 & n43100;
  assign n43102 = pi1156 & ~n43101;
  assign n43103 = ~n43089 & n43102;
  assign n43104 = n43091 & ~n43100;
  assign n43105 = ~pi0211 & ~n43103;
  assign n43106 = ~n43104 & n43105;
  assign n43107 = ~pi0219 & ~n43106;
  assign n43108 = ~n43097 & n43107;
  assign n43109 = pi0263 & ~n43083;
  assign n43110 = ~n43108 & n43109;
  assign n43111 = n40860 & ~n43067;
  assign n43112 = ~n43110 & n43111;
  assign n43113 = ~po1038 & ~n43017;
  assign n43114 = ~n43112 & n43113;
  assign n43115 = n40910 & ~n43016;
  assign n43116 = ~n43114 & n43115;
  assign n43117 = ~pi0230 & ~n42996;
  assign n43118 = ~n43116 & n43117;
  assign n43119 = po1038 & n42990;
  assign n43120 = ~n38578 & n38649;
  assign n43121 = ~pi1156 & ~n43120;
  assign n43122 = n38592 & ~n39112;
  assign n43123 = ~n43121 & n43122;
  assign n43124 = pi1156 & n39854;
  assign n43125 = pi0219 & ~n43124;
  assign n43126 = ~n43123 & n43125;
  assign n43127 = ~n38510 & ~n43123;
  assign n43128 = pi0211 & ~n43127;
  assign n43129 = n42980 & ~n43128;
  assign n43130 = ~po1038 & ~n43126;
  assign n43131 = ~n43129 & n43130;
  assign n43132 = pi0230 & ~n43119;
  assign n43133 = ~n43131 & n43132;
  assign po0420 = ~n43118 & ~n43133;
  assign n43135 = pi1091 & pi1143;
  assign n43136 = ~pi0200 & n43135;
  assign n43137 = ~pi0796 & n40863;
  assign n43138 = pi0264 & ~n40863;
  assign n43139 = ~pi1091 & ~n43137;
  assign n43140 = ~n43138 & n43139;
  assign n43141 = pi0199 & ~n43136;
  assign n43142 = ~n43140 & n43141;
  assign n43143 = pi1091 & pi1141;
  assign n43144 = ~pi0796 & n40885;
  assign n43145 = pi0264 & ~n40885;
  assign n43146 = ~pi1091 & ~n43144;
  assign n43147 = ~n43145 & n43146;
  assign n43148 = ~n43143 & ~n43147;
  assign n43149 = ~pi0200 & ~n43148;
  assign n43150 = pi1091 & pi1142;
  assign n43151 = ~n43147 & ~n43150;
  assign n43152 = pi0200 & ~n43151;
  assign n43153 = ~pi0199 & ~n43149;
  assign n43154 = ~n43152 & n43153;
  assign n43155 = n16479 & ~n43142;
  assign n43156 = ~n43154 & n43155;
  assign n43157 = pi0219 & ~n42455;
  assign n43158 = ~n39410 & ~n43157;
  assign n43159 = ~n43140 & ~n43158;
  assign n43160 = ~pi0211 & ~n43148;
  assign n43161 = pi0211 & ~n43151;
  assign n43162 = ~pi0219 & ~n43160;
  assign n43163 = ~n43161 & n43162;
  assign n43164 = ~n16479 & ~n43159;
  assign n43165 = ~n43163 & n43164;
  assign n43166 = ~n43156 & ~n43165;
  assign n43167 = ~pi0230 & ~n43166;
  assign n43168 = ~pi0211 & pi1141;
  assign n43169 = ~pi0219 & ~n38455;
  assign n43170 = ~n43168 & n43169;
  assign n43171 = ~n39410 & ~n43170;
  assign n43172 = ~n16479 & ~n43171;
  assign n43173 = ~pi0199 & pi1141;
  assign n43174 = n39388 & ~n43173;
  assign n43175 = ~n38444 & ~n43174;
  assign n43176 = n16479 & ~n43175;
  assign n43177 = pi0230 & ~n43172;
  assign n43178 = ~n43176 & n43177;
  assign po0421 = n43167 | n43178;
  assign n43180 = pi1091 & pi1144;
  assign n43181 = ~pi0200 & n43180;
  assign n43182 = ~pi0819 & n40863;
  assign n43183 = pi0265 & ~n40863;
  assign n43184 = ~pi1091 & ~n43182;
  assign n43185 = ~n43183 & n43184;
  assign n43186 = pi0199 & ~n43181;
  assign n43187 = ~n43185 & n43186;
  assign n43188 = ~pi0819 & n40885;
  assign n43189 = pi0265 & ~n40885;
  assign n43190 = ~pi1091 & ~n43188;
  assign n43191 = ~n43189 & n43190;
  assign n43192 = ~n43150 & ~n43191;
  assign n43193 = ~pi0200 & ~n43192;
  assign n43194 = ~n43135 & ~n43191;
  assign n43195 = pi0200 & ~n43194;
  assign n43196 = ~pi0199 & ~n43193;
  assign n43197 = ~n43195 & n43196;
  assign n43198 = n16479 & ~n43187;
  assign n43199 = ~n43197 & n43198;
  assign n43200 = ~n40771 & ~n43157;
  assign n43201 = ~n43185 & ~n43200;
  assign n43202 = ~pi0211 & ~n43192;
  assign n43203 = pi0211 & ~n43194;
  assign n43204 = ~pi0219 & ~n43202;
  assign n43205 = ~n43203 & n43204;
  assign n43206 = ~n16479 & ~n43201;
  assign n43207 = ~n43205 & n43206;
  assign n43208 = ~n43199 & ~n43207;
  assign n43209 = ~pi0230 & ~n43208;
  assign n43210 = ~pi0211 & pi1142;
  assign n43211 = ~pi0219 & ~n38418;
  assign n43212 = ~n43210 & n43211;
  assign n43213 = ~n40771 & ~n43212;
  assign n43214 = ~n16479 & ~n43213;
  assign n43215 = ~n38443 & n40782;
  assign n43216 = ~n38437 & ~n43215;
  assign n43217 = n16479 & ~n43216;
  assign n43218 = pi0230 & ~n43214;
  assign n43219 = ~n43217 & n43218;
  assign po0422 = n43209 | n43219;
  assign n43221 = ~pi0211 & pi1136;
  assign n43222 = pi0219 & ~n43221;
  assign n43223 = pi0211 & ~pi1135;
  assign n43224 = ~n43222 & ~n43223;
  assign n43225 = ~n10844 & n43224;
  assign n43226 = po1038 & n43225;
  assign n43227 = pi0299 & n43225;
  assign n43228 = ~pi0199 & pi1135;
  assign n43229 = pi0200 & ~n43228;
  assign n43230 = pi0199 & pi1136;
  assign n43231 = ~pi0200 & ~n43230;
  assign n43232 = ~pi0299 & ~n43229;
  assign n43233 = ~n43231 & n43232;
  assign n43234 = ~n43227 & ~n43233;
  assign n43235 = ~po1038 & ~n43234;
  assign n43236 = pi0230 & ~n43226;
  assign n43237 = ~n43235 & n43236;
  assign n43238 = ~n43157 & ~n43222;
  assign n43239 = ~pi0266 & ~n40863;
  assign n43240 = ~pi0948 & n40863;
  assign n43241 = ~pi1091 & ~n43239;
  assign n43242 = ~n43240 & n43241;
  assign n43243 = ~n43238 & ~n43242;
  assign n43244 = ~n16479 & ~n43243;
  assign n43245 = ~pi0266 & ~n40885;
  assign n43246 = ~pi0948 & n40885;
  assign n43247 = ~pi1091 & ~n43245;
  assign n43248 = ~n43246 & n43247;
  assign n43249 = ~pi0219 & ~n43248;
  assign n43250 = pi1135 & n42424;
  assign n43251 = n43249 & ~n43250;
  assign n43252 = n43244 & ~n43251;
  assign n43253 = ~pi0199 & ~n43248;
  assign n43254 = pi1091 & pi1136;
  assign n43255 = pi0199 & ~n43242;
  assign n43256 = ~n43254 & n43255;
  assign n43257 = ~n43253 & ~n43256;
  assign n43258 = ~pi0200 & n43257;
  assign n43259 = pi1091 & pi1135;
  assign n43260 = n43253 & ~n43259;
  assign n43261 = pi0200 & ~n43255;
  assign n43262 = ~n43260 & n43261;
  assign n43263 = ~n43258 & ~n43262;
  assign n43264 = n16479 & ~n43263;
  assign n43265 = ~pi0230 & ~n43252;
  assign n43266 = ~n43264 & n43265;
  assign n43267 = ~n43237 & ~n43266;
  assign n43268 = ~pi1134 & ~n43267;
  assign n43269 = n38699 & ~n43230;
  assign n43270 = ~n43229 & ~n43269;
  assign n43271 = n16479 & n43270;
  assign n43272 = ~n16479 & n43224;
  assign n43273 = pi0230 & ~n43271;
  assign n43274 = ~n43272 & n43273;
  assign n43275 = pi1091 & ~n43223;
  assign n43276 = n43249 & ~n43275;
  assign n43277 = n43244 & ~n43276;
  assign n43278 = ~pi0199 & pi1091;
  assign n43279 = ~n43257 & ~n43278;
  assign n43280 = ~pi0200 & ~n43279;
  assign n43281 = ~n43262 & ~n43280;
  assign n43282 = n16479 & ~n43281;
  assign n43283 = ~pi0230 & ~n43277;
  assign n43284 = ~n43282 & n43283;
  assign n43285 = ~n43274 & ~n43284;
  assign n43286 = pi1134 & ~n43285;
  assign po0423 = ~n43268 & ~n43286;
  assign n43288 = pi1155 & ~n42431;
  assign n43289 = ~n42706 & n43288;
  assign n43290 = ~pi1155 & ~n39027;
  assign n43291 = pi1091 & n43290;
  assign n43292 = ~n43289 & ~n43291;
  assign n43293 = ~pi1154 & ~n43292;
  assign n43294 = n42716 & n43288;
  assign n43295 = ~pi1155 & ~n42660;
  assign n43296 = ~n42460 & n43295;
  assign n43297 = ~n43294 & ~n43296;
  assign n43298 = pi1154 & ~n43297;
  assign n43299 = ~pi0219 & ~n43293;
  assign n43300 = ~n43298 & n43299;
  assign n43301 = pi1153 & n38955;
  assign n43302 = n42708 & ~n43301;
  assign n43303 = ~n39668 & n43302;
  assign n43304 = pi1091 & n42928;
  assign n43305 = ~n42430 & n43304;
  assign n43306 = pi1154 & ~n43305;
  assign n43307 = ~pi0299 & n38946;
  assign n43308 = pi1091 & ~n43307;
  assign n43309 = n43306 & n43308;
  assign n43310 = pi0219 & ~n43303;
  assign n43311 = ~n43309 & n43310;
  assign n43312 = ~n43300 & ~n43311;
  assign n43313 = ~pi0211 & ~n43312;
  assign n43314 = pi1155 & n38963;
  assign n43315 = pi1154 & ~n43314;
  assign n43316 = ~pi1155 & ~n38947;
  assign n43317 = ~n38582 & ~n43316;
  assign n43318 = ~n13062 & ~n43317;
  assign n43319 = pi1091 & n43315;
  assign n43320 = ~n43318 & n43319;
  assign n43321 = ~n38701 & ~n40919;
  assign n43322 = n43302 & ~n43321;
  assign n43323 = pi0211 & ~n43322;
  assign n43324 = ~n43320 & n43323;
  assign n43325 = ~n43313 & ~n43324;
  assign n43326 = pi0267 & ~n43325;
  assign n43327 = n38568 & n42448;
  assign n43328 = ~n42685 & ~n43327;
  assign n43329 = ~n43290 & ~n43328;
  assign n43330 = pi0211 & ~pi1154;
  assign n43331 = ~n43329 & n43330;
  assign n43332 = pi1091 & ~pi1155;
  assign n43333 = ~n38947 & n43332;
  assign n43334 = n38488 & ~n43333;
  assign n43335 = ~n43305 & n43334;
  assign n43336 = ~pi1154 & n38545;
  assign n43337 = ~n38670 & ~n43336;
  assign n43338 = ~n38683 & n43337;
  assign n43339 = pi1091 & n43338;
  assign n43340 = ~pi0211 & ~n43339;
  assign n43341 = ~pi0219 & ~n43335;
  assign n43342 = ~n43340 & n43341;
  assign n43343 = n43307 & n43332;
  assign n43344 = n43306 & ~n43343;
  assign n43345 = n42928 & n43315;
  assign n43346 = ~n43344 & ~n43345;
  assign n43347 = pi0211 & ~n43346;
  assign n43348 = pi1154 & ~n43344;
  assign n43349 = ~n38701 & n42708;
  assign n43350 = ~n39667 & n43349;
  assign n43351 = ~pi0211 & ~n43350;
  assign n43352 = ~n43348 & n43351;
  assign n43353 = pi0219 & ~n43347;
  assign n43354 = ~n43352 & n43353;
  assign n43355 = ~n43342 & ~n43354;
  assign n43356 = ~pi0267 & ~n43331;
  assign n43357 = ~n43355 & n43356;
  assign n43358 = ~n43326 & ~n43357;
  assign n43359 = ~po1038 & n43358;
  assign n43360 = ~pi0219 & ~n38488;
  assign n43361 = ~n38497 & n43360;
  assign n43362 = ~n39158 & ~n43361;
  assign n43363 = pi1091 & ~n43362;
  assign n43364 = ~pi0267 & ~pi1091;
  assign n43365 = ~n43363 & ~n43364;
  assign n43366 = po1038 & ~n43365;
  assign n43367 = ~n40910 & ~n43366;
  assign n43368 = ~n43359 & n43367;
  assign n43369 = ~pi0267 & ~n40980;
  assign n43370 = ~n42538 & n43369;
  assign n43371 = pi0267 & n42734;
  assign n43372 = n40859 & ~n43370;
  assign n43373 = ~n43371 & n43372;
  assign n43374 = ~n40859 & n43364;
  assign n43375 = ~n43363 & ~n43374;
  assign n43376 = ~n43373 & n43375;
  assign n43377 = po1038 & ~n43376;
  assign n43378 = ~n40859 & ~n43358;
  assign n43379 = ~n42777 & n42780;
  assign n43380 = n42805 & ~n43379;
  assign n43381 = pi1154 & pi1155;
  assign n43382 = ~n41014 & n43381;
  assign n43383 = ~n42782 & n43382;
  assign n43384 = ~n43380 & ~n43383;
  assign n43385 = pi0211 & ~n43384;
  assign n43386 = pi1153 & n41055;
  assign n43387 = n38487 & ~n42511;
  assign n43388 = ~n43386 & n43387;
  assign n43389 = ~n42761 & n43388;
  assign n43390 = n41039 & n42749;
  assign n43391 = ~pi1155 & ~n43390;
  assign n43392 = ~n43379 & n43391;
  assign n43393 = ~pi0267 & ~n43392;
  assign n43394 = ~n43389 & n43393;
  assign n43395 = ~n43385 & n43394;
  assign n43396 = pi1155 & ~n42583;
  assign n43397 = n41008 & ~n43059;
  assign n43398 = n43396 & ~n43397;
  assign n43399 = ~n42598 & n43398;
  assign n43400 = ~n42501 & ~n42517;
  assign n43401 = n41009 & ~n43400;
  assign n43402 = pi1154 & ~n43401;
  assign n43403 = ~pi1154 & ~n41028;
  assign n43404 = ~n42597 & n43403;
  assign n43405 = ~pi1155 & ~n43404;
  assign n43406 = ~n43402 & n43405;
  assign n43407 = pi0267 & ~n43399;
  assign n43408 = ~n43406 & n43407;
  assign n43409 = ~n43395 & ~n43408;
  assign n43410 = pi0219 & ~n43409;
  assign n43411 = ~pi1155 & ~n42825;
  assign n43412 = ~n43379 & n43411;
  assign n43413 = n41072 & ~n43401;
  assign n43414 = n43070 & ~n43413;
  assign n43415 = pi1154 & ~n43414;
  assign n43416 = ~pi1154 & ~n42497;
  assign n43417 = pi1155 & ~n43416;
  assign n43418 = n41045 & ~n43417;
  assign n43419 = ~n43415 & ~n43418;
  assign n43420 = pi0211 & ~n43412;
  assign n43421 = ~n43419 & n43420;
  assign n43422 = ~n42828 & ~n43386;
  assign n43423 = pi1155 & ~n43422;
  assign n43424 = pi1153 & ~n41116;
  assign n43425 = ~pi1155 & ~n43424;
  assign n43426 = n42605 & n43425;
  assign n43427 = ~pi1154 & ~n43423;
  assign n43428 = ~n43426 & n43427;
  assign n43429 = ~pi1153 & ~n43098;
  assign n43430 = n43425 & ~n43429;
  assign n43431 = pi1154 & ~n43099;
  assign n43432 = ~n43423 & n43431;
  assign n43433 = ~n43430 & n43432;
  assign n43434 = ~pi0211 & ~n43428;
  assign n43435 = ~n43433 & n43434;
  assign n43436 = ~pi0267 & ~n43435;
  assign n43437 = ~n43421 & n43436;
  assign n43438 = ~pi1153 & n41093;
  assign n43439 = ~n41118 & ~n43438;
  assign n43440 = ~pi1155 & n41072;
  assign n43441 = ~n43439 & n43440;
  assign n43442 = n43033 & n43396;
  assign n43443 = pi1154 & ~n43441;
  assign n43444 = ~n43442 & n43443;
  assign n43445 = ~pi1154 & ~n42517;
  assign n43446 = ~n41105 & n43445;
  assign n43447 = ~pi1155 & ~n43446;
  assign n43448 = ~n40988 & n43445;
  assign n43449 = ~n43447 & n43448;
  assign n43450 = ~n43444 & ~n43449;
  assign n43451 = pi0211 & ~n43450;
  assign n43452 = pi1154 & n43439;
  assign n43453 = n43447 & ~n43452;
  assign n43454 = pi1154 & n41008;
  assign n43455 = ~n41091 & ~n42804;
  assign n43456 = pi1155 & ~n43454;
  assign n43457 = ~n43455 & n43456;
  assign n43458 = ~pi0211 & ~n43457;
  assign n43459 = ~n43453 & n43458;
  assign n43460 = pi0267 & ~n43459;
  assign n43461 = ~n43451 & n43460;
  assign n43462 = ~pi0219 & ~n43461;
  assign n43463 = ~n43437 & n43462;
  assign n43464 = ~n43410 & ~n43463;
  assign n43465 = n40859 & ~n43464;
  assign n43466 = ~po1038 & ~n43378;
  assign n43467 = ~n43465 & n43466;
  assign n43468 = n40910 & ~n43377;
  assign n43469 = ~n43467 & n43468;
  assign n43470 = ~pi0230 & ~n43368;
  assign n43471 = ~n43469 & n43470;
  assign n43472 = pi0219 & ~n38963;
  assign n43473 = ~pi1155 & n43301;
  assign n43474 = ~pi1154 & ~n43473;
  assign n43475 = ~n38947 & ~n43474;
  assign n43476 = pi1155 & n39665;
  assign n43477 = ~n43475 & ~n43476;
  assign n43478 = ~n43472 & ~n43477;
  assign n43479 = pi0211 & ~n43478;
  assign n43480 = ~pi0199 & pi1154;
  assign n43481 = pi0200 & ~n43480;
  assign n43482 = ~n38731 & ~n38962;
  assign n43483 = ~n43481 & n43482;
  assign n43484 = ~n38510 & ~n43483;
  assign n43485 = pi0219 & ~n43484;
  assign n43486 = ~pi0219 & n43338;
  assign n43487 = ~pi0211 & ~n43486;
  assign n43488 = ~n43485 & n43487;
  assign n43489 = ~po1038 & ~n43488;
  assign n43490 = ~n43479 & n43489;
  assign n43491 = po1038 & n43362;
  assign n43492 = pi0230 & ~n43491;
  assign n43493 = ~n43490 & n43492;
  assign po0424 = ~n43471 & ~n43493;
  assign n43495 = pi0268 & pi1152;
  assign n43496 = ~pi0211 & ~n16479;
  assign n43497 = ~po1038 & n38568;
  assign n43498 = ~n43496 & ~n43497;
  assign n43499 = ~pi1151 & n43498;
  assign n43500 = ~pi0199 & n16479;
  assign n43501 = ~n40141 & ~n43500;
  assign n43502 = pi1152 & ~n43498;
  assign n43503 = n43501 & ~n43502;
  assign n43504 = pi1150 & ~n43499;
  assign n43505 = ~n43503 & n43504;
  assign n43506 = ~n43495 & n43505;
  assign n43507 = ~pi1151 & n42389;
  assign n43508 = ~po1038 & ~n11448;
  assign n43509 = po1038 & n11446;
  assign n43510 = ~n43508 & ~n43509;
  assign n43511 = pi1151 & ~n43510;
  assign n43512 = ~pi1152 & ~n43511;
  assign n43513 = ~n16479 & n42478;
  assign n43514 = ~po1038 & n38581;
  assign n43515 = ~n43513 & ~n43514;
  assign n43516 = pi1151 & ~n43515;
  assign n43517 = pi1152 & n43516;
  assign n43518 = ~pi1150 & ~n43507;
  assign n43519 = ~n43512 & n43518;
  assign n43520 = ~n43517 & n43519;
  assign n43521 = ~n43506 & ~n43520;
  assign n43522 = pi1091 & ~n43521;
  assign n43523 = pi1152 & n43505;
  assign n43524 = pi1091 & ~n43523;
  assign n43525 = pi0268 & ~n43524;
  assign n43526 = ~n43522 & ~n43525;
  assign n43527 = ~n40909 & ~n43526;
  assign n43528 = ~n42527 & n42572;
  assign n43529 = ~n41012 & n42584;
  assign n43530 = pi0219 & ~n42513;
  assign n43531 = ~n41011 & n43530;
  assign n43532 = ~n43529 & ~n43531;
  assign n43533 = ~po1038 & ~n42505;
  assign n43534 = n43532 & n43533;
  assign n43535 = ~n43528 & ~n43534;
  assign n43536 = ~pi1151 & ~n43535;
  assign n43537 = ~po1038 & ~n42606;
  assign n43538 = pi0219 & n41048;
  assign n43539 = n43537 & ~n43538;
  assign n43540 = n42572 & ~n42733;
  assign n43541 = ~n43539 & ~n43540;
  assign n43542 = pi1151 & ~n43541;
  assign n43543 = ~n43536 & ~n43542;
  assign n43544 = pi0268 & ~n43543;
  assign n43545 = po1038 & ~n42538;
  assign n43546 = ~n42569 & n43545;
  assign n43547 = po1038 & ~n42732;
  assign n43548 = ~n42525 & n43547;
  assign n43549 = n43546 & ~n43548;
  assign n43550 = pi0219 & ~n40994;
  assign n43551 = ~n42548 & ~n43550;
  assign n43552 = ~n40993 & ~n43551;
  assign n43553 = ~po1038 & ~n41026;
  assign n43554 = n43552 & n43553;
  assign n43555 = ~n43549 & ~n43554;
  assign n43556 = ~pi1151 & n43555;
  assign n43557 = ~n40874 & ~n43541;
  assign n43558 = pi0219 & po1038;
  assign n43559 = ~n40868 & n43558;
  assign n43560 = ~n41032 & n43537;
  assign n43561 = ~n42534 & ~n43559;
  assign n43562 = ~n43560 & n43561;
  assign n43563 = ~n43557 & ~n43562;
  assign n43564 = pi1151 & n43563;
  assign n43565 = ~pi0268 & ~n43564;
  assign n43566 = ~n43556 & n43565;
  assign n43567 = ~n43544 & ~n43566;
  assign n43568 = ~pi1152 & ~n43567;
  assign n43569 = ~n42527 & n43547;
  assign n43570 = ~n41062 & ~n42599;
  assign n43571 = ~n43532 & ~n43570;
  assign n43572 = ~po1038 & ~n43571;
  assign n43573 = ~n40868 & ~n42587;
  assign n43574 = n43572 & ~n43573;
  assign n43575 = ~n43569 & ~n43574;
  assign n43576 = ~pi1151 & ~n43575;
  assign n43577 = ~n40870 & n43533;
  assign n43578 = ~n42733 & n43547;
  assign n43579 = ~n43539 & ~n43578;
  assign n43580 = ~n43577 & n43579;
  assign n43581 = pi1151 & ~n43580;
  assign n43582 = pi0268 & ~n43581;
  assign n43583 = ~n43576 & n43582;
  assign n43584 = ~n42512 & ~n43552;
  assign n43585 = ~po1038 & ~n43584;
  assign n43586 = ~n43546 & ~n43585;
  assign n43587 = ~pi1151 & ~n43586;
  assign n43588 = ~n42528 & n43545;
  assign n43589 = ~pi0219 & n41097;
  assign n43590 = ~n43530 & ~n43589;
  assign n43591 = ~po1038 & ~n43590;
  assign n43592 = ~n43549 & ~n43588;
  assign n43593 = ~n43591 & n43592;
  assign n43594 = pi1151 & ~n43593;
  assign n43595 = ~pi0268 & ~n43594;
  assign n43596 = ~n43587 & n43595;
  assign n43597 = pi1152 & ~n43596;
  assign n43598 = ~n43583 & n43597;
  assign n43599 = ~n43568 & ~n43598;
  assign n43600 = pi1150 & ~n43599;
  assign n43601 = ~n42534 & n43545;
  assign n43602 = ~pi0219 & ~n41045;
  assign n43603 = ~n41002 & ~n43602;
  assign n43604 = n43591 & n43603;
  assign n43605 = ~n43601 & ~n43604;
  assign n43606 = ~pi1151 & ~n43605;
  assign n43607 = ~po1038 & ~n43532;
  assign n43608 = ~n43588 & ~n43607;
  assign n43609 = pi1151 & ~n43608;
  assign n43610 = pi1152 & ~n43606;
  assign n43611 = ~n43609 & n43610;
  assign n43612 = ~pi1151 & n43562;
  assign n43613 = ~n42529 & ~n43559;
  assign n43614 = ~n43572 & n43613;
  assign n43615 = pi1151 & n43614;
  assign n43616 = ~pi1152 & ~n43612;
  assign n43617 = ~n43615 & n43616;
  assign n43618 = ~n43611 & ~n43617;
  assign n43619 = ~pi0268 & ~n43618;
  assign n43620 = pi0219 & ~n42598;
  assign n43621 = ~po1038 & ~n42599;
  assign n43622 = ~n43620 & n43621;
  assign n43623 = ~n43548 & ~n43622;
  assign n43624 = ~pi1151 & n43623;
  assign n43625 = ~n42570 & n43547;
  assign n43626 = ~n42548 & ~n43620;
  assign n43627 = n41102 & ~n43626;
  assign n43628 = ~po1038 & ~n43627;
  assign n43629 = ~n43625 & ~n43628;
  assign n43630 = pi1151 & n43629;
  assign n43631 = pi1152 & ~n43624;
  assign n43632 = ~n43630 & n43631;
  assign n43633 = n40874 & ~n43541;
  assign n43634 = ~pi1151 & ~n43633;
  assign n43635 = ~po1038 & ~n42553;
  assign n43636 = ~n42548 & n43635;
  assign n43637 = ~n42573 & ~n43636;
  assign n43638 = pi1151 & n43637;
  assign n43639 = ~pi1152 & ~n43634;
  assign n43640 = ~n43638 & n43639;
  assign n43641 = pi0268 & ~n43640;
  assign n43642 = ~n43632 & n43641;
  assign n43643 = ~pi1150 & ~n43642;
  assign n43644 = ~n43619 & n43643;
  assign n43645 = ~n43600 & ~n43644;
  assign n43646 = n40909 & ~n43645;
  assign n43647 = ~pi0230 & ~n43527;
  assign n43648 = ~n43646 & n43647;
  assign n43649 = pi0230 & ~n43505;
  assign n43650 = ~n43520 & n43649;
  assign po0425 = ~n43648 & ~n43650;
  assign n43652 = ~pi0199 & pi1137;
  assign n43653 = pi0200 & ~n43652;
  assign n43654 = pi0199 & pi1138;
  assign n43655 = ~pi0199 & pi1136;
  assign n43656 = ~pi0200 & ~n43654;
  assign n43657 = ~n43655 & n43656;
  assign n43658 = ~n43653 & ~n43657;
  assign n43659 = n16479 & ~n43658;
  assign n43660 = ~pi0211 & pi1138;
  assign n43661 = pi0219 & n43660;
  assign n43662 = pi0211 & pi1137;
  assign n43663 = ~n43221 & ~n43662;
  assign n43664 = ~pi0219 & ~n43663;
  assign n43665 = ~n43661 & ~n43664;
  assign n43666 = ~n16479 & n43665;
  assign n43667 = ~n43659 & ~n43666;
  assign n43668 = pi0230 & ~n43667;
  assign n43669 = ~pi0200 & n43254;
  assign n43670 = pi1137 & n40951;
  assign n43671 = ~n43669 & ~n43670;
  assign n43672 = n43500 & n43671;
  assign n43673 = pi1091 & ~n43663;
  assign n43674 = n40141 & ~n43673;
  assign n43675 = ~n43672 & ~n43674;
  assign n43676 = ~pi0817 & n40885;
  assign n43677 = pi0269 & ~n40885;
  assign n43678 = ~pi1091 & ~n43676;
  assign n43679 = ~n43677 & n43678;
  assign n43680 = ~n43675 & ~n43679;
  assign n43681 = ~pi0817 & n40863;
  assign n43682 = pi0269 & ~n40863;
  assign n43683 = ~pi1091 & ~n43681;
  assign n43684 = ~n43682 & n43683;
  assign n43685 = pi1138 & n42455;
  assign n43686 = pi0219 & ~n16479;
  assign n43687 = ~n43685 & n43686;
  assign n43688 = ~pi0200 & pi1091;
  assign n43689 = pi1138 & n43688;
  assign n43690 = pi0199 & ~n43689;
  assign n43691 = n16479 & n43690;
  assign n43692 = ~n43687 & ~n43691;
  assign n43693 = ~n43684 & ~n43692;
  assign n43694 = ~n43680 & ~n43693;
  assign n43695 = ~pi0230 & ~n43694;
  assign po0426 = ~n43668 & ~n43695;
  assign n43697 = ~pi0805 & n40863;
  assign n43698 = pi0270 & ~n40863;
  assign n43699 = ~pi1091 & ~n43697;
  assign n43700 = ~n43698 & n43699;
  assign n43701 = n42455 & n43168;
  assign n43702 = n43686 & ~n43701;
  assign n43703 = ~pi0200 & n43143;
  assign n43704 = pi0199 & ~n43703;
  assign n43705 = n16479 & n43704;
  assign n43706 = ~n43702 & ~n43705;
  assign n43707 = ~n43700 & ~n43706;
  assign n43708 = ~pi0805 & n40885;
  assign n43709 = pi0270 & ~n40885;
  assign n43710 = ~pi1091 & ~n43708;
  assign n43711 = ~n43709 & n43710;
  assign n43712 = ~pi0211 & pi1139;
  assign n43713 = pi0211 & pi1140;
  assign n43714 = ~n43712 & ~n43713;
  assign n43715 = pi1091 & ~n43714;
  assign n43716 = n40141 & ~n43715;
  assign n43717 = pi1091 & pi1140;
  assign n43718 = pi0200 & n43717;
  assign n43719 = pi1139 & n43688;
  assign n43720 = ~n43718 & ~n43719;
  assign n43721 = n43500 & n43720;
  assign n43722 = ~n43716 & ~n43721;
  assign n43723 = ~n43711 & ~n43722;
  assign n43724 = ~pi0230 & ~n43707;
  assign n43725 = ~n43723 & n43724;
  assign n43726 = pi0219 & ~n43168;
  assign n43727 = ~pi0219 & n43714;
  assign n43728 = ~n43726 & ~n43727;
  assign n43729 = ~n16479 & ~n43728;
  assign n43730 = ~pi0199 & pi1140;
  assign n43731 = pi0200 & ~n43730;
  assign n43732 = pi0199 & pi1141;
  assign n43733 = ~pi0199 & pi1139;
  assign n43734 = ~pi0200 & ~n43732;
  assign n43735 = ~n43733 & n43734;
  assign n43736 = ~n43731 & ~n43735;
  assign n43737 = n16479 & ~n43736;
  assign n43738 = pi0230 & ~n43729;
  assign n43739 = ~n43737 & n43738;
  assign po0427 = n43725 | n43739;
  assign n43741 = ~pi0211 & pi1147;
  assign n43742 = n42444 & n43741;
  assign n43743 = ~pi0271 & ~n40866;
  assign n43744 = ~n40871 & ~n43743;
  assign n43745 = pi0219 & ~n43744;
  assign n43746 = ~pi1091 & ~n40887;
  assign n43747 = pi0271 & ~n43746;
  assign n43748 = ~pi0271 & ~n40888;
  assign n43749 = ~n43747 & ~n43748;
  assign n43750 = pi1091 & pi1146;
  assign n43751 = ~n43749 & ~n43750;
  assign n43752 = ~pi0211 & n43750;
  assign n43753 = ~n43751 & ~n43752;
  assign n43754 = pi1091 & n39412;
  assign n43755 = ~pi0219 & ~n43754;
  assign n43756 = ~n43753 & n43755;
  assign n43757 = ~n43745 & ~n43756;
  assign n43758 = ~n16479 & ~n43742;
  assign n43759 = ~n43757 & n43758;
  assign n43760 = pi0199 & ~n43744;
  assign n43761 = ~pi0199 & n43751;
  assign n43762 = ~n43760 & ~n43761;
  assign n43763 = pi0200 & ~n43762;
  assign n43764 = pi1147 & n40931;
  assign n43765 = pi1091 & pi1145;
  assign n43766 = ~pi0199 & ~n43765;
  assign n43767 = ~n43749 & n43766;
  assign n43768 = ~n43760 & ~n43767;
  assign n43769 = ~pi0200 & ~n43764;
  assign n43770 = ~n43768 & n43769;
  assign n43771 = ~n43763 & ~n43770;
  assign n43772 = n16479 & ~n43771;
  assign n43773 = ~n43759 & ~n43772;
  assign n43774 = ~pi0230 & ~n43773;
  assign n43775 = pi1147 & n42386;
  assign n43776 = ~n40225 & ~n40235;
  assign n43777 = ~pi0219 & ~n43776;
  assign n43778 = ~pi0200 & ~n39393;
  assign n43779 = n40339 & ~n43778;
  assign n43780 = ~n43775 & ~n43777;
  assign n43781 = ~n43779 & n43780;
  assign n43782 = ~po1038 & ~n43781;
  assign n43783 = pi0219 & ~n43741;
  assign n43784 = ~n39412 & n41531;
  assign n43785 = ~n43783 & ~n43784;
  assign n43786 = po1038 & n43785;
  assign n43787 = pi0230 & ~n43786;
  assign n43788 = ~n43782 & n43787;
  assign po0428 = ~n43774 & ~n43788;
  assign n43790 = po1038 & n10844;
  assign n43791 = ~n13065 & ~n43790;
  assign n43792 = ~pi1150 & n43791;
  assign n43793 = ~n43498 & ~n43792;
  assign n43794 = ~pi1149 & ~n43793;
  assign n43795 = pi1149 & ~pi1150;
  assign n43796 = ~n43498 & ~n43795;
  assign n43797 = n43501 & ~n43796;
  assign n43798 = ~n43794 & ~n43797;
  assign n43799 = pi1091 & ~n43798;
  assign n43800 = pi1148 & ~n43799;
  assign n43801 = pi1150 & ~n42389;
  assign n43802 = ~pi1149 & ~n43801;
  assign n43803 = pi1091 & n43802;
  assign n43804 = ~n16479 & n42712;
  assign n43805 = ~po1038 & n40936;
  assign n43806 = ~n43804 & ~n43805;
  assign n43807 = ~pi1150 & n43806;
  assign n43808 = pi1091 & ~n43515;
  assign n43809 = pi1150 & ~n43808;
  assign n43810 = pi1149 & ~n43807;
  assign n43811 = ~n43809 & n43810;
  assign n43812 = ~pi1148 & ~n43803;
  assign n43813 = ~n43811 & n43812;
  assign n43814 = ~pi0283 & ~n43800;
  assign n43815 = ~n43813 & n43814;
  assign n43816 = ~pi1150 & ~n43633;
  assign n43817 = pi1150 & n43623;
  assign n43818 = ~pi1149 & ~n43816;
  assign n43819 = ~n43817 & n43818;
  assign n43820 = pi1150 & n43629;
  assign n43821 = ~pi1150 & n43637;
  assign n43822 = pi1149 & ~n43821;
  assign n43823 = ~n43820 & n43822;
  assign n43824 = ~n43819 & ~n43823;
  assign n43825 = ~pi1148 & ~n43824;
  assign n43826 = ~pi1150 & n43541;
  assign n43827 = pi1150 & n43580;
  assign n43828 = pi1149 & ~n43826;
  assign n43829 = ~n43827 & n43828;
  assign n43830 = ~pi1150 & n43535;
  assign n43831 = pi1150 & n43575;
  assign n43832 = ~pi1149 & ~n43830;
  assign n43833 = ~n43831 & n43832;
  assign n43834 = ~n43829 & ~n43833;
  assign n43835 = pi1148 & ~n43834;
  assign n43836 = pi0283 & ~n43825;
  assign n43837 = ~n43835 & n43836;
  assign n43838 = pi0272 & ~n43815;
  assign n43839 = ~n43837 & n43838;
  assign n43840 = ~pi1150 & ~n43563;
  assign n43841 = pi1150 & ~n43593;
  assign n43842 = pi1149 & ~n43840;
  assign n43843 = ~n43841 & n43842;
  assign n43844 = pi1150 & ~n43586;
  assign n43845 = ~pi1150 & ~n43555;
  assign n43846 = ~pi1149 & ~n43845;
  assign n43847 = ~n43844 & n43846;
  assign n43848 = ~n43843 & ~n43847;
  assign n43849 = pi1148 & ~n43848;
  assign n43850 = pi1150 & n43605;
  assign n43851 = ~pi1150 & ~n43562;
  assign n43852 = ~pi1149 & ~n43851;
  assign n43853 = ~n43850 & n43852;
  assign n43854 = ~pi1150 & ~n43614;
  assign n43855 = pi1150 & n43608;
  assign n43856 = pi1149 & ~n43855;
  assign n43857 = ~n43854 & n43856;
  assign n43858 = ~pi1148 & ~n43853;
  assign n43859 = ~n43857 & n43858;
  assign n43860 = ~n43849 & ~n43859;
  assign n43861 = pi0283 & ~n43860;
  assign n43862 = ~po1038 & n38550;
  assign n43863 = ~n40141 & ~n43862;
  assign n43864 = ~n43496 & n43863;
  assign n43865 = pi1150 & ~n43864;
  assign n43866 = pi1149 & ~n43865;
  assign n43867 = n43501 & n43866;
  assign n43868 = pi1148 & ~n43794;
  assign n43869 = ~n43867 & n43868;
  assign n43870 = pi1091 & n43869;
  assign n43871 = ~pi1148 & ~n43802;
  assign n43872 = ~pi1150 & ~n43510;
  assign n43873 = pi1150 & n43515;
  assign n43874 = pi1149 & ~n43872;
  assign n43875 = ~n43873 & n43874;
  assign n43876 = pi1091 & ~n43875;
  assign n43877 = n43871 & n43876;
  assign n43878 = ~pi0283 & ~n43877;
  assign n43879 = ~n43870 & n43878;
  assign n43880 = ~pi0272 & ~n43879;
  assign n43881 = ~n43861 & n43880;
  assign n43882 = ~pi0230 & ~n43839;
  assign n43883 = ~n43881 & n43882;
  assign n43884 = pi1149 & ~n43515;
  assign n43885 = ~n43866 & ~n43884;
  assign n43886 = ~n43872 & ~n43885;
  assign n43887 = n43871 & ~n43886;
  assign n43888 = pi0230 & ~n43869;
  assign n43889 = ~n43887 & n43888;
  assign po0429 = ~n43883 & ~n43889;
  assign n43891 = ~pi0273 & ~n40867;
  assign n43892 = ~n40873 & ~n43891;
  assign n43893 = pi0219 & ~n43892;
  assign n43894 = ~pi0273 & ~n40889;
  assign n43895 = n40891 & ~n43894;
  assign n43896 = ~pi0219 & ~n43752;
  assign n43897 = ~n43895 & n43896;
  assign n43898 = ~n43893 & ~n43897;
  assign n43899 = po1038 & n43898;
  assign n43900 = pi0299 & n43898;
  assign n43901 = pi0199 & ~n43892;
  assign n43902 = ~pi0200 & n43750;
  assign n43903 = ~pi0199 & ~n43902;
  assign n43904 = ~n43895 & n43903;
  assign n43905 = ~pi0299 & ~n43901;
  assign n43906 = ~n43904 & n43905;
  assign n43907 = ~n43900 & ~n43906;
  assign n43908 = ~n11447 & ~n41041;
  assign n43909 = pi1091 & ~n43908;
  assign n43910 = n43907 & ~n43909;
  assign n43911 = ~po1038 & ~n43910;
  assign n43912 = pi1091 & n42573;
  assign n43913 = ~n43911 & ~n43912;
  assign n43914 = pi1147 & ~n43913;
  assign n43915 = n40447 & ~n43907;
  assign n43916 = ~pi1148 & ~n43915;
  assign n43917 = pi1091 & n38519;
  assign n43918 = ~n43898 & ~n43917;
  assign n43919 = pi0299 & ~n43918;
  assign n43920 = n40932 & ~n43763;
  assign n43921 = ~n43906 & ~n43920;
  assign n43922 = ~n43919 & n43921;
  assign n43923 = ~po1038 & ~n43922;
  assign n43924 = n40080 & n42444;
  assign n43925 = pi1148 & ~n43924;
  assign n43926 = ~n43923 & n43925;
  assign n43927 = ~n43916 & ~n43926;
  assign n43928 = ~n43899 & ~n43927;
  assign n43929 = ~n43914 & n43928;
  assign n43930 = ~pi0230 & ~n43929;
  assign n43931 = pi1146 & ~n41404;
  assign n43932 = ~n43791 & n43931;
  assign n43933 = ~pi0211 & ~n40234;
  assign n43934 = n40141 & ~n43933;
  assign n43935 = ~pi1146 & n10809;
  assign n43936 = n43500 & ~n43935;
  assign n43937 = ~n43934 & ~n43936;
  assign n43938 = pi1147 & ~n43937;
  assign n43939 = ~pi1148 & ~n43932;
  assign n43940 = ~n43938 & n43939;
  assign n43941 = ~pi0199 & pi1147;
  assign n43942 = pi0200 & ~n43941;
  assign n43943 = ~n43935 & ~n43942;
  assign n43944 = n16479 & n43943;
  assign n43945 = ~pi1146 & n10844;
  assign n43946 = pi1147 & n40141;
  assign n43947 = ~n43496 & ~n43946;
  assign n43948 = ~n43945 & ~n43947;
  assign n43949 = pi1148 & ~n43944;
  assign n43950 = ~n43948 & n43949;
  assign n43951 = pi0230 & ~n43940;
  assign n43952 = ~n43950 & n43951;
  assign po0430 = n43930 | n43952;
  assign n43954 = ~pi0200 & n43765;
  assign n43955 = ~pi0659 & n40863;
  assign n43956 = pi0274 & ~n40863;
  assign n43957 = ~pi1091 & ~n43955;
  assign n43958 = ~n43956 & n43957;
  assign n43959 = pi0199 & ~n43954;
  assign n43960 = ~n43958 & n43959;
  assign n43961 = ~pi0659 & n40885;
  assign n43962 = pi0274 & ~n40885;
  assign n43963 = ~pi1091 & ~n43961;
  assign n43964 = ~n43962 & n43963;
  assign n43965 = ~n43180 & ~n43964;
  assign n43966 = pi0200 & ~n43965;
  assign n43967 = ~n43135 & ~n43964;
  assign n43968 = ~pi0200 & ~n43967;
  assign n43969 = ~pi0199 & ~n43966;
  assign n43970 = ~n43968 & n43969;
  assign n43971 = n16479 & ~n43960;
  assign n43972 = ~n43970 & n43971;
  assign n43973 = pi0211 & ~n43965;
  assign n43974 = ~pi0211 & ~n43967;
  assign n43975 = ~pi0219 & ~n43973;
  assign n43976 = ~n43974 & n43975;
  assign n43977 = pi0219 & ~n43754;
  assign n43978 = ~n43958 & n43977;
  assign n43979 = ~n16479 & ~n43978;
  assign n43980 = ~n43976 & n43979;
  assign n43981 = ~pi0230 & ~n43972;
  assign n43982 = ~n43980 & n43981;
  assign n43983 = ~n38508 & ~n40225;
  assign n43984 = ~pi0219 & ~n38425;
  assign n43985 = ~n39413 & n43984;
  assign n43986 = ~n43983 & ~n43985;
  assign n43987 = ~n38436 & n40332;
  assign n43988 = n40788 & ~n43987;
  assign n43989 = ~n43986 & ~n43988;
  assign n43990 = ~po1038 & ~n43989;
  assign n43991 = ~n40221 & ~n43985;
  assign n43992 = pi0230 & ~n43990;
  assign n43993 = ~n43991 & n43992;
  assign po0431 = ~n43982 & ~n43993;
  assign n43995 = pi1151 & ~n43498;
  assign n43996 = pi1149 & n43501;
  assign n43997 = ~n43995 & n43996;
  assign n43998 = ~pi1149 & n43516;
  assign n43999 = ~n43997 & ~n43998;
  assign n44000 = pi1150 & ~n43999;
  assign n44001 = ~pi1151 & n43791;
  assign n44002 = pi1149 & ~n43498;
  assign n44003 = ~n44001 & n44002;
  assign n44004 = ~pi1149 & pi1151;
  assign n44005 = ~n42389 & n44004;
  assign n44006 = ~pi1150 & ~n44005;
  assign n44007 = ~n44003 & n44006;
  assign n44008 = ~n44000 & ~n44007;
  assign n44009 = pi1091 & ~n44008;
  assign n44010 = ~pi1151 & n41484;
  assign n44011 = ~n43806 & n44010;
  assign n44012 = ~n44009 & ~n44011;
  assign n44013 = pi0275 & ~n44012;
  assign n44014 = n43498 & n43795;
  assign n44015 = n40607 & ~n42389;
  assign n44016 = ~pi1151 & n43510;
  assign n44017 = pi1150 & ~n44016;
  assign n44018 = ~n43516 & n44017;
  assign n44019 = ~pi1149 & ~n44015;
  assign n44020 = ~n44018 & n44019;
  assign n44021 = ~n43997 & ~n44014;
  assign n44022 = ~n44020 & n44021;
  assign n44023 = pi1091 & n44022;
  assign n44024 = ~pi0275 & ~n44023;
  assign n44025 = ~n40908 & ~n44024;
  assign n44026 = ~n44013 & n44025;
  assign n44027 = ~pi1150 & n43605;
  assign n44028 = pi1151 & ~n43855;
  assign n44029 = ~n44027 & n44028;
  assign n44030 = pi1150 & ~n43614;
  assign n44031 = ~pi1151 & ~n43851;
  assign n44032 = ~n44030 & n44031;
  assign n44033 = ~n44029 & ~n44032;
  assign n44034 = ~pi0275 & ~n44033;
  assign n44035 = pi1150 & n43637;
  assign n44036 = ~n43816 & ~n44035;
  assign n44037 = ~pi1151 & ~n44036;
  assign n44038 = ~pi1150 & n43623;
  assign n44039 = ~n43820 & ~n44038;
  assign n44040 = pi1151 & ~n44039;
  assign n44041 = pi0275 & ~n44037;
  assign n44042 = ~n44040 & n44041;
  assign n44043 = ~pi1149 & ~n44042;
  assign n44044 = ~n44034 & n44043;
  assign n44045 = pi1150 & ~n43563;
  assign n44046 = ~pi1151 & ~n44045;
  assign n44047 = ~n43845 & n44046;
  assign n44048 = ~pi1150 & ~n43586;
  assign n44049 = pi1151 & ~n43841;
  assign n44050 = ~n44048 & n44049;
  assign n44051 = ~pi0275 & ~n44047;
  assign n44052 = ~n44050 & n44051;
  assign n44053 = pi1151 & ~n43575;
  assign n44054 = ~pi1150 & ~n43536;
  assign n44055 = ~n44053 & n44054;
  assign n44056 = ~pi1151 & ~n43541;
  assign n44057 = pi1150 & ~n44056;
  assign n44058 = ~n43581 & n44057;
  assign n44059 = pi0275 & ~n44058;
  assign n44060 = ~n44055 & n44059;
  assign n44061 = pi1149 & ~n44052;
  assign n44062 = ~n44060 & n44061;
  assign n44063 = n40908 & ~n44044;
  assign n44064 = ~n44062 & n44063;
  assign n44065 = ~n44026 & ~n44064;
  assign n44066 = ~pi0230 & ~n44065;
  assign n44067 = pi0230 & n44022;
  assign po0432 = n44066 | n44067;
  assign n44069 = ~pi0276 & ~n40886;
  assign n44070 = n43746 & ~n44069;
  assign n44071 = ~n38419 & ~n40210;
  assign n44072 = pi1091 & ~n44071;
  assign n44073 = n40141 & ~n44072;
  assign n44074 = pi1145 & n40951;
  assign n44075 = ~n43181 & ~n44074;
  assign n44076 = n43500 & n44075;
  assign n44077 = ~n44073 & ~n44076;
  assign n44078 = ~n44070 & ~n44077;
  assign n44079 = ~pi0276 & ~n40864;
  assign n44080 = n40870 & ~n44079;
  assign n44081 = n43686 & ~n43752;
  assign n44082 = pi0199 & ~n43902;
  assign n44083 = n16479 & n44082;
  assign n44084 = ~n44081 & ~n44083;
  assign n44085 = ~n44080 & ~n44084;
  assign n44086 = ~pi0230 & ~n44078;
  assign n44087 = ~n44085 & n44086;
  assign n44088 = ~n38434 & n41294;
  assign n44089 = ~n40330 & ~n44088;
  assign n44090 = n16479 & ~n44089;
  assign n44091 = ~pi0219 & ~n44071;
  assign n44092 = pi1146 & n38519;
  assign n44093 = ~n44091 & ~n44092;
  assign n44094 = ~n16479 & n44093;
  assign n44095 = pi0230 & ~n44090;
  assign n44096 = ~n44094 & n44095;
  assign po0433 = n44087 | n44096;
  assign n44098 = ~pi0200 & n43150;
  assign n44099 = ~pi0820 & n40863;
  assign n44100 = pi0277 & ~n40863;
  assign n44101 = ~pi1091 & ~n44099;
  assign n44102 = ~n44100 & n44101;
  assign n44103 = pi0199 & ~n44098;
  assign n44104 = ~n44102 & n44103;
  assign n44105 = ~pi0820 & n40885;
  assign n44106 = pi0277 & ~n40885;
  assign n44107 = ~pi1091 & ~n44105;
  assign n44108 = ~n44106 & n44107;
  assign n44109 = ~n43717 & ~n44108;
  assign n44110 = ~pi0200 & ~n44109;
  assign n44111 = ~n43143 & ~n44108;
  assign n44112 = pi0200 & ~n44111;
  assign n44113 = ~pi0199 & ~n44110;
  assign n44114 = ~n44112 & n44113;
  assign n44115 = n16479 & ~n44104;
  assign n44116 = ~n44114 & n44115;
  assign n44117 = pi0219 & ~n43210;
  assign n44118 = ~n43157 & ~n44117;
  assign n44119 = ~n44102 & ~n44118;
  assign n44120 = ~pi0211 & ~n44109;
  assign n44121 = pi0211 & ~n44111;
  assign n44122 = ~pi0219 & ~n44120;
  assign n44123 = ~n44121 & n44122;
  assign n44124 = ~n16479 & ~n44119;
  assign n44125 = ~n44123 & n44124;
  assign n44126 = ~n44116 & ~n44125;
  assign n44127 = ~pi0230 & ~n44126;
  assign n44128 = pi0211 & pi1141;
  assign n44129 = ~pi0211 & pi1140;
  assign n44130 = ~pi0219 & ~n44128;
  assign n44131 = ~n44129 & n44130;
  assign n44132 = ~n44117 & ~n44131;
  assign n44133 = ~n16479 & ~n44132;
  assign n44134 = n38433 & ~n43730;
  assign n44135 = pi0200 & ~n43173;
  assign n44136 = ~n44134 & ~n44135;
  assign n44137 = n16479 & ~n44136;
  assign n44138 = pi0230 & ~n44133;
  assign n44139 = ~n44137 & n44138;
  assign po0434 = n44127 | n44139;
  assign n44141 = ~pi0278 & ~n40863;
  assign n44142 = ~pi0976 & n40863;
  assign n44143 = ~pi1091 & ~n44141;
  assign n44144 = ~n44142 & n44143;
  assign n44145 = pi0199 & ~n44144;
  assign n44146 = pi1091 & ~pi1132;
  assign n44147 = pi0976 & n40885;
  assign n44148 = pi0278 & ~n40885;
  assign n44149 = ~pi1091 & ~n44147;
  assign n44150 = ~n44148 & n44149;
  assign n44151 = ~n44146 & ~n44150;
  assign n44152 = ~pi0199 & ~n44151;
  assign n44153 = ~n44145 & ~n44152;
  assign n44154 = ~pi0200 & ~n44153;
  assign n44155 = pi1091 & ~pi1133;
  assign n44156 = ~n44150 & ~n44155;
  assign n44157 = ~pi0199 & ~n44156;
  assign n44158 = ~n44145 & ~n44157;
  assign n44159 = pi0200 & ~n44158;
  assign n44160 = ~pi0299 & ~n44159;
  assign n44161 = ~n44154 & n44160;
  assign n44162 = pi0219 & ~n44144;
  assign n44163 = pi0211 & ~pi1133;
  assign n44164 = ~pi0211 & ~pi1132;
  assign n44165 = ~n44163 & ~n44164;
  assign n44166 = pi1091 & ~n44165;
  assign n44167 = ~n44150 & ~n44166;
  assign n44168 = ~pi0219 & ~n44167;
  assign n44169 = ~n44162 & ~n44168;
  assign n44170 = pi0299 & n44169;
  assign n44171 = ~n44161 & ~n44170;
  assign n44172 = ~po1038 & ~n44171;
  assign n44173 = po1038 & n44169;
  assign n44174 = ~pi0230 & ~n44173;
  assign n44175 = ~n44172 & n44174;
  assign n44176 = n39374 & n44165;
  assign n44177 = ~pi0199 & pi1132;
  assign n44178 = ~pi0200 & ~n44177;
  assign n44179 = ~pi0199 & pi1133;
  assign n44180 = pi0200 & ~n44179;
  assign n44181 = ~pi0299 & ~n44180;
  assign n44182 = ~n44178 & n44181;
  assign n44183 = n38508 & n44165;
  assign n44184 = ~n44182 & ~n44183;
  assign n44185 = ~po1038 & ~n44184;
  assign n44186 = pi0230 & ~n44176;
  assign n44187 = ~n44185 & n44186;
  assign n44188 = ~n44175 & ~n44187;
  assign n44189 = ~pi1134 & ~n44188;
  assign n44190 = n10809 & ~n44177;
  assign n44191 = n44181 & ~n44190;
  assign n44192 = ~n42627 & ~n44183;
  assign n44193 = ~n44191 & n44192;
  assign n44194 = ~po1038 & ~n44193;
  assign n44195 = ~pi0219 & ~n44165;
  assign n44196 = ~n40081 & ~n44195;
  assign n44197 = pi0230 & ~n44194;
  assign n44198 = ~n44196 & n44197;
  assign n44199 = ~n40931 & n44154;
  assign n44200 = n44160 & ~n44199;
  assign n44201 = n13062 & n42455;
  assign n44202 = ~n44170 & ~n44201;
  assign n44203 = ~n44200 & n44202;
  assign n44204 = ~po1038 & ~n44203;
  assign n44205 = ~n43924 & n44174;
  assign n44206 = ~n44204 & n44205;
  assign n44207 = ~n44198 & ~n44206;
  assign n44208 = pi1134 & ~n44207;
  assign po0435 = ~n44189 & ~n44208;
  assign n44210 = ~pi0279 & ~n40863;
  assign n44211 = ~pi0958 & n40863;
  assign n44212 = ~pi1091 & ~n44210;
  assign n44213 = ~n44211 & n44212;
  assign n44214 = pi1135 & n43688;
  assign n44215 = ~n44213 & ~n44214;
  assign n44216 = pi0199 & ~n44215;
  assign n44217 = pi0958 & n40885;
  assign n44218 = pi0279 & ~n40885;
  assign n44219 = ~pi1091 & ~n44217;
  assign n44220 = ~n44218 & n44219;
  assign n44221 = ~pi1133 & n43688;
  assign n44222 = ~pi0199 & ~n44221;
  assign n44223 = ~n44220 & n44222;
  assign n44224 = ~n44216 & ~n44223;
  assign n44225 = n16479 & ~n44224;
  assign n44226 = ~n40951 & n44225;
  assign n44227 = ~n42424 & ~n44155;
  assign n44228 = ~n44220 & n44227;
  assign n44229 = ~pi0219 & ~n44228;
  assign n44230 = pi1135 & n42455;
  assign n44231 = pi0219 & ~n44230;
  assign n44232 = ~n44213 & n44231;
  assign n44233 = ~n16479 & ~n44232;
  assign n44234 = ~n44229 & n44233;
  assign n44235 = ~pi0230 & ~n44234;
  assign n44236 = ~n44226 & n44235;
  assign n44237 = pi1135 & n38519;
  assign n44238 = ~pi0211 & ~pi1133;
  assign n44239 = ~pi0219 & ~n44238;
  assign n44240 = ~pi0211 & n44239;
  assign n44241 = ~n44237 & ~n44240;
  assign n44242 = po1038 & ~n44241;
  assign n44243 = pi0199 & pi1135;
  assign n44244 = ~n44179 & ~n44243;
  assign n44245 = n38568 & ~n44244;
  assign n44246 = pi0299 & ~n44241;
  assign n44247 = ~n44245 & ~n44246;
  assign n44248 = ~po1038 & ~n44247;
  assign n44249 = pi0230 & ~n44242;
  assign n44250 = ~n44248 & n44249;
  assign n44251 = ~n44236 & ~n44250;
  assign n44252 = ~pi1134 & ~n44251;
  assign n44253 = ~pi1133 & n10809;
  assign n44254 = ~pi0200 & pi1135;
  assign n44255 = pi0199 & ~n44254;
  assign n44256 = ~n44253 & ~n44255;
  assign n44257 = n16479 & ~n44256;
  assign n44258 = ~n44237 & ~n44239;
  assign n44259 = ~n16479 & n44258;
  assign n44260 = ~n44257 & ~n44259;
  assign n44261 = pi0230 & ~n44260;
  assign n44262 = pi1091 & ~n44238;
  assign n44263 = n40141 & n44262;
  assign n44264 = ~n44225 & ~n44263;
  assign n44265 = n44235 & n44264;
  assign n44266 = ~n44261 & ~n44265;
  assign n44267 = pi1134 & ~n44266;
  assign po0436 = ~n44252 & ~n44267;
  assign n44269 = ~pi0211 & pi1135;
  assign n44270 = pi0211 & pi1136;
  assign n44271 = ~n44269 & ~n44270;
  assign n44272 = pi1091 & n44271;
  assign n44273 = ~pi0280 & ~n40885;
  assign n44274 = pi0914 & n40885;
  assign n44275 = ~pi1091 & ~n44273;
  assign n44276 = ~n44274 & n44275;
  assign n44277 = ~n44272 & ~n44276;
  assign n44278 = ~pi0219 & ~n44277;
  assign n44279 = ~pi0211 & pi1137;
  assign n44280 = pi0219 & ~n44279;
  assign n44281 = ~n43157 & ~n44280;
  assign n44282 = ~pi0914 & n40863;
  assign n44283 = pi0280 & ~n40863;
  assign n44284 = ~pi1091 & ~n44282;
  assign n44285 = ~n44283 & n44284;
  assign n44286 = ~n44281 & ~n44285;
  assign n44287 = ~n44278 & ~n44286;
  assign n44288 = ~n16479 & ~n44287;
  assign n44289 = pi1137 & n43688;
  assign n44290 = ~n44285 & ~n44289;
  assign n44291 = pi0199 & ~n44290;
  assign n44292 = pi0200 & pi1136;
  assign n44293 = pi1091 & ~n44254;
  assign n44294 = ~n44292 & n44293;
  assign n44295 = ~pi0199 & ~n44294;
  assign n44296 = ~n44276 & n44295;
  assign n44297 = n16479 & ~n44291;
  assign n44298 = ~n44296 & n44297;
  assign n44299 = ~n44288 & ~n44298;
  assign n44300 = ~pi0230 & ~n44299;
  assign n44301 = pi0200 & ~n43655;
  assign n44302 = pi0199 & pi1137;
  assign n44303 = ~pi0200 & ~n43228;
  assign n44304 = ~n44302 & n44303;
  assign n44305 = ~n44301 & ~n44304;
  assign n44306 = n16479 & n44305;
  assign n44307 = ~pi0219 & n44271;
  assign n44308 = ~n44280 & ~n44307;
  assign n44309 = ~n16479 & n44308;
  assign n44310 = pi0230 & ~n44306;
  assign n44311 = ~n44309 & n44310;
  assign po0437 = ~n44300 & ~n44311;
  assign n44313 = ~pi0199 & pi1138;
  assign n44314 = pi0200 & ~n44313;
  assign n44315 = pi0199 & pi1139;
  assign n44316 = ~pi0200 & ~n43652;
  assign n44317 = ~n44315 & n44316;
  assign n44318 = ~n44314 & ~n44317;
  assign n44319 = n16479 & ~n44318;
  assign n44320 = pi0219 & n43712;
  assign n44321 = pi0211 & pi1138;
  assign n44322 = ~n44279 & ~n44321;
  assign n44323 = ~pi0219 & ~n44322;
  assign n44324 = ~n44320 & ~n44323;
  assign n44325 = ~n16479 & n44324;
  assign n44326 = ~n44319 & ~n44325;
  assign n44327 = pi0230 & ~n44326;
  assign n44328 = ~pi0830 & n40885;
  assign n44329 = pi0281 & ~n40885;
  assign n44330 = ~pi1091 & ~n44328;
  assign n44331 = ~n44329 & n44330;
  assign n44332 = pi1091 & ~n44322;
  assign n44333 = n40141 & ~n44332;
  assign n44334 = pi1138 & n40951;
  assign n44335 = ~n44289 & ~n44334;
  assign n44336 = n43500 & n44335;
  assign n44337 = ~n44333 & ~n44336;
  assign n44338 = ~n44331 & ~n44337;
  assign n44339 = ~pi0830 & n40863;
  assign n44340 = pi0281 & ~n40863;
  assign n44341 = ~pi1091 & ~n44339;
  assign n44342 = ~n44340 & n44341;
  assign n44343 = pi1139 & n42455;
  assign n44344 = n43686 & ~n44343;
  assign n44345 = pi0199 & ~n43719;
  assign n44346 = n16479 & n44345;
  assign n44347 = ~n44344 & ~n44346;
  assign n44348 = ~n44342 & ~n44347;
  assign n44349 = ~n44338 & ~n44348;
  assign n44350 = ~pi0230 & ~n44349;
  assign po0438 = ~n44327 & ~n44350;
  assign n44352 = pi0200 & ~n43733;
  assign n44353 = pi0199 & pi1140;
  assign n44354 = ~pi0200 & ~n44313;
  assign n44355 = ~n44353 & n44354;
  assign n44356 = ~n44352 & ~n44355;
  assign n44357 = n16479 & ~n44356;
  assign n44358 = pi0219 & n44129;
  assign n44359 = pi0211 & pi1139;
  assign n44360 = ~n43660 & ~n44359;
  assign n44361 = ~pi0219 & ~n44360;
  assign n44362 = ~n44358 & ~n44361;
  assign n44363 = ~n16479 & n44362;
  assign n44364 = ~n44357 & ~n44363;
  assign n44365 = pi0230 & ~n44364;
  assign n44366 = ~pi0836 & n40885;
  assign n44367 = pi0282 & ~n40885;
  assign n44368 = ~pi1091 & ~n44366;
  assign n44369 = ~n44367 & n44368;
  assign n44370 = pi1091 & ~n44360;
  assign n44371 = n40141 & ~n44370;
  assign n44372 = pi1139 & n40951;
  assign n44373 = ~n43689 & ~n44372;
  assign n44374 = n43500 & n44373;
  assign n44375 = ~n44371 & ~n44374;
  assign n44376 = ~n44369 & ~n44375;
  assign n44377 = ~pi0836 & n40863;
  assign n44378 = pi0282 & ~n40863;
  assign n44379 = ~pi1091 & ~n44377;
  assign n44380 = ~n44378 & n44379;
  assign n44381 = pi1140 & n42455;
  assign n44382 = n43686 & ~n44381;
  assign n44383 = ~pi0200 & n43717;
  assign n44384 = pi0199 & ~n44383;
  assign n44385 = n16479 & n44384;
  assign n44386 = ~n44382 & ~n44385;
  assign n44387 = ~n44380 & ~n44386;
  assign n44388 = ~n44376 & ~n44387;
  assign n44389 = ~pi0230 & ~n44388;
  assign po0439 = ~n44365 & ~n44389;
  assign n44391 = pi1147 & ~n43791;
  assign n44392 = pi1149 & ~n42389;
  assign n44393 = ~n44391 & ~n44392;
  assign n44394 = ~pi1148 & ~n44393;
  assign n44395 = n43884 & ~n44391;
  assign n44396 = pi1147 & ~n43501;
  assign n44397 = ~pi1149 & n43510;
  assign n44398 = ~n44396 & n44397;
  assign n44399 = pi1148 & ~n44395;
  assign n44400 = ~n44398 & n44399;
  assign n44401 = pi0230 & ~n44394;
  assign n44402 = ~n44400 & n44401;
  assign n44403 = ~pi1147 & n43637;
  assign n44404 = pi1147 & n43541;
  assign n44405 = pi1148 & ~n44404;
  assign n44406 = ~n44403 & n44405;
  assign n44407 = pi1147 & n43535;
  assign n44408 = ~pi1147 & ~n43633;
  assign n44409 = ~pi1148 & ~n44408;
  assign n44410 = ~n44407 & n44409;
  assign n44411 = ~pi1149 & ~n44406;
  assign n44412 = ~n44410 & n44411;
  assign n44413 = ~pi1147 & n43629;
  assign n44414 = pi1147 & n43580;
  assign n44415 = pi1148 & ~n44414;
  assign n44416 = ~n44413 & n44415;
  assign n44417 = ~pi1147 & n43623;
  assign n44418 = pi1147 & n43575;
  assign n44419 = ~pi1148 & ~n44417;
  assign n44420 = ~n44418 & n44419;
  assign n44421 = pi1149 & ~n44416;
  assign n44422 = ~n44420 & n44421;
  assign n44423 = pi0283 & ~n44412;
  assign n44424 = ~n44422 & n44423;
  assign n44425 = ~pi1147 & n43605;
  assign n44426 = pi1147 & n43586;
  assign n44427 = pi1149 & ~n44425;
  assign n44428 = ~n44426 & n44427;
  assign n44429 = ~pi1147 & ~n43562;
  assign n44430 = pi1147 & n43555;
  assign n44431 = ~pi1149 & ~n44429;
  assign n44432 = ~n44430 & n44431;
  assign n44433 = ~pi1148 & ~n44432;
  assign n44434 = ~n44428 & n44433;
  assign n44435 = ~pi1147 & n43608;
  assign n44436 = pi1147 & n43593;
  assign n44437 = pi1149 & ~n44436;
  assign n44438 = ~n44435 & n44437;
  assign n44439 = pi1147 & n43563;
  assign n44440 = ~pi1147 & ~n43614;
  assign n44441 = ~pi1149 & ~n44439;
  assign n44442 = ~n44440 & n44441;
  assign n44443 = pi1148 & ~n44438;
  assign n44444 = ~n44442 & n44443;
  assign n44445 = ~pi0283 & ~n44434;
  assign n44446 = ~n44444 & n44445;
  assign n44447 = ~pi0230 & ~n44424;
  assign n44448 = ~n44446 & n44447;
  assign po0440 = ~n44402 & ~n44448;
  assign n44450 = ~pi0284 & ~n42902;
  assign n44451 = pi1143 & n42902;
  assign n44452 = ~n40143 & n44451;
  assign po0441 = n44450 | n44452;
  assign n44454 = n2572 & ~n10399;
  assign n44455 = ~n7420 & n44454;
  assign n44456 = pi0286 & n44455;
  assign n44457 = pi0288 & pi0289;
  assign n44458 = n44456 & n44457;
  assign n44459 = pi0285 & n44458;
  assign n44460 = pi0285 & n44454;
  assign n44461 = ~n44458 & ~n44460;
  assign n44462 = ~po1038 & ~n44459;
  assign n44463 = ~n44461 & n44462;
  assign n44464 = ~po1038 & n44458;
  assign n44465 = ~pi0286 & n7420;
  assign n44466 = ~pi0288 & n44465;
  assign n44467 = ~pi0289 & n44466;
  assign n44468 = pi0285 & ~n44467;
  assign n44469 = ~n44464 & n44468;
  assign n44470 = ~n44463 & ~n44469;
  assign po0442 = ~pi0793 & ~n44470;
  assign n44472 = ~pi0288 & ~n7424;
  assign n44473 = n7420 & n44472;
  assign n44474 = pi0286 & ~n44473;
  assign n44475 = ~pi0286 & n44473;
  assign n44476 = po1038 & ~n44474;
  assign n44477 = ~n44475 & n44476;
  assign n44478 = n7420 & ~n44454;
  assign n44479 = pi0286 & ~n44478;
  assign n44480 = ~n44454 & n44465;
  assign n44481 = ~n44479 & ~n44480;
  assign n44482 = n44472 & ~n44481;
  assign n44483 = ~pi0286 & ~n44455;
  assign n44484 = pi0288 & ~n44456;
  assign n44485 = ~n44483 & n44484;
  assign n44486 = ~po1038 & ~n44482;
  assign n44487 = ~n44485 & n44486;
  assign n44488 = ~pi0793 & ~n44477;
  assign po0443 = ~n44487 & n44488;
  assign n44490 = ~pi0287 & pi0457;
  assign po0444 = ~pi0332 & ~n44490;
  assign n44492 = pi0288 & ~n7420;
  assign n44493 = ~n44473 & ~n44492;
  assign po0637 = ~po1038 & n44454;
  assign n44495 = ~n44493 & po0637;
  assign n44496 = n44493 & ~po0637;
  assign n44497 = ~pi0793 & ~n44495;
  assign po0445 = ~n44496 & n44497;
  assign n44499 = pi0289 & ~n44466;
  assign n44500 = pi0285 & ~pi0289;
  assign n44501 = n44466 & n44500;
  assign n44502 = po1038 & ~n44499;
  assign n44503 = ~n44501 & n44502;
  assign n44504 = ~pi0289 & n44484;
  assign n44505 = n44480 & n44500;
  assign n44506 = pi0289 & ~n44480;
  assign n44507 = ~pi0288 & ~n44505;
  assign n44508 = ~n44506 & n44507;
  assign n44509 = ~n44458 & ~n44504;
  assign n44510 = ~n44508 & n44509;
  assign n44511 = ~po1038 & ~n44510;
  assign n44512 = ~pi0793 & ~n44503;
  assign po0446 = ~n44511 & n44512;
  assign n44514 = ~pi0290 & pi0476;
  assign n44515 = ~pi0476 & ~pi1048;
  assign po0447 = ~n44514 & ~n44515;
  assign n44517 = ~pi0291 & pi0476;
  assign n44518 = ~pi0476 & ~pi1049;
  assign po0448 = ~n44517 & ~n44518;
  assign n44520 = ~pi0292 & pi0476;
  assign n44521 = ~pi0476 & ~pi1084;
  assign po0449 = ~n44520 & ~n44521;
  assign n44523 = ~pi0293 & pi0476;
  assign n44524 = ~pi0476 & ~pi1059;
  assign po0450 = ~n44523 & ~n44524;
  assign n44526 = ~pi0294 & pi0476;
  assign n44527 = ~pi0476 & ~pi1072;
  assign po0451 = ~n44526 & ~n44527;
  assign n44529 = ~pi0295 & pi0476;
  assign n44530 = ~pi0476 & ~pi1053;
  assign po0452 = ~n44529 & ~n44530;
  assign n44532 = ~pi0296 & pi0476;
  assign n44533 = ~pi0476 & ~pi1037;
  assign po0453 = ~n44532 & ~n44533;
  assign n44535 = ~pi0297 & pi0476;
  assign n44536 = ~pi0476 & ~pi1044;
  assign po0454 = ~n44535 & ~n44536;
  assign n44538 = ~pi0478 & pi1044;
  assign n44539 = pi0298 & pi0478;
  assign po0455 = n44538 | n44539;
  assign n44541 = pi0054 & n2521;
  assign n44542 = ~pi0054 & n13153;
  assign n44543 = n13411 & n44542;
  assign n44544 = ~n44541 & ~n44543;
  assign n44545 = n2621 & n8880;
  assign n44546 = ~n44544 & n44545;
  assign n44547 = ~pi0039 & ~n44546;
  assign po0456 = ~n11263 & ~n44547;
  assign n44549 = pi0057 & ~pi0059;
  assign n44550 = n10068 & n44549;
  assign n44551 = ~pi0312 & n44550;
  assign n44552 = pi0300 & ~n44551;
  assign n44553 = ~pi0300 & n44551;
  assign n44554 = ~pi0055 & ~n44553;
  assign po0457 = n44552 | ~n44554;
  assign n44556 = ~pi0301 & n44554;
  assign n44557 = ~pi0055 & pi0301;
  assign n44558 = n44553 & n44557;
  assign po0458 = n44556 | n44558;
  assign n44560 = n5836 & ~po1038;
  assign n44561 = ~pi0222 & ~pi0223;
  assign n44562 = pi0937 & ~n44561;
  assign n44563 = pi0273 & n3351;
  assign n44564 = ~n44562 & ~n44563;
  assign n44565 = n44560 & n44564;
  assign n44566 = ~n2603 & n44565;
  assign n44567 = n3449 & ~n16479;
  assign n44568 = ~n44565 & ~n44567;
  assign n44569 = pi0237 & ~n44568;
  assign n44570 = n5780 & ~n16479;
  assign n44571 = ~n44560 & ~n44570;
  assign n44572 = ~pi1148 & n44571;
  assign n44573 = ~pi0215 & n3310;
  assign n44574 = ~pi0273 & n44573;
  assign n44575 = pi0833 & n7570;
  assign n44576 = ~pi0937 & n44575;
  assign n44577 = ~n44574 & ~n44576;
  assign n44578 = ~n16479 & ~n44577;
  assign n44579 = ~n44566 & ~n44578;
  assign n44580 = ~n44569 & n44579;
  assign po0459 = ~n44572 & n44580;
  assign n44582 = ~pi0478 & pi1049;
  assign n44583 = pi0303 & pi0478;
  assign po0460 = n44582 | n44583;
  assign n44585 = ~pi0478 & pi1048;
  assign n44586 = pi0304 & pi0478;
  assign po0461 = n44585 | n44586;
  assign n44588 = ~pi0478 & pi1084;
  assign n44589 = pi0305 & pi0478;
  assign po0462 = n44588 | n44589;
  assign n44591 = ~pi0478 & pi1059;
  assign n44592 = pi0306 & pi0478;
  assign po0463 = n44591 | n44592;
  assign n44594 = ~pi0478 & pi1053;
  assign n44595 = pi0307 & pi0478;
  assign po0464 = n44594 | n44595;
  assign n44597 = ~pi0478 & pi1037;
  assign n44598 = pi0308 & pi0478;
  assign po0465 = n44597 | n44598;
  assign n44600 = ~pi0478 & pi1072;
  assign n44601 = pi0309 & pi0478;
  assign po0466 = n44600 | n44601;
  assign n44603 = pi1147 & n44571;
  assign n44604 = pi0222 & ~pi0934;
  assign n44605 = ~pi0271 & n3351;
  assign n44606 = ~n44604 & ~n44605;
  assign n44607 = n44560 & n44606;
  assign n44608 = ~n3448 & n44570;
  assign n44609 = pi0934 & ~n2526;
  assign n44610 = pi0271 & n3310;
  assign n44611 = ~n44609 & ~n44610;
  assign n44612 = n44608 & ~n44611;
  assign n44613 = ~n44567 & ~n44607;
  assign n44614 = ~n44612 & n44613;
  assign n44615 = ~n44603 & n44614;
  assign n44616 = ~pi0233 & ~n44615;
  assign n44617 = n2604 & n16479;
  assign n44618 = n44560 & ~n44606;
  assign n44619 = n44570 & n44611;
  assign n44620 = pi1147 & ~n44617;
  assign n44621 = ~n44618 & n44620;
  assign n44622 = ~n44619 & n44621;
  assign n44623 = ~n2603 & n44560;
  assign n44624 = ~n44608 & ~n44623;
  assign n44625 = ~pi1147 & ~n44624;
  assign n44626 = ~n44614 & n44625;
  assign n44627 = ~n44622 & ~n44626;
  assign n44628 = pi0233 & ~n44627;
  assign po0467 = n44616 | n44628;
  assign n44630 = ~pi0055 & ~pi0311;
  assign n44631 = ~n44558 & ~n44630;
  assign n44632 = ~pi0311 & n44558;
  assign po0468 = ~n44631 & ~n44632;
  assign n44634 = pi0312 & ~n44550;
  assign n44635 = ~n44551 & ~n44634;
  assign po0469 = ~pi0055 & ~n44635;
  assign n44637 = ~n10388 & ~n13446;
  assign n44638 = po0740 & ~n13453;
  assign n44639 = n10166 & ~n44638;
  assign po0634 = n44637 | ~n44639;
  assign n44641 = ~pi0954 & po0634;
  assign n44642 = pi0313 & pi0954;
  assign po0470 = ~n44641 & ~n44642;
  assign n44644 = n6323 & n8880;
  assign n44645 = n14440 & ~n44644;
  assign n44646 = pi0039 & ~n15297;
  assign n44647 = ~pi0039 & ~n14514;
  assign n44648 = n2608 & ~n44646;
  assign n44649 = ~n44647 & n44648;
  assign n44650 = ~n15333 & ~n44649;
  assign n44651 = n2534 & n10163;
  assign n44652 = ~n44650 & n44651;
  assign n44653 = ~n44645 & ~n44652;
  assign n44654 = n14432 & n14433;
  assign po0471 = ~n44653 & n44654;
  assign n44656 = ~pi0340 & n44454;
  assign n44657 = ~po1038 & n44656;
  assign n44658 = pi0315 & ~n44657;
  assign n44659 = pi1080 & n44657;
  assign po0472 = n44658 | n44659;
  assign n44661 = pi0316 & ~n44657;
  assign n44662 = pi1047 & n44657;
  assign po0473 = n44661 | n44662;
  assign n44664 = ~pi0330 & po0637;
  assign n44665 = pi0317 & ~n44664;
  assign n44666 = pi1078 & n44664;
  assign po0474 = n44665 | n44666;
  assign n44668 = ~pi0341 & n44454;
  assign n44669 = ~po1038 & n44668;
  assign n44670 = pi0318 & ~n44669;
  assign n44671 = pi1074 & n44669;
  assign po0475 = n44670 | n44671;
  assign n44673 = pi0319 & ~n44669;
  assign n44674 = pi1072 & n44669;
  assign po0476 = n44673 | n44674;
  assign n44676 = pi0320 & ~n44657;
  assign n44677 = pi1048 & n44657;
  assign po0477 = n44676 | n44677;
  assign n44679 = pi0321 & ~n44657;
  assign n44680 = pi1058 & n44657;
  assign po0478 = n44679 | n44680;
  assign n44682 = pi0322 & ~n44657;
  assign n44683 = pi1051 & n44657;
  assign po0479 = n44682 | n44683;
  assign n44685 = pi0323 & ~n44657;
  assign n44686 = pi1065 & n44657;
  assign po0480 = n44685 | n44686;
  assign n44688 = pi0324 & ~n44669;
  assign n44689 = pi1086 & n44669;
  assign po0481 = n44688 | n44689;
  assign n44691 = pi0325 & ~n44669;
  assign n44692 = pi1063 & n44669;
  assign po0482 = n44691 | n44692;
  assign n44694 = pi0326 & ~n44669;
  assign n44695 = pi1057 & n44669;
  assign po0483 = n44694 | n44695;
  assign n44697 = pi0327 & ~n44657;
  assign n44698 = pi1040 & n44657;
  assign po0484 = n44697 | n44698;
  assign n44700 = pi0328 & ~n44669;
  assign n44701 = pi1058 & n44669;
  assign po0485 = n44700 | n44701;
  assign n44703 = pi0329 & ~n44669;
  assign n44704 = pi1043 & n44669;
  assign po0486 = n44703 | n44704;
  assign n44706 = pi1092 & ~n2930;
  assign n44707 = po1038 & n44706;
  assign n44708 = ~pi0330 & n44707;
  assign n44709 = ~po1038 & n44706;
  assign n44710 = ~pi0330 & ~n44454;
  assign n44711 = ~n44656 & ~n44710;
  assign n44712 = n44709 & ~n44711;
  assign po0487 = n44708 | n44712;
  assign n44714 = ~pi0331 & n44707;
  assign n44715 = ~pi0331 & ~n44454;
  assign n44716 = ~n44668 & ~n44715;
  assign n44717 = n44709 & ~n44716;
  assign po0488 = n44714 | n44717;
  assign n44719 = n11002 & n13166;
  assign n44720 = ~n11002 & ~n13102;
  assign n44721 = n7445 & ~n44720;
  assign n44722 = ~pi0070 & ~n44721;
  assign n44723 = pi0332 & n9117;
  assign n44724 = ~n44722 & n44723;
  assign n44725 = ~n44719 & ~n44724;
  assign n44726 = ~pi0039 & ~n44725;
  assign n44727 = pi0039 & n10368;
  assign n44728 = ~pi0038 & ~n44727;
  assign n44729 = ~n44726 & n44728;
  assign po0489 = n38269 & ~n44729;
  assign n44731 = pi0333 & ~n44669;
  assign n44732 = pi1040 & n44669;
  assign po0490 = n44731 | n44732;
  assign n44734 = pi0334 & ~n44669;
  assign n44735 = pi1065 & n44669;
  assign po0491 = n44734 | n44735;
  assign n44737 = pi0335 & ~n44669;
  assign n44738 = pi1069 & n44669;
  assign po0492 = n44737 | n44738;
  assign n44740 = pi0336 & ~n44664;
  assign n44741 = pi1070 & n44664;
  assign po0493 = n44740 | n44741;
  assign n44743 = pi0337 & ~n44664;
  assign n44744 = pi1044 & n44664;
  assign po0494 = n44743 | n44744;
  assign n44746 = pi0338 & ~n44664;
  assign n44747 = pi1072 & n44664;
  assign po0495 = n44746 | n44747;
  assign n44749 = pi0339 & ~n44664;
  assign n44750 = pi1086 & n44664;
  assign po0496 = n44749 | n44750;
  assign n44752 = pi0340 & n44707;
  assign n44753 = ~pi0340 & ~n44454;
  assign n44754 = ~pi0331 & n44454;
  assign n44755 = n44709 & ~n44753;
  assign n44756 = ~n44754 & n44755;
  assign po0497 = ~n44752 & ~n44756;
  assign n44758 = ~pi0341 & ~po0637;
  assign n44759 = ~n44664 & ~n44758;
  assign po0498 = n44706 & ~n44759;
  assign n44761 = pi0342 & ~n44657;
  assign n44762 = pi1049 & n44657;
  assign po0499 = n44761 | n44762;
  assign n44764 = pi0343 & ~n44657;
  assign n44765 = pi1062 & n44657;
  assign po0500 = n44764 | n44765;
  assign n44767 = pi0344 & ~n44657;
  assign n44768 = pi1069 & n44657;
  assign po0501 = n44767 | n44768;
  assign n44770 = pi0345 & ~n44657;
  assign n44771 = pi1039 & n44657;
  assign po0502 = n44770 | n44771;
  assign n44773 = pi0346 & ~n44657;
  assign n44774 = pi1067 & n44657;
  assign po0503 = n44773 | n44774;
  assign n44776 = pi0347 & ~n44657;
  assign n44777 = pi1055 & n44657;
  assign po0504 = n44776 | n44777;
  assign n44779 = pi0348 & ~n44657;
  assign n44780 = pi1087 & n44657;
  assign po0505 = n44779 | n44780;
  assign n44782 = pi0349 & ~n44657;
  assign n44783 = pi1043 & n44657;
  assign po0506 = n44782 | n44783;
  assign n44785 = pi0350 & ~n44657;
  assign n44786 = pi1035 & n44657;
  assign po0507 = n44785 | n44786;
  assign n44788 = pi0351 & ~n44657;
  assign n44789 = pi1079 & n44657;
  assign po0508 = n44788 | n44789;
  assign n44791 = pi0352 & ~n44657;
  assign n44792 = pi1078 & n44657;
  assign po0509 = n44791 | n44792;
  assign n44794 = pi0353 & ~n44657;
  assign n44795 = pi1063 & n44657;
  assign po0510 = n44794 | n44795;
  assign n44797 = pi0354 & ~n44657;
  assign n44798 = pi1045 & n44657;
  assign po0511 = n44797 | n44798;
  assign n44800 = pi0355 & ~n44657;
  assign n44801 = pi1084 & n44657;
  assign po0512 = n44800 | n44801;
  assign n44803 = pi0356 & ~n44657;
  assign n44804 = pi1081 & n44657;
  assign po0513 = n44803 | n44804;
  assign n44806 = pi0357 & ~n44657;
  assign n44807 = pi1076 & n44657;
  assign po0514 = n44806 | n44807;
  assign n44809 = pi0358 & ~n44657;
  assign n44810 = pi1071 & n44657;
  assign po0515 = n44809 | n44810;
  assign n44812 = pi0359 & ~n44657;
  assign n44813 = pi1068 & n44657;
  assign po0516 = n44812 | n44813;
  assign n44815 = pi0360 & ~n44657;
  assign n44816 = pi1042 & n44657;
  assign po0517 = n44815 | n44816;
  assign n44818 = pi0361 & ~n44657;
  assign n44819 = pi1059 & n44657;
  assign po0518 = n44818 | n44819;
  assign n44821 = pi0362 & ~n44657;
  assign n44822 = pi1070 & n44657;
  assign po0519 = n44821 | n44822;
  assign n44824 = pi0363 & ~n44664;
  assign n44825 = pi1049 & n44664;
  assign po0520 = n44824 | n44825;
  assign n44827 = pi0364 & ~n44664;
  assign n44828 = pi1062 & n44664;
  assign po0521 = n44827 | n44828;
  assign n44830 = pi0365 & ~n44664;
  assign n44831 = pi1065 & n44664;
  assign po0522 = n44830 | n44831;
  assign n44833 = pi0366 & ~n44664;
  assign n44834 = pi1069 & n44664;
  assign po0523 = n44833 | n44834;
  assign n44836 = pi0367 & ~n44664;
  assign n44837 = pi1039 & n44664;
  assign po0524 = n44836 | n44837;
  assign n44839 = pi0368 & ~n44664;
  assign n44840 = pi1067 & n44664;
  assign po0525 = n44839 | n44840;
  assign n44842 = pi0369 & ~n44664;
  assign n44843 = pi1080 & n44664;
  assign po0526 = n44842 | n44843;
  assign n44845 = pi0370 & ~n44664;
  assign n44846 = pi1055 & n44664;
  assign po0527 = n44845 | n44846;
  assign n44848 = pi0371 & ~n44664;
  assign n44849 = pi1051 & n44664;
  assign po0528 = n44848 | n44849;
  assign n44851 = pi0372 & ~n44664;
  assign n44852 = pi1048 & n44664;
  assign po0529 = n44851 | n44852;
  assign n44854 = pi0373 & ~n44664;
  assign n44855 = pi1087 & n44664;
  assign po0530 = n44854 | n44855;
  assign n44857 = pi0374 & ~n44664;
  assign n44858 = pi1035 & n44664;
  assign po0531 = n44857 | n44858;
  assign n44860 = pi0375 & ~n44664;
  assign n44861 = pi1047 & n44664;
  assign po0532 = n44860 | n44861;
  assign n44863 = pi0376 & ~n44664;
  assign n44864 = pi1079 & n44664;
  assign po0533 = n44863 | n44864;
  assign n44866 = pi0377 & ~n44664;
  assign n44867 = pi1074 & n44664;
  assign po0534 = n44866 | n44867;
  assign n44869 = pi0378 & ~n44664;
  assign n44870 = pi1063 & n44664;
  assign po0535 = n44869 | n44870;
  assign n44872 = pi0379 & ~n44664;
  assign n44873 = pi1045 & n44664;
  assign po0536 = n44872 | n44873;
  assign n44875 = pi0380 & ~n44664;
  assign n44876 = pi1084 & n44664;
  assign po0537 = n44875 | n44876;
  assign n44878 = pi0381 & ~n44664;
  assign n44879 = pi1081 & n44664;
  assign po0538 = n44878 | n44879;
  assign n44881 = pi0382 & ~n44664;
  assign n44882 = pi1076 & n44664;
  assign po0539 = n44881 | n44882;
  assign n44884 = pi0383 & ~n44664;
  assign n44885 = pi1071 & n44664;
  assign po0540 = n44884 | n44885;
  assign n44887 = pi0384 & ~n44664;
  assign n44888 = pi1068 & n44664;
  assign po0541 = n44887 | n44888;
  assign n44890 = pi0385 & ~n44664;
  assign n44891 = pi1042 & n44664;
  assign po0542 = n44890 | n44891;
  assign n44893 = pi0386 & ~n44664;
  assign n44894 = pi1059 & n44664;
  assign po0543 = n44893 | n44894;
  assign n44896 = pi0387 & ~n44664;
  assign n44897 = pi1053 & n44664;
  assign po0544 = n44896 | n44897;
  assign n44899 = pi0388 & ~n44664;
  assign n44900 = pi1037 & n44664;
  assign po0545 = n44899 | n44900;
  assign n44902 = pi0389 & ~n44664;
  assign n44903 = pi1036 & n44664;
  assign po0546 = n44902 | n44903;
  assign n44905 = pi0390 & ~n44669;
  assign n44906 = pi1049 & n44669;
  assign po0547 = n44905 | n44906;
  assign n44908 = pi0391 & ~n44669;
  assign n44909 = pi1062 & n44669;
  assign po0548 = n44908 | n44909;
  assign n44911 = pi0392 & ~n44669;
  assign n44912 = pi1039 & n44669;
  assign po0549 = n44911 | n44912;
  assign n44914 = pi0393 & ~n44669;
  assign n44915 = pi1067 & n44669;
  assign po0550 = n44914 | n44915;
  assign n44917 = pi0394 & ~n44669;
  assign n44918 = pi1080 & n44669;
  assign po0551 = n44917 | n44918;
  assign n44920 = pi0395 & ~n44669;
  assign n44921 = pi1055 & n44669;
  assign po0552 = n44920 | n44921;
  assign n44923 = pi0396 & ~n44669;
  assign n44924 = pi1051 & n44669;
  assign po0553 = n44923 | n44924;
  assign n44926 = pi0397 & ~n44669;
  assign n44927 = pi1048 & n44669;
  assign po0554 = n44926 | n44927;
  assign n44929 = pi0398 & ~n44669;
  assign n44930 = pi1087 & n44669;
  assign po0555 = n44929 | n44930;
  assign n44932 = pi0399 & ~n44669;
  assign n44933 = pi1047 & n44669;
  assign po0556 = n44932 | n44933;
  assign n44935 = pi0400 & ~n44669;
  assign n44936 = pi1035 & n44669;
  assign po0557 = n44935 | n44936;
  assign n44938 = pi0401 & ~n44669;
  assign n44939 = pi1079 & n44669;
  assign po0558 = n44938 | n44939;
  assign n44941 = pi0402 & ~n44669;
  assign n44942 = pi1078 & n44669;
  assign po0559 = n44941 | n44942;
  assign n44944 = pi0403 & ~n44669;
  assign n44945 = pi1045 & n44669;
  assign po0560 = n44944 | n44945;
  assign n44947 = pi0404 & ~n44669;
  assign n44948 = pi1084 & n44669;
  assign po0561 = n44947 | n44948;
  assign n44950 = pi0405 & ~n44669;
  assign n44951 = pi1081 & n44669;
  assign po0562 = n44950 | n44951;
  assign n44953 = pi0406 & ~n44669;
  assign n44954 = pi1076 & n44669;
  assign po0563 = n44953 | n44954;
  assign n44956 = pi0407 & ~n44669;
  assign n44957 = pi1071 & n44669;
  assign po0564 = n44956 | n44957;
  assign n44959 = pi0408 & ~n44669;
  assign n44960 = pi1068 & n44669;
  assign po0565 = n44959 | n44960;
  assign n44962 = pi0409 & ~n44669;
  assign n44963 = pi1042 & n44669;
  assign po0566 = n44962 | n44963;
  assign n44965 = pi0410 & ~n44669;
  assign n44966 = pi1059 & n44669;
  assign po0567 = n44965 | n44966;
  assign n44968 = pi0411 & ~n44669;
  assign n44969 = pi1053 & n44669;
  assign po0568 = n44968 | n44969;
  assign n44971 = pi0412 & ~n44669;
  assign n44972 = pi1037 & n44669;
  assign po0569 = n44971 | n44972;
  assign n44974 = pi0413 & ~n44669;
  assign n44975 = pi1036 & n44669;
  assign po0570 = n44974 | n44975;
  assign n44977 = ~po1038 & n44754;
  assign n44978 = pi0414 & ~n44977;
  assign n44979 = pi1049 & n44977;
  assign po0571 = n44978 | n44979;
  assign n44981 = pi0415 & ~n44977;
  assign n44982 = pi1062 & n44977;
  assign po0572 = n44981 | n44982;
  assign n44984 = pi0416 & ~n44977;
  assign n44985 = pi1069 & n44977;
  assign po0573 = n44984 | n44985;
  assign n44987 = pi0417 & ~n44977;
  assign n44988 = pi1039 & n44977;
  assign po0574 = n44987 | n44988;
  assign n44990 = pi0418 & ~n44977;
  assign n44991 = pi1067 & n44977;
  assign po0575 = n44990 | n44991;
  assign n44993 = pi0419 & ~n44977;
  assign n44994 = pi1080 & n44977;
  assign po0576 = n44993 | n44994;
  assign n44996 = pi0420 & ~n44977;
  assign n44997 = pi1055 & n44977;
  assign po0577 = n44996 | n44997;
  assign n44999 = pi0421 & ~n44977;
  assign n45000 = pi1051 & n44977;
  assign po0578 = n44999 | n45000;
  assign n45002 = pi0422 & ~n44977;
  assign n45003 = pi1048 & n44977;
  assign po0579 = n45002 | n45003;
  assign n45005 = pi0423 & ~n44977;
  assign n45006 = pi1087 & n44977;
  assign po0580 = n45005 | n45006;
  assign n45008 = pi0424 & ~n44977;
  assign n45009 = pi1047 & n44977;
  assign po0581 = n45008 | n45009;
  assign n45011 = pi0425 & ~n44977;
  assign n45012 = pi1035 & n44977;
  assign po0582 = n45011 | n45012;
  assign n45014 = pi0426 & ~n44977;
  assign n45015 = pi1079 & n44977;
  assign po0583 = n45014 | n45015;
  assign n45017 = pi0427 & ~n44977;
  assign n45018 = pi1078 & n44977;
  assign po0584 = n45017 | n45018;
  assign n45020 = pi0428 & ~n44977;
  assign n45021 = pi1045 & n44977;
  assign po0585 = n45020 | n45021;
  assign n45023 = pi0429 & ~n44977;
  assign n45024 = pi1084 & n44977;
  assign po0586 = n45023 | n45024;
  assign n45026 = pi0430 & ~n44977;
  assign n45027 = pi1076 & n44977;
  assign po0587 = n45026 | n45027;
  assign n45029 = pi0431 & ~n44977;
  assign n45030 = pi1071 & n44977;
  assign po0588 = n45029 | n45030;
  assign n45032 = pi0432 & ~n44977;
  assign n45033 = pi1068 & n44977;
  assign po0589 = n45032 | n45033;
  assign n45035 = pi0433 & ~n44977;
  assign n45036 = pi1042 & n44977;
  assign po0590 = n45035 | n45036;
  assign n45038 = pi0434 & ~n44977;
  assign n45039 = pi1059 & n44977;
  assign po0591 = n45038 | n45039;
  assign n45041 = pi0435 & ~n44977;
  assign n45042 = pi1053 & n44977;
  assign po0592 = n45041 | n45042;
  assign n45044 = pi0436 & ~n44977;
  assign n45045 = pi1037 & n44977;
  assign po0593 = n45044 | n45045;
  assign n45047 = pi0437 & ~n44977;
  assign n45048 = pi1070 & n44977;
  assign po0594 = n45047 | n45048;
  assign n45050 = pi0438 & ~n44977;
  assign n45051 = pi1036 & n44977;
  assign po0595 = n45050 | n45051;
  assign n45053 = pi0439 & ~n44664;
  assign n45054 = pi1057 & n44664;
  assign po0596 = n45053 | n45054;
  assign n45056 = pi0440 & ~n44664;
  assign n45057 = pi1043 & n44664;
  assign po0597 = n45056 | n45057;
  assign n45059 = pi0441 & ~n44657;
  assign n45060 = pi1044 & n44657;
  assign po0598 = n45059 | n45060;
  assign n45062 = pi0442 & ~n44664;
  assign n45063 = pi1058 & n44664;
  assign po0599 = n45062 | n45063;
  assign n45065 = pi0443 & ~n44977;
  assign n45066 = pi1044 & n44977;
  assign po0600 = n45065 | n45066;
  assign n45068 = pi0444 & ~n44977;
  assign n45069 = pi1072 & n44977;
  assign po0601 = n45068 | n45069;
  assign n45071 = pi0445 & ~n44977;
  assign n45072 = pi1081 & n44977;
  assign po0602 = n45071 | n45072;
  assign n45074 = pi0446 & ~n44977;
  assign n45075 = pi1086 & n44977;
  assign po0603 = n45074 | n45075;
  assign n45077 = pi0447 & ~n44664;
  assign n45078 = pi1040 & n44664;
  assign po0604 = n45077 | n45078;
  assign n45080 = pi0448 & ~n44977;
  assign n45081 = pi1074 & n44977;
  assign po0605 = n45080 | n45081;
  assign n45083 = pi0449 & ~n44977;
  assign n45084 = pi1057 & n44977;
  assign po0606 = n45083 | n45084;
  assign n45086 = pi0450 & ~n44657;
  assign n45087 = pi1036 & n44657;
  assign po0607 = n45086 | n45087;
  assign n45089 = pi0451 & ~n44977;
  assign n45090 = pi1063 & n44977;
  assign po0608 = n45089 | n45090;
  assign n45092 = pi0452 & ~n44657;
  assign n45093 = pi1053 & n44657;
  assign po0609 = n45092 | n45093;
  assign n45095 = pi0453 & ~n44977;
  assign n45096 = pi1040 & n44977;
  assign po0610 = n45095 | n45096;
  assign n45098 = pi0454 & ~n44977;
  assign n45099 = pi1043 & n44977;
  assign po0611 = n45098 | n45099;
  assign n45101 = pi0455 & ~n44657;
  assign n45102 = pi1037 & n44657;
  assign po0612 = n45101 | n45102;
  assign n45104 = pi0456 & ~n44669;
  assign n45105 = pi1044 & n44669;
  assign po0613 = n45104 | n45105;
  assign n45107 = pi0594 & pi0600;
  assign n45108 = pi0597 & n45107;
  assign n45109 = pi0601 & n45108;
  assign n45110 = ~pi0804 & ~pi0810;
  assign n45111 = ~pi0595 & n45110;
  assign n45112 = ~pi0599 & pi0810;
  assign n45113 = pi0596 & ~n45112;
  assign n45114 = pi0804 & ~n45113;
  assign n45115 = pi0595 & pi0815;
  assign n45116 = ~n45114 & n45115;
  assign n45117 = ~n45111 & ~n45116;
  assign n45118 = n45109 & ~n45117;
  assign n45119 = pi0600 & ~pi0810;
  assign n45120 = pi0804 & ~n45119;
  assign n45121 = ~pi0601 & ~n45110;
  assign n45122 = ~pi0815 & ~n45120;
  assign n45123 = ~n45121 & n45122;
  assign n45124 = ~n45118 & ~n45123;
  assign n45125 = pi0605 & ~n45124;
  assign n45126 = pi0990 & n45107;
  assign n45127 = ~pi0815 & n45120;
  assign n45128 = n45126 & n45127;
  assign n45129 = ~n45125 & ~n45128;
  assign po0614 = pi0821 & ~n45129;
  assign n45131 = pi0458 & ~n44657;
  assign n45132 = pi1072 & n44657;
  assign po0615 = n45131 | n45132;
  assign n45134 = pi0459 & ~n44977;
  assign n45135 = pi1058 & n44977;
  assign po0616 = n45134 | n45135;
  assign n45137 = pi0460 & ~n44657;
  assign n45138 = pi1086 & n44657;
  assign po0617 = n45137 | n45138;
  assign n45140 = pi0461 & ~n44657;
  assign n45141 = pi1057 & n44657;
  assign po0618 = n45140 | n45141;
  assign n45143 = pi0462 & ~n44657;
  assign n45144 = pi1074 & n44657;
  assign po0619 = n45143 | n45144;
  assign n45146 = pi0463 & ~n44669;
  assign n45147 = pi1070 & n44669;
  assign po0620 = n45146 | n45147;
  assign n45149 = pi0464 & ~n44977;
  assign n45150 = pi1065 & n44977;
  assign po0621 = n45149 | n45150;
  assign n45152 = ~pi0299 & n44561;
  assign n45153 = ~n11423 & ~n45152;
  assign n45154 = ~n11396 & ~n11399;
  assign n45155 = ~pi0243 & ~n45154;
  assign n45156 = ~pi0243 & pi1157;
  assign n45157 = ~n45153 & ~n45156;
  assign n45158 = ~n45155 & n45157;
  assign n45159 = ~n3471 & ~n11424;
  assign n45160 = pi0926 & n45156;
  assign n45161 = ~n45159 & n45160;
  assign n45162 = ~n5836 & ~n5854;
  assign n45163 = pi0926 & ~n45162;
  assign n45164 = pi1157 & n45162;
  assign n45165 = ~n45155 & ~n45163;
  assign n45166 = ~n45164 & n45165;
  assign n45167 = ~n45158 & ~n45161;
  assign n45168 = ~n45166 & n45167;
  assign n45169 = ~po1038 & ~n45168;
  assign n45170 = ~pi0243 & n44573;
  assign n45171 = pi0926 & n44575;
  assign n45172 = pi1157 & ~n5780;
  assign n45173 = po1038 & ~n45170;
  assign n45174 = ~n45171 & ~n45172;
  assign n45175 = n45173 & n45174;
  assign po0622 = ~n45169 & ~n45175;
  assign n45177 = po1038 & ~n44573;
  assign n45178 = ~po1038 & n45154;
  assign n45179 = ~n45177 & ~n45178;
  assign n45180 = ~pi0943 & ~n45179;
  assign n45181 = ~n44571 & n45180;
  assign n45182 = pi0943 & n44624;
  assign n45183 = ~n45180 & ~n45182;
  assign n45184 = ~pi1151 & ~n45183;
  assign n45185 = ~po1038 & ~n45153;
  assign n45186 = n2526 & po1038;
  assign n45187 = ~n45185 & ~n45186;
  assign n45188 = ~pi0275 & ~n45187;
  assign n45189 = ~n44567 & ~n44617;
  assign n45190 = pi0943 & pi1151;
  assign n45191 = ~n45189 & n45190;
  assign n45192 = ~n45181 & ~n45188;
  assign n45193 = ~n45191 & n45192;
  assign po0623 = ~n45184 & n45193;
  assign n45195 = pi0040 & ~pi0287;
  assign n45196 = n42346 & n45195;
  assign n45197 = po0950 & n45196;
  assign n45198 = ~n10165 & ~n45197;
  assign n45199 = ~pi0102 & ~n13381;
  assign n45200 = n8897 & n10162;
  assign n45201 = n16847 & n45200;
  assign n45202 = ~n45199 & n45201;
  assign n45203 = n16845 & n45202;
  assign n45204 = n45196 & ~n45203;
  assign n45205 = ~n45196 & n45203;
  assign n45206 = ~n45204 & ~n45205;
  assign n45207 = n7490 & ~n45206;
  assign n45208 = ~n6277 & ~n45206;
  assign n45209 = n6277 & n45203;
  assign n45210 = ~n45208 & ~n45209;
  assign n45211 = ~n7490 & ~n45210;
  assign n45212 = pi1091 & ~n45207;
  assign n45213 = ~n45211 & n45212;
  assign n45214 = ~pi1093 & ~n45210;
  assign n45215 = ~n7417 & ~n45206;
  assign n45216 = n7417 & n45203;
  assign n45217 = ~n45215 & ~n45216;
  assign n45218 = pi1093 & ~n45217;
  assign n45219 = ~pi1091 & ~n45214;
  assign n45220 = ~n45218 & n45219;
  assign n45221 = ~n45213 & ~n45220;
  assign n45222 = n2610 & n44644;
  assign n45223 = ~n45221 & n45222;
  assign po0624 = ~n45198 & ~n45223;
  assign n45225 = n10200 & n11337;
  assign n45226 = pi0038 & ~pi0039;
  assign n45227 = n10197 & n45226;
  assign n45228 = n8962 & n45227;
  assign n45229 = pi0468 & ~n45228;
  assign po0625 = n45225 | n45229;
  assign n45231 = ~pi0263 & ~n45154;
  assign n45232 = ~pi0263 & pi1156;
  assign n45233 = ~n45153 & ~n45232;
  assign n45234 = ~n45231 & n45233;
  assign n45235 = pi0942 & n45232;
  assign n45236 = ~n45159 & n45235;
  assign n45237 = pi0942 & ~n45162;
  assign n45238 = pi1156 & n45162;
  assign n45239 = ~n45231 & ~n45237;
  assign n45240 = ~n45238 & n45239;
  assign n45241 = ~n45234 & ~n45236;
  assign n45242 = ~n45240 & n45241;
  assign n45243 = ~po1038 & ~n45242;
  assign n45244 = pi1156 & ~n5780;
  assign n45245 = pi0942 & n44575;
  assign n45246 = ~pi0263 & n44573;
  assign n45247 = po1038 & ~n45246;
  assign n45248 = ~n45244 & ~n45245;
  assign n45249 = n45247 & n45248;
  assign po0626 = ~n45243 & ~n45249;
  assign n45251 = pi0267 & ~n45154;
  assign n45252 = pi0267 & pi1155;
  assign n45253 = ~n45153 & ~n45252;
  assign n45254 = ~n45251 & n45253;
  assign n45255 = pi0925 & n45252;
  assign n45256 = ~n45159 & n45255;
  assign n45257 = pi0925 & ~n45162;
  assign n45258 = pi1155 & n45162;
  assign n45259 = ~n45251 & ~n45257;
  assign n45260 = ~n45258 & n45259;
  assign n45261 = ~n45254 & ~n45256;
  assign n45262 = ~n45260 & n45261;
  assign n45263 = ~po1038 & ~n45262;
  assign n45264 = pi1155 & ~n5780;
  assign n45265 = pi0925 & n44575;
  assign n45266 = pi0267 & n44573;
  assign n45267 = po1038 & ~n45266;
  assign n45268 = ~n45264 & ~n45265;
  assign n45269 = n45267 & n45268;
  assign po0627 = ~n45263 & ~n45269;
  assign n45271 = pi0253 & ~n45154;
  assign n45272 = pi0253 & pi1153;
  assign n45273 = ~n45153 & ~n45272;
  assign n45274 = ~n45271 & n45273;
  assign n45275 = pi0941 & n45272;
  assign n45276 = ~n45159 & n45275;
  assign n45277 = pi0941 & ~n45162;
  assign n45278 = pi1153 & n45162;
  assign n45279 = ~n45271 & ~n45277;
  assign n45280 = ~n45278 & n45279;
  assign n45281 = ~n45274 & ~n45276;
  assign n45282 = ~n45280 & n45281;
  assign n45283 = ~po1038 & ~n45282;
  assign n45284 = pi1153 & ~n5780;
  assign n45285 = pi0941 & n44575;
  assign n45286 = pi0253 & n44573;
  assign n45287 = po1038 & ~n45286;
  assign n45288 = ~n45284 & ~n45285;
  assign n45289 = n45287 & n45288;
  assign po0628 = ~n45283 & ~n45289;
  assign n45291 = pi0254 & ~n45154;
  assign n45292 = pi0254 & pi1154;
  assign n45293 = ~n45153 & ~n45292;
  assign n45294 = ~n45291 & n45293;
  assign n45295 = pi0923 & n45292;
  assign n45296 = ~n45159 & n45295;
  assign n45297 = pi0923 & ~n45162;
  assign n45298 = pi1154 & n45162;
  assign n45299 = ~n45291 & ~n45297;
  assign n45300 = ~n45298 & n45299;
  assign n45301 = ~n45294 & ~n45296;
  assign n45302 = ~n45300 & n45301;
  assign n45303 = ~po1038 & ~n45302;
  assign n45304 = pi1154 & ~n5780;
  assign n45305 = pi0923 & n44575;
  assign n45306 = pi0254 & n44573;
  assign n45307 = po1038 & ~n45306;
  assign n45308 = ~n45304 & ~n45305;
  assign n45309 = n45307 & n45308;
  assign po0629 = ~n45303 & ~n45309;
  assign n45311 = ~pi0922 & ~n45179;
  assign n45312 = ~n44571 & n45311;
  assign n45313 = pi0922 & n44624;
  assign n45314 = ~n45311 & ~n45313;
  assign n45315 = ~pi1152 & ~n45314;
  assign n45316 = ~pi0268 & ~n45187;
  assign n45317 = pi0922 & pi1152;
  assign n45318 = ~n45189 & n45317;
  assign n45319 = ~n45312 & ~n45316;
  assign n45320 = ~n45318 & n45319;
  assign po0630 = ~n45315 & n45320;
  assign n45322 = ~pi0931 & ~n45179;
  assign n45323 = ~n44571 & n45322;
  assign n45324 = pi0931 & n44624;
  assign n45325 = ~n45322 & ~n45324;
  assign n45326 = ~pi1150 & ~n45325;
  assign n45327 = ~pi0272 & ~n45187;
  assign n45328 = pi0931 & pi1150;
  assign n45329 = ~n45189 & n45328;
  assign n45330 = ~n45323 & ~n45327;
  assign n45331 = ~n45329 & n45330;
  assign po0631 = ~n45326 & n45331;
  assign n45333 = ~pi0936 & ~n45179;
  assign n45334 = ~n44571 & n45333;
  assign n45335 = pi0936 & n44624;
  assign n45336 = ~n45333 & ~n45335;
  assign n45337 = ~pi1149 & ~n45336;
  assign n45338 = ~pi0283 & ~n45187;
  assign n45339 = pi0936 & pi1149;
  assign n45340 = ~n45189 & n45339;
  assign n45341 = ~n45334 & ~n45338;
  assign n45342 = ~n45340 & n45341;
  assign po0632 = ~n45337 & n45342;
  assign n45344 = pi0071 & n43509;
  assign n45345 = pi0071 & ~n11448;
  assign n45346 = n11448 & n13052;
  assign n45347 = n10150 & ~n11448;
  assign n45348 = n10147 & n45347;
  assign n45349 = ~n45346 & ~n45348;
  assign n45350 = n2572 & n10162;
  assign n45351 = ~n45349 & n45350;
  assign n45352 = n13050 & n45351;
  assign n45353 = ~n45345 & ~n45352;
  assign n45354 = ~po1038 & ~n45353;
  assign po0633 = n45344 | n45354;
  assign po0635 = pi0071 & ~n43791;
  assign n45357 = pi0481 & ~n34775;
  assign n45358 = pi0248 & n34775;
  assign po0638 = n45357 | n45358;
  assign n45360 = pi0482 & ~n34791;
  assign n45361 = pi0249 & n34791;
  assign po0639 = n45360 | n45361;
  assign n45363 = pi0483 & ~n34915;
  assign n45364 = pi0242 & n34915;
  assign po0640 = n45363 | n45364;
  assign n45366 = pi0484 & ~n34915;
  assign n45367 = pi0249 & n34915;
  assign po0641 = n45366 | n45367;
  assign n45369 = pi0485 & ~n36111;
  assign n45370 = pi0234 & n36111;
  assign po0642 = n45369 | n45370;
  assign n45372 = pi0486 & ~n36111;
  assign n45373 = pi0244 & n36111;
  assign po0643 = n45372 | n45373;
  assign n45375 = pi0487 & ~n34775;
  assign n45376 = pi0246 & n34775;
  assign po0644 = n45375 | n45376;
  assign n45378 = pi0488 & ~n34775;
  assign n45379 = ~pi0239 & n34775;
  assign po0645 = ~n45378 & ~n45379;
  assign n45381 = pi0489 & ~n36111;
  assign n45382 = pi0242 & n36111;
  assign po0646 = n45381 | n45382;
  assign n45384 = pi0490 & ~n34915;
  assign n45385 = pi0241 & n34915;
  assign po0647 = n45384 | n45385;
  assign n45387 = pi0491 & ~n34915;
  assign n45388 = pi0238 & n34915;
  assign po0648 = n45387 | n45388;
  assign n45390 = pi0492 & ~n34915;
  assign n45391 = pi0240 & n34915;
  assign po0649 = n45390 | n45391;
  assign n45393 = pi0493 & ~n34915;
  assign n45394 = pi0244 & n34915;
  assign po0650 = n45393 | n45394;
  assign n45396 = pi0494 & ~n34915;
  assign n45397 = ~pi0239 & n34915;
  assign po0651 = ~n45396 & ~n45397;
  assign n45399 = pi0495 & ~n34915;
  assign n45400 = pi0235 & n34915;
  assign po0652 = n45399 | n45400;
  assign n45402 = pi0496 & ~n34907;
  assign n45403 = pi0249 & n34907;
  assign po0653 = n45402 | n45403;
  assign n45405 = pi0497 & ~n34907;
  assign n45406 = ~pi0239 & n34907;
  assign po0654 = ~n45405 & ~n45406;
  assign n45408 = pi0498 & ~n34791;
  assign n45409 = pi0238 & n34791;
  assign po0655 = n45408 | n45409;
  assign n45411 = pi0499 & ~n34907;
  assign n45412 = pi0246 & n34907;
  assign po0656 = n45411 | n45412;
  assign n45414 = pi0500 & ~n34907;
  assign n45415 = pi0241 & n34907;
  assign po0657 = n45414 | n45415;
  assign n45417 = pi0501 & ~n34907;
  assign n45418 = pi0248 & n34907;
  assign po0658 = n45417 | n45418;
  assign n45420 = pi0502 & ~n34907;
  assign n45421 = pi0247 & n34907;
  assign po0659 = n45420 | n45421;
  assign n45423 = pi0503 & ~n34907;
  assign n45424 = pi0245 & n34907;
  assign po0660 = n45423 | n45424;
  assign n45426 = pi0504 & ~n34900;
  assign n45427 = pi0242 & n34900;
  assign po0661 = n45426 | n45427;
  assign n45429 = ~n6326 & n16479;
  assign n45430 = ~n34895 & ~n45429;
  assign n45431 = ~pi0234 & n45430;
  assign n45432 = n34907 & n45431;
  assign n45433 = pi0505 & ~n45432;
  assign n45434 = pi0234 & n34899;
  assign n45435 = ~pi0505 & n34778;
  assign n45436 = n45434 & n45435;
  assign po0662 = n45433 | n45436;
  assign n45438 = pi0506 & ~n34900;
  assign n45439 = pi0241 & n34900;
  assign po0663 = n45438 | n45439;
  assign n45441 = pi0507 & ~n34900;
  assign n45442 = pi0238 & n34900;
  assign po0664 = n45441 | n45442;
  assign n45444 = pi0508 & ~n34900;
  assign n45445 = pi0247 & n34900;
  assign po0665 = n45444 | n45445;
  assign n45447 = pi0509 & ~n34900;
  assign n45448 = pi0245 & n34900;
  assign po0666 = n45447 | n45448;
  assign n45450 = pi0510 & ~n34775;
  assign n45451 = pi0242 & n34775;
  assign po0667 = n45450 | n45451;
  assign n45453 = n6584 & ~po1038;
  assign n45454 = ~n34769 & ~n45453;
  assign n45455 = ~pi0234 & n45454;
  assign n45456 = n34775 & ~n45455;
  assign n45457 = pi0511 & ~n34775;
  assign po0668 = n45456 | n45457;
  assign n45459 = pi0512 & ~n34775;
  assign n45460 = pi0235 & n34775;
  assign po0669 = n45459 | n45460;
  assign n45462 = pi0513 & ~n34775;
  assign n45463 = pi0244 & n34775;
  assign po0670 = n45462 | n45463;
  assign n45465 = pi0514 & ~n34775;
  assign n45466 = pi0245 & n34775;
  assign po0671 = n45465 | n45466;
  assign n45468 = pi0515 & ~n34775;
  assign n45469 = pi0240 & n34775;
  assign po0672 = n45468 | n45469;
  assign n45471 = pi0516 & ~n34775;
  assign n45472 = pi0247 & n34775;
  assign po0673 = n45471 | n45472;
  assign n45474 = pi0517 & ~n34775;
  assign n45475 = pi0238 & n34775;
  assign po0674 = n45474 | n45475;
  assign n45477 = n34783 & n45455;
  assign n45478 = pi0518 & ~n45477;
  assign n45479 = pi0234 & n34774;
  assign n45480 = ~pi0518 & n34778;
  assign n45481 = n45479 & n45480;
  assign po0675 = n45478 | n45481;
  assign n45483 = pi0519 & ~n34783;
  assign n45484 = ~pi0239 & n34783;
  assign po0676 = ~n45483 & ~n45484;
  assign n45486 = pi0520 & ~n34783;
  assign n45487 = pi0246 & n34783;
  assign po0677 = n45486 | n45487;
  assign n45489 = pi0521 & ~n34783;
  assign n45490 = pi0248 & n34783;
  assign po0678 = n45489 | n45490;
  assign n45492 = pi0522 & ~n34783;
  assign n45493 = pi0238 & n34783;
  assign po0679 = n45492 | n45493;
  assign n45495 = n36139 & n45455;
  assign n45496 = pi0523 & ~n45495;
  assign n45497 = ~pi0523 & n34910;
  assign n45498 = n45479 & n45497;
  assign po0680 = n45496 | n45498;
  assign n45500 = pi0524 & ~n36139;
  assign n45501 = ~pi0239 & n36139;
  assign po0681 = ~n45500 & ~n45501;
  assign n45503 = pi0525 & ~n36139;
  assign n45504 = pi0245 & n36139;
  assign po0682 = n45503 | n45504;
  assign n45506 = pi0526 & ~n36139;
  assign n45507 = pi0246 & n36139;
  assign po0683 = n45506 | n45507;
  assign n45509 = pi0527 & ~n36139;
  assign n45510 = pi0247 & n36139;
  assign po0684 = n45509 | n45510;
  assign n45512 = pi0528 & ~n36139;
  assign n45513 = pi0249 & n36139;
  assign po0685 = n45512 | n45513;
  assign n45515 = pi0529 & ~n36139;
  assign n45516 = pi0238 & n36139;
  assign po0686 = n45515 | n45516;
  assign n45518 = pi0530 & ~n36139;
  assign n45519 = pi0240 & n36139;
  assign po0687 = n45518 | n45519;
  assign n45521 = pi0531 & ~n34791;
  assign n45522 = pi0235 & n34791;
  assign po0688 = n45521 | n45522;
  assign n45524 = pi0532 & ~n34791;
  assign n45525 = pi0247 & n34791;
  assign po0689 = n45524 | n45525;
  assign n45527 = pi0533 & ~n34900;
  assign n45528 = pi0235 & n34900;
  assign po0690 = n45527 | n45528;
  assign n45530 = pi0534 & ~n34900;
  assign n45531 = ~pi0239 & n34900;
  assign po0691 = ~n45530 & ~n45531;
  assign n45533 = pi0535 & ~n34900;
  assign n45534 = pi0240 & n34900;
  assign po0692 = n45533 | n45534;
  assign n45536 = pi0536 & ~n34900;
  assign n45537 = pi0246 & n34900;
  assign po0693 = n45536 | n45537;
  assign n45539 = pi0537 & ~n34900;
  assign n45540 = pi0248 & n34900;
  assign po0694 = n45539 | n45540;
  assign n45542 = pi0538 & ~n34900;
  assign n45543 = pi0249 & n34900;
  assign po0695 = n45542 | n45543;
  assign n45545 = pi0539 & ~n34907;
  assign n45546 = pi0242 & n34907;
  assign po0696 = n45545 | n45546;
  assign n45548 = pi0540 & ~n34907;
  assign n45549 = pi0235 & n34907;
  assign po0697 = n45548 | n45549;
  assign n45551 = pi0541 & ~n34907;
  assign n45552 = pi0244 & n34907;
  assign po0698 = n45551 | n45552;
  assign n45554 = pi0542 & ~n34907;
  assign n45555 = pi0240 & n34907;
  assign po0699 = n45554 | n45555;
  assign n45557 = pi0543 & ~n34907;
  assign n45558 = pi0238 & n34907;
  assign po0700 = n45557 | n45558;
  assign n45560 = n34915 & n45431;
  assign n45561 = pi0544 & ~n45560;
  assign n45562 = ~pi0544 & n34910;
  assign n45563 = n45434 & n45562;
  assign po0701 = n45561 | n45563;
  assign n45565 = pi0545 & ~n34915;
  assign n45566 = pi0245 & n34915;
  assign po0702 = n45565 | n45566;
  assign n45568 = pi0546 & ~n34915;
  assign n45569 = pi0246 & n34915;
  assign po0703 = n45568 | n45569;
  assign n45571 = pi0547 & ~n34915;
  assign n45572 = pi0247 & n34915;
  assign po0704 = n45571 | n45572;
  assign n45574 = pi0548 & ~n34915;
  assign n45575 = pi0248 & n34915;
  assign po0705 = n45574 | n45575;
  assign n45577 = pi0549 & ~n36111;
  assign n45578 = pi0235 & n36111;
  assign po0706 = n45577 | n45578;
  assign n45580 = pi0550 & ~n36111;
  assign n45581 = ~pi0239 & n36111;
  assign po0707 = ~n45580 & ~n45581;
  assign n45583 = pi0551 & ~n36111;
  assign n45584 = pi0240 & n36111;
  assign po0708 = n45583 | n45584;
  assign n45586 = pi0552 & ~n36111;
  assign n45587 = pi0247 & n36111;
  assign po0709 = n45586 | n45587;
  assign n45589 = pi0553 & ~n36111;
  assign n45590 = pi0241 & n36111;
  assign po0710 = n45589 | n45590;
  assign n45592 = pi0554 & ~n36111;
  assign n45593 = pi0248 & n36111;
  assign po0711 = n45592 | n45593;
  assign n45595 = pi0555 & ~n36111;
  assign n45596 = pi0249 & n36111;
  assign po0712 = n45595 | n45596;
  assign n45598 = pi0556 & ~n34791;
  assign n45599 = pi0242 & n34791;
  assign po0713 = n45598 | n45599;
  assign n45601 = n34900 & n45431;
  assign n45602 = pi0557 & ~n45601;
  assign n45603 = ~pi0557 & n34583;
  assign n45604 = n45434 & n45603;
  assign po0714 = n45602 | n45604;
  assign n45606 = pi0558 & ~n34900;
  assign n45607 = pi0244 & n34900;
  assign po0715 = n45606 | n45607;
  assign n45609 = pi0559 & ~n34775;
  assign n45610 = pi0241 & n34775;
  assign po0716 = n45609 | n45610;
  assign n45612 = pi0560 & ~n34791;
  assign n45613 = pi0240 & n34791;
  assign po0717 = n45612 | n45613;
  assign n45615 = pi0561 & ~n34783;
  assign n45616 = pi0247 & n34783;
  assign po0718 = n45615 | n45616;
  assign n45618 = pi0562 & ~n34791;
  assign n45619 = pi0241 & n34791;
  assign po0719 = n45618 | n45619;
  assign n45621 = pi0563 & ~n36111;
  assign n45622 = pi0246 & n36111;
  assign po0720 = n45621 | n45622;
  assign n45624 = pi0564 & ~n34791;
  assign n45625 = pi0246 & n34791;
  assign po0721 = n45624 | n45625;
  assign n45627 = pi0565 & ~n34791;
  assign n45628 = pi0248 & n34791;
  assign po0722 = n45627 | n45628;
  assign n45630 = pi0566 & ~n34791;
  assign n45631 = pi0244 & n34791;
  assign po0723 = n45630 | n45631;
  assign n45633 = ~pi0567 & pi1092;
  assign n45634 = ~pi1093 & n45633;
  assign n45635 = pi0603 & ~n17117;
  assign n45636 = n17182 & ~n20225;
  assign n45637 = ~n20235 & n45636;
  assign n45638 = n45635 & n45637;
  assign n45639 = ~pi0789 & ~n45634;
  assign n45640 = ~n45638 & n45639;
  assign n45641 = ~pi0619 & n45638;
  assign n45642 = ~n45634 & ~n45641;
  assign n45643 = ~pi1159 & ~n45642;
  assign n45644 = pi0619 & n45638;
  assign n45645 = ~n45634 & ~n45644;
  assign n45646 = pi1159 & ~n45645;
  assign n45647 = pi0789 & ~n45643;
  assign n45648 = ~n45646 & n45647;
  assign n45649 = ~n45640 & ~n45648;
  assign n45650 = pi0680 & n16826;
  assign n45651 = ~n19146 & n45650;
  assign n45652 = ~n45634 & ~n45651;
  assign n45653 = n19150 & ~n45652;
  assign n45654 = ~n16634 & n45648;
  assign n45655 = n45653 & ~n45654;
  assign n45656 = ~n45649 & ~n45655;
  assign n45657 = n17970 & ~n45656;
  assign n45658 = n35357 & n45649;
  assign n45659 = ~n16635 & n45653;
  assign n45660 = pi0641 & n45659;
  assign n45661 = ~n45634 & ~n45660;
  assign n45662 = n17865 & ~n45661;
  assign n45663 = ~pi0641 & n45659;
  assign n45664 = ~n45634 & ~n45663;
  assign n45665 = n17866 & ~n45664;
  assign n45666 = ~n45662 & ~n45665;
  assign n45667 = ~n45658 & n45666;
  assign n45668 = pi0788 & ~n45667;
  assign n45669 = ~n45657 & ~n45668;
  assign n45670 = ~n20364 & ~n45669;
  assign n45671 = n19151 & ~n45652;
  assign n45672 = pi0628 & n45671;
  assign n45673 = ~n45634 & ~n45672;
  assign n45674 = pi1156 & ~n45673;
  assign n45675 = ~n17969 & n45649;
  assign n45676 = n17969 & n45634;
  assign n45677 = ~n45675 & ~n45676;
  assign n45678 = n17854 & ~n45677;
  assign n45679 = ~pi0629 & ~n45674;
  assign n45680 = ~n45678 & n45679;
  assign n45681 = ~pi0628 & n45671;
  assign n45682 = ~n45634 & ~n45681;
  assign n45683 = ~pi1156 & ~n45682;
  assign n45684 = n17853 & ~n45677;
  assign n45685 = pi0629 & ~n45683;
  assign n45686 = ~n45684 & n45685;
  assign n45687 = pi0792 & ~n45680;
  assign n45688 = ~n45686 & n45687;
  assign n45689 = ~n45670 & ~n45688;
  assign n45690 = ~pi0647 & ~n45689;
  assign n45691 = ~n17779 & ~n45677;
  assign n45692 = n17779 & n45634;
  assign n45693 = ~n45691 & ~n45692;
  assign n45694 = pi0647 & ~n45693;
  assign n45695 = ~pi1157 & ~n45694;
  assign n45696 = ~n45690 & n45695;
  assign n45697 = ~n19142 & n45671;
  assign n45698 = pi0647 & n45697;
  assign n45699 = pi1157 & ~n45634;
  assign n45700 = ~n45698 & n45699;
  assign n45701 = ~pi0630 & ~n45700;
  assign n45702 = ~n45696 & n45701;
  assign n45703 = pi0647 & ~n45689;
  assign n45704 = ~pi0647 & ~n45693;
  assign n45705 = pi1157 & ~n45704;
  assign n45706 = ~n45703 & n45705;
  assign n45707 = ~pi0647 & n45697;
  assign n45708 = ~pi1157 & ~n45634;
  assign n45709 = ~n45707 & n45708;
  assign n45710 = pi0630 & ~n45709;
  assign n45711 = ~n45706 & n45710;
  assign n45712 = ~n45702 & ~n45711;
  assign n45713 = pi0787 & ~n45712;
  assign n45714 = ~pi0787 & ~n45689;
  assign n45715 = ~n45713 & ~n45714;
  assign n45716 = ~pi0790 & ~n45715;
  assign n45717 = ~n19342 & n45697;
  assign n45718 = ~n45634 & ~n45717;
  assign n45719 = pi0644 & ~n45718;
  assign n45720 = ~pi0644 & ~n45715;
  assign n45721 = ~pi0715 & ~n45719;
  assign n45722 = ~n45720 & n45721;
  assign n45723 = ~n17804 & n45691;
  assign n45724 = ~pi0644 & n45723;
  assign n45725 = pi0715 & ~n45634;
  assign n45726 = ~n45724 & n45725;
  assign n45727 = ~n45722 & ~n45726;
  assign n45728 = ~pi1160 & ~n45727;
  assign n45729 = pi0644 & n45723;
  assign n45730 = ~n45634 & ~n45729;
  assign n45731 = ~pi0715 & ~n45730;
  assign n45732 = ~pi0644 & n45718;
  assign n45733 = pi0644 & n45715;
  assign n45734 = pi0715 & ~n45732;
  assign n45735 = ~n45733 & n45734;
  assign n45736 = pi1160 & ~n45731;
  assign n45737 = ~n45735 & n45736;
  assign n45738 = pi0790 & ~n45737;
  assign n45739 = ~n45728 & n45738;
  assign n45740 = ~n45716 & ~n45739;
  assign n45741 = pi0230 & ~n45740;
  assign n45742 = ~pi0230 & n45633;
  assign po0724 = n45741 | n45742;
  assign n45744 = pi0568 & ~n34791;
  assign n45745 = pi0245 & n34791;
  assign po0725 = n45744 | n45745;
  assign n45747 = pi0569 & ~n34791;
  assign n45748 = ~pi0239 & n34791;
  assign po0726 = ~n45747 & ~n45748;
  assign n45750 = n34791 & n45455;
  assign n45751 = pi0570 & ~n45750;
  assign n45752 = ~pi0570 & n34786;
  assign n45753 = n45479 & n45752;
  assign po0727 = n45751 | n45753;
  assign n45755 = pi0571 & ~n36139;
  assign n45756 = pi0241 & n36139;
  assign po0728 = n45755 | n45756;
  assign n45758 = pi0572 & ~n36139;
  assign n45759 = pi0244 & n36139;
  assign po0729 = n45758 | n45759;
  assign n45761 = pi0573 & ~n36139;
  assign n45762 = pi0242 & n36139;
  assign po0730 = n45761 | n45762;
  assign n45764 = pi0574 & ~n34783;
  assign n45765 = pi0241 & n34783;
  assign po0731 = n45764 | n45765;
  assign n45767 = pi0575 & ~n36139;
  assign n45768 = pi0235 & n36139;
  assign po0732 = n45767 | n45768;
  assign n45770 = pi0576 & ~n36139;
  assign n45771 = pi0248 & n36139;
  assign po0733 = n45770 | n45771;
  assign n45773 = pi0577 & ~n36111;
  assign n45774 = pi0238 & n36111;
  assign po0734 = n45773 | n45774;
  assign n45776 = pi0578 & ~n34783;
  assign n45777 = pi0249 & n34783;
  assign po0735 = n45776 | n45777;
  assign n45779 = pi0579 & ~n34775;
  assign n45780 = pi0249 & n34775;
  assign po0736 = n45779 | n45780;
  assign n45782 = pi0580 & ~n36111;
  assign n45783 = pi0245 & n36111;
  assign po0737 = n45782 | n45783;
  assign n45785 = pi0581 & ~n34783;
  assign n45786 = pi0235 & n34783;
  assign po0738 = n45785 | n45786;
  assign n45788 = pi0582 & ~n34783;
  assign n45789 = pi0240 & n34783;
  assign po0739 = n45788 | n45789;
  assign n45791 = pi0584 & ~n34783;
  assign n45792 = pi0245 & n34783;
  assign po0741 = n45791 | n45792;
  assign n45794 = pi0585 & ~n34783;
  assign n45795 = pi0244 & n34783;
  assign po0742 = n45794 | n45795;
  assign n45797 = pi0586 & ~n34783;
  assign n45798 = pi0242 & n34783;
  assign po0743 = n45797 | n45798;
  assign n45800 = ~pi0230 & pi0587;
  assign n45801 = pi0230 & n17168;
  assign n45802 = ~n20225 & n45801;
  assign n45803 = ~n35575 & n45802;
  assign n45804 = n20237 & n45803;
  assign n45805 = n30797 & n45804;
  assign po0744 = n45800 | n45805;
  assign n45807 = ~pi0123 & n12373;
  assign n45808 = ~pi0588 & ~n45807;
  assign n45809 = ~pi0591 & n45807;
  assign n45810 = n44706 & ~n45808;
  assign po0745 = ~n45809 & n45810;
  assign n45812 = ~pi0204 & n45430;
  assign n45813 = ~pi0201 & n45454;
  assign n45814 = pi0233 & ~n45812;
  assign n45815 = ~n45813 & n45814;
  assign n45816 = ~pi0205 & n45430;
  assign n45817 = ~pi0202 & n45454;
  assign n45818 = ~pi0233 & ~n45816;
  assign n45819 = ~n45817 & n45818;
  assign n45820 = ~n45815 & ~n45819;
  assign n45821 = pi0237 & ~n45820;
  assign n45822 = ~pi0206 & n45430;
  assign n45823 = ~pi0220 & n45454;
  assign n45824 = pi0233 & ~n45822;
  assign n45825 = ~n45823 & n45824;
  assign n45826 = ~pi0218 & n45430;
  assign n45827 = ~pi0203 & n45454;
  assign n45828 = ~pi0233 & ~n45826;
  assign n45829 = ~n45827 & n45828;
  assign n45830 = ~n45825 & ~n45829;
  assign n45831 = ~pi0237 & ~n45830;
  assign po0746 = ~n45821 & ~n45831;
  assign n45833 = pi0588 & n45807;
  assign n45834 = pi0590 & ~n45807;
  assign n45835 = n44706 & ~n45833;
  assign po0747 = n45834 | ~n45835;
  assign n45837 = ~pi0591 & ~n45807;
  assign n45838 = ~pi0592 & n45807;
  assign n45839 = n44706 & ~n45837;
  assign po0748 = ~n45838 & n45839;
  assign n45841 = ~pi0592 & ~n45807;
  assign n45842 = ~pi0590 & n45807;
  assign n45843 = n44706 & ~n45841;
  assign po0749 = ~n45842 & n45843;
  assign n45845 = pi0234 & n45454;
  assign n45846 = pi0518 & ~n45845;
  assign n45847 = pi0246 & ~pi0520;
  assign n45848 = ~pi0246 & pi0520;
  assign n45849 = pi0249 & ~pi0578;
  assign n45850 = ~pi0249 & pi0578;
  assign n45851 = pi0248 & ~pi0521;
  assign n45852 = ~pi0248 & pi0521;
  assign n45853 = pi0241 & pi0574;
  assign n45854 = ~pi0241 & ~pi0574;
  assign n45855 = ~n45853 & ~n45854;
  assign n45856 = ~pi0518 & ~n45455;
  assign n45857 = ~n45847 & ~n45848;
  assign n45858 = ~n45849 & ~n45850;
  assign n45859 = ~n45851 & ~n45852;
  assign n45860 = n45858 & n45859;
  assign n45861 = ~n45855 & n45857;
  assign n45862 = n45860 & n45861;
  assign n45863 = ~n45846 & n45862;
  assign n45864 = ~n45856 & n45863;
  assign n45865 = pi0582 & n45864;
  assign n45866 = pi0240 & ~n45865;
  assign n45867 = ~pi0582 & n45864;
  assign n45868 = ~pi0240 & ~n45867;
  assign n45869 = ~n45866 & ~n45868;
  assign n45870 = ~pi0239 & pi0519;
  assign n45871 = pi0239 & ~pi0519;
  assign n45872 = ~n45870 & ~n45871;
  assign n45873 = n45869 & ~n45872;
  assign n45874 = pi0242 & pi0586;
  assign n45875 = ~pi0242 & ~pi0586;
  assign n45876 = ~n45874 & ~n45875;
  assign n45877 = n45873 & ~n45876;
  assign n45878 = pi0235 & pi0581;
  assign n45879 = ~pi0235 & ~pi0581;
  assign n45880 = ~n45878 & ~n45879;
  assign n45881 = n45877 & ~n45880;
  assign n45882 = pi0585 & n45881;
  assign n45883 = pi0244 & ~n45882;
  assign n45884 = ~pi0585 & n45881;
  assign n45885 = ~pi0244 & ~n45884;
  assign n45886 = ~n45883 & ~n45885;
  assign n45887 = pi0584 & n45886;
  assign n45888 = pi0245 & ~n45887;
  assign n45889 = ~pi0584 & n45886;
  assign n45890 = ~pi0245 & ~n45889;
  assign n45891 = ~n45888 & ~n45890;
  assign n45892 = ~pi0247 & ~pi0561;
  assign n45893 = pi0247 & pi0561;
  assign n45894 = ~n45892 & ~n45893;
  assign n45895 = n45891 & ~n45894;
  assign n45896 = pi0238 & n45895;
  assign n45897 = pi0240 & pi0542;
  assign n45898 = ~pi0240 & ~pi0542;
  assign n45899 = ~n45897 & ~n45898;
  assign n45900 = ~pi0248 & ~pi0501;
  assign n45901 = pi0248 & pi0501;
  assign n45902 = ~n45900 & ~n45901;
  assign n45903 = pi0234 & n45430;
  assign n45904 = pi0505 & ~n45903;
  assign n45905 = ~pi0505 & ~n45431;
  assign n45906 = pi0249 & ~pi0496;
  assign n45907 = ~pi0249 & pi0496;
  assign n45908 = ~pi0246 & ~pi0499;
  assign n45909 = pi0246 & pi0499;
  assign n45910 = ~n45908 & ~n45909;
  assign n45911 = ~n45906 & ~n45907;
  assign n45912 = ~n45902 & n45911;
  assign n45913 = ~n45910 & n45912;
  assign n45914 = ~n45904 & n45913;
  assign n45915 = ~n45905 & n45914;
  assign n45916 = ~pi0241 & ~pi0500;
  assign n45917 = pi0241 & pi0500;
  assign n45918 = ~n45916 & ~n45917;
  assign n45919 = n45915 & ~n45918;
  assign n45920 = ~n45899 & n45919;
  assign n45921 = pi0497 & n45920;
  assign n45922 = ~pi0239 & ~n45921;
  assign n45923 = ~pi0497 & n45920;
  assign n45924 = pi0239 & ~n45923;
  assign n45925 = ~n45922 & ~n45924;
  assign n45926 = pi0539 & n45925;
  assign n45927 = pi0242 & ~n45926;
  assign n45928 = ~pi0539 & n45925;
  assign n45929 = ~pi0242 & ~n45928;
  assign n45930 = ~n45927 & ~n45929;
  assign n45931 = pi0540 & n45930;
  assign n45932 = pi0235 & ~n45931;
  assign n45933 = ~pi0540 & n45930;
  assign n45934 = ~pi0235 & ~n45933;
  assign n45935 = ~n45932 & ~n45934;
  assign n45936 = pi0244 & pi0541;
  assign n45937 = ~pi0244 & ~pi0541;
  assign n45938 = ~n45936 & ~n45937;
  assign n45939 = n45935 & ~n45938;
  assign n45940 = pi0245 & pi0503;
  assign n45941 = ~pi0245 & ~pi0503;
  assign n45942 = ~n45940 & ~n45941;
  assign n45943 = n45939 & ~n45942;
  assign n45944 = ~pi0502 & n45943;
  assign n45945 = ~pi0247 & ~n45944;
  assign n45946 = pi0502 & n45943;
  assign n45947 = pi0247 & ~n45946;
  assign n45948 = ~n45945 & ~n45947;
  assign n45949 = ~pi0238 & n45948;
  assign n45950 = pi0522 & ~n45896;
  assign n45951 = ~n45949 & n45950;
  assign n45952 = ~n45892 & ~n45945;
  assign n45953 = pi0502 & ~n45891;
  assign n45954 = ~pi0500 & n45919;
  assign n45955 = n45915 & n45917;
  assign n45956 = ~n45864 & ~n45955;
  assign n45957 = ~n45954 & n45956;
  assign n45958 = ~pi0582 & ~n45957;
  assign n45959 = pi0582 & n45919;
  assign n45960 = ~pi0240 & ~n45959;
  assign n45961 = ~n45958 & n45960;
  assign n45962 = ~n45866 & ~n45961;
  assign n45963 = ~pi0542 & ~n45962;
  assign n45964 = pi0582 & ~n45957;
  assign n45965 = ~pi0582 & n45919;
  assign n45966 = pi0240 & ~n45965;
  assign n45967 = ~n45964 & n45966;
  assign n45968 = ~n45868 & ~n45967;
  assign n45969 = pi0542 & ~n45968;
  assign n45970 = ~n45963 & ~n45969;
  assign n45971 = ~pi0497 & n45970;
  assign n45972 = pi0497 & n45869;
  assign n45973 = pi0239 & ~n45972;
  assign n45974 = ~n45971 & n45973;
  assign n45975 = ~n45922 & ~n45974;
  assign n45976 = ~pi0519 & ~n45975;
  assign n45977 = pi0497 & n45970;
  assign n45978 = ~pi0497 & n45869;
  assign n45979 = ~pi0239 & ~n45978;
  assign n45980 = ~n45977 & n45979;
  assign n45981 = ~n45924 & ~n45980;
  assign n45982 = pi0519 & ~n45981;
  assign n45983 = ~n45976 & ~n45982;
  assign n45984 = ~pi0539 & n45983;
  assign n45985 = pi0539 & n45873;
  assign n45986 = ~pi0242 & ~n45985;
  assign n45987 = ~n45984 & n45986;
  assign n45988 = ~n45927 & ~n45987;
  assign n45989 = ~pi0586 & ~n45988;
  assign n45990 = pi0539 & n45983;
  assign n45991 = ~pi0539 & n45873;
  assign n45992 = pi0242 & ~n45991;
  assign n45993 = ~n45990 & n45992;
  assign n45994 = ~n45929 & ~n45993;
  assign n45995 = pi0586 & ~n45994;
  assign n45996 = ~n45989 & ~n45995;
  assign n45997 = ~pi0540 & n45996;
  assign n45998 = pi0540 & n45877;
  assign n45999 = ~pi0235 & ~n45998;
  assign n46000 = ~n45997 & n45999;
  assign n46001 = ~n45932 & ~n46000;
  assign n46002 = ~pi0581 & ~n46001;
  assign n46003 = pi0540 & n45996;
  assign n46004 = ~pi0540 & n45877;
  assign n46005 = pi0235 & ~n46004;
  assign n46006 = ~n46003 & n46005;
  assign n46007 = ~n45934 & ~n46006;
  assign n46008 = pi0581 & ~n46007;
  assign n46009 = ~n46002 & ~n46008;
  assign n46010 = ~pi0585 & n46009;
  assign n46011 = pi0585 & n45935;
  assign n46012 = ~pi0244 & ~n46011;
  assign n46013 = ~n46010 & n46012;
  assign n46014 = ~n45883 & ~n46013;
  assign n46015 = ~pi0541 & ~n46014;
  assign n46016 = pi0585 & n46009;
  assign n46017 = ~pi0585 & n45935;
  assign n46018 = pi0244 & ~n46017;
  assign n46019 = ~n46016 & n46018;
  assign n46020 = ~n45885 & ~n46019;
  assign n46021 = pi0541 & ~n46020;
  assign n46022 = ~n46015 & ~n46021;
  assign n46023 = ~pi0584 & n46022;
  assign n46024 = pi0584 & n45939;
  assign n46025 = ~pi0245 & ~n46024;
  assign n46026 = ~n46023 & n46025;
  assign n46027 = ~n45888 & ~n46026;
  assign n46028 = ~pi0503 & ~n46027;
  assign n46029 = pi0584 & n46022;
  assign n46030 = ~pi0584 & n45939;
  assign n46031 = pi0245 & ~n46030;
  assign n46032 = ~n46029 & n46031;
  assign n46033 = ~n45890 & ~n46032;
  assign n46034 = pi0503 & ~n46033;
  assign n46035 = ~n46028 & ~n46034;
  assign n46036 = ~pi0502 & ~n46035;
  assign n46037 = ~pi0561 & ~n45953;
  assign n46038 = ~n46036 & n46037;
  assign n46039 = ~n45952 & ~n46038;
  assign n46040 = ~n45893 & ~n45947;
  assign n46041 = ~pi0502 & ~n45891;
  assign n46042 = pi0502 & ~n46035;
  assign n46043 = pi0561 & ~n46041;
  assign n46044 = ~n46042 & n46043;
  assign n46045 = ~n46040 & ~n46044;
  assign n46046 = ~n46039 & ~n46045;
  assign n46047 = ~pi0238 & n46046;
  assign n46048 = ~pi0522 & ~n46047;
  assign n46049 = ~pi0543 & ~n45951;
  assign n46050 = ~n46048 & n46049;
  assign n46051 = ~pi0238 & n45895;
  assign n46052 = pi0238 & n45948;
  assign n46053 = ~pi0522 & ~n46051;
  assign n46054 = ~n46052 & n46053;
  assign n46055 = pi0238 & n46046;
  assign n46056 = pi0522 & ~n46055;
  assign n46057 = pi0543 & ~n46054;
  assign n46058 = ~n46056 & n46057;
  assign n46059 = ~n46050 & ~n46058;
  assign n46060 = ~pi0233 & ~n46059;
  assign n46061 = pi0246 & pi0536;
  assign n46062 = ~pi0246 & ~pi0536;
  assign n46063 = ~n46061 & ~n46062;
  assign n46064 = ~pi0557 & ~n45431;
  assign n46065 = pi0557 & ~n45903;
  assign n46066 = ~n46063 & ~n46064;
  assign n46067 = ~n46065 & n46066;
  assign n46068 = ~pi0538 & n46067;
  assign n46069 = ~pi0249 & ~n46068;
  assign n46070 = pi0538 & n46067;
  assign n46071 = pi0249 & ~n46070;
  assign n46072 = ~n46069 & ~n46071;
  assign n46073 = ~pi0537 & n46072;
  assign n46074 = ~pi0248 & ~n46073;
  assign n46075 = pi0537 & n46072;
  assign n46076 = pi0248 & ~n46075;
  assign n46077 = ~n46074 & ~n46076;
  assign n46078 = pi0241 & pi0506;
  assign n46079 = ~pi0241 & ~pi0506;
  assign n46080 = ~n46078 & ~n46079;
  assign n46081 = n46077 & ~n46080;
  assign n46082 = pi0240 & pi0535;
  assign n46083 = ~pi0240 & ~pi0535;
  assign n46084 = ~n46082 & ~n46083;
  assign n46085 = n46081 & ~n46084;
  assign n46086 = pi0534 & n46085;
  assign n46087 = ~pi0239 & ~n46086;
  assign n46088 = ~pi0534 & n46085;
  assign n46089 = pi0239 & ~n46088;
  assign n46090 = ~n46087 & ~n46089;
  assign n46091 = pi0504 & n46090;
  assign n46092 = pi0242 & ~n46091;
  assign n46093 = ~pi0504 & n46090;
  assign n46094 = ~pi0242 & ~n46093;
  assign n46095 = ~n46092 & ~n46094;
  assign n46096 = pi0533 & n46095;
  assign n46097 = pi0235 & ~n46096;
  assign n46098 = ~pi0533 & n46095;
  assign n46099 = ~pi0235 & ~n46098;
  assign n46100 = ~n46097 & ~n46099;
  assign n46101 = pi0558 & n46100;
  assign n46102 = pi0244 & ~n46101;
  assign n46103 = ~pi0558 & n46100;
  assign n46104 = ~pi0244 & ~n46103;
  assign n46105 = ~n46102 & ~n46104;
  assign n46106 = pi0509 & n46105;
  assign n46107 = pi0245 & ~n46106;
  assign n46108 = ~pi0509 & n46105;
  assign n46109 = ~pi0245 & ~n46108;
  assign n46110 = ~n46107 & ~n46109;
  assign n46111 = pi0508 & n46110;
  assign n46112 = pi0247 & ~n46111;
  assign n46113 = ~pi0508 & n46110;
  assign n46114 = ~pi0247 & ~n46113;
  assign n46115 = ~n46112 & ~n46114;
  assign n46116 = ~pi0238 & n46115;
  assign n46117 = pi0248 & pi0481;
  assign n46118 = ~pi0248 & ~pi0481;
  assign n46119 = ~n46117 & ~n46118;
  assign n46120 = pi0246 & pi0487;
  assign n46121 = ~pi0246 & ~pi0487;
  assign n46122 = ~n46120 & ~n46121;
  assign n46123 = ~pi0511 & ~n45455;
  assign n46124 = pi0511 & ~n45845;
  assign n46125 = ~n46122 & ~n46123;
  assign n46126 = ~n46124 & n46125;
  assign n46127 = ~pi0249 & ~pi0579;
  assign n46128 = pi0249 & pi0579;
  assign n46129 = ~n46127 & ~n46128;
  assign n46130 = n46126 & ~n46129;
  assign n46131 = ~n46119 & n46130;
  assign n46132 = pi0559 & n46131;
  assign n46133 = pi0241 & ~n46132;
  assign n46134 = ~pi0559 & n46131;
  assign n46135 = ~pi0241 & ~n46134;
  assign n46136 = ~n46133 & ~n46135;
  assign n46137 = pi0515 & n46136;
  assign n46138 = pi0240 & ~n46137;
  assign n46139 = ~pi0515 & n46136;
  assign n46140 = ~pi0240 & ~n46139;
  assign n46141 = ~n46138 & ~n46140;
  assign n46142 = ~pi0239 & pi0488;
  assign n46143 = pi0239 & ~pi0488;
  assign n46144 = ~n46142 & ~n46143;
  assign n46145 = n46141 & ~n46144;
  assign n46146 = pi0242 & pi0510;
  assign n46147 = ~pi0242 & ~pi0510;
  assign n46148 = ~n46146 & ~n46147;
  assign n46149 = n46145 & ~n46148;
  assign n46150 = pi0235 & pi0512;
  assign n46151 = ~pi0235 & ~pi0512;
  assign n46152 = ~n46150 & ~n46151;
  assign n46153 = n46149 & ~n46152;
  assign n46154 = pi0244 & pi0513;
  assign n46155 = ~pi0244 & ~pi0513;
  assign n46156 = ~n46154 & ~n46155;
  assign n46157 = n46153 & ~n46156;
  assign n46158 = pi0245 & pi0514;
  assign n46159 = ~pi0245 & ~pi0514;
  assign n46160 = ~n46158 & ~n46159;
  assign n46161 = n46157 & ~n46160;
  assign n46162 = pi0247 & pi0516;
  assign n46163 = ~pi0247 & ~pi0516;
  assign n46164 = ~n46162 & ~n46163;
  assign n46165 = n46161 & ~n46164;
  assign n46166 = pi0238 & n46165;
  assign n46167 = pi0517 & ~n46166;
  assign n46168 = ~n46116 & n46167;
  assign n46169 = ~pi0579 & ~n46130;
  assign n46170 = ~n46069 & n46126;
  assign n46171 = pi0579 & ~n46170;
  assign n46172 = ~n46169 & ~n46171;
  assign n46173 = ~n46072 & ~n46172;
  assign n46174 = ~pi0537 & ~n46173;
  assign n46175 = pi0537 & n46130;
  assign n46176 = ~pi0248 & ~n46175;
  assign n46177 = ~n46174 & n46176;
  assign n46178 = ~n46076 & ~n46177;
  assign n46179 = ~pi0481 & ~n46178;
  assign n46180 = pi0537 & ~n46173;
  assign n46181 = ~pi0537 & n46130;
  assign n46182 = pi0248 & ~n46181;
  assign n46183 = ~n46180 & n46182;
  assign n46184 = ~n46074 & ~n46183;
  assign n46185 = pi0481 & ~n46184;
  assign n46186 = ~n46179 & ~n46185;
  assign n46187 = ~pi0559 & n46186;
  assign n46188 = pi0559 & n46077;
  assign n46189 = ~pi0241 & ~n46188;
  assign n46190 = ~n46187 & n46189;
  assign n46191 = ~n46133 & ~n46190;
  assign n46192 = ~pi0506 & ~n46191;
  assign n46193 = pi0559 & n46186;
  assign n46194 = ~pi0559 & n46077;
  assign n46195 = pi0241 & ~n46194;
  assign n46196 = ~n46193 & n46195;
  assign n46197 = ~n46135 & ~n46196;
  assign n46198 = pi0506 & ~n46197;
  assign n46199 = ~n46192 & ~n46198;
  assign n46200 = ~pi0515 & n46199;
  assign n46201 = pi0515 & n46081;
  assign n46202 = ~pi0240 & ~n46201;
  assign n46203 = ~n46200 & n46202;
  assign n46204 = ~n46138 & ~n46203;
  assign n46205 = ~pi0535 & ~n46204;
  assign n46206 = pi0515 & n46199;
  assign n46207 = ~pi0515 & n46081;
  assign n46208 = pi0240 & ~n46207;
  assign n46209 = ~n46206 & n46208;
  assign n46210 = ~n46140 & ~n46209;
  assign n46211 = pi0535 & ~n46210;
  assign n46212 = ~n46205 & ~n46211;
  assign n46213 = ~pi0534 & n46212;
  assign n46214 = pi0534 & n46141;
  assign n46215 = pi0239 & ~n46214;
  assign n46216 = ~n46213 & n46215;
  assign n46217 = ~n46087 & ~n46216;
  assign n46218 = ~pi0488 & ~n46217;
  assign n46219 = pi0534 & n46212;
  assign n46220 = ~pi0534 & n46141;
  assign n46221 = ~pi0239 & ~n46220;
  assign n46222 = ~n46219 & n46221;
  assign n46223 = ~n46089 & ~n46222;
  assign n46224 = pi0488 & ~n46223;
  assign n46225 = ~n46218 & ~n46224;
  assign n46226 = ~pi0504 & n46225;
  assign n46227 = pi0504 & n46145;
  assign n46228 = ~pi0242 & ~n46227;
  assign n46229 = ~n46226 & n46228;
  assign n46230 = ~n46092 & ~n46229;
  assign n46231 = ~pi0510 & ~n46230;
  assign n46232 = pi0504 & n46225;
  assign n46233 = ~pi0504 & n46145;
  assign n46234 = pi0242 & ~n46233;
  assign n46235 = ~n46232 & n46234;
  assign n46236 = ~n46094 & ~n46235;
  assign n46237 = pi0510 & ~n46236;
  assign n46238 = ~n46231 & ~n46237;
  assign n46239 = ~pi0533 & n46238;
  assign n46240 = pi0533 & n46149;
  assign n46241 = ~pi0235 & ~n46240;
  assign n46242 = ~n46239 & n46241;
  assign n46243 = ~n46097 & ~n46242;
  assign n46244 = ~pi0512 & ~n46243;
  assign n46245 = pi0533 & n46238;
  assign n46246 = ~pi0533 & n46149;
  assign n46247 = pi0235 & ~n46246;
  assign n46248 = ~n46245 & n46247;
  assign n46249 = ~n46099 & ~n46248;
  assign n46250 = pi0512 & ~n46249;
  assign n46251 = ~n46244 & ~n46250;
  assign n46252 = ~pi0558 & n46251;
  assign n46253 = pi0558 & n46153;
  assign n46254 = ~pi0244 & ~n46253;
  assign n46255 = ~n46252 & n46254;
  assign n46256 = ~n46102 & ~n46255;
  assign n46257 = ~pi0513 & ~n46256;
  assign n46258 = pi0558 & n46251;
  assign n46259 = ~pi0558 & n46153;
  assign n46260 = pi0244 & ~n46259;
  assign n46261 = ~n46258 & n46260;
  assign n46262 = ~n46104 & ~n46261;
  assign n46263 = pi0513 & ~n46262;
  assign n46264 = ~n46257 & ~n46263;
  assign n46265 = ~pi0509 & n46264;
  assign n46266 = pi0509 & n46157;
  assign n46267 = ~pi0245 & ~n46266;
  assign n46268 = ~n46265 & n46267;
  assign n46269 = ~n46107 & ~n46268;
  assign n46270 = ~pi0514 & ~n46269;
  assign n46271 = pi0509 & n46264;
  assign n46272 = ~pi0509 & n46157;
  assign n46273 = pi0245 & ~n46272;
  assign n46274 = ~n46271 & n46273;
  assign n46275 = ~n46109 & ~n46274;
  assign n46276 = pi0514 & ~n46275;
  assign n46277 = ~n46270 & ~n46276;
  assign n46278 = ~pi0508 & n46277;
  assign n46279 = pi0508 & n46161;
  assign n46280 = ~pi0247 & ~n46279;
  assign n46281 = ~n46278 & n46280;
  assign n46282 = ~n46112 & ~n46281;
  assign n46283 = ~pi0516 & ~n46282;
  assign n46284 = pi0508 & n46277;
  assign n46285 = ~pi0508 & n46161;
  assign n46286 = pi0247 & ~n46285;
  assign n46287 = ~n46284 & n46286;
  assign n46288 = ~n46114 & ~n46287;
  assign n46289 = pi0516 & ~n46288;
  assign n46290 = ~n46283 & ~n46289;
  assign n46291 = ~pi0238 & n46290;
  assign n46292 = ~pi0517 & ~n46291;
  assign n46293 = ~pi0507 & ~n46168;
  assign n46294 = ~n46292 & n46293;
  assign n46295 = pi0238 & n46115;
  assign n46296 = ~pi0238 & n46165;
  assign n46297 = ~pi0517 & ~n46296;
  assign n46298 = ~n46295 & n46297;
  assign n46299 = pi0238 & n46290;
  assign n46300 = pi0517 & ~n46299;
  assign n46301 = pi0507 & ~n46298;
  assign n46302 = ~n46300 & n46301;
  assign n46303 = ~n46294 & ~n46302;
  assign n46304 = pi0233 & ~n46303;
  assign n46305 = pi0237 & ~n46060;
  assign n46306 = ~n46304 & n46305;
  assign n46307 = ~pi0240 & ~pi0492;
  assign n46308 = pi0240 & pi0492;
  assign n46309 = ~n46307 & ~n46308;
  assign n46310 = pi0241 & pi0490;
  assign n46311 = ~pi0241 & ~pi0490;
  assign n46312 = ~n46310 & ~n46311;
  assign n46313 = pi0248 & pi0548;
  assign n46314 = ~pi0248 & ~pi0548;
  assign n46315 = ~n46313 & ~n46314;
  assign n46316 = pi0249 & pi0484;
  assign n46317 = ~pi0249 & ~pi0484;
  assign n46318 = ~n46316 & ~n46317;
  assign n46319 = pi0246 & pi0546;
  assign n46320 = ~pi0246 & ~pi0546;
  assign n46321 = ~n46319 & ~n46320;
  assign n46322 = ~pi0544 & ~n45431;
  assign n46323 = pi0544 & ~n45903;
  assign n46324 = ~n46315 & ~n46318;
  assign n46325 = ~n46321 & n46324;
  assign n46326 = ~n46322 & n46325;
  assign n46327 = ~n46323 & n46326;
  assign n46328 = ~n46312 & n46327;
  assign n46329 = ~n46309 & n46328;
  assign n46330 = pi0494 & n46329;
  assign n46331 = ~pi0239 & ~n46330;
  assign n46332 = ~pi0494 & n46329;
  assign n46333 = pi0239 & ~n46332;
  assign n46334 = ~n46331 & ~n46333;
  assign n46335 = pi0483 & n46334;
  assign n46336 = pi0242 & ~n46335;
  assign n46337 = ~pi0483 & n46334;
  assign n46338 = ~pi0242 & ~n46337;
  assign n46339 = ~n46336 & ~n46338;
  assign n46340 = pi0495 & n46339;
  assign n46341 = pi0235 & ~n46340;
  assign n46342 = ~pi0495 & n46339;
  assign n46343 = ~pi0235 & ~n46342;
  assign n46344 = ~n46341 & ~n46343;
  assign n46345 = pi0244 & pi0493;
  assign n46346 = ~pi0244 & ~pi0493;
  assign n46347 = ~n46345 & ~n46346;
  assign n46348 = n46344 & ~n46347;
  assign n46349 = pi0545 & n46348;
  assign n46350 = pi0245 & ~n46349;
  assign n46351 = ~pi0545 & n46348;
  assign n46352 = ~pi0245 & ~n46351;
  assign n46353 = ~n46350 & ~n46352;
  assign n46354 = pi0547 & n46353;
  assign n46355 = pi0247 & ~n46354;
  assign n46356 = ~pi0547 & n46353;
  assign n46357 = ~pi0247 & ~n46356;
  assign n46358 = ~n46355 & ~n46357;
  assign n46359 = ~pi0238 & n46358;
  assign n46360 = pi0523 & ~n45845;
  assign n46361 = pi0248 & pi0576;
  assign n46362 = ~pi0248 & ~pi0576;
  assign n46363 = ~n46361 & ~n46362;
  assign n46364 = pi0249 & pi0528;
  assign n46365 = ~pi0249 & ~pi0528;
  assign n46366 = ~n46364 & ~n46365;
  assign n46367 = pi0246 & pi0526;
  assign n46368 = ~pi0246 & ~pi0526;
  assign n46369 = ~n46367 & ~n46368;
  assign n46370 = ~pi0523 & ~n45455;
  assign n46371 = ~n46363 & ~n46366;
  assign n46372 = ~n46369 & n46371;
  assign n46373 = ~n46360 & n46372;
  assign n46374 = ~n46370 & n46373;
  assign n46375 = pi0571 & n46374;
  assign n46376 = pi0241 & ~n46375;
  assign n46377 = ~pi0571 & n46374;
  assign n46378 = ~pi0241 & ~n46377;
  assign n46379 = ~n46376 & ~n46378;
  assign n46380 = ~pi0530 & n46379;
  assign n46381 = ~pi0240 & ~n46380;
  assign n46382 = pi0530 & n46379;
  assign n46383 = pi0240 & ~n46382;
  assign n46384 = ~n46381 & ~n46383;
  assign n46385 = ~pi0239 & pi0524;
  assign n46386 = pi0239 & ~pi0524;
  assign n46387 = ~n46385 & ~n46386;
  assign n46388 = n46384 & ~n46387;
  assign n46389 = pi0242 & pi0573;
  assign n46390 = ~pi0242 & ~pi0573;
  assign n46391 = ~n46389 & ~n46390;
  assign n46392 = n46388 & ~n46391;
  assign n46393 = pi0235 & pi0575;
  assign n46394 = ~pi0235 & ~pi0575;
  assign n46395 = ~n46393 & ~n46394;
  assign n46396 = n46392 & ~n46395;
  assign n46397 = pi0572 & n46396;
  assign n46398 = pi0244 & ~n46397;
  assign n46399 = ~pi0572 & n46396;
  assign n46400 = ~pi0244 & ~n46399;
  assign n46401 = ~n46398 & ~n46400;
  assign n46402 = pi0245 & pi0525;
  assign n46403 = ~pi0245 & ~pi0525;
  assign n46404 = ~n46402 & ~n46403;
  assign n46405 = n46401 & ~n46404;
  assign n46406 = pi0247 & pi0527;
  assign n46407 = ~pi0247 & ~pi0527;
  assign n46408 = ~n46406 & ~n46407;
  assign n46409 = n46405 & ~n46408;
  assign n46410 = pi0238 & n46409;
  assign n46411 = pi0529 & ~n46410;
  assign n46412 = ~n46359 & n46411;
  assign n46413 = ~n46307 & ~n46381;
  assign n46414 = pi0530 & ~n46328;
  assign n46415 = ~pi0241 & ~n46327;
  assign n46416 = ~n46377 & n46415;
  assign n46417 = ~n46376 & ~n46416;
  assign n46418 = ~pi0490 & ~n46417;
  assign n46419 = pi0241 & ~n46327;
  assign n46420 = ~n46375 & n46419;
  assign n46421 = ~n46378 & ~n46420;
  assign n46422 = pi0490 & ~n46421;
  assign n46423 = ~n46418 & ~n46422;
  assign n46424 = ~pi0530 & ~n46423;
  assign n46425 = ~pi0492 & ~n46414;
  assign n46426 = ~n46424 & n46425;
  assign n46427 = ~n46413 & ~n46426;
  assign n46428 = ~n46308 & ~n46383;
  assign n46429 = ~pi0530 & ~n46328;
  assign n46430 = pi0530 & ~n46423;
  assign n46431 = pi0492 & ~n46429;
  assign n46432 = ~n46430 & n46431;
  assign n46433 = ~n46428 & ~n46432;
  assign n46434 = ~n46427 & ~n46433;
  assign n46435 = ~pi0494 & n46434;
  assign n46436 = pi0494 & n46384;
  assign n46437 = pi0239 & ~n46436;
  assign n46438 = ~n46435 & n46437;
  assign n46439 = ~n46331 & ~n46438;
  assign n46440 = ~pi0524 & ~n46439;
  assign n46441 = pi0494 & n46434;
  assign n46442 = ~pi0494 & n46384;
  assign n46443 = ~pi0239 & ~n46442;
  assign n46444 = ~n46441 & n46443;
  assign n46445 = ~n46333 & ~n46444;
  assign n46446 = pi0524 & ~n46445;
  assign n46447 = ~n46440 & ~n46446;
  assign n46448 = ~pi0483 & n46447;
  assign n46449 = pi0483 & n46388;
  assign n46450 = ~pi0242 & ~n46449;
  assign n46451 = ~n46448 & n46450;
  assign n46452 = ~n46336 & ~n46451;
  assign n46453 = ~pi0573 & ~n46452;
  assign n46454 = pi0483 & n46447;
  assign n46455 = ~pi0483 & n46388;
  assign n46456 = pi0242 & ~n46455;
  assign n46457 = ~n46454 & n46456;
  assign n46458 = ~n46338 & ~n46457;
  assign n46459 = pi0573 & ~n46458;
  assign n46460 = ~n46453 & ~n46459;
  assign n46461 = ~pi0495 & n46460;
  assign n46462 = pi0495 & n46392;
  assign n46463 = ~pi0235 & ~n46462;
  assign n46464 = ~n46461 & n46463;
  assign n46465 = ~n46341 & ~n46464;
  assign n46466 = ~pi0575 & ~n46465;
  assign n46467 = pi0495 & n46460;
  assign n46468 = ~pi0495 & n46392;
  assign n46469 = pi0235 & ~n46468;
  assign n46470 = ~n46467 & n46469;
  assign n46471 = ~n46343 & ~n46470;
  assign n46472 = pi0575 & ~n46471;
  assign n46473 = ~n46466 & ~n46472;
  assign n46474 = ~pi0572 & n46473;
  assign n46475 = pi0572 & n46344;
  assign n46476 = ~pi0244 & ~n46475;
  assign n46477 = ~n46474 & n46476;
  assign n46478 = ~n46398 & ~n46477;
  assign n46479 = ~pi0493 & ~n46478;
  assign n46480 = pi0572 & n46473;
  assign n46481 = ~pi0572 & n46344;
  assign n46482 = pi0244 & ~n46481;
  assign n46483 = ~n46480 & n46482;
  assign n46484 = ~n46400 & ~n46483;
  assign n46485 = pi0493 & ~n46484;
  assign n46486 = ~n46479 & ~n46485;
  assign n46487 = ~pi0545 & n46486;
  assign n46488 = pi0545 & n46401;
  assign n46489 = ~pi0245 & ~n46488;
  assign n46490 = ~n46487 & n46489;
  assign n46491 = ~n46350 & ~n46490;
  assign n46492 = ~pi0525 & ~n46491;
  assign n46493 = pi0545 & n46486;
  assign n46494 = ~pi0545 & n46401;
  assign n46495 = pi0245 & ~n46494;
  assign n46496 = ~n46493 & n46495;
  assign n46497 = ~n46352 & ~n46496;
  assign n46498 = pi0525 & ~n46497;
  assign n46499 = ~n46492 & ~n46498;
  assign n46500 = ~pi0547 & n46499;
  assign n46501 = pi0547 & n46405;
  assign n46502 = ~pi0247 & ~n46501;
  assign n46503 = ~n46500 & n46502;
  assign n46504 = ~n46355 & ~n46503;
  assign n46505 = ~pi0527 & ~n46504;
  assign n46506 = pi0547 & n46499;
  assign n46507 = ~pi0547 & n46405;
  assign n46508 = pi0247 & ~n46507;
  assign n46509 = ~n46506 & n46508;
  assign n46510 = ~n46357 & ~n46509;
  assign n46511 = pi0527 & ~n46510;
  assign n46512 = ~n46505 & ~n46511;
  assign n46513 = ~pi0238 & n46512;
  assign n46514 = ~pi0529 & ~n46513;
  assign n46515 = ~pi0491 & ~n46412;
  assign n46516 = ~n46514 & n46515;
  assign n46517 = pi0238 & n46358;
  assign n46518 = ~pi0238 & n46409;
  assign n46519 = ~pi0529 & ~n46518;
  assign n46520 = ~n46517 & n46519;
  assign n46521 = pi0238 & n46512;
  assign n46522 = pi0529 & ~n46521;
  assign n46523 = pi0491 & ~n46520;
  assign n46524 = ~n46522 & n46523;
  assign n46525 = ~n46516 & ~n46524;
  assign n46526 = pi0233 & ~n46525;
  assign n46527 = pi0485 & ~n45903;
  assign n46528 = pi0240 & pi0551;
  assign n46529 = ~pi0240 & ~pi0551;
  assign n46530 = ~n46528 & ~n46529;
  assign n46531 = pi0249 & ~pi0555;
  assign n46532 = ~pi0249 & pi0555;
  assign n46533 = pi0241 & ~pi0553;
  assign n46534 = ~pi0241 & pi0553;
  assign n46535 = pi0248 & ~pi0554;
  assign n46536 = ~pi0248 & pi0554;
  assign n46537 = ~pi0246 & pi0563;
  assign n46538 = pi0246 & ~pi0563;
  assign n46539 = ~pi0485 & ~n45431;
  assign n46540 = ~n46531 & ~n46532;
  assign n46541 = ~n46533 & ~n46534;
  assign n46542 = ~n46535 & ~n46536;
  assign n46543 = ~n46537 & ~n46538;
  assign n46544 = n46542 & n46543;
  assign n46545 = n46540 & n46541;
  assign n46546 = ~n46530 & n46545;
  assign n46547 = n46544 & n46546;
  assign n46548 = ~n46527 & n46547;
  assign n46549 = ~n46539 & n46548;
  assign n46550 = pi0550 & n46549;
  assign n46551 = ~pi0239 & ~n46550;
  assign n46552 = ~pi0550 & n46549;
  assign n46553 = pi0239 & ~n46552;
  assign n46554 = ~n46551 & ~n46553;
  assign n46555 = ~pi0489 & n46554;
  assign n46556 = ~pi0242 & ~n46555;
  assign n46557 = pi0489 & n46554;
  assign n46558 = pi0242 & ~n46557;
  assign n46559 = ~n46556 & ~n46558;
  assign n46560 = pi0549 & n46559;
  assign n46561 = pi0235 & ~n46560;
  assign n46562 = ~pi0549 & n46559;
  assign n46563 = ~pi0235 & ~n46562;
  assign n46564 = ~n46561 & ~n46563;
  assign n46565 = pi0486 & n46564;
  assign n46566 = pi0244 & ~n46565;
  assign n46567 = ~pi0486 & n46564;
  assign n46568 = ~pi0244 & ~n46567;
  assign n46569 = ~n46566 & ~n46568;
  assign n46570 = pi0245 & pi0580;
  assign n46571 = ~pi0245 & ~pi0580;
  assign n46572 = ~n46570 & ~n46571;
  assign n46573 = n46569 & ~n46572;
  assign n46574 = pi0552 & n46573;
  assign n46575 = pi0247 & ~n46574;
  assign n46576 = ~pi0552 & n46573;
  assign n46577 = ~pi0247 & ~n46576;
  assign n46578 = ~n46575 & ~n46577;
  assign n46579 = pi0238 & n46578;
  assign n46580 = ~pi0242 & ~pi0556;
  assign n46581 = pi0242 & pi0556;
  assign n46582 = ~n46580 & ~n46581;
  assign n46583 = pi0246 & ~pi0564;
  assign n46584 = pi0570 & ~n45845;
  assign n46585 = ~pi0246 & pi0564;
  assign n46586 = pi0249 & ~pi0482;
  assign n46587 = ~pi0249 & pi0482;
  assign n46588 = pi0241 & pi0562;
  assign n46589 = ~pi0241 & ~pi0562;
  assign n46590 = ~n46588 & ~n46589;
  assign n46591 = ~pi0570 & ~n45455;
  assign n46592 = ~n46585 & ~n46586;
  assign n46593 = ~n46587 & n46592;
  assign n46594 = ~n46590 & n46593;
  assign n46595 = ~n46584 & n46594;
  assign n46596 = ~n46591 & n46595;
  assign n46597 = pi0248 & ~pi0565;
  assign n46598 = ~pi0248 & pi0565;
  assign n46599 = ~n46597 & ~n46598;
  assign n46600 = pi0240 & pi0560;
  assign n46601 = ~pi0240 & ~pi0560;
  assign n46602 = ~n46600 & ~n46601;
  assign n46603 = ~n46583 & n46599;
  assign n46604 = ~n46602 & n46603;
  assign n46605 = n46596 & n46604;
  assign n46606 = ~pi0240 & ~n46605;
  assign n46607 = pi0560 & ~n46583;
  assign n46608 = n46599 & n46607;
  assign n46609 = n46596 & n46608;
  assign n46610 = pi0240 & ~n46609;
  assign n46611 = ~n46606 & ~n46610;
  assign n46612 = ~pi0239 & pi0569;
  assign n46613 = pi0239 & ~pi0569;
  assign n46614 = ~n46612 & ~n46613;
  assign n46615 = n46611 & ~n46614;
  assign n46616 = ~n46582 & n46615;
  assign n46617 = pi0235 & pi0531;
  assign n46618 = ~pi0235 & ~pi0531;
  assign n46619 = ~n46617 & ~n46618;
  assign n46620 = n46616 & ~n46619;
  assign n46621 = pi0244 & pi0566;
  assign n46622 = ~pi0244 & ~pi0566;
  assign n46623 = ~n46621 & ~n46622;
  assign n46624 = n46620 & ~n46623;
  assign n46625 = pi0568 & n46624;
  assign n46626 = pi0245 & ~n46625;
  assign n46627 = ~pi0568 & n46624;
  assign n46628 = ~pi0245 & ~n46627;
  assign n46629 = ~n46626 & ~n46628;
  assign n46630 = pi0247 & pi0532;
  assign n46631 = ~pi0247 & ~pi0532;
  assign n46632 = ~n46630 & ~n46631;
  assign n46633 = n46629 & ~n46632;
  assign n46634 = ~pi0238 & n46633;
  assign n46635 = pi0577 & ~n46634;
  assign n46636 = ~n46579 & n46635;
  assign n46637 = ~n46556 & ~n46580;
  assign n46638 = pi0489 & ~n46615;
  assign n46639 = n46605 & n46613;
  assign n46640 = pi0569 & ~n46553;
  assign n46641 = n46611 & n46640;
  assign n46642 = ~n46554 & ~n46639;
  assign n46643 = ~n46641 & n46642;
  assign n46644 = ~pi0489 & n46643;
  assign n46645 = ~pi0556 & ~n46638;
  assign n46646 = ~n46644 & n46645;
  assign n46647 = ~n46637 & ~n46646;
  assign n46648 = ~n46558 & ~n46581;
  assign n46649 = ~pi0489 & ~n46615;
  assign n46650 = pi0489 & n46643;
  assign n46651 = pi0556 & ~n46649;
  assign n46652 = ~n46650 & n46651;
  assign n46653 = ~n46648 & ~n46652;
  assign n46654 = ~n46647 & ~n46653;
  assign n46655 = ~pi0549 & n46654;
  assign n46656 = pi0549 & n46616;
  assign n46657 = ~pi0235 & ~n46656;
  assign n46658 = ~n46655 & n46657;
  assign n46659 = ~n46561 & ~n46658;
  assign n46660 = ~pi0531 & ~n46659;
  assign n46661 = pi0549 & n46654;
  assign n46662 = ~pi0549 & n46616;
  assign n46663 = pi0235 & ~n46662;
  assign n46664 = ~n46661 & n46663;
  assign n46665 = ~n46563 & ~n46664;
  assign n46666 = pi0531 & ~n46665;
  assign n46667 = ~n46660 & ~n46666;
  assign n46668 = ~pi0486 & n46667;
  assign n46669 = pi0486 & n46620;
  assign n46670 = ~pi0244 & ~n46669;
  assign n46671 = ~n46668 & n46670;
  assign n46672 = ~n46566 & ~n46671;
  assign n46673 = ~pi0566 & ~n46672;
  assign n46674 = pi0486 & n46667;
  assign n46675 = ~pi0486 & n46620;
  assign n46676 = pi0244 & ~n46675;
  assign n46677 = ~n46674 & n46676;
  assign n46678 = ~n46568 & ~n46677;
  assign n46679 = pi0566 & ~n46678;
  assign n46680 = ~n46673 & ~n46679;
  assign n46681 = ~pi0568 & n46680;
  assign n46682 = pi0568 & n46569;
  assign n46683 = ~pi0245 & ~n46682;
  assign n46684 = ~n46681 & n46683;
  assign n46685 = ~n46626 & ~n46684;
  assign n46686 = ~pi0580 & ~n46685;
  assign n46687 = pi0568 & n46680;
  assign n46688 = ~pi0568 & n46569;
  assign n46689 = pi0245 & ~n46688;
  assign n46690 = ~n46687 & n46689;
  assign n46691 = ~n46628 & ~n46690;
  assign n46692 = pi0580 & ~n46691;
  assign n46693 = ~n46686 & ~n46692;
  assign n46694 = ~pi0552 & n46693;
  assign n46695 = pi0552 & n46629;
  assign n46696 = ~pi0247 & ~n46695;
  assign n46697 = ~n46694 & n46696;
  assign n46698 = ~n46575 & ~n46697;
  assign n46699 = ~pi0532 & ~n46698;
  assign n46700 = pi0552 & n46693;
  assign n46701 = ~pi0552 & n46629;
  assign n46702 = pi0247 & ~n46701;
  assign n46703 = ~n46700 & n46702;
  assign n46704 = ~n46577 & ~n46703;
  assign n46705 = pi0532 & ~n46704;
  assign n46706 = ~n46699 & ~n46705;
  assign n46707 = ~pi0238 & n46706;
  assign n46708 = ~pi0577 & ~n46707;
  assign n46709 = ~pi0498 & ~n46636;
  assign n46710 = ~n46708 & n46709;
  assign n46711 = ~pi0238 & n46578;
  assign n46712 = pi0238 & n46633;
  assign n46713 = ~pi0577 & ~n46712;
  assign n46714 = ~n46711 & n46713;
  assign n46715 = pi0238 & n46706;
  assign n46716 = pi0577 & ~n46715;
  assign n46717 = pi0498 & ~n46714;
  assign n46718 = ~n46716 & n46717;
  assign n46719 = ~n46710 & ~n46718;
  assign n46720 = ~pi0233 & ~n46719;
  assign n46721 = ~pi0237 & ~n46720;
  assign n46722 = ~n46526 & n46721;
  assign po0750 = ~n46306 & ~n46722;
  assign n46724 = ~pi0806 & n45126;
  assign n46725 = ~pi0332 & ~pi0806;
  assign n46726 = pi0990 & n46725;
  assign n46727 = pi0600 & n46726;
  assign n46728 = ~pi0332 & pi0594;
  assign n46729 = ~n46727 & ~n46728;
  assign po0751 = ~n46724 & ~n46729;
  assign n46731 = pi0605 & ~pi0806;
  assign n46732 = n45109 & n46731;
  assign n46733 = ~pi0595 & ~n46732;
  assign n46734 = pi0595 & n46732;
  assign n46735 = ~pi0332 & ~n46733;
  assign po0752 = ~n46734 & n46735;
  assign n46737 = ~pi0332 & pi0596;
  assign n46738 = pi0595 & n45108;
  assign n46739 = n46726 & n46738;
  assign n46740 = ~n46737 & ~n46739;
  assign n46741 = pi0596 & n46739;
  assign po0753 = ~n46740 & ~n46741;
  assign n46743 = ~pi0597 & ~n46724;
  assign n46744 = pi0597 & n46724;
  assign n46745 = ~pi0332 & ~n46743;
  assign po0754 = ~n46744 & n46745;
  assign n46747 = ~pi0882 & ~po1038;
  assign n46748 = pi0947 & n46747;
  assign n46749 = pi0598 & ~n46748;
  assign n46750 = pi0740 & pi0780;
  assign n46751 = n6192 & n46750;
  assign po0755 = n46749 | n46751;
  assign n46753 = ~pi0332 & pi0599;
  assign n46754 = ~n46741 & ~n46753;
  assign n46755 = pi0599 & n46741;
  assign po0756 = ~n46754 & ~n46755;
  assign n46757 = ~pi0332 & pi0600;
  assign n46758 = ~n46726 & ~n46757;
  assign po0757 = ~n46727 & ~n46758;
  assign n46760 = ~pi0806 & ~pi0989;
  assign n46761 = ~pi0601 & pi0806;
  assign n46762 = ~pi0332 & ~n46760;
  assign po0758 = ~n46761 & n46762;
  assign n46764 = ~pi0230 & pi0602;
  assign n46765 = ~pi0715 & ~pi1160;
  assign n46766 = pi0715 & pi1160;
  assign n46767 = pi0790 & ~n46765;
  assign n46768 = ~n46766 & n46767;
  assign n46769 = pi0230 & n16644;
  assign n46770 = ~n17856 & n46769;
  assign n46771 = ~n19146 & ~n19342;
  assign n46772 = ~n46768 & n46771;
  assign n46773 = n46770 & n46772;
  assign n46774 = n19151 & n46773;
  assign po0759 = n46764 | n46774;
  assign n46776 = pi0871 & pi0966;
  assign n46777 = pi0872 & pi0966;
  assign n46778 = pi0832 & ~pi1100;
  assign n46779 = ~pi0980 & pi1038;
  assign n46780 = pi1060 & n46779;
  assign n46781 = pi0952 & ~pi1061;
  assign n46782 = n46780 & n46781;
  assign n46783 = n46778 & n46782;
  assign po0897 = pi0832 & n46782;
  assign n46785 = ~pi0603 & ~po0897;
  assign n46786 = ~pi0966 & ~n46783;
  assign n46787 = ~n46785 & n46786;
  assign n46788 = ~n46776 & ~n46777;
  assign po0760 = n46787 | ~n46788;
  assign n46790 = pi0823 & n16657;
  assign n46791 = ~pi0779 & n46790;
  assign n46792 = ~pi0299 & pi0983;
  assign n46793 = pi0907 & n46792;
  assign n46794 = pi0604 & ~n46793;
  assign n46795 = ~n46790 & n46794;
  assign po0761 = n46791 | n46795;
  assign n46797 = ~pi0605 & ~n46725;
  assign n46798 = ~pi0332 & ~n46731;
  assign po0762 = ~n46797 & n46798;
  assign n46800 = ~pi0606 & ~po0897;
  assign n46801 = ~pi1104 & po0897;
  assign n46802 = ~n46800 & ~n46801;
  assign n46803 = ~pi0966 & ~n46802;
  assign n46804 = ~pi0837 & pi0966;
  assign po0763 = ~n46803 & ~n46804;
  assign n46806 = ~pi0607 & ~po0897;
  assign n46807 = ~pi1107 & po0897;
  assign n46808 = ~pi0966 & ~n46806;
  assign po0764 = ~n46807 & n46808;
  assign n46810 = ~pi0608 & ~po0897;
  assign n46811 = ~pi1116 & po0897;
  assign n46812 = ~pi0966 & ~n46810;
  assign po0765 = ~n46811 & n46812;
  assign n46814 = ~pi0609 & ~po0897;
  assign n46815 = ~pi1118 & po0897;
  assign n46816 = ~pi0966 & ~n46814;
  assign po0766 = ~n46815 & n46816;
  assign n46818 = ~pi0610 & ~po0897;
  assign n46819 = ~pi1113 & po0897;
  assign n46820 = ~pi0966 & ~n46818;
  assign po0767 = ~n46819 & n46820;
  assign n46822 = ~pi0611 & ~po0897;
  assign n46823 = ~pi1114 & po0897;
  assign n46824 = ~pi0966 & ~n46822;
  assign po0768 = ~n46823 & n46824;
  assign n46826 = ~pi0612 & ~po0897;
  assign n46827 = ~pi1111 & po0897;
  assign n46828 = ~pi0966 & ~n46826;
  assign po0769 = ~n46827 & n46828;
  assign n46830 = ~pi0613 & ~po0897;
  assign n46831 = ~pi1115 & po0897;
  assign n46832 = ~pi0966 & ~n46830;
  assign po0770 = ~n46831 & n46832;
  assign n46834 = ~pi0614 & ~po0897;
  assign n46835 = ~pi1102 & po0897;
  assign n46836 = ~pi0966 & ~n46834;
  assign n46837 = ~n46835 & n46836;
  assign po0771 = n46776 | n46837;
  assign n46839 = pi0907 & n46747;
  assign n46840 = ~pi0615 & ~n46839;
  assign n46841 = pi0779 & pi0797;
  assign n46842 = n6195 & n46841;
  assign po0772 = n46840 | n46842;
  assign n46844 = ~pi0616 & ~po0897;
  assign n46845 = ~pi1101 & po0897;
  assign n46846 = ~pi0966 & ~n46844;
  assign n46847 = ~n46845 & n46846;
  assign po0773 = n46777 | n46847;
  assign n46849 = ~pi0617 & ~po0897;
  assign n46850 = ~pi1105 & po0897;
  assign n46851 = ~n46849 & ~n46850;
  assign n46852 = ~pi0966 & ~n46851;
  assign n46853 = ~pi0850 & pi0966;
  assign po0774 = ~n46852 & ~n46853;
  assign n46855 = ~pi0618 & ~po0897;
  assign n46856 = ~pi1117 & po0897;
  assign n46857 = ~pi0966 & ~n46855;
  assign po0775 = ~n46856 & n46857;
  assign n46859 = ~pi0619 & ~po0897;
  assign n46860 = ~pi1122 & po0897;
  assign n46861 = ~pi0966 & ~n46859;
  assign po0776 = ~n46860 & n46861;
  assign n46863 = ~pi0620 & ~po0897;
  assign n46864 = ~pi1112 & po0897;
  assign n46865 = ~pi0966 & ~n46863;
  assign po0777 = ~n46864 & n46865;
  assign n46867 = ~pi0621 & ~po0897;
  assign n46868 = ~pi1108 & po0897;
  assign n46869 = ~pi0966 & ~n46867;
  assign po0778 = ~n46868 & n46869;
  assign n46871 = ~pi0622 & ~po0897;
  assign n46872 = ~pi1109 & po0897;
  assign n46873 = ~pi0966 & ~n46871;
  assign po0779 = ~n46872 & n46873;
  assign n46875 = ~pi0623 & ~po0897;
  assign n46876 = ~pi1106 & po0897;
  assign n46877 = ~pi0966 & ~n46875;
  assign po0780 = ~n46876 & n46877;
  assign n46879 = pi0831 & n17167;
  assign n46880 = ~pi0780 & n46879;
  assign n46881 = pi0947 & n46792;
  assign n46882 = pi0624 & ~n46881;
  assign n46883 = ~n46879 & n46882;
  assign po0781 = n46880 | n46883;
  assign n46885 = pi0832 & ~pi0973;
  assign n46886 = ~pi1054 & pi1066;
  assign n46887 = pi1088 & n46886;
  assign n46888 = n46885 & n46887;
  assign po0954 = ~pi0953 & n46888;
  assign n46890 = ~pi0625 & ~po0954;
  assign n46891 = ~pi1116 & po0954;
  assign n46892 = ~pi0962 & ~n46890;
  assign po0782 = ~n46891 & n46892;
  assign n46894 = ~pi0626 & ~po0897;
  assign n46895 = ~pi1121 & po0897;
  assign n46896 = ~pi0966 & ~n46894;
  assign po0783 = ~n46895 & n46896;
  assign n46898 = ~pi0627 & ~po0954;
  assign n46899 = ~pi1117 & po0954;
  assign n46900 = ~pi0962 & ~n46898;
  assign po0784 = ~n46899 & n46900;
  assign n46902 = ~pi0628 & ~po0954;
  assign n46903 = ~pi1119 & po0954;
  assign n46904 = ~pi0962 & ~n46902;
  assign po0785 = ~n46903 & n46904;
  assign n46906 = ~pi0629 & ~po0897;
  assign n46907 = ~pi1119 & po0897;
  assign n46908 = ~pi0966 & ~n46906;
  assign po0786 = ~n46907 & n46908;
  assign n46910 = ~pi0630 & ~po0897;
  assign n46911 = ~pi1120 & po0897;
  assign n46912 = ~pi0966 & ~n46910;
  assign po0787 = ~n46911 & n46912;
  assign n46914 = ~pi1113 & po0954;
  assign n46915 = pi0631 & ~po0954;
  assign n46916 = ~pi0962 & ~n46914;
  assign po0788 = ~n46915 & n46916;
  assign n46918 = ~pi1115 & po0954;
  assign n46919 = pi0632 & ~po0954;
  assign n46920 = ~pi0962 & ~n46918;
  assign po0789 = ~n46919 & n46920;
  assign n46922 = ~pi0633 & ~po0897;
  assign n46923 = ~pi1110 & po0897;
  assign n46924 = ~pi0966 & ~n46922;
  assign po0790 = ~n46923 & n46924;
  assign n46926 = ~pi0634 & ~po0954;
  assign n46927 = ~pi1110 & po0954;
  assign n46928 = ~pi0962 & ~n46926;
  assign po0791 = ~n46927 & n46928;
  assign n46930 = ~pi1112 & po0954;
  assign n46931 = pi0635 & ~po0954;
  assign n46932 = ~pi0962 & ~n46930;
  assign po0792 = ~n46931 & n46932;
  assign n46934 = ~pi0636 & ~po0897;
  assign n46935 = ~pi1127 & po0897;
  assign n46936 = ~pi0966 & ~n46934;
  assign po0793 = ~n46935 & n46936;
  assign n46938 = ~pi0637 & ~po0954;
  assign n46939 = ~pi1105 & po0954;
  assign n46940 = ~pi0962 & ~n46938;
  assign po0794 = ~n46939 & n46940;
  assign n46942 = ~pi0638 & ~po0954;
  assign n46943 = ~pi1107 & po0954;
  assign n46944 = ~pi0962 & ~n46942;
  assign po0795 = ~n46943 & n46944;
  assign n46946 = ~pi0639 & ~po0954;
  assign n46947 = ~pi1109 & po0954;
  assign n46948 = ~pi0962 & ~n46946;
  assign po0796 = ~n46947 & n46948;
  assign n46950 = ~pi0640 & ~po0897;
  assign n46951 = ~pi1128 & po0897;
  assign n46952 = ~pi0966 & ~n46950;
  assign po0797 = ~n46951 & n46952;
  assign n46954 = ~pi0641 & ~po0954;
  assign n46955 = ~pi1121 & po0954;
  assign n46956 = ~pi0962 & ~n46954;
  assign po0798 = ~n46955 & n46956;
  assign n46958 = ~pi0642 & ~po0897;
  assign n46959 = ~pi1103 & po0897;
  assign n46960 = ~pi0966 & ~n46958;
  assign po0799 = ~n46959 & n46960;
  assign n46962 = ~pi0643 & ~po0954;
  assign n46963 = ~pi1104 & po0954;
  assign n46964 = ~pi0962 & ~n46962;
  assign po0800 = ~n46963 & n46964;
  assign n46966 = ~pi0644 & ~po0897;
  assign n46967 = ~pi1123 & po0897;
  assign n46968 = ~pi0966 & ~n46966;
  assign po0801 = ~n46967 & n46968;
  assign n46970 = ~pi0645 & ~po0897;
  assign n46971 = ~pi1125 & po0897;
  assign n46972 = ~pi0966 & ~n46970;
  assign po0802 = ~n46971 & n46972;
  assign n46974 = ~pi1114 & po0954;
  assign n46975 = pi0646 & ~po0954;
  assign n46976 = ~pi0962 & ~n46974;
  assign po0803 = ~n46975 & n46976;
  assign n46978 = ~pi0647 & ~po0954;
  assign n46979 = ~pi1120 & po0954;
  assign n46980 = ~pi0962 & ~n46978;
  assign po0804 = ~n46979 & n46980;
  assign n46982 = ~pi0648 & ~po0954;
  assign n46983 = ~pi1122 & po0954;
  assign n46984 = ~pi0962 & ~n46982;
  assign po0805 = ~n46983 & n46984;
  assign n46986 = ~pi1126 & po0954;
  assign n46987 = pi0649 & ~po0954;
  assign n46988 = ~pi0962 & ~n46986;
  assign po0806 = ~n46987 & n46988;
  assign n46990 = ~pi1127 & po0954;
  assign n46991 = pi0650 & ~po0954;
  assign n46992 = ~pi0962 & ~n46990;
  assign po0807 = ~n46991 & n46992;
  assign n46994 = ~pi0651 & ~po0897;
  assign n46995 = ~pi1130 & po0897;
  assign n46996 = ~pi0966 & ~n46994;
  assign po0808 = ~n46995 & n46996;
  assign n46998 = ~pi0652 & ~po0897;
  assign n46999 = ~pi1131 & po0897;
  assign n47000 = ~pi0966 & ~n46998;
  assign po0809 = ~n46999 & n47000;
  assign n47002 = ~pi0653 & ~po0897;
  assign n47003 = ~pi1129 & po0897;
  assign n47004 = ~pi0966 & ~n47002;
  assign po0810 = ~n47003 & n47004;
  assign n47006 = ~pi1130 & po0954;
  assign n47007 = pi0654 & ~po0954;
  assign n47008 = ~pi0962 & ~n47006;
  assign po0811 = ~n47007 & n47008;
  assign n47010 = ~pi1124 & po0954;
  assign n47011 = pi0655 & ~po0954;
  assign n47012 = ~pi0962 & ~n47010;
  assign po0812 = ~n47011 & n47012;
  assign n47014 = ~pi0656 & ~po0897;
  assign n47015 = ~pi1126 & po0897;
  assign n47016 = ~pi0966 & ~n47014;
  assign po0813 = ~n47015 & n47016;
  assign n47018 = ~pi1131 & po0954;
  assign n47019 = pi0657 & ~po0954;
  assign n47020 = ~pi0962 & ~n47018;
  assign po0814 = ~n47019 & n47020;
  assign n47022 = ~pi0658 & ~po0897;
  assign n47023 = ~pi1124 & po0897;
  assign n47024 = ~pi0966 & ~n47022;
  assign po0815 = ~n47023 & n47024;
  assign n47026 = pi0266 & pi0992;
  assign n47027 = ~pi0280 & n47026;
  assign n47028 = ~pi0269 & n47027;
  assign n47029 = ~pi0281 & n47028;
  assign n47030 = ~pi0270 & ~pi0277;
  assign n47031 = ~pi0282 & n47030;
  assign n47032 = n47029 & n47031;
  assign n47033 = ~pi0264 & n47032;
  assign n47034 = ~pi0265 & n47033;
  assign po0959 = ~pi0274 & n47034;
  assign n47036 = pi0274 & ~n47034;
  assign po0816 = ~po0959 & ~n47036;
  assign n47038 = ~pi0660 & ~po0954;
  assign n47039 = ~pi1118 & po0954;
  assign n47040 = ~pi0962 & ~n47038;
  assign po0817 = ~n47039 & n47040;
  assign n47042 = ~pi0661 & ~po0954;
  assign n47043 = ~pi1101 & po0954;
  assign n47044 = ~pi0962 & ~n47042;
  assign po0818 = ~n47043 & n47044;
  assign n47046 = ~pi0662 & ~po0954;
  assign n47047 = ~pi1102 & po0954;
  assign n47048 = ~pi0962 & ~n47046;
  assign po0819 = ~n47047 & n47048;
  assign n47050 = ~pi0223 & ~pi0224;
  assign n47051 = ~pi0199 & ~pi0257;
  assign n47052 = pi0199 & ~pi1065;
  assign n47053 = ~n47050 & ~n47051;
  assign n47054 = ~n47052 & n47053;
  assign n47055 = ~pi0592 & n8041;
  assign n47056 = pi0464 & n47055;
  assign n47057 = pi0588 & ~n47056;
  assign n47058 = ~pi0591 & pi0592;
  assign n47059 = pi0365 & n47058;
  assign n47060 = pi0334 & pi0591;
  assign n47061 = ~pi0592 & n47060;
  assign n47062 = ~n47059 & ~n47061;
  assign n47063 = ~pi0590 & ~n47062;
  assign n47064 = pi0590 & ~pi0591;
  assign n47065 = ~pi0592 & n47064;
  assign n47066 = pi0323 & n47065;
  assign n47067 = ~pi0588 & ~n47066;
  assign n47068 = ~n47063 & n47067;
  assign n47069 = n47050 & ~n47057;
  assign n47070 = ~n47068 & n47069;
  assign n47071 = ~n47054 & ~n47070;
  assign n47072 = n7643 & ~n47071;
  assign n47073 = ~pi1137 & ~pi1138;
  assign n47074 = ~pi1134 & n47073;
  assign n47075 = ~pi0784 & ~pi1136;
  assign n47076 = ~pi0634 & pi1136;
  assign n47077 = pi1135 & ~n47075;
  assign n47078 = ~n47076 & n47077;
  assign n47079 = ~pi0815 & ~pi1136;
  assign n47080 = ~pi0633 & pi1136;
  assign n47081 = ~pi1135 & ~n47079;
  assign n47082 = ~n47080 & n47081;
  assign n47083 = ~n47078 & ~n47082;
  assign n47084 = n47074 & ~n47083;
  assign n47085 = pi1135 & n47073;
  assign n47086 = pi1136 & ~n47085;
  assign n47087 = ~pi0766 & n47086;
  assign n47088 = ~pi0855 & ~pi1136;
  assign n47089 = ~pi0700 & pi1135;
  assign n47090 = pi1135 & ~pi1136;
  assign n47091 = pi1134 & n47073;
  assign n47092 = ~n47090 & n47091;
  assign n47093 = ~n47088 & ~n47089;
  assign n47094 = n47092 & n47093;
  assign n47095 = ~n47087 & n47094;
  assign n47096 = ~n47084 & ~n47095;
  assign n47097 = ~n7643 & ~n47096;
  assign po0820 = n47072 | n47097;
  assign n47099 = pi0429 & n47055;
  assign n47100 = pi0588 & ~n47099;
  assign n47101 = ~pi0590 & pi0591;
  assign n47102 = pi0404 & n47101;
  assign n47103 = ~pi0590 & pi0592;
  assign n47104 = ~pi0588 & ~n47103;
  assign n47105 = ~n47102 & n47104;
  assign n47106 = pi0380 & ~pi0591;
  assign n47107 = pi0592 & ~n47106;
  assign n47108 = ~n47105 & ~n47107;
  assign n47109 = pi0355 & n47065;
  assign n47110 = ~n47108 & ~n47109;
  assign n47111 = n47050 & ~n47100;
  assign n47112 = ~n47110 & n47111;
  assign n47113 = ~pi0199 & ~pi0292;
  assign n47114 = pi0199 & ~pi1084;
  assign n47115 = ~n47050 & ~n47113;
  assign n47116 = ~n47114 & n47115;
  assign n47117 = ~n47112 & ~n47116;
  assign n47118 = n7643 & ~n47117;
  assign n47119 = ~pi1135 & ~pi1136;
  assign n47120 = pi0872 & n47119;
  assign n47121 = ~pi0772 & ~pi1135;
  assign n47122 = ~pi0727 & pi1135;
  assign n47123 = pi1136 & ~n47121;
  assign n47124 = ~n47122 & n47123;
  assign n47125 = pi1134 & ~n47120;
  assign n47126 = ~n47124 & n47125;
  assign n47127 = ~n7643 & n47073;
  assign n47128 = pi0614 & ~pi1135;
  assign n47129 = pi0662 & pi1135;
  assign n47130 = pi1136 & ~n47128;
  assign n47131 = ~n47129 & n47130;
  assign n47132 = pi0811 & ~pi1135;
  assign n47133 = pi0785 & pi1135;
  assign n47134 = ~pi1136 & ~n47132;
  assign n47135 = ~n47133 & n47134;
  assign n47136 = ~n47131 & ~n47135;
  assign n47137 = ~pi1134 & ~n47136;
  assign n47138 = ~n47126 & n47127;
  assign n47139 = ~n47137 & n47138;
  assign po0821 = n47118 | n47139;
  assign n47141 = ~pi0665 & ~po0954;
  assign n47142 = ~pi1108 & po0954;
  assign n47143 = ~pi0962 & ~n47141;
  assign po0822 = ~n47142 & n47143;
  assign n47145 = ~pi0607 & ~pi1135;
  assign n47146 = ~pi0638 & pi1135;
  assign n47147 = pi1136 & ~n47145;
  assign n47148 = ~n47146 & n47147;
  assign n47149 = ~pi0790 & pi1135;
  assign n47150 = pi0799 & ~pi1135;
  assign n47151 = ~pi1136 & ~n47149;
  assign n47152 = ~n47150 & n47151;
  assign n47153 = ~n47148 & ~n47152;
  assign n47154 = n47074 & ~n47153;
  assign n47155 = ~pi0764 & n47086;
  assign n47156 = ~pi0691 & pi1135;
  assign n47157 = ~pi0873 & ~pi1136;
  assign n47158 = ~n47156 & ~n47157;
  assign n47159 = n47092 & n47158;
  assign n47160 = ~n47155 & n47159;
  assign n47161 = ~n47154 & ~n47160;
  assign n47162 = ~n7643 & ~n47161;
  assign n47163 = ~pi0199 & ~pi0297;
  assign n47164 = pi0199 & ~pi1044;
  assign n47165 = ~n47050 & ~n47163;
  assign n47166 = ~n47164 & n47165;
  assign n47167 = pi0443 & n47055;
  assign n47168 = pi0588 & ~n47167;
  assign n47169 = pi0456 & n47101;
  assign n47170 = n47104 & ~n47169;
  assign n47171 = pi0337 & ~pi0591;
  assign n47172 = pi0592 & ~n47171;
  assign n47173 = ~n47170 & ~n47172;
  assign n47174 = pi0441 & n47065;
  assign n47175 = ~n47173 & ~n47174;
  assign n47176 = n47050 & ~n47168;
  assign n47177 = ~n47175 & n47176;
  assign n47178 = ~n47166 & ~n47177;
  assign n47179 = n7643 & ~n47178;
  assign po0823 = n47162 | n47179;
  assign n47181 = pi0444 & n47055;
  assign n47182 = pi0588 & ~n47181;
  assign n47183 = pi0319 & n47101;
  assign n47184 = n47104 & ~n47183;
  assign n47185 = pi0338 & ~pi0591;
  assign n47186 = pi0592 & ~n47185;
  assign n47187 = ~n47184 & ~n47186;
  assign n47188 = pi0458 & n47065;
  assign n47189 = ~n47187 & ~n47188;
  assign n47190 = n47050 & ~n47182;
  assign n47191 = ~n47189 & n47190;
  assign n47192 = ~pi0199 & ~pi0294;
  assign n47193 = pi0199 & ~pi1072;
  assign n47194 = ~n47050 & ~n47192;
  assign n47195 = ~n47193 & n47194;
  assign n47196 = ~n47191 & ~n47195;
  assign n47197 = n7643 & ~n47196;
  assign n47198 = pi0871 & n47119;
  assign n47199 = ~pi0763 & ~pi1135;
  assign n47200 = ~pi0699 & pi1135;
  assign n47201 = pi1136 & ~n47199;
  assign n47202 = ~n47200 & n47201;
  assign n47203 = pi1134 & ~n47198;
  assign n47204 = ~n47202 & n47203;
  assign n47205 = pi0792 & ~pi1136;
  assign n47206 = pi0681 & pi1136;
  assign n47207 = pi1135 & ~n47205;
  assign n47208 = ~n47206 & n47207;
  assign n47209 = ~pi0809 & ~pi1136;
  assign n47210 = pi0642 & pi1136;
  assign n47211 = ~pi1135 & ~n47209;
  assign n47212 = ~n47210 & n47211;
  assign n47213 = ~n47208 & ~n47212;
  assign n47214 = ~pi1134 & ~n47213;
  assign n47215 = n47127 & ~n47204;
  assign n47216 = ~n47214 & n47215;
  assign po0824 = n47197 | n47216;
  assign n47218 = ~pi0603 & ~pi1135;
  assign n47219 = ~pi0680 & pi1135;
  assign n47220 = pi1136 & ~n47218;
  assign n47221 = ~n47219 & n47220;
  assign n47222 = ~pi0981 & ~pi1135;
  assign n47223 = ~pi0778 & pi1135;
  assign n47224 = ~pi1136 & ~n47222;
  assign n47225 = ~n47223 & n47224;
  assign n47226 = ~n47221 & ~n47225;
  assign n47227 = n47074 & ~n47226;
  assign n47228 = ~pi0759 & n47086;
  assign n47229 = ~pi0696 & pi1135;
  assign n47230 = ~pi0837 & ~pi1136;
  assign n47231 = ~n47229 & ~n47230;
  assign n47232 = n47092 & n47231;
  assign n47233 = ~n47228 & n47232;
  assign n47234 = ~n47227 & ~n47233;
  assign n47235 = ~n7643 & ~n47234;
  assign n47236 = ~pi0199 & ~pi0291;
  assign n47237 = pi0199 & ~pi1049;
  assign n47238 = ~n47050 & ~n47236;
  assign n47239 = ~n47237 & n47238;
  assign n47240 = pi0414 & n47055;
  assign n47241 = pi0588 & ~n47240;
  assign n47242 = pi0390 & n47101;
  assign n47243 = n47104 & ~n47242;
  assign n47244 = pi0363 & ~pi0591;
  assign n47245 = pi0592 & ~n47244;
  assign n47246 = ~n47243 & ~n47245;
  assign n47247 = pi0342 & n47065;
  assign n47248 = ~n47246 & ~n47247;
  assign n47249 = n47050 & ~n47241;
  assign n47250 = ~n47248 & n47249;
  assign n47251 = ~n47239 & ~n47250;
  assign n47252 = n7643 & ~n47251;
  assign po0825 = n47235 | n47252;
  assign n47254 = ~pi1125 & po0954;
  assign n47255 = pi0669 & ~po0954;
  assign n47256 = ~pi0962 & ~n47254;
  assign po0826 = ~n47255 & n47256;
  assign n47258 = ~pi0199 & ~pi0258;
  assign n47259 = pi0199 & ~pi1062;
  assign n47260 = ~n47050 & ~n47258;
  assign n47261 = ~n47259 & n47260;
  assign n47262 = pi0415 & n47055;
  assign n47263 = pi0588 & ~n47262;
  assign n47264 = pi0364 & n47058;
  assign n47265 = pi0391 & pi0591;
  assign n47266 = ~pi0592 & n47265;
  assign n47267 = ~n47264 & ~n47266;
  assign n47268 = ~pi0590 & ~n47267;
  assign n47269 = pi0343 & n47065;
  assign n47270 = ~pi0588 & ~n47269;
  assign n47271 = ~n47268 & n47270;
  assign n47272 = n47050 & ~n47263;
  assign n47273 = ~n47271 & n47272;
  assign n47274 = ~n47261 & ~n47273;
  assign n47275 = n7643 & ~n47274;
  assign n47276 = pi0723 & pi1135;
  assign n47277 = ~pi0852 & ~pi1136;
  assign n47278 = pi0745 & n47086;
  assign n47279 = ~n47276 & ~n47277;
  assign n47280 = n47092 & n47279;
  assign n47281 = ~n47278 & n47280;
  assign n47282 = pi0695 & pi1135;
  assign n47283 = pi1136 & n47073;
  assign n47284 = ~pi0612 & ~pi1135;
  assign n47285 = ~pi1134 & ~n47282;
  assign n47286 = ~n47284 & n47285;
  assign n47287 = n47283 & n47286;
  assign n47288 = ~n47281 & ~n47287;
  assign n47289 = ~n7643 & ~n47288;
  assign po0827 = n47275 | n47289;
  assign n47291 = ~pi0199 & ~pi0261;
  assign n47292 = pi0199 & ~pi1040;
  assign n47293 = ~n47050 & ~n47291;
  assign n47294 = ~n47292 & n47293;
  assign n47295 = pi0453 & n47055;
  assign n47296 = pi0588 & ~n47295;
  assign n47297 = pi0447 & n47058;
  assign n47298 = pi0333 & pi0591;
  assign n47299 = ~pi0592 & n47298;
  assign n47300 = ~n47297 & ~n47299;
  assign n47301 = ~pi0590 & ~n47300;
  assign n47302 = pi0327 & n47065;
  assign n47303 = ~pi0588 & ~n47302;
  assign n47304 = ~n47301 & n47303;
  assign n47305 = n47050 & ~n47296;
  assign n47306 = ~n47304 & n47305;
  assign n47307 = ~n47294 & ~n47306;
  assign n47308 = n7643 & ~n47307;
  assign n47309 = pi0724 & pi1135;
  assign n47310 = ~pi0865 & ~pi1136;
  assign n47311 = pi0741 & n47086;
  assign n47312 = ~n47309 & ~n47310;
  assign n47313 = n47092 & n47312;
  assign n47314 = ~n47311 & n47313;
  assign n47315 = pi0646 & pi1135;
  assign n47316 = ~pi0611 & ~pi1135;
  assign n47317 = ~pi1134 & ~n47315;
  assign n47318 = ~n47316 & n47317;
  assign n47319 = n47283 & n47318;
  assign n47320 = ~n47314 & ~n47319;
  assign n47321 = ~n7643 & ~n47320;
  assign po0828 = n47308 | n47321;
  assign n47323 = ~pi0616 & ~pi1135;
  assign n47324 = ~pi0661 & pi1135;
  assign n47325 = pi1136 & ~n47323;
  assign n47326 = ~n47324 & n47325;
  assign n47327 = ~pi0808 & ~pi1135;
  assign n47328 = ~pi0781 & pi1135;
  assign n47329 = ~pi1136 & ~n47327;
  assign n47330 = ~n47328 & n47329;
  assign n47331 = ~n47326 & ~n47330;
  assign n47332 = n47074 & ~n47331;
  assign n47333 = ~pi0758 & n47086;
  assign n47334 = ~pi0736 & pi1135;
  assign n47335 = ~pi0850 & ~pi1136;
  assign n47336 = ~n47334 & ~n47335;
  assign n47337 = n47092 & n47336;
  assign n47338 = ~n47333 & n47337;
  assign n47339 = ~n47332 & ~n47338;
  assign n47340 = ~n7643 & ~n47339;
  assign n47341 = ~pi0199 & ~pi0290;
  assign n47342 = pi0199 & ~pi1048;
  assign n47343 = ~n47050 & ~n47341;
  assign n47344 = ~n47342 & n47343;
  assign n47345 = pi0422 & n47055;
  assign n47346 = pi0588 & ~n47345;
  assign n47347 = pi0397 & n47101;
  assign n47348 = n47104 & ~n47347;
  assign n47349 = pi0372 & ~pi0591;
  assign n47350 = pi0592 & ~n47349;
  assign n47351 = ~n47348 & ~n47350;
  assign n47352 = pi0320 & n47065;
  assign n47353 = ~n47351 & ~n47352;
  assign n47354 = n47050 & ~n47346;
  assign n47355 = ~n47353 & n47354;
  assign n47356 = ~n47344 & ~n47355;
  assign n47357 = n7643 & ~n47356;
  assign po0829 = n47340 | n47357;
  assign n47359 = ~pi0617 & ~pi1135;
  assign n47360 = ~pi0637 & pi1135;
  assign n47361 = pi1136 & ~n47359;
  assign n47362 = ~n47360 & n47361;
  assign n47363 = ~pi0788 & pi1135;
  assign n47364 = pi0814 & ~pi1135;
  assign n47365 = ~pi1136 & ~n47363;
  assign n47366 = ~n47364 & n47365;
  assign n47367 = ~n47362 & ~n47366;
  assign n47368 = n47074 & ~n47367;
  assign n47369 = ~pi0749 & n47086;
  assign n47370 = ~pi0706 & pi1135;
  assign n47371 = ~pi0866 & ~pi1136;
  assign n47372 = ~n47370 & ~n47371;
  assign n47373 = n47092 & n47372;
  assign n47374 = ~n47369 & n47373;
  assign n47375 = ~n47368 & ~n47374;
  assign n47376 = ~n7643 & ~n47375;
  assign n47377 = ~pi0199 & ~pi0295;
  assign n47378 = pi0199 & ~pi1053;
  assign n47379 = ~n47050 & ~n47377;
  assign n47380 = ~n47378 & n47379;
  assign n47381 = pi0435 & n47055;
  assign n47382 = pi0588 & ~n47381;
  assign n47383 = pi0411 & n47101;
  assign n47384 = n47104 & ~n47383;
  assign n47385 = pi0387 & ~pi0591;
  assign n47386 = pi0592 & ~n47385;
  assign n47387 = ~n47384 & ~n47386;
  assign n47388 = pi0452 & n47065;
  assign n47389 = ~n47387 & ~n47388;
  assign n47390 = n47050 & ~n47382;
  assign n47391 = ~n47389 & n47390;
  assign n47392 = ~n47380 & ~n47391;
  assign n47393 = n7643 & ~n47392;
  assign po0830 = n47376 | n47393;
  assign n47395 = ~pi0199 & ~pi0256;
  assign n47396 = pi0199 & ~pi1070;
  assign n47397 = ~n47050 & ~n47395;
  assign n47398 = ~n47396 & n47397;
  assign n47399 = pi0437 & n47055;
  assign n47400 = pi0588 & ~n47399;
  assign n47401 = pi0336 & n47058;
  assign n47402 = pi0463 & pi0591;
  assign n47403 = ~pi0592 & n47402;
  assign n47404 = ~n47401 & ~n47403;
  assign n47405 = ~pi0590 & ~n47404;
  assign n47406 = pi0362 & n47065;
  assign n47407 = ~pi0588 & ~n47406;
  assign n47408 = ~n47405 & n47407;
  assign n47409 = n47050 & ~n47400;
  assign n47410 = ~n47408 & n47409;
  assign n47411 = ~n47398 & ~n47410;
  assign n47412 = n7643 & ~n47411;
  assign n47413 = pi0859 & n47119;
  assign n47414 = ~pi0743 & ~pi1135;
  assign n47415 = ~pi0735 & pi1135;
  assign n47416 = pi1136 & ~n47414;
  assign n47417 = ~n47415 & n47416;
  assign n47418 = pi1134 & ~n47413;
  assign n47419 = ~n47417 & n47418;
  assign n47420 = pi0622 & ~pi1135;
  assign n47421 = pi0639 & pi1135;
  assign n47422 = pi1136 & ~n47420;
  assign n47423 = ~n47421 & n47422;
  assign n47424 = pi0804 & ~pi1135;
  assign n47425 = pi0783 & pi1135;
  assign n47426 = ~pi1136 & ~n47424;
  assign n47427 = ~n47425 & n47426;
  assign n47428 = ~n47423 & ~n47427;
  assign n47429 = ~pi1134 & ~n47428;
  assign n47430 = n47127 & ~n47419;
  assign n47431 = ~n47429 & n47430;
  assign po0831 = n47412 | n47431;
  assign n47433 = pi0876 & n47119;
  assign n47434 = ~pi0748 & ~pi1135;
  assign n47435 = ~pi0730 & pi1135;
  assign n47436 = pi1136 & ~n47434;
  assign n47437 = ~n47435 & n47436;
  assign n47438 = ~n47433 & ~n47437;
  assign n47439 = n47091 & ~n47438;
  assign n47440 = ~pi0623 & n47086;
  assign n47441 = pi0789 & n47090;
  assign n47442 = ~pi0710 & pi1135;
  assign n47443 = pi1136 & ~n47442;
  assign n47444 = ~pi0803 & ~pi1135;
  assign n47445 = ~n47441 & ~n47444;
  assign n47446 = ~n47443 & n47445;
  assign n47447 = n47074 & ~n47440;
  assign n47448 = ~n47446 & n47447;
  assign n47449 = ~n47439 & ~n47448;
  assign n47450 = ~n7643 & ~n47449;
  assign n47451 = ~pi0199 & ~pi0296;
  assign n47452 = pi0199 & ~pi1037;
  assign n47453 = ~n47050 & ~n47451;
  assign n47454 = ~n47452 & n47453;
  assign n47455 = pi0436 & n47055;
  assign n47456 = pi0588 & ~n47455;
  assign n47457 = pi0412 & n47101;
  assign n47458 = n47104 & ~n47457;
  assign n47459 = pi0388 & ~pi0591;
  assign n47460 = pi0592 & ~n47459;
  assign n47461 = ~n47458 & ~n47460;
  assign n47462 = pi0455 & n47065;
  assign n47463 = ~n47461 & ~n47462;
  assign n47464 = n47050 & ~n47456;
  assign n47465 = ~n47463 & n47464;
  assign n47466 = ~n47454 & ~n47465;
  assign n47467 = n7643 & ~n47466;
  assign po0832 = n47450 | n47467;
  assign n47469 = ~pi0606 & ~pi1135;
  assign n47470 = ~pi0643 & pi1135;
  assign n47471 = pi1136 & ~n47469;
  assign n47472 = ~n47470 & n47471;
  assign n47473 = ~pi0787 & pi1135;
  assign n47474 = pi0812 & ~pi1135;
  assign n47475 = ~pi1136 & ~n47473;
  assign n47476 = ~n47474 & n47475;
  assign n47477 = ~n47472 & ~n47476;
  assign n47478 = n47074 & ~n47477;
  assign n47479 = ~pi0746 & n47086;
  assign n47480 = ~pi0729 & pi1135;
  assign n47481 = ~pi0881 & ~pi1136;
  assign n47482 = ~n47480 & ~n47481;
  assign n47483 = n47092 & n47482;
  assign n47484 = ~n47479 & n47483;
  assign n47485 = ~n47478 & ~n47484;
  assign n47486 = ~n7643 & ~n47485;
  assign n47487 = ~pi0199 & ~pi0293;
  assign n47488 = pi0199 & ~pi1059;
  assign n47489 = ~n47050 & ~n47487;
  assign n47490 = ~n47488 & n47489;
  assign n47491 = pi0434 & n47055;
  assign n47492 = pi0588 & ~n47491;
  assign n47493 = pi0410 & n47101;
  assign n47494 = n47104 & ~n47493;
  assign n47495 = pi0386 & ~pi0591;
  assign n47496 = pi0592 & ~n47495;
  assign n47497 = ~n47494 & ~n47496;
  assign n47498 = pi0361 & n47065;
  assign n47499 = ~n47497 & ~n47498;
  assign n47500 = n47050 & ~n47492;
  assign n47501 = ~n47499 & n47500;
  assign n47502 = ~n47490 & ~n47501;
  assign n47503 = n7643 & ~n47502;
  assign po0833 = n47486 | n47503;
  assign n47505 = ~pi0199 & ~pi0259;
  assign n47506 = pi0199 & ~pi1069;
  assign n47507 = ~n47050 & ~n47505;
  assign n47508 = ~n47506 & n47507;
  assign n47509 = pi0416 & n47055;
  assign n47510 = pi0588 & ~n47509;
  assign n47511 = pi0366 & n47058;
  assign n47512 = pi0335 & pi0591;
  assign n47513 = ~pi0592 & n47512;
  assign n47514 = ~n47511 & ~n47513;
  assign n47515 = ~pi0590 & ~n47514;
  assign n47516 = pi0344 & n47065;
  assign n47517 = ~pi0588 & ~n47516;
  assign n47518 = ~n47515 & n47517;
  assign n47519 = n47050 & ~n47510;
  assign n47520 = ~n47518 & n47519;
  assign n47521 = ~n47508 & ~n47520;
  assign n47522 = n7643 & ~n47521;
  assign n47523 = pi0704 & pi1135;
  assign n47524 = ~pi0870 & ~pi1136;
  assign n47525 = pi0742 & n47086;
  assign n47526 = ~n47523 & ~n47524;
  assign n47527 = n47092 & n47526;
  assign n47528 = ~n47525 & n47527;
  assign n47529 = pi0635 & pi1135;
  assign n47530 = ~pi0620 & ~pi1135;
  assign n47531 = ~pi1134 & ~n47529;
  assign n47532 = ~n47530 & n47531;
  assign n47533 = n47283 & n47532;
  assign n47534 = ~n47528 & ~n47533;
  assign n47535 = ~n7643 & ~n47534;
  assign po0834 = n47522 | n47535;
  assign n47537 = ~pi0199 & ~pi0260;
  assign n47538 = pi0199 & ~pi1067;
  assign n47539 = ~n47050 & ~n47537;
  assign n47540 = ~n47538 & n47539;
  assign n47541 = pi0418 & n47055;
  assign n47542 = pi0588 & ~n47541;
  assign n47543 = pi0368 & n47058;
  assign n47544 = pi0393 & pi0591;
  assign n47545 = ~pi0592 & n47544;
  assign n47546 = ~n47543 & ~n47545;
  assign n47547 = ~pi0590 & ~n47546;
  assign n47548 = pi0346 & n47065;
  assign n47549 = ~pi0588 & ~n47548;
  assign n47550 = ~n47547 & n47549;
  assign n47551 = n47050 & ~n47542;
  assign n47552 = ~n47550 & n47551;
  assign n47553 = ~n47540 & ~n47552;
  assign n47554 = n7643 & ~n47553;
  assign n47555 = pi0688 & pi1135;
  assign n47556 = ~pi0856 & ~pi1136;
  assign n47557 = pi0760 & n47086;
  assign n47558 = ~n47555 & ~n47556;
  assign n47559 = n47092 & n47558;
  assign n47560 = ~n47557 & n47559;
  assign n47561 = pi0632 & pi1135;
  assign n47562 = ~pi0613 & ~pi1135;
  assign n47563 = ~pi1134 & ~n47561;
  assign n47564 = ~n47562 & n47563;
  assign n47565 = n47283 & n47564;
  assign n47566 = ~n47560 & ~n47565;
  assign n47567 = ~n7643 & ~n47566;
  assign po0835 = n47554 | n47567;
  assign n47569 = ~pi0199 & ~pi0255;
  assign n47570 = pi0199 & ~pi1036;
  assign n47571 = ~n47050 & ~n47569;
  assign n47572 = ~n47570 & n47571;
  assign n47573 = pi0438 & n47055;
  assign n47574 = pi0588 & ~n47573;
  assign n47575 = pi0389 & n47058;
  assign n47576 = pi0413 & pi0591;
  assign n47577 = ~pi0592 & n47576;
  assign n47578 = ~n47575 & ~n47577;
  assign n47579 = ~pi0590 & ~n47578;
  assign n47580 = pi0450 & n47065;
  assign n47581 = ~pi0588 & ~n47580;
  assign n47582 = ~n47579 & n47581;
  assign n47583 = n47050 & ~n47574;
  assign n47584 = ~n47582 & n47583;
  assign n47585 = ~n47572 & ~n47584;
  assign n47586 = n7643 & ~n47585;
  assign n47587 = ~pi0791 & ~pi1136;
  assign n47588 = ~pi0665 & pi1136;
  assign n47589 = pi1135 & ~n47587;
  assign n47590 = ~n47588 & n47589;
  assign n47591 = ~pi0810 & ~pi1136;
  assign n47592 = ~pi0621 & pi1136;
  assign n47593 = ~pi1135 & ~n47591;
  assign n47594 = ~n47592 & n47593;
  assign n47595 = ~n47590 & ~n47594;
  assign n47596 = n47074 & ~n47595;
  assign n47597 = ~pi0739 & n47086;
  assign n47598 = ~pi0874 & ~pi1136;
  assign n47599 = ~pi0690 & pi1135;
  assign n47600 = ~n47598 & ~n47599;
  assign n47601 = n47092 & n47600;
  assign n47602 = ~n47597 & n47601;
  assign n47603 = ~n47596 & ~n47602;
  assign n47604 = ~n7643 & ~n47603;
  assign po0836 = n47586 | n47604;
  assign n47606 = ~pi0680 & ~po0954;
  assign n47607 = ~pi1100 & po0954;
  assign n47608 = ~pi0962 & ~n47606;
  assign po0837 = ~n47607 & n47608;
  assign n47610 = ~pi0681 & ~po0954;
  assign n47611 = ~pi1103 & po0954;
  assign n47612 = ~pi0962 & ~n47610;
  assign po0838 = ~n47611 & n47612;
  assign n47614 = ~pi0199 & ~pi0251;
  assign n47615 = pi0199 & ~pi1039;
  assign n47616 = ~n47050 & ~n47614;
  assign n47617 = ~n47615 & n47616;
  assign n47618 = pi0417 & n47055;
  assign n47619 = pi0588 & ~n47618;
  assign n47620 = pi0367 & n47058;
  assign n47621 = pi0392 & pi0591;
  assign n47622 = ~pi0592 & n47621;
  assign n47623 = ~n47620 & ~n47622;
  assign n47624 = ~pi0590 & ~n47623;
  assign n47625 = pi0345 & n47065;
  assign n47626 = ~pi0588 & ~n47625;
  assign n47627 = ~n47624 & n47626;
  assign n47628 = n47050 & ~n47619;
  assign n47629 = ~n47627 & n47628;
  assign n47630 = ~n47617 & ~n47629;
  assign n47631 = n7643 & ~n47630;
  assign n47632 = pi0686 & pi1135;
  assign n47633 = ~pi0848 & ~pi1136;
  assign n47634 = pi0757 & n47086;
  assign n47635 = ~n47632 & ~n47633;
  assign n47636 = n47092 & n47635;
  assign n47637 = ~n47634 & n47636;
  assign n47638 = pi0631 & pi1135;
  assign n47639 = ~pi0610 & ~pi1135;
  assign n47640 = ~pi1134 & ~n47638;
  assign n47641 = ~n47639 & n47640;
  assign n47642 = n47283 & n47641;
  assign n47643 = ~n47637 & ~n47642;
  assign n47644 = ~n7643 & ~n47643;
  assign po0839 = n47631 | n47644;
  assign po0980 = pi0953 & n46888;
  assign n47647 = ~pi1130 & po0980;
  assign n47648 = pi0684 & ~po0980;
  assign n47649 = ~pi0962 & ~n47647;
  assign po0841 = ~n47648 & n47649;
  assign n47651 = pi0590 & ~pi0592;
  assign n47652 = pi0357 & n47651;
  assign n47653 = pi0382 & n47103;
  assign n47654 = ~n47652 & ~n47653;
  assign n47655 = ~pi0591 & ~n47654;
  assign n47656 = pi0406 & ~pi0592;
  assign n47657 = n47101 & n47656;
  assign n47658 = ~n47655 & ~n47657;
  assign n47659 = ~pi0588 & ~n47658;
  assign n47660 = ~pi0591 & ~pi0592;
  assign n47661 = pi0588 & ~pi0590;
  assign n47662 = pi0430 & n47660;
  assign n47663 = n47661 & n47662;
  assign n47664 = ~n47659 & ~n47663;
  assign n47665 = n47050 & ~n47664;
  assign n47666 = pi0199 & ~pi1076;
  assign n47667 = ~n47050 & ~n47666;
  assign n47668 = ~n42880 & n47667;
  assign n47669 = ~n47665 & ~n47668;
  assign n47670 = n7643 & ~n47669;
  assign n47671 = pi0860 & n47119;
  assign n47672 = pi0744 & ~pi1135;
  assign n47673 = pi0728 & pi1135;
  assign n47674 = pi1136 & ~n47672;
  assign n47675 = ~n47673 & n47674;
  assign n47676 = ~n47671 & ~n47675;
  assign n47677 = n47091 & ~n47676;
  assign n47678 = pi1136 & ~n47073;
  assign n47679 = ~pi1134 & ~n47678;
  assign n47680 = ~pi0652 & ~pi1135;
  assign n47681 = pi0657 & pi1135;
  assign n47682 = pi1136 & ~n47680;
  assign n47683 = ~n47681 & n47682;
  assign n47684 = pi0813 & n47073;
  assign n47685 = n47119 & n47684;
  assign n47686 = ~n47683 & ~n47685;
  assign n47687 = n47679 & ~n47686;
  assign n47688 = ~n47677 & ~n47687;
  assign n47689 = ~n7643 & ~n47688;
  assign po0842 = n47670 | n47689;
  assign n47691 = ~pi1113 & po0980;
  assign n47692 = pi0686 & ~po0980;
  assign n47693 = ~pi0962 & ~n47691;
  assign po0843 = ~n47692 & n47693;
  assign n47695 = ~pi0687 & ~po0980;
  assign n47696 = ~pi1127 & po0980;
  assign n47697 = ~pi0962 & ~n47695;
  assign po0844 = ~n47696 & n47697;
  assign n47699 = ~pi1115 & po0980;
  assign n47700 = pi0688 & ~po0980;
  assign n47701 = ~pi0962 & ~n47699;
  assign po0845 = ~n47700 & n47701;
  assign n47703 = pi0351 & n47651;
  assign n47704 = pi0376 & n47103;
  assign n47705 = ~n47703 & ~n47704;
  assign n47706 = ~pi0591 & ~n47705;
  assign n47707 = pi0401 & ~pi0592;
  assign n47708 = n47101 & n47707;
  assign n47709 = ~n47706 & ~n47708;
  assign n47710 = ~pi0588 & ~n47709;
  assign n47711 = pi0426 & n47660;
  assign n47712 = n47661 & n47711;
  assign n47713 = ~n47710 & ~n47712;
  assign n47714 = n47050 & ~n47713;
  assign n47715 = pi0199 & ~pi1079;
  assign n47716 = ~pi0199 & n42849;
  assign n47717 = ~n47050 & ~n47715;
  assign n47718 = ~n47716 & n47717;
  assign n47719 = ~n47714 & ~n47718;
  assign n47720 = n7643 & ~n47719;
  assign n47721 = pi0798 & n47119;
  assign n47722 = ~pi0658 & ~pi1135;
  assign n47723 = pi0655 & pi1135;
  assign n47724 = pi1136 & ~n47722;
  assign n47725 = ~n47723 & n47724;
  assign n47726 = ~n47721 & ~n47725;
  assign n47727 = n47074 & ~n47726;
  assign n47728 = pi0752 & n47086;
  assign n47729 = ~pi0703 & pi1135;
  assign n47730 = ~pi0843 & ~pi1136;
  assign n47731 = ~n47729 & ~n47730;
  assign n47732 = n47092 & n47731;
  assign n47733 = ~n47728 & n47732;
  assign n47734 = ~n47727 & ~n47733;
  assign n47735 = ~n7643 & ~n47734;
  assign po0846 = n47720 | n47735;
  assign n47737 = ~pi0690 & ~po0980;
  assign n47738 = ~pi1108 & po0980;
  assign n47739 = ~pi0962 & ~n47737;
  assign po0847 = ~n47738 & n47739;
  assign n47741 = ~pi0691 & ~po0980;
  assign n47742 = ~pi1107 & po0980;
  assign n47743 = ~pi0962 & ~n47741;
  assign po0848 = ~n47742 & n47743;
  assign n47745 = pi0352 & n47651;
  assign n47746 = pi0317 & n47103;
  assign n47747 = ~n47745 & ~n47746;
  assign n47748 = ~pi0591 & ~n47747;
  assign n47749 = pi0402 & ~pi0592;
  assign n47750 = n47101 & n47749;
  assign n47751 = ~n47748 & ~n47750;
  assign n47752 = ~pi0588 & ~n47751;
  assign n47753 = pi0427 & n47660;
  assign n47754 = n47661 & n47753;
  assign n47755 = ~n47752 & ~n47754;
  assign n47756 = n47050 & ~n47755;
  assign n47757 = pi0199 & ~pi1078;
  assign n47758 = ~pi0199 & n42861;
  assign n47759 = ~n47050 & ~n47757;
  assign n47760 = ~n47758 & n47759;
  assign n47761 = ~n47756 & ~n47760;
  assign n47762 = n7643 & ~n47761;
  assign n47763 = pi0844 & n47119;
  assign n47764 = ~pi0726 & pi1135;
  assign n47765 = pi0770 & ~pi1135;
  assign n47766 = pi1136 & ~n47764;
  assign n47767 = ~n47765 & n47766;
  assign n47768 = pi1134 & ~n47763;
  assign n47769 = ~n47767 & n47768;
  assign n47770 = pi0801 & n47119;
  assign n47771 = ~pi0656 & ~pi1135;
  assign n47772 = pi0649 & pi1135;
  assign n47773 = pi1136 & ~n47771;
  assign n47774 = ~n47772 & n47773;
  assign n47775 = ~pi1134 & ~n47770;
  assign n47776 = ~n47774 & n47775;
  assign n47777 = n47127 & ~n47769;
  assign n47778 = ~n47776 & n47777;
  assign po0849 = n47762 | n47778;
  assign n47780 = ~pi1129 & po0954;
  assign n47781 = pi0693 & ~po0954;
  assign n47782 = ~pi0962 & ~n47780;
  assign po0850 = ~n47781 & n47782;
  assign n47784 = ~pi1128 & po0980;
  assign n47785 = pi0694 & ~po0980;
  assign n47786 = ~pi0962 & ~n47784;
  assign po0851 = ~n47785 & n47786;
  assign n47788 = ~pi1111 & po0954;
  assign n47789 = pi0695 & ~po0954;
  assign n47790 = ~pi0962 & ~n47788;
  assign po0852 = ~n47789 & n47790;
  assign n47792 = ~pi0696 & ~po0980;
  assign n47793 = ~pi1100 & po0980;
  assign n47794 = ~pi0962 & ~n47792;
  assign po0853 = ~n47793 & n47794;
  assign n47796 = ~pi1129 & po0980;
  assign n47797 = pi0697 & ~po0980;
  assign n47798 = ~pi0962 & ~n47796;
  assign po0854 = ~n47797 & n47798;
  assign n47800 = ~pi1116 & po0980;
  assign n47801 = pi0698 & ~po0980;
  assign n47802 = ~pi0962 & ~n47800;
  assign po0855 = ~n47801 & n47802;
  assign n47804 = ~pi0699 & ~po0980;
  assign n47805 = ~pi1103 & po0980;
  assign n47806 = ~pi0962 & ~n47804;
  assign po0856 = ~n47805 & n47806;
  assign n47808 = ~pi0700 & ~po0980;
  assign n47809 = ~pi1110 & po0980;
  assign n47810 = ~pi0962 & ~n47808;
  assign po0857 = ~n47809 & n47810;
  assign n47812 = ~pi1123 & po0980;
  assign n47813 = pi0701 & ~po0980;
  assign n47814 = ~pi0962 & ~n47812;
  assign po0858 = ~n47813 & n47814;
  assign n47816 = ~pi1117 & po0980;
  assign n47817 = pi0702 & ~po0980;
  assign n47818 = ~pi0962 & ~n47816;
  assign po0859 = ~n47817 & n47818;
  assign n47820 = ~pi0703 & ~po0980;
  assign n47821 = ~pi1124 & po0980;
  assign n47822 = ~pi0962 & ~n47820;
  assign po0860 = ~n47821 & n47822;
  assign n47824 = ~pi1112 & po0980;
  assign n47825 = pi0704 & ~po0980;
  assign n47826 = ~pi0962 & ~n47824;
  assign po0861 = ~n47825 & n47826;
  assign n47828 = ~pi0705 & ~po0980;
  assign n47829 = ~pi1125 & po0980;
  assign n47830 = ~pi0962 & ~n47828;
  assign po0862 = ~n47829 & n47830;
  assign n47832 = ~pi0706 & ~po0980;
  assign n47833 = ~pi1105 & po0980;
  assign n47834 = ~pi0962 & ~n47832;
  assign po0863 = ~n47833 & n47834;
  assign n47836 = pi0370 & n47058;
  assign n47837 = pi0395 & pi0591;
  assign n47838 = ~pi0592 & n47837;
  assign n47839 = ~n47836 & ~n47838;
  assign n47840 = ~pi0590 & ~n47839;
  assign n47841 = pi0347 & n47065;
  assign n47842 = ~n47840 & ~n47841;
  assign n47843 = ~pi0588 & n47050;
  assign n47844 = ~n47842 & n47843;
  assign n47845 = pi0199 & ~pi1055;
  assign n47846 = ~pi0200 & ~pi0304;
  assign n47847 = pi0200 & ~pi1048;
  assign n47848 = ~n47846 & ~n47847;
  assign n47849 = ~pi0199 & ~n47848;
  assign n47850 = ~n47050 & ~n47845;
  assign n47851 = ~n47849 & n47850;
  assign n47852 = n47050 & n47055;
  assign n47853 = pi0420 & pi0588;
  assign n47854 = n47852 & n47853;
  assign n47855 = ~n47851 & ~n47854;
  assign n47856 = ~n47844 & n47855;
  assign n47857 = n7643 & ~n47856;
  assign n47858 = ~pi0627 & pi1135;
  assign n47859 = ~pi0618 & ~pi1135;
  assign n47860 = ~pi1134 & ~n47858;
  assign n47861 = ~n47859 & n47860;
  assign n47862 = n47283 & n47861;
  assign n47863 = pi0702 & pi1135;
  assign n47864 = ~pi0847 & ~pi1136;
  assign n47865 = pi0753 & n47086;
  assign n47866 = ~n47863 & ~n47864;
  assign n47867 = n47092 & n47866;
  assign n47868 = ~n47865 & n47867;
  assign n47869 = ~n47862 & ~n47868;
  assign n47870 = ~n7643 & ~n47869;
  assign po0864 = n47857 | n47870;
  assign n47872 = n47050 & n47660;
  assign n47873 = pi0459 & n47661;
  assign n47874 = n47872 & n47873;
  assign n47875 = n47050 & n47058;
  assign n47876 = pi0442 & n47875;
  assign n47877 = ~pi0592 & n47050;
  assign n47878 = pi0328 & pi0591;
  assign n47879 = n47877 & n47878;
  assign n47880 = ~n47876 & ~n47879;
  assign n47881 = ~pi0590 & ~n47880;
  assign n47882 = pi0321 & n47050;
  assign n47883 = n47065 & n47882;
  assign n47884 = ~n47881 & ~n47883;
  assign n47885 = ~pi0588 & ~n47884;
  assign n47886 = pi0199 & ~pi1058;
  assign n47887 = ~pi0200 & ~pi0305;
  assign n47888 = pi0200 & ~pi1084;
  assign n47889 = ~n47887 & ~n47888;
  assign n47890 = ~pi0199 & ~n47889;
  assign n47891 = ~n47050 & ~n47886;
  assign n47892 = ~n47890 & n47891;
  assign n47893 = n7643 & ~n47874;
  assign n47894 = ~n47892 & n47893;
  assign n47895 = ~n47885 & n47894;
  assign n47896 = ~pi0609 & ~pi1135;
  assign n47897 = ~pi0660 & pi1135;
  assign n47898 = ~pi1134 & ~n47896;
  assign n47899 = ~n47897 & n47898;
  assign n47900 = n47283 & n47899;
  assign n47901 = n47073 & ~n47090;
  assign n47902 = pi0709 & pi1135;
  assign n47903 = ~pi0857 & ~pi1136;
  assign n47904 = pi0754 & n47086;
  assign n47905 = pi1134 & ~n47902;
  assign n47906 = ~n47903 & n47905;
  assign n47907 = n47901 & n47906;
  assign n47908 = ~n47904 & n47907;
  assign n47909 = ~n7643 & ~n47900;
  assign n47910 = ~n47908 & n47909;
  assign po0865 = ~n47895 & ~n47910;
  assign n47912 = ~pi1118 & po0980;
  assign n47913 = pi0709 & ~po0980;
  assign n47914 = ~pi0962 & ~n47912;
  assign po0866 = ~n47913 & n47914;
  assign n47916 = ~pi0710 & ~po0954;
  assign n47917 = ~pi1106 & po0954;
  assign n47918 = ~pi0962 & ~n47916;
  assign po0867 = ~n47917 & n47918;
  assign n47920 = pi0373 & n47058;
  assign n47921 = pi0398 & pi0591;
  assign n47922 = ~pi0592 & n47921;
  assign n47923 = ~n47920 & ~n47922;
  assign n47924 = ~pi0590 & ~n47923;
  assign n47925 = pi0348 & n47065;
  assign n47926 = ~n47924 & ~n47925;
  assign n47927 = n47843 & ~n47926;
  assign n47928 = pi0199 & ~pi1087;
  assign n47929 = ~pi0200 & ~pi0306;
  assign n47930 = pi0200 & ~pi1059;
  assign n47931 = ~n47929 & ~n47930;
  assign n47932 = ~pi0199 & ~n47931;
  assign n47933 = ~n47050 & ~n47928;
  assign n47934 = ~n47932 & n47933;
  assign n47935 = pi0423 & pi0588;
  assign n47936 = n47852 & n47935;
  assign n47937 = ~n47934 & ~n47936;
  assign n47938 = ~n47927 & n47937;
  assign n47939 = n7643 & ~n47938;
  assign n47940 = ~pi0647 & pi1135;
  assign n47941 = ~pi0630 & ~pi1135;
  assign n47942 = ~pi1134 & ~n47940;
  assign n47943 = ~n47941 & n47942;
  assign n47944 = n47283 & n47943;
  assign n47945 = pi0725 & pi1135;
  assign n47946 = ~pi0858 & ~pi1136;
  assign n47947 = pi0755 & n47086;
  assign n47948 = ~n47945 & ~n47946;
  assign n47949 = n47092 & n47948;
  assign n47950 = ~n47947 & n47949;
  assign n47951 = ~n47944 & ~n47950;
  assign n47952 = ~n7643 & ~n47951;
  assign po0868 = n47939 | n47952;
  assign n47954 = pi0701 & pi1135;
  assign n47955 = ~pi0842 & ~pi1136;
  assign n47956 = pi0751 & n47086;
  assign n47957 = pi1134 & ~n47954;
  assign n47958 = ~n47955 & n47957;
  assign n47959 = n47901 & n47958;
  assign n47960 = ~n47956 & n47959;
  assign n47961 = ~pi0715 & pi1135;
  assign n47962 = ~pi0644 & ~pi1135;
  assign n47963 = ~pi1134 & ~n47961;
  assign n47964 = ~n47962 & n47963;
  assign n47965 = n47283 & n47964;
  assign n47966 = ~n47960 & ~n47965;
  assign n47967 = ~n7643 & ~n47966;
  assign n47968 = pi0199 & pi1035;
  assign n47969 = pi0298 & n10809;
  assign n47970 = pi1044 & n11444;
  assign n47971 = ~n47050 & ~n47968;
  assign n47972 = ~n47969 & n47971;
  assign n47973 = ~n47970 & n47972;
  assign n47974 = pi0425 & n47660;
  assign n47975 = n47661 & n47974;
  assign n47976 = pi0374 & n47058;
  assign n47977 = pi0400 & pi0591;
  assign n47978 = ~pi0592 & n47977;
  assign n47979 = ~n47976 & ~n47978;
  assign n47980 = ~pi0590 & ~n47979;
  assign n47981 = pi0350 & n47065;
  assign n47982 = ~n47980 & ~n47981;
  assign n47983 = ~pi0588 & ~n47982;
  assign n47984 = n47050 & ~n47975;
  assign n47985 = ~n47983 & n47984;
  assign n47986 = n7643 & ~n47973;
  assign n47987 = ~n47985 & n47986;
  assign po0869 = n47967 | n47987;
  assign n47989 = pi0371 & n47058;
  assign n47990 = pi0396 & pi0591;
  assign n47991 = ~pi0592 & n47990;
  assign n47992 = ~n47989 & ~n47991;
  assign n47993 = ~pi0590 & ~n47992;
  assign n47994 = pi0322 & n47065;
  assign n47995 = ~n47993 & ~n47994;
  assign n47996 = n47843 & ~n47995;
  assign n47997 = pi0199 & ~pi1051;
  assign n47998 = ~pi0200 & ~pi0309;
  assign n47999 = pi0200 & ~pi1072;
  assign n48000 = ~n47998 & ~n47999;
  assign n48001 = ~pi0199 & ~n48000;
  assign n48002 = ~n47050 & ~n47997;
  assign n48003 = ~n48001 & n48002;
  assign n48004 = pi0421 & pi0588;
  assign n48005 = n47852 & n48004;
  assign n48006 = ~n48003 & ~n48005;
  assign n48007 = ~n47996 & n48006;
  assign n48008 = n7643 & ~n48007;
  assign n48009 = ~pi0628 & pi1135;
  assign n48010 = ~pi0629 & ~pi1135;
  assign n48011 = ~pi1134 & ~n48009;
  assign n48012 = ~n48010 & n48011;
  assign n48013 = n47283 & n48012;
  assign n48014 = pi0734 & pi1135;
  assign n48015 = ~pi0854 & ~pi1136;
  assign n48016 = pi0756 & n47086;
  assign n48017 = ~n48014 & ~n48015;
  assign n48018 = n47092 & n48017;
  assign n48019 = ~n48016 & n48018;
  assign n48020 = ~n48013 & ~n48019;
  assign n48021 = ~n7643 & ~n48020;
  assign po0870 = n48008 | n48021;
  assign n48023 = pi0461 & n47651;
  assign n48024 = pi0439 & n47103;
  assign n48025 = ~n48023 & ~n48024;
  assign n48026 = ~pi0591 & ~n48025;
  assign n48027 = pi0326 & ~pi0592;
  assign n48028 = n47101 & n48027;
  assign n48029 = ~n48026 & ~n48028;
  assign n48030 = ~pi0588 & ~n48029;
  assign n48031 = pi0449 & n47660;
  assign n48032 = n47661 & n48031;
  assign n48033 = ~n48030 & ~n48032;
  assign n48034 = n47050 & ~n48033;
  assign n48035 = pi0199 & ~pi1057;
  assign n48036 = ~n47050 & ~n48035;
  assign n48037 = ~n42339 & n48036;
  assign n48038 = ~n48034 & ~n48037;
  assign n48039 = n7643 & ~n48038;
  assign n48040 = pi0867 & n47119;
  assign n48041 = pi0762 & ~pi1135;
  assign n48042 = pi0697 & pi1135;
  assign n48043 = pi1136 & ~n48041;
  assign n48044 = ~n48042 & n48043;
  assign n48045 = ~n48040 & ~n48044;
  assign n48046 = n47091 & ~n48045;
  assign n48047 = ~pi0653 & ~pi1135;
  assign n48048 = pi0693 & pi1135;
  assign n48049 = pi1136 & ~n48047;
  assign n48050 = ~n48048 & n48049;
  assign n48051 = pi0816 & n47073;
  assign n48052 = n47119 & n48051;
  assign n48053 = ~n48050 & ~n48052;
  assign n48054 = n47679 & ~n48053;
  assign n48055 = ~n48046 & ~n48054;
  assign n48056 = ~n7643 & ~n48055;
  assign po0871 = n48039 | n48056;
  assign n48058 = ~pi0715 & ~po0954;
  assign n48059 = ~pi1123 & po0954;
  assign n48060 = ~pi0962 & ~n48058;
  assign po0872 = ~n48059 & n48060;
  assign n48062 = pi0454 & n47661;
  assign n48063 = n47872 & n48062;
  assign n48064 = pi0440 & n47875;
  assign n48065 = pi0329 & pi0591;
  assign n48066 = n47877 & n48065;
  assign n48067 = ~n48064 & ~n48066;
  assign n48068 = ~pi0590 & ~n48067;
  assign n48069 = pi0349 & n47050;
  assign n48070 = n47065 & n48069;
  assign n48071 = ~n48068 & ~n48070;
  assign n48072 = ~pi0588 & ~n48071;
  assign n48073 = pi0199 & ~pi1043;
  assign n48074 = ~pi0200 & ~pi0307;
  assign n48075 = pi0200 & ~pi1053;
  assign n48076 = ~n48074 & ~n48075;
  assign n48077 = ~pi0199 & ~n48076;
  assign n48078 = ~n47050 & ~n48073;
  assign n48079 = ~n48077 & n48078;
  assign n48080 = n7643 & ~n48063;
  assign n48081 = ~n48079 & n48080;
  assign n48082 = ~n48072 & n48081;
  assign n48083 = ~pi0626 & ~pi1135;
  assign n48084 = ~pi0641 & pi1135;
  assign n48085 = ~pi1134 & ~n48083;
  assign n48086 = ~n48084 & n48085;
  assign n48087 = n47283 & n48086;
  assign n48088 = pi0738 & pi1135;
  assign n48089 = ~pi0845 & ~pi1136;
  assign n48090 = pi0761 & n47086;
  assign n48091 = pi1134 & ~n48088;
  assign n48092 = ~n48089 & n48091;
  assign n48093 = n47901 & n48092;
  assign n48094 = ~n48090 & n48093;
  assign n48095 = ~n7643 & ~n48087;
  assign n48096 = ~n48094 & n48095;
  assign po0873 = ~n48082 & ~n48096;
  assign n48098 = pi0318 & pi0591;
  assign n48099 = ~pi0592 & n48098;
  assign n48100 = ~pi0591 & n8468;
  assign n48101 = ~n48099 & ~n48100;
  assign n48102 = ~pi0590 & ~n48101;
  assign n48103 = pi0462 & n47065;
  assign n48104 = ~n48102 & ~n48103;
  assign n48105 = n47843 & ~n48104;
  assign n48106 = pi0199 & ~pi1074;
  assign n48107 = ~pi0199 & n42855;
  assign n48108 = ~n47050 & ~n48106;
  assign n48109 = ~n48107 & n48108;
  assign n48110 = pi0448 & pi0588;
  assign n48111 = n47852 & n48110;
  assign n48112 = ~n48109 & ~n48111;
  assign n48113 = ~n48105 & n48112;
  assign n48114 = n7643 & ~n48113;
  assign n48115 = ~pi0705 & pi1135;
  assign n48116 = pi0768 & n47086;
  assign n48117 = ~pi0839 & ~pi1136;
  assign n48118 = pi1134 & ~n48115;
  assign n48119 = ~n48117 & n48118;
  assign n48120 = n47901 & n48119;
  assign n48121 = ~n48116 & n48120;
  assign n48122 = pi0800 & n47119;
  assign n48123 = ~pi0645 & ~pi1135;
  assign n48124 = pi0669 & pi1135;
  assign n48125 = pi1136 & ~n48123;
  assign n48126 = ~n48124 & n48125;
  assign n48127 = ~n48122 & ~n48126;
  assign n48128 = n47074 & ~n48127;
  assign n48129 = ~n48121 & ~n48128;
  assign n48130 = ~n7643 & ~n48129;
  assign po0874 = n48114 | n48130;
  assign n48132 = pi0419 & n47661;
  assign n48133 = n47872 & n48132;
  assign n48134 = pi0369 & n47875;
  assign n48135 = pi0394 & pi0591;
  assign n48136 = n47877 & n48135;
  assign n48137 = ~n48134 & ~n48136;
  assign n48138 = ~pi0590 & ~n48137;
  assign n48139 = pi0315 & n47050;
  assign n48140 = n47065 & n48139;
  assign n48141 = ~n48138 & ~n48140;
  assign n48142 = ~pi0588 & ~n48141;
  assign n48143 = pi0199 & ~pi1080;
  assign n48144 = ~pi0200 & ~pi0303;
  assign n48145 = pi0200 & ~pi1049;
  assign n48146 = ~n48144 & ~n48145;
  assign n48147 = ~pi0199 & ~n48146;
  assign n48148 = ~n47050 & ~n48143;
  assign n48149 = ~n48147 & n48148;
  assign n48150 = n7643 & ~n48133;
  assign n48151 = ~n48149 & n48150;
  assign n48152 = ~n48142 & n48151;
  assign n48153 = ~pi0608 & ~pi1135;
  assign n48154 = ~pi0625 & pi1135;
  assign n48155 = ~pi1134 & ~n48153;
  assign n48156 = ~n48154 & n48155;
  assign n48157 = n47283 & n48156;
  assign n48158 = pi0698 & pi1135;
  assign n48159 = ~pi0853 & ~pi1136;
  assign n48160 = pi0767 & n47086;
  assign n48161 = pi1134 & ~n48158;
  assign n48162 = ~n48159 & n48161;
  assign n48163 = n47901 & n48162;
  assign n48164 = ~n48160 & n48163;
  assign n48165 = ~n7643 & ~n48157;
  assign n48166 = ~n48164 & n48165;
  assign po0875 = ~n48152 & ~n48166;
  assign n48168 = pi0378 & n47058;
  assign n48169 = pi0325 & pi0591;
  assign n48170 = ~pi0592 & n48169;
  assign n48171 = ~n48168 & ~n48170;
  assign n48172 = ~pi0590 & ~n48171;
  assign n48173 = pi0353 & n47065;
  assign n48174 = ~n48172 & ~n48173;
  assign n48175 = n47843 & ~n48174;
  assign n48176 = pi0199 & ~pi1063;
  assign n48177 = ~pi0199 & n42867;
  assign n48178 = ~n47050 & ~n48176;
  assign n48179 = ~n48177 & n48178;
  assign n48180 = pi0451 & pi0588;
  assign n48181 = n47852 & n48180;
  assign n48182 = ~n48179 & ~n48181;
  assign n48183 = ~n48175 & n48182;
  assign n48184 = n7643 & ~n48183;
  assign n48185 = ~pi0687 & pi1135;
  assign n48186 = pi0774 & n47086;
  assign n48187 = ~pi0868 & ~pi1136;
  assign n48188 = pi1134 & ~n48185;
  assign n48189 = ~n48187 & n48188;
  assign n48190 = n47901 & n48189;
  assign n48191 = ~n48186 & n48190;
  assign n48192 = pi0807 & n47119;
  assign n48193 = ~pi0636 & ~pi1135;
  assign n48194 = pi0650 & pi1135;
  assign n48195 = pi1136 & ~n48193;
  assign n48196 = ~n48194 & n48195;
  assign n48197 = ~n48192 & ~n48196;
  assign n48198 = n47074 & ~n48197;
  assign n48199 = ~n48191 & ~n48198;
  assign n48200 = ~n7643 & ~n48199;
  assign po0876 = n48184 | n48200;
  assign n48202 = pi0356 & n47651;
  assign n48203 = pi0381 & n47103;
  assign n48204 = ~n48202 & ~n48203;
  assign n48205 = ~pi0591 & ~n48204;
  assign n48206 = pi0405 & ~pi0592;
  assign n48207 = n47101 & n48206;
  assign n48208 = ~n48205 & ~n48207;
  assign n48209 = ~pi0588 & ~n48208;
  assign n48210 = pi0445 & n47660;
  assign n48211 = n47661 & n48210;
  assign n48212 = ~n48209 & ~n48211;
  assign n48213 = n47050 & ~n48212;
  assign n48214 = pi0199 & ~pi1081;
  assign n48215 = ~n47050 & ~n48214;
  assign n48216 = ~n42887 & n48215;
  assign n48217 = ~n48213 & ~n48216;
  assign n48218 = n7643 & ~n48217;
  assign n48219 = pi0880 & n47119;
  assign n48220 = pi0750 & ~pi1135;
  assign n48221 = pi0684 & pi1135;
  assign n48222 = pi1136 & ~n48220;
  assign n48223 = ~n48221 & n48222;
  assign n48224 = ~n48219 & ~n48223;
  assign n48225 = n47091 & ~n48224;
  assign n48226 = ~pi0651 & ~pi1135;
  assign n48227 = pi0654 & pi1135;
  assign n48228 = pi1136 & ~n48226;
  assign n48229 = ~n48227 & n48228;
  assign n48230 = pi0794 & n47073;
  assign n48231 = n47119 & n48230;
  assign n48232 = ~n48229 & ~n48231;
  assign n48233 = n47679 & ~n48232;
  assign n48234 = ~n48225 & ~n48233;
  assign n48235 = ~n7643 & ~n48234;
  assign po0877 = n48218 | n48235;
  assign n48237 = pi0721 & ~pi0775;
  assign n48238 = pi0721 & pi0813;
  assign n48239 = ~pi0773 & ~pi0801;
  assign n48240 = pi0773 & pi0801;
  assign n48241 = ~n48239 & ~n48240;
  assign n48242 = ~pi0771 & ~pi0800;
  assign n48243 = pi0771 & pi0800;
  assign n48244 = ~n48242 & ~n48243;
  assign n48245 = ~pi0769 & ~pi0794;
  assign n48246 = pi0769 & pi0794;
  assign n48247 = ~n48245 & ~n48246;
  assign n48248 = ~pi0765 & ~pi0798;
  assign n48249 = pi0765 & pi0798;
  assign n48250 = ~n48248 & ~n48249;
  assign n48251 = pi0807 & ~n48250;
  assign n48252 = pi0747 & n48251;
  assign n48253 = ~pi0747 & ~pi0807;
  assign n48254 = ~n48250 & n48253;
  assign n48255 = ~n48252 & ~n48254;
  assign n48256 = ~n48247 & ~n48255;
  assign n48257 = ~n48244 & n48256;
  assign n48258 = ~n48241 & n48257;
  assign n48259 = n48238 & n48258;
  assign n48260 = ~pi0775 & ~pi0816;
  assign n48261 = pi0775 & pi0816;
  assign n48262 = ~n48260 & ~n48261;
  assign n48263 = n48259 & ~n48262;
  assign n48264 = n48237 & ~n48263;
  assign n48265 = pi0747 & pi0773;
  assign n48266 = pi0769 & n48265;
  assign n48267 = pi0721 & n48266;
  assign n48268 = ~pi0721 & ~n48266;
  assign n48269 = pi0775 & ~n48267;
  assign n48270 = ~n48268 & n48269;
  assign n48271 = ~n48244 & n48251;
  assign n48272 = ~pi0721 & ~pi0813;
  assign n48273 = pi0794 & pi0801;
  assign n48274 = n48272 & n48273;
  assign n48275 = n48271 & n48274;
  assign n48276 = ~n48259 & ~n48275;
  assign n48277 = pi0816 & ~n48276;
  assign n48278 = n48270 & ~n48277;
  assign n48279 = pi0795 & ~n48278;
  assign n48280 = ~pi0945 & pi0988;
  assign n48281 = pi0731 & n48280;
  assign n48282 = ~n48237 & ~n48270;
  assign n48283 = n48281 & ~n48282;
  assign n48284 = ~n48279 & n48283;
  assign n48285 = ~pi0731 & ~pi0795;
  assign n48286 = pi0731 & pi0795;
  assign n48287 = ~n48285 & ~n48286;
  assign n48288 = n48263 & ~n48287;
  assign n48289 = pi0721 & ~n48281;
  assign n48290 = ~n48288 & n48289;
  assign n48291 = ~n48264 & ~n48290;
  assign po0878 = n48284 | ~n48291;
  assign n48293 = pi0379 & n47058;
  assign n48294 = pi0403 & pi0591;
  assign n48295 = ~pi0592 & n48294;
  assign n48296 = ~n48293 & ~n48295;
  assign n48297 = ~pi0590 & ~n48296;
  assign n48298 = pi0354 & n47065;
  assign n48299 = ~n48297 & ~n48298;
  assign n48300 = n47843 & ~n48299;
  assign n48301 = pi0199 & ~pi1045;
  assign n48302 = ~pi0199 & n42873;
  assign n48303 = ~n47050 & ~n48301;
  assign n48304 = ~n48302 & n48303;
  assign n48305 = pi0428 & pi0588;
  assign n48306 = n47852 & n48305;
  assign n48307 = ~n48304 & ~n48306;
  assign n48308 = ~n48300 & n48307;
  assign n48309 = n7643 & ~n48308;
  assign n48310 = ~pi0795 & ~pi1134;
  assign n48311 = ~pi0851 & pi1134;
  assign n48312 = ~pi1136 & ~n48310;
  assign n48313 = ~n48311 & n48312;
  assign n48314 = ~pi0640 & ~pi1134;
  assign n48315 = pi0776 & pi1134;
  assign n48316 = pi1136 & ~n48314;
  assign n48317 = ~n48315 & n48316;
  assign n48318 = ~n48313 & ~n48317;
  assign n48319 = ~pi1135 & ~n48318;
  assign n48320 = pi0694 & pi1134;
  assign n48321 = pi0732 & ~pi1134;
  assign n48322 = pi1135 & pi1136;
  assign n48323 = ~n48320 & n48322;
  assign n48324 = ~n48321 & n48323;
  assign n48325 = ~n48319 & ~n48324;
  assign n48326 = n47127 & ~n48325;
  assign po0879 = n48309 | n48326;
  assign n48328 = ~pi1111 & po0980;
  assign n48329 = pi0723 & ~po0980;
  assign n48330 = ~pi0962 & ~n48328;
  assign po0880 = ~n48329 & n48330;
  assign n48332 = ~pi1114 & po0980;
  assign n48333 = pi0724 & ~po0980;
  assign n48334 = ~pi0962 & ~n48332;
  assign po0881 = ~n48333 & n48334;
  assign n48336 = ~pi1120 & po0980;
  assign n48337 = pi0725 & ~po0980;
  assign n48338 = ~pi0962 & ~n48336;
  assign po0882 = ~n48337 & n48338;
  assign n48340 = ~pi0726 & ~po0980;
  assign n48341 = ~pi1126 & po0980;
  assign n48342 = ~pi0962 & ~n48340;
  assign po0883 = ~n48341 & n48342;
  assign n48344 = ~pi0727 & ~po0980;
  assign n48345 = ~pi1102 & po0980;
  assign n48346 = ~pi0962 & ~n48344;
  assign po0884 = ~n48345 & n48346;
  assign n48348 = ~pi1131 & po0980;
  assign n48349 = pi0728 & ~po0980;
  assign n48350 = ~pi0962 & ~n48348;
  assign po0885 = ~n48349 & n48350;
  assign n48352 = ~pi0729 & ~po0980;
  assign n48353 = ~pi1104 & po0980;
  assign n48354 = ~pi0962 & ~n48352;
  assign po0886 = ~n48353 & n48354;
  assign n48356 = ~pi0730 & ~po0980;
  assign n48357 = ~pi1106 & po0980;
  assign n48358 = ~pi0962 & ~n48356;
  assign po0887 = ~n48357 & n48358;
  assign n48360 = ~n48238 & ~n48272;
  assign n48361 = n48258 & ~n48360;
  assign n48362 = pi0795 & ~n48262;
  assign n48363 = n48361 & n48362;
  assign n48364 = ~n48265 & ~n48363;
  assign n48365 = n48281 & ~n48364;
  assign n48366 = pi0731 & ~n48363;
  assign n48367 = ~n48262 & ~n48360;
  assign n48368 = ~pi0795 & pi0801;
  assign n48369 = ~n48247 & n48368;
  assign n48370 = n48367 & n48369;
  assign n48371 = n48271 & n48370;
  assign n48372 = n48265 & ~n48371;
  assign n48373 = ~pi0731 & ~n48372;
  assign n48374 = n48280 & ~n48373;
  assign n48375 = ~n48366 & ~n48374;
  assign po0888 = ~n48365 & ~n48375;
  assign n48377 = ~pi1128 & po0954;
  assign n48378 = pi0732 & ~po0954;
  assign n48379 = ~pi0962 & ~n48377;
  assign po0889 = ~n48378 & n48379;
  assign n48381 = pi0424 & n47661;
  assign n48382 = n47872 & n48381;
  assign n48383 = pi0375 & n47875;
  assign n48384 = pi0399 & pi0591;
  assign n48385 = n47877 & n48384;
  assign n48386 = ~n48383 & ~n48385;
  assign n48387 = ~pi0590 & ~n48386;
  assign n48388 = pi0316 & n47050;
  assign n48389 = n47065 & n48388;
  assign n48390 = ~n48387 & ~n48389;
  assign n48391 = ~pi0588 & ~n48390;
  assign n48392 = pi0199 & ~pi1047;
  assign n48393 = ~pi0200 & ~pi0308;
  assign n48394 = pi0200 & ~pi1037;
  assign n48395 = ~n48393 & ~n48394;
  assign n48396 = ~pi0199 & ~n48395;
  assign n48397 = ~n47050 & ~n48392;
  assign n48398 = ~n48396 & n48397;
  assign n48399 = n7643 & ~n48382;
  assign n48400 = ~n48398 & n48399;
  assign n48401 = ~n48391 & n48400;
  assign n48402 = ~pi0619 & ~pi1135;
  assign n48403 = ~pi0648 & pi1135;
  assign n48404 = ~pi1134 & ~n48402;
  assign n48405 = ~n48403 & n48404;
  assign n48406 = n47283 & n48405;
  assign n48407 = pi0737 & pi1135;
  assign n48408 = ~pi0838 & ~pi1136;
  assign n48409 = pi0777 & n47086;
  assign n48410 = pi1134 & ~n48407;
  assign n48411 = ~n48408 & n48410;
  assign n48412 = n47901 & n48411;
  assign n48413 = ~n48409 & n48412;
  assign n48414 = ~n7643 & ~n48406;
  assign n48415 = ~n48413 & n48414;
  assign po0890 = ~n48401 & ~n48415;
  assign n48417 = ~pi1119 & po0980;
  assign n48418 = pi0734 & ~po0980;
  assign n48419 = ~pi0962 & ~n48417;
  assign po0891 = ~n48418 & n48419;
  assign n48421 = ~pi0735 & ~po0980;
  assign n48422 = ~pi1109 & po0980;
  assign n48423 = ~pi0962 & ~n48421;
  assign po0892 = ~n48422 & n48423;
  assign n48425 = ~pi0736 & ~po0980;
  assign n48426 = ~pi1101 & po0980;
  assign n48427 = ~pi0962 & ~n48425;
  assign po0893 = ~n48426 & n48427;
  assign n48429 = ~pi1122 & po0980;
  assign n48430 = pi0737 & ~po0980;
  assign n48431 = ~pi0962 & ~n48429;
  assign po0894 = ~n48430 & n48431;
  assign n48433 = ~pi1121 & po0980;
  assign n48434 = pi0738 & ~po0980;
  assign n48435 = ~pi0962 & ~n48433;
  assign po0895 = ~n48434 & n48435;
  assign n48437 = ~pi0952 & ~pi1061;
  assign n48438 = n46780 & n48437;
  assign po0988 = pi0832 & n48438;
  assign n48440 = pi1108 & po0988;
  assign n48441 = pi0739 & ~po0988;
  assign n48442 = ~pi0966 & ~n48440;
  assign po0896 = n48441 | ~n48442;
  assign n48444 = ~pi0741 & ~po0988;
  assign n48445 = pi1114 & po0988;
  assign n48446 = ~pi0966 & ~n48444;
  assign po0898 = n48445 | ~n48446;
  assign n48448 = ~pi0742 & ~po0988;
  assign n48449 = pi1112 & po0988;
  assign n48450 = ~pi0966 & ~n48448;
  assign po0899 = n48449 | ~n48450;
  assign n48452 = pi1109 & po0988;
  assign n48453 = pi0743 & ~po0988;
  assign n48454 = ~pi0966 & ~n48452;
  assign po0900 = n48453 | ~n48454;
  assign n48456 = ~pi0744 & ~po0988;
  assign n48457 = pi1131 & po0988;
  assign n48458 = ~pi0966 & ~n48456;
  assign po0901 = n48457 | ~n48458;
  assign n48460 = ~pi0745 & ~po0988;
  assign n48461 = pi1111 & po0988;
  assign n48462 = ~pi0966 & ~n48460;
  assign po0902 = n48461 | ~n48462;
  assign n48464 = pi1104 & po0988;
  assign n48465 = pi0746 & ~po0988;
  assign n48466 = ~pi0966 & ~n48464;
  assign po0903 = n48465 | ~n48466;
  assign n48468 = pi0773 & n48280;
  assign n48469 = ~pi0747 & ~n48468;
  assign n48470 = n48265 & n48280;
  assign n48471 = ~n48287 & n48367;
  assign n48472 = pi0801 & n48254;
  assign n48473 = ~n48241 & ~n48468;
  assign n48474 = n48251 & n48473;
  assign n48475 = ~n48472 & ~n48474;
  assign n48476 = ~n48244 & ~n48247;
  assign n48477 = n48471 & n48476;
  assign n48478 = ~n48475 & n48477;
  assign n48479 = ~n48469 & ~n48470;
  assign po0904 = ~n48478 & n48479;
  assign n48481 = pi1106 & po0988;
  assign n48482 = pi0748 & ~po0988;
  assign n48483 = ~pi0966 & ~n48481;
  assign po0905 = n48482 | ~n48483;
  assign n48485 = pi1105 & po0988;
  assign n48486 = pi0749 & ~po0988;
  assign n48487 = ~pi0966 & ~n48485;
  assign po0906 = n48486 | ~n48487;
  assign n48489 = ~pi0750 & ~po0988;
  assign n48490 = pi1130 & po0988;
  assign n48491 = ~pi0966 & ~n48489;
  assign po0907 = n48490 | ~n48491;
  assign n48493 = ~pi0751 & ~po0988;
  assign n48494 = pi1123 & po0988;
  assign n48495 = ~pi0966 & ~n48493;
  assign po0908 = n48494 | ~n48495;
  assign n48497 = ~pi0752 & ~po0988;
  assign n48498 = pi1124 & po0988;
  assign n48499 = ~pi0966 & ~n48497;
  assign po0909 = n48498 | ~n48499;
  assign n48501 = ~pi0753 & ~po0988;
  assign n48502 = pi1117 & po0988;
  assign n48503 = ~pi0966 & ~n48501;
  assign po0910 = n48502 | ~n48503;
  assign n48505 = ~pi0754 & ~po0988;
  assign n48506 = pi1118 & po0988;
  assign n48507 = ~pi0966 & ~n48505;
  assign po0911 = n48506 | ~n48507;
  assign n48509 = ~pi0755 & ~po0988;
  assign n48510 = pi1120 & po0988;
  assign n48511 = ~pi0966 & ~n48509;
  assign po0912 = n48510 | ~n48511;
  assign n48513 = ~pi0756 & ~po0988;
  assign n48514 = pi1119 & po0988;
  assign n48515 = ~pi0966 & ~n48513;
  assign po0913 = n48514 | ~n48515;
  assign n48517 = ~pi0757 & ~po0988;
  assign n48518 = pi1113 & po0988;
  assign n48519 = ~pi0966 & ~n48517;
  assign po0914 = n48518 | ~n48519;
  assign n48521 = pi1101 & po0988;
  assign n48522 = pi0758 & ~po0988;
  assign n48523 = ~pi0966 & ~n48521;
  assign po0915 = n48522 | ~n48523;
  assign n48525 = ~pi0759 & ~po0988;
  assign n48526 = n46778 & n48438;
  assign n48527 = ~n48525 & ~n48526;
  assign po0916 = pi0966 | n48527;
  assign n48529 = ~pi0760 & ~po0988;
  assign n48530 = pi1115 & po0988;
  assign n48531 = ~pi0966 & ~n48529;
  assign po0917 = n48530 | ~n48531;
  assign n48533 = ~pi0761 & ~po0988;
  assign n48534 = pi1121 & po0988;
  assign n48535 = ~pi0966 & ~n48533;
  assign po0918 = n48534 | ~n48535;
  assign n48537 = ~pi0762 & ~po0988;
  assign n48538 = pi1129 & po0988;
  assign n48539 = ~pi0966 & ~n48537;
  assign po0919 = n48538 | ~n48539;
  assign n48541 = pi1103 & po0988;
  assign n48542 = pi0763 & ~po0988;
  assign n48543 = ~pi0966 & ~n48541;
  assign po0920 = n48542 | ~n48543;
  assign n48545 = pi1107 & po0988;
  assign n48546 = pi0764 & ~po0988;
  assign n48547 = ~pi0966 & ~n48545;
  assign po0921 = n48546 | ~n48547;
  assign po0978 = n48258 & n48471;
  assign n48550 = pi0765 & ~po0978;
  assign n48551 = pi0945 & ~n48550;
  assign n48552 = ~n48259 & ~n48272;
  assign n48553 = ~pi0765 & ~n48243;
  assign n48554 = ~n48246 & n48553;
  assign n48555 = ~n48252 & n48554;
  assign n48556 = n48239 & ~n48555;
  assign n48557 = ~n48240 & ~n48556;
  assign n48558 = n48257 & ~n48557;
  assign n48559 = ~pi0721 & ~n48558;
  assign n48560 = n48260 & ~n48559;
  assign n48561 = ~n48552 & n48560;
  assign n48562 = n48261 & n48361;
  assign n48563 = ~pi0765 & ~n48562;
  assign n48564 = ~n48561 & n48563;
  assign n48565 = ~pi0795 & ~n48564;
  assign n48566 = ~pi0731 & ~n48565;
  assign n48567 = ~pi0795 & n48566;
  assign n48568 = pi0765 & ~n48567;
  assign n48569 = ~n48366 & ~n48566;
  assign n48570 = ~n48568 & ~n48569;
  assign n48571 = ~pi0945 & ~n48570;
  assign po0922 = ~n48551 & ~n48571;
  assign n48573 = pi1110 & po0988;
  assign n48574 = pi0766 & ~po0988;
  assign n48575 = ~pi0966 & ~n48573;
  assign po0923 = n48574 | ~n48575;
  assign n48577 = ~pi0767 & ~po0988;
  assign n48578 = pi1116 & po0988;
  assign n48579 = ~pi0966 & ~n48577;
  assign po0924 = n48578 | ~n48579;
  assign n48581 = ~pi0768 & ~po0988;
  assign n48582 = pi1125 & po0988;
  assign n48583 = ~pi0966 & ~n48581;
  assign po0925 = n48582 | ~n48583;
  assign n48585 = pi0794 & ~n48241;
  assign n48586 = ~n48244 & n48585;
  assign n48587 = n48367 & n48586;
  assign n48588 = ~n48255 & n48587;
  assign n48589 = ~pi0775 & n48588;
  assign n48590 = ~n48562 & ~n48589;
  assign n48591 = pi0795 & ~n48590;
  assign n48592 = pi0775 & n48265;
  assign n48593 = pi0769 & ~n48592;
  assign n48594 = ~pi0769 & n48592;
  assign n48595 = ~n48593 & ~n48594;
  assign n48596 = n48281 & ~n48595;
  assign n48597 = ~n48591 & n48596;
  assign n48598 = ~n48287 & n48588;
  assign n48599 = pi0769 & ~n48281;
  assign n48600 = ~n48598 & n48599;
  assign po0926 = n48597 | n48600;
  assign n48602 = ~pi0770 & ~po0988;
  assign n48603 = pi1126 & po0988;
  assign n48604 = ~pi0966 & ~n48602;
  assign po0927 = n48603 | ~n48604;
  assign n48606 = ~n48261 & ~n48560;
  assign n48607 = n48285 & ~n48606;
  assign n48608 = ~n48262 & n48286;
  assign n48609 = ~n48607 & ~n48608;
  assign po0963 = n48361 & ~n48609;
  assign n48611 = ~pi0945 & pi0987;
  assign n48612 = ~po0963 & n48611;
  assign n48613 = pi0771 & pi0945;
  assign n48614 = ~po0978 & n48613;
  assign po0928 = n48612 | n48614;
  assign n48616 = pi1102 & po0988;
  assign n48617 = pi0772 & ~po0988;
  assign n48618 = ~pi0966 & ~n48616;
  assign po0929 = n48617 | ~n48618;
  assign n48620 = ~pi0801 & n48257;
  assign n48621 = po0963 & n48620;
  assign n48622 = n48280 & ~n48621;
  assign n48623 = pi0801 & ~n48471;
  assign n48624 = n48258 & ~n48623;
  assign n48625 = pi0773 & ~n48624;
  assign n48626 = ~n48622 & ~n48625;
  assign po0930 = ~n48468 & ~n48626;
  assign n48628 = ~pi0774 & ~po0988;
  assign n48629 = pi1127 & po0988;
  assign n48630 = ~pi0966 & ~n48628;
  assign po0931 = n48629 | ~n48630;
  assign n48632 = pi0775 & ~po0978;
  assign n48633 = pi0731 & ~pi0945;
  assign n48634 = pi0765 & pi0771;
  assign n48635 = n48265 & n48634;
  assign n48636 = pi0795 & pi0800;
  assign n48637 = pi0801 & ~pi0816;
  assign n48638 = n48636 & n48637;
  assign n48639 = ~n48360 & n48638;
  assign n48640 = n48256 & n48639;
  assign n48641 = n48635 & ~n48640;
  assign n48642 = ~pi0775 & ~n48641;
  assign n48643 = n48633 & ~n48642;
  assign n48644 = ~n48632 & ~n48643;
  assign n48645 = ~n48363 & ~n48635;
  assign n48646 = pi0775 & n48633;
  assign n48647 = ~n48645 & n48646;
  assign po0932 = ~n48644 & ~n48647;
  assign n48649 = ~pi0776 & ~po0988;
  assign n48650 = pi1128 & po0988;
  assign n48651 = ~pi0966 & ~n48649;
  assign po0933 = n48650 | ~n48651;
  assign n48653 = ~pi0777 & ~po0988;
  assign n48654 = pi1122 & po0988;
  assign n48655 = ~pi0966 & ~n48653;
  assign po0934 = n48654 | ~n48655;
  assign n48657 = pi0832 & pi0956;
  assign n48658 = ~pi1046 & ~pi1083;
  assign n48659 = pi1085 & n48658;
  assign n48660 = n48657 & n48659;
  assign n48661 = ~pi0968 & n48660;
  assign n48662 = pi0778 & ~n48661;
  assign n48663 = pi1100 & n48661;
  assign po0935 = n48662 | n48663;
  assign po0936 = ~pi0779 | n46839;
  assign po0937 = ~pi0780 | n46748;
  assign n48667 = pi0781 & ~n48661;
  assign n48668 = pi1101 & n48661;
  assign po0938 = n48667 | n48668;
  assign n48670 = ~n42345 & ~n46792;
  assign po0939 = n46747 | ~n48670;
  assign n48672 = pi0783 & ~n48661;
  assign n48673 = pi1109 & n48661;
  assign po0940 = n48672 | n48673;
  assign n48675 = pi0784 & ~n48661;
  assign n48676 = pi1110 & n48661;
  assign po0941 = n48675 | n48676;
  assign n48678 = pi0785 & ~n48661;
  assign n48679 = pi1102 & n48661;
  assign po0942 = n48678 | n48679;
  assign n48681 = pi0024 & ~pi0954;
  assign n48682 = pi0786 & pi0954;
  assign po0943 = ~n48681 & ~n48682;
  assign n48684 = pi0787 & ~n48661;
  assign n48685 = pi1104 & n48661;
  assign po0944 = n48684 | n48685;
  assign n48687 = pi0788 & ~n48661;
  assign n48688 = pi1105 & n48661;
  assign po0945 = n48687 | n48688;
  assign n48690 = pi0789 & ~n48661;
  assign n48691 = pi1106 & n48661;
  assign po0946 = n48690 | n48691;
  assign n48693 = pi0790 & ~n48661;
  assign n48694 = pi1107 & n48661;
  assign po0947 = n48693 | n48694;
  assign n48696 = pi0791 & ~n48661;
  assign n48697 = pi1108 & n48661;
  assign po0948 = n48696 | n48697;
  assign n48699 = pi0792 & ~n48661;
  assign n48700 = pi1103 & n48661;
  assign po0949 = n48699 | n48700;
  assign n48702 = pi0968 & n48660;
  assign n48703 = pi0794 & ~n48702;
  assign n48704 = pi1130 & n48702;
  assign po0951 = n48703 | n48704;
  assign n48706 = pi0795 & ~n48702;
  assign n48707 = pi1128 & n48702;
  assign po0952 = n48706 | n48707;
  assign n48709 = pi0266 & ~pi0269;
  assign n48710 = pi0278 & pi0279;
  assign n48711 = ~pi0280 & n48710;
  assign n48712 = n48709 & n48711;
  assign n48713 = ~pi0281 & n48712;
  assign n48714 = n47031 & n48713;
  assign n48715 = pi0264 & ~n48714;
  assign n48716 = ~pi0264 & n48714;
  assign po0953 = ~n48715 & ~n48716;
  assign n48718 = pi0798 & ~n48702;
  assign n48719 = pi1124 & n48702;
  assign po0955 = n48718 | n48719;
  assign n48721 = pi0799 & ~n48702;
  assign n48722 = ~pi1107 & n48702;
  assign po0956 = ~n48721 & ~n48722;
  assign n48724 = pi0800 & ~n48702;
  assign n48725 = pi1125 & n48702;
  assign po0957 = n48724 | n48725;
  assign n48727 = pi0801 & ~n48702;
  assign n48728 = pi1126 & n48702;
  assign po0958 = n48727 | n48728;
  assign n48730 = pi0803 & ~n48702;
  assign n48731 = ~pi1106 & n48702;
  assign po0960 = ~n48730 & ~n48731;
  assign n48733 = pi0804 & ~n48702;
  assign n48734 = pi1109 & n48702;
  assign po0961 = n48733 | n48734;
  assign n48736 = ~pi0282 & n47029;
  assign n48737 = ~pi0270 & n48736;
  assign n48738 = pi0270 & ~n48736;
  assign po0962 = ~n48737 & ~n48738;
  assign n48740 = pi0807 & ~n48702;
  assign n48741 = pi1127 & n48702;
  assign po0964 = n48740 | n48741;
  assign n48743 = pi0808 & ~n48702;
  assign n48744 = pi1101 & n48702;
  assign po0965 = n48743 | n48744;
  assign n48746 = pi0809 & ~n48702;
  assign n48747 = ~pi1103 & n48702;
  assign po0966 = ~n48746 & ~n48747;
  assign n48749 = pi0810 & ~n48702;
  assign n48750 = pi1108 & n48702;
  assign po0967 = n48749 | n48750;
  assign n48752 = pi0811 & ~n48702;
  assign n48753 = pi1102 & n48702;
  assign po0968 = n48752 | n48753;
  assign n48755 = pi0812 & ~n48702;
  assign n48756 = ~pi1104 & n48702;
  assign po0969 = ~n48755 & ~n48756;
  assign n48758 = pi0813 & ~n48702;
  assign n48759 = pi1131 & n48702;
  assign po0970 = n48758 | n48759;
  assign n48761 = pi0814 & ~n48702;
  assign n48762 = ~pi1105 & n48702;
  assign po0971 = ~n48761 & ~n48762;
  assign n48764 = pi0815 & ~n48702;
  assign n48765 = pi1110 & n48702;
  assign po0972 = n48764 | n48765;
  assign n48767 = pi0816 & ~n48702;
  assign n48768 = pi1129 & n48702;
  assign po0973 = n48767 | n48768;
  assign n48770 = pi0269 & ~n47027;
  assign po0974 = ~n47028 & ~n48770;
  assign n48772 = n7643 & n14172;
  assign po0975 = n14025 | n48772;
  assign n48774 = pi0265 & ~n47033;
  assign po0976 = ~n47034 & ~n48774;
  assign n48776 = pi0277 & ~n48737;
  assign po0977 = ~n47032 & ~n48776;
  assign po0979 = ~pi0811 & ~pi0893;
  assign n48779 = ~pi0982 & ~n10074;
  assign n48780 = n7626 & n7643;
  assign n48781 = ~n48779 & ~n48780;
  assign po0981 = n2932 & ~n48781;
  assign n48783 = pi0123 & n2604;
  assign n48784 = pi1131 & ~n48783;
  assign n48785 = pi1127 & ~n48783;
  assign n48786 = ~n48784 & ~n48785;
  assign n48787 = ~pi0825 & n48783;
  assign n48788 = n48786 & ~n48787;
  assign n48789 = pi1131 & n48785;
  assign n48790 = ~n48788 & ~n48789;
  assign n48791 = pi1124 & ~pi1130;
  assign n48792 = ~pi1124 & pi1130;
  assign n48793 = ~n48791 & ~n48792;
  assign n48794 = ~pi1128 & ~pi1129;
  assign n48795 = pi1128 & pi1129;
  assign n48796 = ~n48794 & ~n48795;
  assign n48797 = ~pi1125 & ~pi1126;
  assign n48798 = pi1125 & pi1126;
  assign n48799 = ~n48797 & ~n48798;
  assign n48800 = n48796 & ~n48799;
  assign n48801 = ~n48796 & n48799;
  assign n48802 = ~n48800 & ~n48801;
  assign n48803 = n48793 & n48802;
  assign n48804 = ~n48793 & ~n48802;
  assign n48805 = ~n48803 & ~n48804;
  assign n48806 = ~n48790 & ~n48805;
  assign n48807 = pi0825 & n48783;
  assign n48808 = n48786 & ~n48807;
  assign n48809 = ~n48789 & n48805;
  assign n48810 = ~n48808 & n48809;
  assign po0982 = ~n48806 & ~n48810;
  assign n48812 = pi1123 & ~n48783;
  assign n48813 = pi1122 & ~n48783;
  assign n48814 = ~n48812 & ~n48813;
  assign n48815 = ~pi0826 & n48783;
  assign n48816 = n48814 & ~n48815;
  assign n48817 = pi1123 & n48813;
  assign n48818 = ~n48816 & ~n48817;
  assign n48819 = pi1118 & ~pi1119;
  assign n48820 = ~pi1118 & pi1119;
  assign n48821 = ~n48819 & ~n48820;
  assign n48822 = ~pi1120 & ~pi1121;
  assign n48823 = pi1120 & pi1121;
  assign n48824 = ~n48822 & ~n48823;
  assign n48825 = ~pi1116 & ~pi1117;
  assign n48826 = pi1116 & pi1117;
  assign n48827 = ~n48825 & ~n48826;
  assign n48828 = n48824 & ~n48827;
  assign n48829 = ~n48824 & n48827;
  assign n48830 = ~n48828 & ~n48829;
  assign n48831 = n48821 & n48830;
  assign n48832 = ~n48821 & ~n48830;
  assign n48833 = ~n48831 & ~n48832;
  assign n48834 = ~n48818 & ~n48833;
  assign n48835 = pi0826 & n48783;
  assign n48836 = n48814 & ~n48835;
  assign n48837 = ~n48817 & n48833;
  assign n48838 = ~n48836 & n48837;
  assign po0983 = ~n48834 & ~n48838;
  assign n48840 = pi1100 & ~n48783;
  assign n48841 = pi1107 & ~n48783;
  assign n48842 = ~n48840 & ~n48841;
  assign n48843 = ~pi0827 & n48783;
  assign n48844 = n48842 & ~n48843;
  assign n48845 = pi1100 & n48841;
  assign n48846 = ~n48844 & ~n48845;
  assign n48847 = pi1103 & ~pi1105;
  assign n48848 = ~pi1103 & pi1105;
  assign n48849 = ~n48847 & ~n48848;
  assign n48850 = ~pi1101 & ~pi1102;
  assign n48851 = pi1101 & pi1102;
  assign n48852 = ~n48850 & ~n48851;
  assign n48853 = ~pi1104 & ~pi1106;
  assign n48854 = pi1104 & pi1106;
  assign n48855 = ~n48853 & ~n48854;
  assign n48856 = n48852 & ~n48855;
  assign n48857 = ~n48852 & n48855;
  assign n48858 = ~n48856 & ~n48857;
  assign n48859 = n48849 & n48858;
  assign n48860 = ~n48849 & ~n48858;
  assign n48861 = ~n48859 & ~n48860;
  assign n48862 = ~n48846 & ~n48861;
  assign n48863 = pi0827 & n48783;
  assign n48864 = n48842 & ~n48863;
  assign n48865 = ~n48845 & n48861;
  assign n48866 = ~n48864 & n48865;
  assign po0984 = ~n48862 & ~n48866;
  assign n48868 = pi1115 & ~n48783;
  assign n48869 = pi1114 & ~n48783;
  assign n48870 = ~n48868 & ~n48869;
  assign n48871 = ~pi0828 & n48783;
  assign n48872 = n48870 & ~n48871;
  assign n48873 = pi1115 & n48869;
  assign n48874 = ~n48872 & ~n48873;
  assign n48875 = pi1110 & ~pi1111;
  assign n48876 = ~pi1110 & pi1111;
  assign n48877 = ~n48875 & ~n48876;
  assign n48878 = ~pi1112 & ~pi1113;
  assign n48879 = pi1112 & pi1113;
  assign n48880 = ~n48878 & ~n48879;
  assign n48881 = ~pi1108 & ~pi1109;
  assign n48882 = pi1108 & pi1109;
  assign n48883 = ~n48881 & ~n48882;
  assign n48884 = n48880 & ~n48883;
  assign n48885 = ~n48880 & n48883;
  assign n48886 = ~n48884 & ~n48885;
  assign n48887 = n48877 & n48886;
  assign n48888 = ~n48877 & ~n48886;
  assign n48889 = ~n48887 & ~n48888;
  assign n48890 = ~n48874 & ~n48889;
  assign n48891 = pi0828 & n48783;
  assign n48892 = n48870 & ~n48891;
  assign n48893 = ~n48873 & n48889;
  assign n48894 = ~n48892 & n48893;
  assign po0985 = ~n48890 & ~n48894;
  assign n48896 = n2930 & n7643;
  assign n48897 = pi0951 & ~n48896;
  assign po0986 = pi1092 & ~n48897;
  assign n48899 = pi0281 & ~n48712;
  assign po0987 = ~n48713 & ~n48899;
  assign n48901 = ~pi0832 & pi1091;
  assign n48902 = pi1162 & n48901;
  assign po0989 = n8874 & n48902;
  assign n48904 = pi0833 & ~n2926;
  assign po0990 = n16887 | n48904;
  assign po0991 = pi0946 & n2926;
  assign n48907 = pi0282 & ~n47029;
  assign po0992 = ~n48736 & ~n48907;
  assign n48909 = ~pi0955 & pi1049;
  assign n48910 = pi0837 & pi0955;
  assign po0993 = n48909 | n48910;
  assign n48912 = ~pi0955 & pi1047;
  assign n48913 = pi0838 & pi0955;
  assign po0994 = n48912 | n48913;
  assign n48915 = ~pi0955 & pi1074;
  assign n48916 = pi0839 & pi0955;
  assign po0995 = n48915 | n48916;
  assign n48918 = pi0840 & ~n2926;
  assign n48919 = pi1196 & n2926;
  assign po0996 = n48918 | n48919;
  assign po0997 = ~pi0033 & n8979;
  assign n48922 = ~pi0955 & pi1035;
  assign n48923 = pi0842 & pi0955;
  assign po0998 = n48922 | n48923;
  assign n48925 = ~pi0955 & pi1079;
  assign n48926 = pi0843 & pi0955;
  assign po0999 = n48925 | n48926;
  assign n48928 = ~pi0955 & pi1078;
  assign n48929 = pi0844 & pi0955;
  assign po1000 = n48928 | n48929;
  assign n48931 = ~pi0955 & pi1043;
  assign n48932 = pi0845 & pi0955;
  assign po1001 = n48931 | n48932;
  assign n48934 = pi0846 & ~n42902;
  assign n48935 = pi1134 & n42902;
  assign po1002 = n48934 | n48935;
  assign n48937 = ~pi0955 & pi1055;
  assign n48938 = pi0847 & pi0955;
  assign po1003 = n48937 | n48938;
  assign n48940 = ~pi0955 & pi1039;
  assign n48941 = pi0848 & pi0955;
  assign po1004 = n48940 | n48941;
  assign n48943 = pi0849 & ~n2926;
  assign n48944 = pi1198 & n2926;
  assign po1005 = n48943 | n48944;
  assign n48946 = ~pi0955 & pi1048;
  assign n48947 = pi0850 & pi0955;
  assign po1006 = n48946 | n48947;
  assign n48949 = ~pi0955 & pi1045;
  assign n48950 = pi0851 & pi0955;
  assign po1007 = n48949 | n48950;
  assign n48952 = ~pi0955 & pi1062;
  assign n48953 = pi0852 & pi0955;
  assign po1008 = n48952 | n48953;
  assign n48955 = ~pi0955 & pi1080;
  assign n48956 = pi0853 & pi0955;
  assign po1009 = n48955 | n48956;
  assign n48958 = ~pi0955 & pi1051;
  assign n48959 = pi0854 & pi0955;
  assign po1010 = n48958 | n48959;
  assign n48961 = ~pi0955 & pi1065;
  assign n48962 = pi0855 & pi0955;
  assign po1011 = n48961 | n48962;
  assign n48964 = ~pi0955 & pi1067;
  assign n48965 = pi0856 & pi0955;
  assign po1012 = n48964 | n48965;
  assign n48967 = ~pi0955 & pi1058;
  assign n48968 = pi0857 & pi0955;
  assign po1013 = n48967 | n48968;
  assign n48970 = ~pi0955 & pi1087;
  assign n48971 = pi0858 & pi0955;
  assign po1014 = n48970 | n48971;
  assign n48973 = ~pi0955 & pi1070;
  assign n48974 = pi0859 & pi0955;
  assign po1015 = n48973 | n48974;
  assign n48976 = ~pi0955 & pi1076;
  assign n48977 = pi0860 & pi0955;
  assign po1016 = n48976 | n48977;
  assign n48979 = pi1093 & pi1141;
  assign n48980 = pi0861 & ~pi1093;
  assign n48981 = ~n48979 & ~n48980;
  assign n48982 = ~pi0228 & ~n48981;
  assign n48983 = ~pi0123 & ~pi1141;
  assign n48984 = pi0123 & ~pi0861;
  assign n48985 = pi0228 & ~n48983;
  assign n48986 = ~n48984 & n48985;
  assign po1017 = n48982 | n48986;
  assign n48988 = pi0862 & ~n42902;
  assign n48989 = pi1139 & n42902;
  assign po1018 = n48988 | n48989;
  assign n48991 = pi0863 & ~n2926;
  assign n48992 = pi1199 & n2926;
  assign po1019 = n48991 | n48992;
  assign n48994 = pi0864 & ~n2926;
  assign n48995 = pi1197 & n2926;
  assign po1020 = n48994 | n48995;
  assign n48997 = ~pi0955 & pi1040;
  assign n48998 = pi0865 & pi0955;
  assign po1021 = n48997 | n48998;
  assign n49000 = ~pi0955 & pi1053;
  assign n49001 = pi0866 & pi0955;
  assign po1022 = n49000 | n49001;
  assign n49003 = ~pi0955 & pi1057;
  assign n49004 = pi0867 & pi0955;
  assign po1023 = n49003 | n49004;
  assign n49006 = ~pi0955 & pi1063;
  assign n49007 = pi0868 & pi0955;
  assign po1024 = n49006 | n49007;
  assign n49009 = pi1093 & pi1140;
  assign n49010 = pi0869 & ~pi1093;
  assign n49011 = ~n49009 & ~n49010;
  assign n49012 = ~pi0228 & ~n49011;
  assign n49013 = ~pi0123 & ~pi1140;
  assign n49014 = pi0123 & ~pi0869;
  assign n49015 = pi0228 & ~n49013;
  assign n49016 = ~n49014 & n49015;
  assign po1025 = n49012 | n49016;
  assign n49018 = ~pi0955 & pi1069;
  assign n49019 = pi0870 & pi0955;
  assign po1026 = n49018 | n49019;
  assign n49021 = ~pi0955 & pi1072;
  assign n49022 = pi0871 & pi0955;
  assign po1027 = n49021 | n49022;
  assign n49024 = ~pi0955 & pi1084;
  assign n49025 = pi0872 & pi0955;
  assign po1028 = n49024 | n49025;
  assign n49027 = ~pi0955 & pi1044;
  assign n49028 = pi0873 & pi0955;
  assign po1029 = n49027 | n49028;
  assign n49030 = ~pi0955 & pi1036;
  assign n49031 = pi0874 & pi0955;
  assign po1030 = n49030 | n49031;
  assign n49033 = pi1093 & ~pi1136;
  assign n49034 = ~pi0875 & ~pi1093;
  assign n49035 = ~n49033 & ~n49034;
  assign n49036 = ~pi0228 & ~n49035;
  assign n49037 = ~pi0123 & pi1136;
  assign n49038 = pi0123 & pi0875;
  assign n49039 = pi0228 & ~n49037;
  assign n49040 = ~n49038 & n49039;
  assign po1031 = ~n49036 & ~n49040;
  assign n49042 = ~pi0955 & pi1037;
  assign n49043 = pi0876 & pi0955;
  assign po1032 = n49042 | n49043;
  assign n49045 = pi1093 & pi1138;
  assign n49046 = pi0877 & ~pi1093;
  assign n49047 = ~n49045 & ~n49046;
  assign n49048 = ~pi0228 & ~n49047;
  assign n49049 = ~pi0123 & ~pi1138;
  assign n49050 = pi0123 & ~pi0877;
  assign n49051 = pi0228 & ~n49049;
  assign n49052 = ~n49050 & n49051;
  assign po1033 = n49048 | n49052;
  assign n49054 = pi1093 & pi1137;
  assign n49055 = pi0878 & ~pi1093;
  assign n49056 = ~n49054 & ~n49055;
  assign n49057 = ~pi0228 & ~n49056;
  assign n49058 = ~pi0123 & ~pi1137;
  assign n49059 = pi0123 & ~pi0878;
  assign n49060 = pi0228 & ~n49058;
  assign n49061 = ~n49059 & n49060;
  assign po1034 = n49057 | n49061;
  assign n49063 = pi1093 & pi1135;
  assign n49064 = pi0879 & ~pi1093;
  assign n49065 = ~n49063 & ~n49064;
  assign n49066 = ~pi0228 & ~n49065;
  assign n49067 = ~pi0123 & ~pi1135;
  assign n49068 = pi0123 & ~pi0879;
  assign n49069 = pi0228 & ~n49067;
  assign n49070 = ~n49068 & n49069;
  assign po1035 = n49066 | n49070;
  assign n49072 = ~pi0955 & pi1081;
  assign n49073 = pi0880 & pi0955;
  assign po1036 = n49072 | n49073;
  assign n49075 = ~pi0955 & pi1059;
  assign n49076 = pi0881 & pi0955;
  assign po1037 = n49075 | n49076;
  assign n49078 = ~pi0883 & n48783;
  assign po1039 = n48841 | n49078;
  assign n49080 = pi1124 & ~n48783;
  assign n49081 = ~pi0884 & n48783;
  assign po1040 = n49080 | n49081;
  assign n49083 = pi1125 & ~n48783;
  assign n49084 = ~pi0885 & n48783;
  assign po1041 = n49083 | n49084;
  assign n49086 = pi1109 & ~n48783;
  assign n49087 = ~pi0886 & n48783;
  assign po1042 = n49086 | n49087;
  assign n49089 = ~pi0887 & n48783;
  assign po1043 = n48840 | n49089;
  assign n49091 = pi1120 & ~n48783;
  assign n49092 = ~pi0888 & n48783;
  assign po1044 = n49091 | n49092;
  assign n49094 = pi1103 & ~n48783;
  assign n49095 = ~pi0889 & n48783;
  assign po1045 = n49094 | n49095;
  assign n49097 = pi1126 & ~n48783;
  assign n49098 = ~pi0890 & n48783;
  assign po1046 = n49097 | n49098;
  assign n49100 = pi1116 & ~n48783;
  assign n49101 = ~pi0891 & n48783;
  assign po1047 = n49100 | n49101;
  assign n49103 = pi1101 & ~n48783;
  assign n49104 = ~pi0892 & n48783;
  assign po1048 = n49103 | n49104;
  assign n49106 = pi1119 & ~n48783;
  assign n49107 = ~pi0894 & n48783;
  assign po1050 = n49106 | n49107;
  assign n49109 = pi1113 & ~n48783;
  assign n49110 = ~pi0895 & n48783;
  assign po1051 = n49109 | n49110;
  assign n49112 = pi1118 & ~n48783;
  assign n49113 = ~pi0896 & n48783;
  assign po1052 = n49112 | n49113;
  assign n49115 = pi1129 & ~n48783;
  assign n49116 = ~pi0898 & n48783;
  assign po1054 = n49115 | n49116;
  assign n49118 = ~pi0899 & n48783;
  assign po1055 = n48868 | n49118;
  assign n49120 = pi1110 & ~n48783;
  assign n49121 = ~pi0900 & n48783;
  assign po1056 = n49120 | n49121;
  assign n49123 = pi1111 & ~n48783;
  assign n49124 = ~pi0902 & n48783;
  assign po1058 = n49123 | n49124;
  assign n49126 = pi1121 & ~n48783;
  assign n49127 = ~pi0903 & n48783;
  assign po1059 = n49126 | n49127;
  assign n49129 = ~pi0904 & n48783;
  assign po1060 = n48785 | n49129;
  assign n49131 = ~pi0905 & n48783;
  assign po1061 = n48784 | n49131;
  assign n49133 = pi1128 & ~n48783;
  assign n49134 = ~pi0906 & n48783;
  assign po1062 = n49133 | n49134;
  assign n49136 = ~pi0782 & ~pi0907;
  assign n49137 = ~pi0624 & ~pi0979;
  assign n49138 = ~pi0598 & pi0979;
  assign n49139 = pi0782 & ~n49137;
  assign n49140 = ~n49138 & n49139;
  assign n49141 = ~pi0604 & ~pi0979;
  assign n49142 = pi0615 & pi0979;
  assign n49143 = ~n49141 & ~n49142;
  assign n49144 = pi0782 & ~n49143;
  assign n49145 = ~n49136 & ~n49140;
  assign po1063 = ~n49144 & n49145;
  assign n49147 = ~pi0908 & n48783;
  assign po1064 = n48813 | n49147;
  assign n49149 = pi1105 & ~n48783;
  assign n49150 = ~pi0909 & n48783;
  assign po1065 = n49149 | n49150;
  assign n49152 = pi1117 & ~n48783;
  assign n49153 = ~pi0910 & n48783;
  assign po1066 = n49152 | n49153;
  assign n49155 = pi1130 & ~n48783;
  assign n49156 = ~pi0911 & n48783;
  assign po1067 = n49155 | n49156;
  assign n49158 = ~pi0912 & n48783;
  assign po1068 = n48869 | n49158;
  assign n49160 = pi1106 & ~n48783;
  assign n49161 = ~pi0913 & n48783;
  assign po1069 = n49160 | n49161;
  assign n49163 = pi0280 & ~n47026;
  assign po1070 = ~n47027 & ~n49163;
  assign n49165 = pi1108 & ~n48783;
  assign n49166 = ~pi0915 & n48783;
  assign po1071 = n49165 | n49166;
  assign n49168 = ~pi0916 & n48783;
  assign po1072 = n48812 | n49168;
  assign n49170 = pi1112 & ~n48783;
  assign n49171 = ~pi0917 & n48783;
  assign po1073 = n49170 | n49171;
  assign n49173 = pi1104 & ~n48783;
  assign n49174 = ~pi0918 & n48783;
  assign po1074 = n49173 | n49174;
  assign n49176 = pi1102 & ~n48783;
  assign n49177 = ~pi0919 & n48783;
  assign po1075 = n49176 | n49177;
  assign n49179 = pi1093 & pi1139;
  assign n49180 = pi0920 & ~pi1093;
  assign po1076 = n49179 | n49180;
  assign n49182 = pi0921 & ~pi1093;
  assign po1077 = n49009 | n49182;
  assign n49184 = ~pi0922 & ~pi1093;
  assign n49185 = pi1093 & ~pi1152;
  assign po1078 = ~n49184 & ~n49185;
  assign n49187 = ~pi0923 & ~pi1093;
  assign n49188 = pi1093 & ~pi1154;
  assign po1079 = ~n49187 & ~n49188;
  assign n49190 = ~pi0300 & pi0301;
  assign n49191 = pi0311 & ~pi0312;
  assign po1080 = n49190 & n49191;
  assign n49193 = ~pi0925 & ~pi1093;
  assign n49194 = pi1093 & ~pi1155;
  assign po1081 = ~n49193 & ~n49194;
  assign n49196 = ~pi0926 & ~pi1093;
  assign n49197 = pi1093 & ~pi1157;
  assign po1082 = ~n49196 & ~n49197;
  assign n49199 = ~pi0927 & ~pi1093;
  assign n49200 = pi1093 & ~pi1145;
  assign po1083 = ~n49199 & ~n49200;
  assign n49202 = ~pi0928 & ~pi1093;
  assign po1084 = ~n49033 & ~n49202;
  assign n49204 = ~pi0929 & ~pi1093;
  assign n49205 = pi1093 & ~pi1144;
  assign po1085 = ~n49204 & ~n49205;
  assign n49207 = ~pi0930 & ~pi1093;
  assign n49208 = pi1093 & ~pi1134;
  assign po1086 = ~n49207 & ~n49208;
  assign n49210 = ~pi0931 & ~pi1093;
  assign n49211 = pi1093 & ~pi1150;
  assign po1087 = ~n49210 & ~n49211;
  assign n49213 = pi0932 & ~pi1093;
  assign po1088 = n42891 | n49213;
  assign n49215 = pi0933 & ~pi1093;
  assign po1089 = n49054 | n49215;
  assign n49217 = ~pi0934 & ~pi1093;
  assign n49218 = pi1093 & ~pi1147;
  assign po1090 = ~n49217 & ~n49218;
  assign n49220 = pi0935 & ~pi1093;
  assign po1091 = n48979 | n49220;
  assign n49222 = ~pi0936 & ~pi1093;
  assign n49223 = pi1093 & ~pi1149;
  assign po1092 = ~n49222 & ~n49223;
  assign n49225 = ~pi0937 & ~pi1093;
  assign n49226 = pi1093 & ~pi1148;
  assign po1093 = ~n49225 & ~n49226;
  assign n49228 = pi0938 & ~pi1093;
  assign po1094 = n49063 | n49228;
  assign n49230 = ~pi0939 & ~pi1093;
  assign n49231 = pi1093 & ~pi1146;
  assign po1095 = ~n49230 & ~n49231;
  assign n49233 = pi0940 & ~pi1093;
  assign po1096 = n49045 | n49233;
  assign n49235 = ~pi0941 & ~pi1093;
  assign n49236 = pi1093 & ~pi1153;
  assign po1097 = ~n49235 & ~n49236;
  assign n49238 = ~pi0942 & ~pi1093;
  assign n49239 = pi1093 & ~pi1156;
  assign po1098 = ~n49238 & ~n49239;
  assign n49241 = ~pi0943 & ~pi1093;
  assign n49242 = pi1093 & ~pi1151;
  assign po1099 = ~n49241 & ~n49242;
  assign n49244 = pi1093 & pi1143;
  assign n49245 = pi0944 & ~pi1093;
  assign po1100 = n49244 | n49245;
  assign po1102 = pi0230 & n2926;
  assign n49248 = ~pi0782 & pi0947;
  assign po1103 = n49140 | n49248;
  assign n49250 = ~pi0266 & ~pi0992;
  assign po1104 = ~n47026 & ~n49250;
  assign n49252 = ~pi0313 & ~pi0954;
  assign n49253 = pi0949 & pi0954;
  assign po1105 = n49252 | n49253;
  assign po1107 = ~n7626 & n14271;
  assign n49256 = pi0957 & pi1092;
  assign po1112 = pi0031 | n49256;
  assign po1115 = ~pi0782 & pi0960;
  assign po1116 = ~pi0230 & pi0961;
  assign po1118 = ~pi0782 & pi0963;
  assign po1122 = ~pi0230 & pi0967;
  assign po1124 = ~pi0230 & pi0969;
  assign po1125 = ~pi0782 & pi0970;
  assign po1126 = ~pi0230 & pi0971;
  assign po1127 = ~pi0782 & pi0972;
  assign po1128 = ~pi0230 & pi0974;
  assign po1129 = ~pi0782 & pi0975;
  assign po1131 = ~pi0230 & pi0977;
  assign po1132 = ~pi0782 & pi0978;
  assign po1133 = pi0598 | ~pi0615;
  assign po1135 = pi0824 & pi1092;
  assign po1137 = pi0604 | pi0624;
  assign po0166 = 1'b1;
  assign po0170 = ~pi1090;
  assign po1110 = ~pi0954;
  assign po1130 = ~pi0278;
  assign po1146 = ~pi0915;
  assign po1147 = ~pi0825;
  assign po1148 = ~pi0826;
  assign po1149 = ~pi0913;
  assign po1150 = ~pi0894;
  assign po1151 = ~pi0905;
  assign po1153 = ~pi0890;
  assign po1155 = ~pi0906;
  assign po1156 = ~pi0896;
  assign po1157 = ~pi0909;
  assign po1158 = ~pi0911;
  assign po1159 = ~pi0908;
  assign po1160 = ~pi0891;
  assign po1161 = ~pi0902;
  assign po1162 = ~pi0903;
  assign po1163 = ~pi0883;
  assign po1164 = ~pi0888;
  assign po1165 = ~pi0919;
  assign po1166 = ~pi0886;
  assign po1167 = ~pi0912;
  assign po1168 = ~pi0895;
  assign po1169 = ~pi0916;
  assign po1170 = ~pi0889;
  assign po1171 = ~pi0900;
  assign po1172 = ~pi0885;
  assign po1173 = ~pi0904;
  assign po1174 = ~pi0899;
  assign po1175 = ~pi0918;
  assign po1176 = ~pi0898;
  assign po1177 = ~pi0917;
  assign po1178 = ~pi0827;
  assign po1179 = ~pi0887;
  assign po1180 = ~pi0884;
  assign po1181 = ~pi0910;
  assign po1182 = ~pi0828;
  assign po1183 = ~pi0892;
  assign po0000 = pi0668;
  assign po0001 = pi0672;
  assign po0002 = pi0664;
  assign po0003 = pi0667;
  assign po0004 = pi0676;
  assign po0005 = pi0673;
  assign po0006 = pi0675;
  assign po0007 = pi0666;
  assign po0008 = pi0679;
  assign po0009 = pi0674;
  assign po0010 = pi0663;
  assign po0011 = pi0670;
  assign po0012 = pi0677;
  assign po0013 = pi0682;
  assign po0014 = pi0671;
  assign po0015 = pi0678;
  assign po0016 = pi0718;
  assign po0017 = pi0707;
  assign po0018 = pi0708;
  assign po0019 = pi0713;
  assign po0020 = pi0711;
  assign po0021 = pi0716;
  assign po0022 = pi0733;
  assign po0023 = pi0712;
  assign po0024 = pi0689;
  assign po0025 = pi0717;
  assign po0026 = pi0692;
  assign po0027 = pi0719;
  assign po0028 = pi0722;
  assign po0029 = pi0714;
  assign po0030 = pi0720;
  assign po0031 = pi0685;
  assign po0032 = pi0837;
  assign po0033 = pi0850;
  assign po0034 = pi0872;
  assign po0035 = pi0871;
  assign po0036 = pi0881;
  assign po0037 = pi0866;
  assign po0038 = pi0876;
  assign po0039 = pi0873;
  assign po0040 = pi0874;
  assign po0041 = pi0859;
  assign po0042 = pi0855;
  assign po0043 = pi0852;
  assign po0044 = pi0870;
  assign po0045 = pi0848;
  assign po0046 = pi0865;
  assign po0047 = pi0856;
  assign po0048 = pi0853;
  assign po0049 = pi0847;
  assign po0050 = pi0857;
  assign po0051 = pi0854;
  assign po0052 = pi0858;
  assign po0053 = pi0845;
  assign po0054 = pi0838;
  assign po0055 = pi0842;
  assign po0056 = pi0843;
  assign po0057 = pi0839;
  assign po0058 = pi0844;
  assign po0059 = pi0868;
  assign po0060 = pi0851;
  assign po0061 = pi0867;
  assign po0062 = pi0880;
  assign po0063 = pi0860;
  assign po0064 = pi1030;
  assign po0065 = pi1034;
  assign po0066 = pi1015;
  assign po0067 = pi1020;
  assign po0068 = pi1025;
  assign po0069 = pi1005;
  assign po0070 = pi0996;
  assign po0071 = pi1012;
  assign po0072 = pi0993;
  assign po0073 = pi1016;
  assign po0074 = pi1021;
  assign po0075 = pi1010;
  assign po0076 = pi1027;
  assign po0077 = pi1018;
  assign po0078 = pi1017;
  assign po0079 = pi1024;
  assign po0080 = pi1009;
  assign po0081 = pi1032;
  assign po0082 = pi1003;
  assign po0083 = pi0997;
  assign po0084 = pi1013;
  assign po0085 = pi1011;
  assign po0086 = pi1008;
  assign po0087 = pi1019;
  assign po0088 = pi1031;
  assign po0089 = pi1022;
  assign po0090 = pi1000;
  assign po0091 = pi1023;
  assign po0092 = pi1002;
  assign po0093 = pi1026;
  assign po0094 = pi1006;
  assign po0095 = pi0998;
  assign po0096 = pi0031;
  assign po0097 = pi0080;
  assign po0098 = pi0893;
  assign po0099 = pi0467;
  assign po0100 = pi0078;
  assign po0101 = pi0112;
  assign po0102 = pi0013;
  assign po0103 = pi0025;
  assign po0104 = pi0226;
  assign po0105 = pi0127;
  assign po0106 = pi0822;
  assign po0107 = pi0808;
  assign po0108 = pi0227;
  assign po0109 = pi0477;
  assign po0110 = pi0834;
  assign po0111 = pi0229;
  assign po0112 = pi0012;
  assign po0113 = pi0011;
  assign po0114 = pi0010;
  assign po0115 = pi0009;
  assign po0116 = pi0008;
  assign po0117 = pi0007;
  assign po0118 = pi0006;
  assign po0119 = pi0005;
  assign po0120 = pi0004;
  assign po0121 = pi0003;
  assign po0122 = pi0000;
  assign po0123 = pi0002;
  assign po0124 = pi0001;
  assign po0125 = pi0310;
  assign po0126 = pi0302;
  assign po0127 = pi0475;
  assign po0128 = pi0474;
  assign po0129 = pi0466;
  assign po0130 = pi0473;
  assign po0131 = pi0471;
  assign po0132 = pi0472;
  assign po0133 = pi0470;
  assign po0134 = pi0469;
  assign po0135 = pi0465;
  assign po0136 = pi1028;
  assign po0137 = pi1033;
  assign po0138 = pi0995;
  assign po0139 = pi0994;
  assign po0140 = pi0028;
  assign po0141 = pi0027;
  assign po0142 = pi0026;
  assign po0143 = pi0029;
  assign po0144 = pi0015;
  assign po0145 = pi0014;
  assign po0146 = pi0021;
  assign po0147 = pi0020;
  assign po0148 = pi0019;
  assign po0149 = pi0018;
  assign po0150 = pi0017;
  assign po0151 = pi0016;
  assign po0152 = pi1096;
  assign po0168 = pi0228;
  assign po0169 = pi0022;
  assign po0179 = pi1089;
  assign po0180 = pi0023;
  assign po0181 = po0167;
  assign po0188 = pi0037;
  assign po0263 = pi0117;
  assign po0285 = pi0131;
  assign po0386 = pi0232;
  assign po0388 = pi0236;
  assign po0636 = pi0583;
  assign po1053 = pi0067;
  assign po1108 = pi1134;
  assign po1109 = pi0964;
  assign po1111 = pi0965;
  assign po1113 = pi0991;
  assign po1114 = pi0985;
  assign po1117 = pi1014;
  assign po1119 = pi1029;
  assign po1120 = pi1004;
  assign po1121 = pi1007;
  assign po1123 = pi1135;
  assign po1134 = pi1064;
  assign po1136 = pi0299;
  assign po1138 = pi1075;
  assign po1139 = pi1052;
  assign po1140 = pi0771;
  assign po1141 = pi0765;
  assign po1142 = pi0605;
  assign po1143 = pi0601;
  assign po1144 = pi0278;
  assign po1145 = pi0279;
  assign po1152 = pi1095;
  assign po1154 = pi1094;
  assign po1184 = pi1187;
  assign po1185 = pi1172;
  assign po1186 = pi1170;
  assign po1187 = pi1138;
  assign po1188 = pi1177;
  assign po1189 = pi1178;
  assign po1190 = pi0863;
  assign po1191 = pi1203;
  assign po1192 = pi1185;
  assign po1193 = pi1171;
  assign po1194 = pi1192;
  assign po1195 = pi1137;
  assign po1196 = pi1186;
  assign po1197 = pi1165;
  assign po1198 = pi1164;
  assign po1199 = pi1098;
  assign po1200 = pi1183;
  assign po1201 = pi0230;
  assign po1202 = pi1169;
  assign po1203 = pi1136;
  assign po1204 = pi1181;
  assign po1205 = pi0849;
  assign po1206 = pi1193;
  assign po1207 = pi1182;
  assign po1208 = pi1168;
  assign po1209 = pi1175;
  assign po1210 = pi1191;
  assign po1211 = pi1099;
  assign po1212 = pi1174;
  assign po1213 = pi1179;
  assign po1214 = pi1202;
  assign po1215 = pi1176;
  assign po1216 = pi1173;
  assign po1217 = pi1201;
  assign po1218 = pi1167;
  assign po1219 = pi0840;
  assign po1220 = pi1189;
  assign po1221 = pi1195;
  assign po1222 = pi0864;
  assign po1223 = pi1190;
  assign po1224 = pi1188;
  assign po1225 = pi1180;
  assign po1226 = pi1194;
  assign po1227 = pi1097;
  assign po1228 = pi1166;
  assign po1229 = pi1200;
  assign po1230 = pi1184;
endmodule


