module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] , \shift[2] ,
    \shift[3] , \shift[4] , \shift[5] , \shift[6] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] ,
    \shift[2] , \shift[3] , \shift[4] , \shift[5] , \shift[6] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ;
  wire n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
    n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
    n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
    n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
    n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
    n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
    n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
    n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
    n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
    n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
    n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
    n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
    n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
    n695, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
    n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
    n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
    n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
    n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
    n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
    n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
    n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
    n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
    n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
    n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
    n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
    n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
    n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
    n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
    n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
    n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
    n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
    n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
    n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
    n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
    n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
    n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
    n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
    n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1789,
    n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
    n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
    n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
    n1860, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
    n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
    n1931, n1932, n1933, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
    n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
    n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
    n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
    n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2008, n2009, n2010, n2011, n2012,
    n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
    n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
    n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
    n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
    n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
    n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
    n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
    n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
    n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
    n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
    n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2154,
    n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
    n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
    n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
    n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
    n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
    n2225, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
    n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
    n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
    n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
    n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
    n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
    n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
    n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2373, n2374, n2375, n2376, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
    n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
    n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
    n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
    n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2519,
    n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
    n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
    n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
    n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
    n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2609, n2610, n2611,
    n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
    n2622, n2623, n2624, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
    n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
    n2654, n2655, n2656, n2657, n2658, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
    n2675, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
    n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2728,
    n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
    n2760, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
    n2792, n2793, n2794, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2813,
    n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2830, n2831, n2832, n2833, n2834,
    n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
    n2845, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
    n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2864, n2865, n2866,
    n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
    n2877, n2878, n2879, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
    n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
    n2909, n2910, n2911, n2912, n2913, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2949, n2950, n2951,
    n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
    n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2983,
    n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
    n2994, n2995, n2996, n2997, n2998, n3000, n3001, n3002, n3003, n3004,
    n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
    n3015, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3034, n3035, n3036,
    n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
    n3047, n3048, n3049, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3068,
    n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3085, n3086, n3087, n3088, n3089,
    n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
    n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3119, n3120, n3121,
    n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
    n3132, n3133, n3134, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
    n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
    n3164, n3165, n3166, n3167, n3168, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
    n3185, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3204, n3205, n3206,
    n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
    n3217, n3218, n3219, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
    n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3238,
    n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
    n3270, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
    n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3289, n3290, n3291,
    n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
    n3302, n3303, n3304, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
    n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3323,
    n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
    n3334, n3335, n3336, n3337, n3338, n3340, n3341, n3342, n3343, n3344,
    n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
    n3355, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
    n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3374, n3375, n3376,
    n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
    n3387, n3388, n3389, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3408,
    n3409, n3411, n3412, n3414, n3415, n3417, n3418, n3420, n3421, n3423,
    n3424, n3426, n3427, n3429, n3430, n3432, n3433, n3435, n3436, n3438,
    n3439, n3441, n3442, n3444, n3445, n3447, n3448, n3450, n3451, n3453,
    n3454, n3456, n3457, n3459, n3460, n3462, n3463, n3465, n3466, n3468,
    n3469, n3471, n3472, n3474, n3475, n3477, n3478, n3480, n3481, n3483,
    n3484, n3486, n3487, n3489, n3490, n3492, n3493, n3495, n3496, n3498,
    n3499, n3501, n3502, n3504, n3505, n3507, n3508, n3510, n3511, n3513,
    n3514, n3516, n3517, n3519, n3520, n3522, n3523, n3525, n3526, n3528,
    n3529, n3531, n3532, n3534, n3535, n3537, n3538, n3540, n3541, n3543,
    n3544, n3546, n3547, n3549, n3550, n3552, n3553, n3555, n3556, n3558,
    n3559, n3561, n3562, n3564, n3565, n3567, n3568, n3570, n3571, n3573,
    n3574, n3576, n3577, n3579, n3580, n3582, n3583, n3585, n3586, n3588,
    n3589, n3591, n3592, n3594, n3595, n3597, n3598;
  assign n264 = \a[77]  & \shift[0] ;
  assign n265 = \shift[1]  & n264;
  assign n266 = \a[78]  & ~\shift[0] ;
  assign n267 = \shift[1]  & n266;
  assign n268 = ~n265 & ~n267;
  assign n269 = \a[80]  & ~\shift[0] ;
  assign n270 = ~\shift[1]  & n269;
  assign n271 = \a[79]  & \shift[0] ;
  assign n272 = ~\shift[1]  & n271;
  assign n273 = ~n270 & ~n272;
  assign n274 = n268 & n273;
  assign n275 = ~\shift[2]  & ~\shift[3] ;
  assign n276 = ~n274 & n275;
  assign n277 = \a[73]  & \shift[0] ;
  assign n278 = \shift[1]  & n277;
  assign n279 = \a[74]  & ~\shift[0] ;
  assign n280 = \shift[1]  & n279;
  assign n281 = ~n278 & ~n280;
  assign n282 = \a[76]  & ~\shift[0] ;
  assign n283 = ~\shift[1]  & n282;
  assign n284 = \a[75]  & \shift[0] ;
  assign n285 = ~\shift[1]  & n284;
  assign n286 = ~n283 & ~n285;
  assign n287 = n281 & n286;
  assign n288 = \shift[2]  & ~\shift[3] ;
  assign n289 = ~n287 & n288;
  assign n290 = ~n276 & ~n289;
  assign n291 = \a[65]  & \shift[0] ;
  assign n292 = \shift[1]  & n291;
  assign n293 = \a[66]  & ~\shift[0] ;
  assign n294 = \shift[1]  & n293;
  assign n295 = ~n292 & ~n294;
  assign n296 = \a[68]  & ~\shift[0] ;
  assign n297 = ~\shift[1]  & n296;
  assign n298 = \a[67]  & \shift[0] ;
  assign n299 = ~\shift[1]  & n298;
  assign n300 = ~n297 & ~n299;
  assign n301 = n295 & n300;
  assign n302 = \shift[2]  & \shift[3] ;
  assign n303 = ~n301 & n302;
  assign n304 = \a[69]  & \shift[0] ;
  assign n305 = \shift[1]  & n304;
  assign n306 = \a[70]  & ~\shift[0] ;
  assign n307 = \shift[1]  & n306;
  assign n308 = ~n305 & ~n307;
  assign n309 = \a[72]  & ~\shift[0] ;
  assign n310 = ~\shift[1]  & n309;
  assign n311 = \a[71]  & \shift[0] ;
  assign n312 = ~\shift[1]  & n311;
  assign n313 = ~n310 & ~n312;
  assign n314 = n308 & n313;
  assign n315 = ~\shift[2]  & \shift[3] ;
  assign n316 = ~n314 & n315;
  assign n317 = ~n303 & ~n316;
  assign n318 = n290 & n317;
  assign n319 = \shift[4]  & \shift[5] ;
  assign n320 = ~n318 & n319;
  assign n321 = \a[93]  & \shift[0] ;
  assign n322 = \shift[1]  & n321;
  assign n323 = \a[94]  & ~\shift[0] ;
  assign n324 = \shift[1]  & n323;
  assign n325 = ~n322 & ~n324;
  assign n326 = \a[96]  & ~\shift[0] ;
  assign n327 = ~\shift[1]  & n326;
  assign n328 = \a[95]  & \shift[0] ;
  assign n329 = ~\shift[1]  & n328;
  assign n330 = ~n327 & ~n329;
  assign n331 = n325 & n330;
  assign n332 = n275 & ~n331;
  assign n333 = \a[89]  & \shift[0] ;
  assign n334 = \shift[1]  & n333;
  assign n335 = \a[90]  & ~\shift[0] ;
  assign n336 = \shift[1]  & n335;
  assign n337 = ~n334 & ~n336;
  assign n338 = \a[92]  & ~\shift[0] ;
  assign n339 = ~\shift[1]  & n338;
  assign n340 = \a[91]  & \shift[0] ;
  assign n341 = ~\shift[1]  & n340;
  assign n342 = ~n339 & ~n341;
  assign n343 = n337 & n342;
  assign n344 = n288 & ~n343;
  assign n345 = ~n332 & ~n344;
  assign n346 = \a[81]  & \shift[0] ;
  assign n347 = \shift[1]  & n346;
  assign n348 = \a[82]  & ~\shift[0] ;
  assign n349 = \shift[1]  & n348;
  assign n350 = ~n347 & ~n349;
  assign n351 = \a[84]  & ~\shift[0] ;
  assign n352 = ~\shift[1]  & n351;
  assign n353 = \a[83]  & \shift[0] ;
  assign n354 = ~\shift[1]  & n353;
  assign n355 = ~n352 & ~n354;
  assign n356 = n350 & n355;
  assign n357 = n302 & ~n356;
  assign n358 = \a[85]  & \shift[0] ;
  assign n359 = \shift[1]  & n358;
  assign n360 = \a[86]  & ~\shift[0] ;
  assign n361 = \shift[1]  & n360;
  assign n362 = ~n359 & ~n361;
  assign n363 = \a[88]  & ~\shift[0] ;
  assign n364 = ~\shift[1]  & n363;
  assign n365 = \a[87]  & \shift[0] ;
  assign n366 = ~\shift[1]  & n365;
  assign n367 = ~n364 & ~n366;
  assign n368 = n362 & n367;
  assign n369 = n315 & ~n368;
  assign n370 = ~n357 & ~n369;
  assign n371 = n345 & n370;
  assign n372 = ~\shift[4]  & \shift[5] ;
  assign n373 = ~n371 & n372;
  assign n374 = ~n320 & ~n373;
  assign n375 = \a[125]  & \shift[0] ;
  assign n376 = \shift[1]  & n375;
  assign n377 = \a[126]  & ~\shift[0] ;
  assign n378 = \shift[1]  & n377;
  assign n379 = ~n376 & ~n378;
  assign n380 = \a[0]  & ~\shift[0] ;
  assign n381 = ~\shift[1]  & n380;
  assign n382 = \a[127]  & \shift[0] ;
  assign n383 = ~\shift[1]  & n382;
  assign n384 = ~n381 & ~n383;
  assign n385 = n379 & n384;
  assign n386 = n275 & ~n385;
  assign n387 = \a[121]  & \shift[0] ;
  assign n388 = \shift[1]  & n387;
  assign n389 = \a[122]  & ~\shift[0] ;
  assign n390 = \shift[1]  & n389;
  assign n391 = ~n388 & ~n390;
  assign n392 = \a[124]  & ~\shift[0] ;
  assign n393 = ~\shift[1]  & n392;
  assign n394 = \a[123]  & \shift[0] ;
  assign n395 = ~\shift[1]  & n394;
  assign n396 = ~n393 & ~n395;
  assign n397 = n391 & n396;
  assign n398 = n288 & ~n397;
  assign n399 = ~n386 & ~n398;
  assign n400 = \a[113]  & \shift[0] ;
  assign n401 = \shift[1]  & n400;
  assign n402 = \a[114]  & ~\shift[0] ;
  assign n403 = \shift[1]  & n402;
  assign n404 = ~n401 & ~n403;
  assign n405 = \a[116]  & ~\shift[0] ;
  assign n406 = ~\shift[1]  & n405;
  assign n407 = \a[115]  & \shift[0] ;
  assign n408 = ~\shift[1]  & n407;
  assign n409 = ~n406 & ~n408;
  assign n410 = n404 & n409;
  assign n411 = n302 & ~n410;
  assign n412 = \a[117]  & \shift[0] ;
  assign n413 = \shift[1]  & n412;
  assign n414 = \a[118]  & ~\shift[0] ;
  assign n415 = \shift[1]  & n414;
  assign n416 = ~n413 & ~n415;
  assign n417 = \a[120]  & ~\shift[0] ;
  assign n418 = ~\shift[1]  & n417;
  assign n419 = \a[119]  & \shift[0] ;
  assign n420 = ~\shift[1]  & n419;
  assign n421 = ~n418 & ~n420;
  assign n422 = n416 & n421;
  assign n423 = n315 & ~n422;
  assign n424 = ~n411 & ~n423;
  assign n425 = n399 & n424;
  assign n426 = ~\shift[4]  & ~\shift[5] ;
  assign n427 = ~n425 & n426;
  assign n428 = \a[109]  & \shift[0] ;
  assign n429 = \shift[1]  & n428;
  assign n430 = \a[110]  & ~\shift[0] ;
  assign n431 = \shift[1]  & n430;
  assign n432 = ~n429 & ~n431;
  assign n433 = \a[112]  & ~\shift[0] ;
  assign n434 = ~\shift[1]  & n433;
  assign n435 = \a[111]  & \shift[0] ;
  assign n436 = ~\shift[1]  & n435;
  assign n437 = ~n434 & ~n436;
  assign n438 = n432 & n437;
  assign n439 = n275 & ~n438;
  assign n440 = \a[105]  & \shift[0] ;
  assign n441 = \shift[1]  & n440;
  assign n442 = \a[106]  & ~\shift[0] ;
  assign n443 = \shift[1]  & n442;
  assign n444 = ~n441 & ~n443;
  assign n445 = \a[108]  & ~\shift[0] ;
  assign n446 = ~\shift[1]  & n445;
  assign n447 = \a[107]  & \shift[0] ;
  assign n448 = ~\shift[1]  & n447;
  assign n449 = ~n446 & ~n448;
  assign n450 = n444 & n449;
  assign n451 = n288 & ~n450;
  assign n452 = ~n439 & ~n451;
  assign n453 = \a[97]  & \shift[0] ;
  assign n454 = \shift[1]  & n453;
  assign n455 = \a[98]  & ~\shift[0] ;
  assign n456 = \shift[1]  & n455;
  assign n457 = ~n454 & ~n456;
  assign n458 = \a[100]  & ~\shift[0] ;
  assign n459 = ~\shift[1]  & n458;
  assign n460 = \a[99]  & \shift[0] ;
  assign n461 = ~\shift[1]  & n460;
  assign n462 = ~n459 & ~n461;
  assign n463 = n457 & n462;
  assign n464 = n302 & ~n463;
  assign n465 = \a[101]  & \shift[0] ;
  assign n466 = \shift[1]  & n465;
  assign n467 = \a[102]  & ~\shift[0] ;
  assign n468 = \shift[1]  & n467;
  assign n469 = ~n466 & ~n468;
  assign n470 = \a[104]  & ~\shift[0] ;
  assign n471 = ~\shift[1]  & n470;
  assign n472 = \a[103]  & \shift[0] ;
  assign n473 = ~\shift[1]  & n472;
  assign n474 = ~n471 & ~n473;
  assign n475 = n469 & n474;
  assign n476 = n315 & ~n475;
  assign n477 = ~n464 & ~n476;
  assign n478 = n452 & n477;
  assign n479 = \shift[4]  & ~\shift[5] ;
  assign n480 = ~n478 & n479;
  assign n481 = ~n427 & ~n480;
  assign n482 = n374 & n481;
  assign n483 = ~\shift[6]  & ~n482;
  assign n484 = \a[13]  & \shift[0] ;
  assign n485 = \shift[1]  & n484;
  assign n486 = \a[14]  & ~\shift[0] ;
  assign n487 = \shift[1]  & n486;
  assign n488 = ~n485 & ~n487;
  assign n489 = \a[16]  & ~\shift[0] ;
  assign n490 = ~\shift[1]  & n489;
  assign n491 = \a[15]  & \shift[0] ;
  assign n492 = ~\shift[1]  & n491;
  assign n493 = ~n490 & ~n492;
  assign n494 = n488 & n493;
  assign n495 = n275 & ~n494;
  assign n496 = \a[9]  & \shift[0] ;
  assign n497 = \shift[1]  & n496;
  assign n498 = \a[10]  & ~\shift[0] ;
  assign n499 = \shift[1]  & n498;
  assign n500 = ~n497 & ~n499;
  assign n501 = \a[12]  & ~\shift[0] ;
  assign n502 = ~\shift[1]  & n501;
  assign n503 = \a[11]  & \shift[0] ;
  assign n504 = ~\shift[1]  & n503;
  assign n505 = ~n502 & ~n504;
  assign n506 = n500 & n505;
  assign n507 = n288 & ~n506;
  assign n508 = ~n495 & ~n507;
  assign n509 = \a[1]  & \shift[0] ;
  assign n510 = \shift[1]  & n509;
  assign n511 = \a[2]  & ~\shift[0] ;
  assign n512 = \shift[1]  & n511;
  assign n513 = ~n510 & ~n512;
  assign n514 = \a[4]  & ~\shift[0] ;
  assign n515 = ~\shift[1]  & n514;
  assign n516 = \a[3]  & \shift[0] ;
  assign n517 = ~\shift[1]  & n516;
  assign n518 = ~n515 & ~n517;
  assign n519 = n513 & n518;
  assign n520 = n302 & ~n519;
  assign n521 = \a[5]  & \shift[0] ;
  assign n522 = \shift[1]  & n521;
  assign n523 = \a[6]  & ~\shift[0] ;
  assign n524 = \shift[1]  & n523;
  assign n525 = ~n522 & ~n524;
  assign n526 = \a[8]  & ~\shift[0] ;
  assign n527 = ~\shift[1]  & n526;
  assign n528 = \a[7]  & \shift[0] ;
  assign n529 = ~\shift[1]  & n528;
  assign n530 = ~n527 & ~n529;
  assign n531 = n525 & n530;
  assign n532 = n315 & ~n531;
  assign n533 = ~n520 & ~n532;
  assign n534 = n508 & n533;
  assign n535 = n319 & ~n534;
  assign n536 = \a[29]  & \shift[0] ;
  assign n537 = \shift[1]  & n536;
  assign n538 = \a[30]  & ~\shift[0] ;
  assign n539 = \shift[1]  & n538;
  assign n540 = ~n537 & ~n539;
  assign n541 = \a[32]  & ~\shift[0] ;
  assign n542 = ~\shift[1]  & n541;
  assign n543 = \a[31]  & \shift[0] ;
  assign n544 = ~\shift[1]  & n543;
  assign n545 = ~n542 & ~n544;
  assign n546 = n540 & n545;
  assign n547 = n275 & ~n546;
  assign n548 = \a[25]  & \shift[0] ;
  assign n549 = \shift[1]  & n548;
  assign n550 = \a[26]  & ~\shift[0] ;
  assign n551 = \shift[1]  & n550;
  assign n552 = ~n549 & ~n551;
  assign n553 = \a[28]  & ~\shift[0] ;
  assign n554 = ~\shift[1]  & n553;
  assign n555 = \a[27]  & \shift[0] ;
  assign n556 = ~\shift[1]  & n555;
  assign n557 = ~n554 & ~n556;
  assign n558 = n552 & n557;
  assign n559 = n288 & ~n558;
  assign n560 = ~n547 & ~n559;
  assign n561 = \a[17]  & \shift[0] ;
  assign n562 = \shift[1]  & n561;
  assign n563 = \a[18]  & ~\shift[0] ;
  assign n564 = \shift[1]  & n563;
  assign n565 = ~n562 & ~n564;
  assign n566 = \a[20]  & ~\shift[0] ;
  assign n567 = ~\shift[1]  & n566;
  assign n568 = \a[19]  & \shift[0] ;
  assign n569 = ~\shift[1]  & n568;
  assign n570 = ~n567 & ~n569;
  assign n571 = n565 & n570;
  assign n572 = n302 & ~n571;
  assign n573 = \a[21]  & \shift[0] ;
  assign n574 = \shift[1]  & n573;
  assign n575 = \a[22]  & ~\shift[0] ;
  assign n576 = \shift[1]  & n575;
  assign n577 = ~n574 & ~n576;
  assign n578 = \a[24]  & ~\shift[0] ;
  assign n579 = ~\shift[1]  & n578;
  assign n580 = \a[23]  & \shift[0] ;
  assign n581 = ~\shift[1]  & n580;
  assign n582 = ~n579 & ~n581;
  assign n583 = n577 & n582;
  assign n584 = n315 & ~n583;
  assign n585 = ~n572 & ~n584;
  assign n586 = n560 & n585;
  assign n587 = n372 & ~n586;
  assign n588 = ~n535 & ~n587;
  assign n589 = \a[61]  & \shift[0] ;
  assign n590 = \shift[1]  & n589;
  assign n591 = \a[62]  & ~\shift[0] ;
  assign n592 = \shift[1]  & n591;
  assign n593 = ~n590 & ~n592;
  assign n594 = \a[64]  & ~\shift[0] ;
  assign n595 = ~\shift[1]  & n594;
  assign n596 = \a[63]  & \shift[0] ;
  assign n597 = ~\shift[1]  & n596;
  assign n598 = ~n595 & ~n597;
  assign n599 = n593 & n598;
  assign n600 = n275 & ~n599;
  assign n601 = \a[57]  & \shift[0] ;
  assign n602 = \shift[1]  & n601;
  assign n603 = \a[58]  & ~\shift[0] ;
  assign n604 = \shift[1]  & n603;
  assign n605 = ~n602 & ~n604;
  assign n606 = \a[60]  & ~\shift[0] ;
  assign n607 = ~\shift[1]  & n606;
  assign n608 = \a[59]  & \shift[0] ;
  assign n609 = ~\shift[1]  & n608;
  assign n610 = ~n607 & ~n609;
  assign n611 = n605 & n610;
  assign n612 = n288 & ~n611;
  assign n613 = ~n600 & ~n612;
  assign n614 = \a[49]  & \shift[0] ;
  assign n615 = \shift[1]  & n614;
  assign n616 = \a[50]  & ~\shift[0] ;
  assign n617 = \shift[1]  & n616;
  assign n618 = ~n615 & ~n617;
  assign n619 = \a[52]  & ~\shift[0] ;
  assign n620 = ~\shift[1]  & n619;
  assign n621 = \a[51]  & \shift[0] ;
  assign n622 = ~\shift[1]  & n621;
  assign n623 = ~n620 & ~n622;
  assign n624 = n618 & n623;
  assign n625 = n302 & ~n624;
  assign n626 = \a[53]  & \shift[0] ;
  assign n627 = \shift[1]  & n626;
  assign n628 = \a[54]  & ~\shift[0] ;
  assign n629 = \shift[1]  & n628;
  assign n630 = ~n627 & ~n629;
  assign n631 = \a[56]  & ~\shift[0] ;
  assign n632 = ~\shift[1]  & n631;
  assign n633 = \a[55]  & \shift[0] ;
  assign n634 = ~\shift[1]  & n633;
  assign n635 = ~n632 & ~n634;
  assign n636 = n630 & n635;
  assign n637 = n315 & ~n636;
  assign n638 = ~n625 & ~n637;
  assign n639 = n613 & n638;
  assign n640 = n426 & ~n639;
  assign n641 = \a[45]  & \shift[0] ;
  assign n642 = \shift[1]  & n641;
  assign n643 = \a[46]  & ~\shift[0] ;
  assign n644 = \shift[1]  & n643;
  assign n645 = ~n642 & ~n644;
  assign n646 = \a[48]  & ~\shift[0] ;
  assign n647 = ~\shift[1]  & n646;
  assign n648 = \a[47]  & \shift[0] ;
  assign n649 = ~\shift[1]  & n648;
  assign n650 = ~n647 & ~n649;
  assign n651 = n645 & n650;
  assign n652 = n275 & ~n651;
  assign n653 = \a[41]  & \shift[0] ;
  assign n654 = \shift[1]  & n653;
  assign n655 = \a[42]  & ~\shift[0] ;
  assign n656 = \shift[1]  & n655;
  assign n657 = ~n654 & ~n656;
  assign n658 = \a[44]  & ~\shift[0] ;
  assign n659 = ~\shift[1]  & n658;
  assign n660 = \a[43]  & \shift[0] ;
  assign n661 = ~\shift[1]  & n660;
  assign n662 = ~n659 & ~n661;
  assign n663 = n657 & n662;
  assign n664 = n288 & ~n663;
  assign n665 = ~n652 & ~n664;
  assign n666 = \a[33]  & \shift[0] ;
  assign n667 = \shift[1]  & n666;
  assign n668 = \a[34]  & ~\shift[0] ;
  assign n669 = \shift[1]  & n668;
  assign n670 = ~n667 & ~n669;
  assign n671 = \a[36]  & ~\shift[0] ;
  assign n672 = ~\shift[1]  & n671;
  assign n673 = \a[35]  & \shift[0] ;
  assign n674 = ~\shift[1]  & n673;
  assign n675 = ~n672 & ~n674;
  assign n676 = n670 & n675;
  assign n677 = n302 & ~n676;
  assign n678 = \a[40]  & ~\shift[0] ;
  assign n679 = ~\shift[1]  & n678;
  assign n680 = \a[37]  & \shift[0] ;
  assign n681 = \shift[1]  & n680;
  assign n682 = ~n679 & ~n681;
  assign n683 = \a[39]  & \shift[0] ;
  assign n684 = ~\shift[1]  & n683;
  assign n685 = \a[38]  & ~\shift[0] ;
  assign n686 = \shift[1]  & n685;
  assign n687 = ~n684 & ~n686;
  assign n688 = n682 & n687;
  assign n689 = n315 & ~n688;
  assign n690 = ~n677 & ~n689;
  assign n691 = n665 & n690;
  assign n692 = n479 & ~n691;
  assign n693 = ~n640 & ~n692;
  assign n694 = n588 & n693;
  assign n695 = \shift[6]  & ~n694;
  assign \result[0]  = n483 | n695;
  assign n697 = \a[81]  & ~\shift[0] ;
  assign n698 = ~\shift[1]  & n697;
  assign n699 = \a[78]  & \shift[0] ;
  assign n700 = \shift[1]  & n699;
  assign n701 = ~n698 & ~n700;
  assign n702 = \a[80]  & \shift[0] ;
  assign n703 = ~\shift[1]  & n702;
  assign n704 = \a[79]  & ~\shift[0] ;
  assign n705 = \shift[1]  & n704;
  assign n706 = ~n703 & ~n705;
  assign n707 = n701 & n706;
  assign n708 = n275 & ~n707;
  assign n709 = \a[77]  & ~\shift[0] ;
  assign n710 = ~\shift[1]  & n709;
  assign n711 = \a[74]  & \shift[0] ;
  assign n712 = \shift[1]  & n711;
  assign n713 = ~n710 & ~n712;
  assign n714 = \a[76]  & \shift[0] ;
  assign n715 = ~\shift[1]  & n714;
  assign n716 = \a[75]  & ~\shift[0] ;
  assign n717 = \shift[1]  & n716;
  assign n718 = ~n715 & ~n717;
  assign n719 = n713 & n718;
  assign n720 = n288 & ~n719;
  assign n721 = ~n708 & ~n720;
  assign n722 = \a[69]  & ~\shift[0] ;
  assign n723 = ~\shift[1]  & n722;
  assign n724 = \a[66]  & \shift[0] ;
  assign n725 = \shift[1]  & n724;
  assign n726 = ~n723 & ~n725;
  assign n727 = \a[68]  & \shift[0] ;
  assign n728 = ~\shift[1]  & n727;
  assign n729 = \a[67]  & ~\shift[0] ;
  assign n730 = \shift[1]  & n729;
  assign n731 = ~n728 & ~n730;
  assign n732 = n726 & n731;
  assign n733 = n302 & ~n732;
  assign n734 = \a[73]  & ~\shift[0] ;
  assign n735 = ~\shift[1]  & n734;
  assign n736 = \a[70]  & \shift[0] ;
  assign n737 = \shift[1]  & n736;
  assign n738 = ~n735 & ~n737;
  assign n739 = \a[72]  & \shift[0] ;
  assign n740 = ~\shift[1]  & n739;
  assign n741 = \a[71]  & ~\shift[0] ;
  assign n742 = \shift[1]  & n741;
  assign n743 = ~n740 & ~n742;
  assign n744 = n738 & n743;
  assign n745 = n315 & ~n744;
  assign n746 = ~n733 & ~n745;
  assign n747 = n721 & n746;
  assign n748 = n319 & ~n747;
  assign n749 = \a[97]  & ~\shift[0] ;
  assign n750 = ~\shift[1]  & n749;
  assign n751 = \a[94]  & \shift[0] ;
  assign n752 = \shift[1]  & n751;
  assign n753 = ~n750 & ~n752;
  assign n754 = \a[96]  & \shift[0] ;
  assign n755 = ~\shift[1]  & n754;
  assign n756 = \a[95]  & ~\shift[0] ;
  assign n757 = \shift[1]  & n756;
  assign n758 = ~n755 & ~n757;
  assign n759 = n753 & n758;
  assign n760 = n275 & ~n759;
  assign n761 = \a[93]  & ~\shift[0] ;
  assign n762 = ~\shift[1]  & n761;
  assign n763 = \a[90]  & \shift[0] ;
  assign n764 = \shift[1]  & n763;
  assign n765 = ~n762 & ~n764;
  assign n766 = \a[92]  & \shift[0] ;
  assign n767 = ~\shift[1]  & n766;
  assign n768 = \a[91]  & ~\shift[0] ;
  assign n769 = \shift[1]  & n768;
  assign n770 = ~n767 & ~n769;
  assign n771 = n765 & n770;
  assign n772 = n288 & ~n771;
  assign n773 = ~n760 & ~n772;
  assign n774 = \a[85]  & ~\shift[0] ;
  assign n775 = ~\shift[1]  & n774;
  assign n776 = \a[82]  & \shift[0] ;
  assign n777 = \shift[1]  & n776;
  assign n778 = ~n775 & ~n777;
  assign n779 = \a[84]  & \shift[0] ;
  assign n780 = ~\shift[1]  & n779;
  assign n781 = \a[83]  & ~\shift[0] ;
  assign n782 = \shift[1]  & n781;
  assign n783 = ~n780 & ~n782;
  assign n784 = n778 & n783;
  assign n785 = n302 & ~n784;
  assign n786 = \a[89]  & ~\shift[0] ;
  assign n787 = ~\shift[1]  & n786;
  assign n788 = \a[86]  & \shift[0] ;
  assign n789 = \shift[1]  & n788;
  assign n790 = ~n787 & ~n789;
  assign n791 = \a[88]  & \shift[0] ;
  assign n792 = ~\shift[1]  & n791;
  assign n793 = \a[87]  & ~\shift[0] ;
  assign n794 = \shift[1]  & n793;
  assign n795 = ~n792 & ~n794;
  assign n796 = n790 & n795;
  assign n797 = n315 & ~n796;
  assign n798 = ~n785 & ~n797;
  assign n799 = n773 & n798;
  assign n800 = n372 & ~n799;
  assign n801 = ~n748 & ~n800;
  assign n802 = \a[1]  & ~\shift[0] ;
  assign n803 = ~\shift[1]  & n802;
  assign n804 = \a[126]  & \shift[0] ;
  assign n805 = \shift[1]  & n804;
  assign n806 = ~n803 & ~n805;
  assign n807 = \a[0]  & \shift[0] ;
  assign n808 = ~\shift[1]  & n807;
  assign n809 = \a[127]  & ~\shift[0] ;
  assign n810 = \shift[1]  & n809;
  assign n811 = ~n808 & ~n810;
  assign n812 = n806 & n811;
  assign n813 = n275 & ~n812;
  assign n814 = \a[125]  & ~\shift[0] ;
  assign n815 = ~\shift[1]  & n814;
  assign n816 = \a[122]  & \shift[0] ;
  assign n817 = \shift[1]  & n816;
  assign n818 = ~n815 & ~n817;
  assign n819 = \a[124]  & \shift[0] ;
  assign n820 = ~\shift[1]  & n819;
  assign n821 = \a[123]  & ~\shift[0] ;
  assign n822 = \shift[1]  & n821;
  assign n823 = ~n820 & ~n822;
  assign n824 = n818 & n823;
  assign n825 = n288 & ~n824;
  assign n826 = ~n813 & ~n825;
  assign n827 = \a[117]  & ~\shift[0] ;
  assign n828 = ~\shift[1]  & n827;
  assign n829 = \a[114]  & \shift[0] ;
  assign n830 = \shift[1]  & n829;
  assign n831 = ~n828 & ~n830;
  assign n832 = \a[116]  & \shift[0] ;
  assign n833 = ~\shift[1]  & n832;
  assign n834 = \a[115]  & ~\shift[0] ;
  assign n835 = \shift[1]  & n834;
  assign n836 = ~n833 & ~n835;
  assign n837 = n831 & n836;
  assign n838 = n302 & ~n837;
  assign n839 = \a[121]  & ~\shift[0] ;
  assign n840 = ~\shift[1]  & n839;
  assign n841 = \a[118]  & \shift[0] ;
  assign n842 = \shift[1]  & n841;
  assign n843 = ~n840 & ~n842;
  assign n844 = \a[120]  & \shift[0] ;
  assign n845 = ~\shift[1]  & n844;
  assign n846 = \a[119]  & ~\shift[0] ;
  assign n847 = \shift[1]  & n846;
  assign n848 = ~n845 & ~n847;
  assign n849 = n843 & n848;
  assign n850 = n315 & ~n849;
  assign n851 = ~n838 & ~n850;
  assign n852 = n826 & n851;
  assign n853 = n426 & ~n852;
  assign n854 = \a[113]  & ~\shift[0] ;
  assign n855 = ~\shift[1]  & n854;
  assign n856 = \a[110]  & \shift[0] ;
  assign n857 = \shift[1]  & n856;
  assign n858 = ~n855 & ~n857;
  assign n859 = \a[112]  & \shift[0] ;
  assign n860 = ~\shift[1]  & n859;
  assign n861 = \a[111]  & ~\shift[0] ;
  assign n862 = \shift[1]  & n861;
  assign n863 = ~n860 & ~n862;
  assign n864 = n858 & n863;
  assign n865 = n275 & ~n864;
  assign n866 = \a[109]  & ~\shift[0] ;
  assign n867 = ~\shift[1]  & n866;
  assign n868 = \a[106]  & \shift[0] ;
  assign n869 = \shift[1]  & n868;
  assign n870 = ~n867 & ~n869;
  assign n871 = \a[108]  & \shift[0] ;
  assign n872 = ~\shift[1]  & n871;
  assign n873 = \a[107]  & ~\shift[0] ;
  assign n874 = \shift[1]  & n873;
  assign n875 = ~n872 & ~n874;
  assign n876 = n870 & n875;
  assign n877 = n288 & ~n876;
  assign n878 = ~n865 & ~n877;
  assign n879 = \a[101]  & ~\shift[0] ;
  assign n880 = ~\shift[1]  & n879;
  assign n881 = \a[98]  & \shift[0] ;
  assign n882 = \shift[1]  & n881;
  assign n883 = ~n880 & ~n882;
  assign n884 = \a[100]  & \shift[0] ;
  assign n885 = ~\shift[1]  & n884;
  assign n886 = \a[99]  & ~\shift[0] ;
  assign n887 = \shift[1]  & n886;
  assign n888 = ~n885 & ~n887;
  assign n889 = n883 & n888;
  assign n890 = n302 & ~n889;
  assign n891 = \a[105]  & ~\shift[0] ;
  assign n892 = ~\shift[1]  & n891;
  assign n893 = \a[102]  & \shift[0] ;
  assign n894 = \shift[1]  & n893;
  assign n895 = ~n892 & ~n894;
  assign n896 = \a[104]  & \shift[0] ;
  assign n897 = ~\shift[1]  & n896;
  assign n898 = \a[103]  & ~\shift[0] ;
  assign n899 = \shift[1]  & n898;
  assign n900 = ~n897 & ~n899;
  assign n901 = n895 & n900;
  assign n902 = n315 & ~n901;
  assign n903 = ~n890 & ~n902;
  assign n904 = n878 & n903;
  assign n905 = n479 & ~n904;
  assign n906 = ~n853 & ~n905;
  assign n907 = n801 & n906;
  assign n908 = ~\shift[6]  & ~n907;
  assign n909 = \a[65]  & ~\shift[0] ;
  assign n910 = ~\shift[1]  & n909;
  assign n911 = \a[62]  & \shift[0] ;
  assign n912 = \shift[1]  & n911;
  assign n913 = ~n910 & ~n912;
  assign n914 = \a[64]  & \shift[0] ;
  assign n915 = ~\shift[1]  & n914;
  assign n916 = \a[63]  & ~\shift[0] ;
  assign n917 = \shift[1]  & n916;
  assign n918 = ~n915 & ~n917;
  assign n919 = n913 & n918;
  assign n920 = n275 & ~n919;
  assign n921 = \a[61]  & ~\shift[0] ;
  assign n922 = ~\shift[1]  & n921;
  assign n923 = \a[58]  & \shift[0] ;
  assign n924 = \shift[1]  & n923;
  assign n925 = ~n922 & ~n924;
  assign n926 = \a[60]  & \shift[0] ;
  assign n927 = ~\shift[1]  & n926;
  assign n928 = \a[59]  & ~\shift[0] ;
  assign n929 = \shift[1]  & n928;
  assign n930 = ~n927 & ~n929;
  assign n931 = n925 & n930;
  assign n932 = n288 & ~n931;
  assign n933 = ~n920 & ~n932;
  assign n934 = \a[53]  & ~\shift[0] ;
  assign n935 = ~\shift[1]  & n934;
  assign n936 = \a[50]  & \shift[0] ;
  assign n937 = \shift[1]  & n936;
  assign n938 = ~n935 & ~n937;
  assign n939 = \a[52]  & \shift[0] ;
  assign n940 = ~\shift[1]  & n939;
  assign n941 = \a[51]  & ~\shift[0] ;
  assign n942 = \shift[1]  & n941;
  assign n943 = ~n940 & ~n942;
  assign n944 = n938 & n943;
  assign n945 = n302 & ~n944;
  assign n946 = \a[57]  & ~\shift[0] ;
  assign n947 = ~\shift[1]  & n946;
  assign n948 = \a[54]  & \shift[0] ;
  assign n949 = \shift[1]  & n948;
  assign n950 = ~n947 & ~n949;
  assign n951 = \a[56]  & \shift[0] ;
  assign n952 = ~\shift[1]  & n951;
  assign n953 = \a[55]  & ~\shift[0] ;
  assign n954 = \shift[1]  & n953;
  assign n955 = ~n952 & ~n954;
  assign n956 = n950 & n955;
  assign n957 = n315 & ~n956;
  assign n958 = ~n945 & ~n957;
  assign n959 = n933 & n958;
  assign n960 = n426 & ~n959;
  assign n961 = \a[17]  & ~\shift[0] ;
  assign n962 = ~\shift[1]  & n961;
  assign n963 = \a[14]  & \shift[0] ;
  assign n964 = \shift[1]  & n963;
  assign n965 = ~n962 & ~n964;
  assign n966 = \a[16]  & \shift[0] ;
  assign n967 = ~\shift[1]  & n966;
  assign n968 = \a[15]  & ~\shift[0] ;
  assign n969 = \shift[1]  & n968;
  assign n970 = ~n967 & ~n969;
  assign n971 = n965 & n970;
  assign n972 = n275 & ~n971;
  assign n973 = \a[13]  & ~\shift[0] ;
  assign n974 = ~\shift[1]  & n973;
  assign n975 = \a[10]  & \shift[0] ;
  assign n976 = \shift[1]  & n975;
  assign n977 = ~n974 & ~n976;
  assign n978 = \a[12]  & \shift[0] ;
  assign n979 = ~\shift[1]  & n978;
  assign n980 = \a[11]  & ~\shift[0] ;
  assign n981 = \shift[1]  & n980;
  assign n982 = ~n979 & ~n981;
  assign n983 = n977 & n982;
  assign n984 = n288 & ~n983;
  assign n985 = ~n972 & ~n984;
  assign n986 = \a[5]  & ~\shift[0] ;
  assign n987 = ~\shift[1]  & n986;
  assign n988 = \a[2]  & \shift[0] ;
  assign n989 = \shift[1]  & n988;
  assign n990 = ~n987 & ~n989;
  assign n991 = \a[4]  & \shift[0] ;
  assign n992 = ~\shift[1]  & n991;
  assign n993 = \a[3]  & ~\shift[0] ;
  assign n994 = \shift[1]  & n993;
  assign n995 = ~n992 & ~n994;
  assign n996 = n990 & n995;
  assign n997 = n302 & ~n996;
  assign n998 = \a[9]  & ~\shift[0] ;
  assign n999 = ~\shift[1]  & n998;
  assign n1000 = \a[6]  & \shift[0] ;
  assign n1001 = \shift[1]  & n1000;
  assign n1002 = ~n999 & ~n1001;
  assign n1003 = \a[8]  & \shift[0] ;
  assign n1004 = ~\shift[1]  & n1003;
  assign n1005 = \a[7]  & ~\shift[0] ;
  assign n1006 = \shift[1]  & n1005;
  assign n1007 = ~n1004 & ~n1006;
  assign n1008 = n1002 & n1007;
  assign n1009 = n315 & ~n1008;
  assign n1010 = ~n997 & ~n1009;
  assign n1011 = n985 & n1010;
  assign n1012 = n319 & ~n1011;
  assign n1013 = ~n960 & ~n1012;
  assign n1014 = \a[49]  & ~\shift[0] ;
  assign n1015 = ~\shift[1]  & n1014;
  assign n1016 = \a[46]  & \shift[0] ;
  assign n1017 = \shift[1]  & n1016;
  assign n1018 = ~n1015 & ~n1017;
  assign n1019 = \a[48]  & \shift[0] ;
  assign n1020 = ~\shift[1]  & n1019;
  assign n1021 = \a[47]  & ~\shift[0] ;
  assign n1022 = \shift[1]  & n1021;
  assign n1023 = ~n1020 & ~n1022;
  assign n1024 = n1018 & n1023;
  assign n1025 = n275 & ~n1024;
  assign n1026 = \a[42]  & \shift[0] ;
  assign n1027 = \shift[1]  & n1026;
  assign n1028 = \a[43]  & ~\shift[0] ;
  assign n1029 = \shift[1]  & n1028;
  assign n1030 = ~n1027 & ~n1029;
  assign n1031 = \a[45]  & ~\shift[0] ;
  assign n1032 = ~\shift[1]  & n1031;
  assign n1033 = \a[44]  & \shift[0] ;
  assign n1034 = ~\shift[1]  & n1033;
  assign n1035 = ~n1032 & ~n1034;
  assign n1036 = n1030 & n1035;
  assign n1037 = n288 & ~n1036;
  assign n1038 = ~n1025 & ~n1037;
  assign n1039 = \a[37]  & ~\shift[0] ;
  assign n1040 = ~\shift[1]  & n1039;
  assign n1041 = \a[34]  & \shift[0] ;
  assign n1042 = \shift[1]  & n1041;
  assign n1043 = ~n1040 & ~n1042;
  assign n1044 = \a[36]  & \shift[0] ;
  assign n1045 = ~\shift[1]  & n1044;
  assign n1046 = \a[35]  & ~\shift[0] ;
  assign n1047 = \shift[1]  & n1046;
  assign n1048 = ~n1045 & ~n1047;
  assign n1049 = n1043 & n1048;
  assign n1050 = n302 & ~n1049;
  assign n1051 = \a[41]  & ~\shift[0] ;
  assign n1052 = ~\shift[1]  & n1051;
  assign n1053 = \a[40]  & \shift[0] ;
  assign n1054 = ~\shift[1]  & n1053;
  assign n1055 = ~n1052 & ~n1054;
  assign n1056 = \a[39]  & ~\shift[0] ;
  assign n1057 = \shift[1]  & n1056;
  assign n1058 = \a[38]  & \shift[0] ;
  assign n1059 = \shift[1]  & n1058;
  assign n1060 = ~n1057 & ~n1059;
  assign n1061 = n1055 & n1060;
  assign n1062 = n315 & ~n1061;
  assign n1063 = ~n1050 & ~n1062;
  assign n1064 = n1038 & n1063;
  assign n1065 = n479 & ~n1064;
  assign n1066 = \a[33]  & ~\shift[0] ;
  assign n1067 = ~\shift[1]  & n1066;
  assign n1068 = \a[30]  & \shift[0] ;
  assign n1069 = \shift[1]  & n1068;
  assign n1070 = ~n1067 & ~n1069;
  assign n1071 = \a[32]  & \shift[0] ;
  assign n1072 = ~\shift[1]  & n1071;
  assign n1073 = \a[31]  & ~\shift[0] ;
  assign n1074 = \shift[1]  & n1073;
  assign n1075 = ~n1072 & ~n1074;
  assign n1076 = n1070 & n1075;
  assign n1077 = n275 & ~n1076;
  assign n1078 = \a[29]  & ~\shift[0] ;
  assign n1079 = ~\shift[1]  & n1078;
  assign n1080 = \a[26]  & \shift[0] ;
  assign n1081 = \shift[1]  & n1080;
  assign n1082 = ~n1079 & ~n1081;
  assign n1083 = \a[28]  & \shift[0] ;
  assign n1084 = ~\shift[1]  & n1083;
  assign n1085 = \a[27]  & ~\shift[0] ;
  assign n1086 = \shift[1]  & n1085;
  assign n1087 = ~n1084 & ~n1086;
  assign n1088 = n1082 & n1087;
  assign n1089 = n288 & ~n1088;
  assign n1090 = ~n1077 & ~n1089;
  assign n1091 = \a[21]  & ~\shift[0] ;
  assign n1092 = ~\shift[1]  & n1091;
  assign n1093 = \a[18]  & \shift[0] ;
  assign n1094 = \shift[1]  & n1093;
  assign n1095 = ~n1092 & ~n1094;
  assign n1096 = \a[20]  & \shift[0] ;
  assign n1097 = ~\shift[1]  & n1096;
  assign n1098 = \a[19]  & ~\shift[0] ;
  assign n1099 = \shift[1]  & n1098;
  assign n1100 = ~n1097 & ~n1099;
  assign n1101 = n1095 & n1100;
  assign n1102 = n302 & ~n1101;
  assign n1103 = \a[25]  & ~\shift[0] ;
  assign n1104 = ~\shift[1]  & n1103;
  assign n1105 = \a[22]  & \shift[0] ;
  assign n1106 = \shift[1]  & n1105;
  assign n1107 = ~n1104 & ~n1106;
  assign n1108 = \a[24]  & \shift[0] ;
  assign n1109 = ~\shift[1]  & n1108;
  assign n1110 = \a[23]  & ~\shift[0] ;
  assign n1111 = \shift[1]  & n1110;
  assign n1112 = ~n1109 & ~n1111;
  assign n1113 = n1107 & n1112;
  assign n1114 = n315 & ~n1113;
  assign n1115 = ~n1102 & ~n1114;
  assign n1116 = n1090 & n1115;
  assign n1117 = n372 & ~n1116;
  assign n1118 = ~n1065 & ~n1117;
  assign n1119 = n1013 & n1118;
  assign n1120 = \shift[6]  & ~n1119;
  assign \result[1]  = n908 | n1120;
  assign n1122 = ~\shift[1]  & n346;
  assign n1123 = ~\shift[1]  & n348;
  assign n1124 = ~n1122 & ~n1123;
  assign n1125 = \shift[1]  & n269;
  assign n1126 = \shift[1]  & n271;
  assign n1127 = ~n1125 & ~n1126;
  assign n1128 = n1124 & n1127;
  assign n1129 = n275 & ~n1128;
  assign n1130 = ~\shift[1]  & n264;
  assign n1131 = ~\shift[1]  & n266;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = \shift[1]  & n282;
  assign n1134 = \shift[1]  & n284;
  assign n1135 = ~n1133 & ~n1134;
  assign n1136 = n1132 & n1135;
  assign n1137 = n288 & ~n1136;
  assign n1138 = ~n1129 & ~n1137;
  assign n1139 = ~\shift[1]  & n304;
  assign n1140 = ~\shift[1]  & n306;
  assign n1141 = ~n1139 & ~n1140;
  assign n1142 = \shift[1]  & n296;
  assign n1143 = \shift[1]  & n298;
  assign n1144 = ~n1142 & ~n1143;
  assign n1145 = n1141 & n1144;
  assign n1146 = n302 & ~n1145;
  assign n1147 = ~\shift[1]  & n277;
  assign n1148 = ~\shift[1]  & n279;
  assign n1149 = ~n1147 & ~n1148;
  assign n1150 = \shift[1]  & n309;
  assign n1151 = \shift[1]  & n311;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = n1149 & n1152;
  assign n1154 = n315 & ~n1153;
  assign n1155 = ~n1146 & ~n1154;
  assign n1156 = n1138 & n1155;
  assign n1157 = n319 & ~n1156;
  assign n1158 = ~\shift[1]  & n453;
  assign n1159 = ~\shift[1]  & n455;
  assign n1160 = ~n1158 & ~n1159;
  assign n1161 = \shift[1]  & n326;
  assign n1162 = \shift[1]  & n328;
  assign n1163 = ~n1161 & ~n1162;
  assign n1164 = n1160 & n1163;
  assign n1165 = n275 & ~n1164;
  assign n1166 = ~\shift[1]  & n321;
  assign n1167 = ~\shift[1]  & n323;
  assign n1168 = ~n1166 & ~n1167;
  assign n1169 = \shift[1]  & n338;
  assign n1170 = \shift[1]  & n340;
  assign n1171 = ~n1169 & ~n1170;
  assign n1172 = n1168 & n1171;
  assign n1173 = n288 & ~n1172;
  assign n1174 = ~n1165 & ~n1173;
  assign n1175 = ~\shift[1]  & n358;
  assign n1176 = ~\shift[1]  & n360;
  assign n1177 = ~n1175 & ~n1176;
  assign n1178 = \shift[1]  & n351;
  assign n1179 = \shift[1]  & n353;
  assign n1180 = ~n1178 & ~n1179;
  assign n1181 = n1177 & n1180;
  assign n1182 = n302 & ~n1181;
  assign n1183 = ~\shift[1]  & n333;
  assign n1184 = ~\shift[1]  & n335;
  assign n1185 = ~n1183 & ~n1184;
  assign n1186 = \shift[1]  & n363;
  assign n1187 = \shift[1]  & n365;
  assign n1188 = ~n1186 & ~n1187;
  assign n1189 = n1185 & n1188;
  assign n1190 = n315 & ~n1189;
  assign n1191 = ~n1182 & ~n1190;
  assign n1192 = n1174 & n1191;
  assign n1193 = n372 & ~n1192;
  assign n1194 = ~n1157 & ~n1193;
  assign n1195 = ~\shift[1]  & n509;
  assign n1196 = ~\shift[1]  & n511;
  assign n1197 = ~n1195 & ~n1196;
  assign n1198 = \shift[1]  & n380;
  assign n1199 = \shift[1]  & n382;
  assign n1200 = ~n1198 & ~n1199;
  assign n1201 = n1197 & n1200;
  assign n1202 = n275 & ~n1201;
  assign n1203 = ~\shift[1]  & n375;
  assign n1204 = ~\shift[1]  & n377;
  assign n1205 = ~n1203 & ~n1204;
  assign n1206 = \shift[1]  & n392;
  assign n1207 = \shift[1]  & n394;
  assign n1208 = ~n1206 & ~n1207;
  assign n1209 = n1205 & n1208;
  assign n1210 = n288 & ~n1209;
  assign n1211 = ~n1202 & ~n1210;
  assign n1212 = ~\shift[1]  & n412;
  assign n1213 = ~\shift[1]  & n414;
  assign n1214 = ~n1212 & ~n1213;
  assign n1215 = \shift[1]  & n405;
  assign n1216 = \shift[1]  & n407;
  assign n1217 = ~n1215 & ~n1216;
  assign n1218 = n1214 & n1217;
  assign n1219 = n302 & ~n1218;
  assign n1220 = ~\shift[1]  & n387;
  assign n1221 = ~\shift[1]  & n389;
  assign n1222 = ~n1220 & ~n1221;
  assign n1223 = \shift[1]  & n417;
  assign n1224 = \shift[1]  & n419;
  assign n1225 = ~n1223 & ~n1224;
  assign n1226 = n1222 & n1225;
  assign n1227 = n315 & ~n1226;
  assign n1228 = ~n1219 & ~n1227;
  assign n1229 = n1211 & n1228;
  assign n1230 = n426 & ~n1229;
  assign n1231 = ~\shift[1]  & n400;
  assign n1232 = ~\shift[1]  & n402;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = \shift[1]  & n433;
  assign n1235 = \shift[1]  & n435;
  assign n1236 = ~n1234 & ~n1235;
  assign n1237 = n1233 & n1236;
  assign n1238 = n275 & ~n1237;
  assign n1239 = ~\shift[1]  & n428;
  assign n1240 = ~\shift[1]  & n430;
  assign n1241 = ~n1239 & ~n1240;
  assign n1242 = \shift[1]  & n445;
  assign n1243 = \shift[1]  & n447;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = n1241 & n1244;
  assign n1246 = n288 & ~n1245;
  assign n1247 = ~n1238 & ~n1246;
  assign n1248 = ~\shift[1]  & n465;
  assign n1249 = ~\shift[1]  & n467;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = \shift[1]  & n458;
  assign n1252 = \shift[1]  & n460;
  assign n1253 = ~n1251 & ~n1252;
  assign n1254 = n1250 & n1253;
  assign n1255 = n302 & ~n1254;
  assign n1256 = ~\shift[1]  & n440;
  assign n1257 = ~\shift[1]  & n442;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = \shift[1]  & n470;
  assign n1260 = \shift[1]  & n472;
  assign n1261 = ~n1259 & ~n1260;
  assign n1262 = n1258 & n1261;
  assign n1263 = n315 & ~n1262;
  assign n1264 = ~n1255 & ~n1263;
  assign n1265 = n1247 & n1264;
  assign n1266 = n479 & ~n1265;
  assign n1267 = ~n1230 & ~n1266;
  assign n1268 = n1194 & n1267;
  assign n1269 = ~\shift[6]  & ~n1268;
  assign n1270 = ~\shift[1]  & n291;
  assign n1271 = ~\shift[1]  & n293;
  assign n1272 = ~n1270 & ~n1271;
  assign n1273 = \shift[1]  & n594;
  assign n1274 = \shift[1]  & n596;
  assign n1275 = ~n1273 & ~n1274;
  assign n1276 = n1272 & n1275;
  assign n1277 = n275 & ~n1276;
  assign n1278 = ~\shift[1]  & n589;
  assign n1279 = ~\shift[1]  & n591;
  assign n1280 = ~n1278 & ~n1279;
  assign n1281 = \shift[1]  & n606;
  assign n1282 = \shift[1]  & n608;
  assign n1283 = ~n1281 & ~n1282;
  assign n1284 = n1280 & n1283;
  assign n1285 = n288 & ~n1284;
  assign n1286 = ~n1277 & ~n1285;
  assign n1287 = ~\shift[1]  & n626;
  assign n1288 = ~\shift[1]  & n628;
  assign n1289 = ~n1287 & ~n1288;
  assign n1290 = \shift[1]  & n619;
  assign n1291 = \shift[1]  & n621;
  assign n1292 = ~n1290 & ~n1291;
  assign n1293 = n1289 & n1292;
  assign n1294 = n302 & ~n1293;
  assign n1295 = ~\shift[1]  & n601;
  assign n1296 = ~\shift[1]  & n603;
  assign n1297 = ~n1295 & ~n1296;
  assign n1298 = \shift[1]  & n631;
  assign n1299 = \shift[1]  & n633;
  assign n1300 = ~n1298 & ~n1299;
  assign n1301 = n1297 & n1300;
  assign n1302 = n315 & ~n1301;
  assign n1303 = ~n1294 & ~n1302;
  assign n1304 = n1286 & n1303;
  assign n1305 = n426 & ~n1304;
  assign n1306 = ~\shift[1]  & n561;
  assign n1307 = ~\shift[1]  & n563;
  assign n1308 = ~n1306 & ~n1307;
  assign n1309 = \shift[1]  & n489;
  assign n1310 = \shift[1]  & n491;
  assign n1311 = ~n1309 & ~n1310;
  assign n1312 = n1308 & n1311;
  assign n1313 = n275 & ~n1312;
  assign n1314 = ~\shift[1]  & n484;
  assign n1315 = ~\shift[1]  & n486;
  assign n1316 = ~n1314 & ~n1315;
  assign n1317 = \shift[1]  & n501;
  assign n1318 = \shift[1]  & n503;
  assign n1319 = ~n1317 & ~n1318;
  assign n1320 = n1316 & n1319;
  assign n1321 = n288 & ~n1320;
  assign n1322 = ~n1313 & ~n1321;
  assign n1323 = ~\shift[1]  & n521;
  assign n1324 = ~\shift[1]  & n523;
  assign n1325 = ~n1323 & ~n1324;
  assign n1326 = \shift[1]  & n514;
  assign n1327 = \shift[1]  & n516;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = n1325 & n1328;
  assign n1330 = n302 & ~n1329;
  assign n1331 = ~\shift[1]  & n496;
  assign n1332 = ~\shift[1]  & n498;
  assign n1333 = ~n1331 & ~n1332;
  assign n1334 = \shift[1]  & n526;
  assign n1335 = \shift[1]  & n528;
  assign n1336 = ~n1334 & ~n1335;
  assign n1337 = n1333 & n1336;
  assign n1338 = n315 & ~n1337;
  assign n1339 = ~n1330 & ~n1338;
  assign n1340 = n1322 & n1339;
  assign n1341 = n319 & ~n1340;
  assign n1342 = ~n1305 & ~n1341;
  assign n1343 = ~\shift[1]  & n614;
  assign n1344 = ~\shift[1]  & n616;
  assign n1345 = ~n1343 & ~n1344;
  assign n1346 = \shift[1]  & n646;
  assign n1347 = \shift[1]  & n648;
  assign n1348 = ~n1346 & ~n1347;
  assign n1349 = n1345 & n1348;
  assign n1350 = n275 & ~n1349;
  assign n1351 = \shift[1]  & n660;
  assign n1352 = \shift[1]  & n658;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = ~\shift[1]  & n643;
  assign n1355 = ~\shift[1]  & n641;
  assign n1356 = ~n1354 & ~n1355;
  assign n1357 = n1353 & n1356;
  assign n1358 = n288 & ~n1357;
  assign n1359 = ~n1350 & ~n1358;
  assign n1360 = ~\shift[1]  & n680;
  assign n1361 = ~\shift[1]  & n685;
  assign n1362 = ~n1360 & ~n1361;
  assign n1363 = \shift[1]  & n671;
  assign n1364 = \shift[1]  & n673;
  assign n1365 = ~n1363 & ~n1364;
  assign n1366 = n1362 & n1365;
  assign n1367 = n302 & ~n1366;
  assign n1368 = ~\shift[1]  & n653;
  assign n1369 = ~\shift[1]  & n655;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = \shift[1]  & n683;
  assign n1372 = \shift[1]  & n678;
  assign n1373 = ~n1371 & ~n1372;
  assign n1374 = n1370 & n1373;
  assign n1375 = n315 & ~n1374;
  assign n1376 = ~n1367 & ~n1375;
  assign n1377 = n1359 & n1376;
  assign n1378 = n479 & ~n1377;
  assign n1379 = ~\shift[1]  & n666;
  assign n1380 = ~\shift[1]  & n668;
  assign n1381 = ~n1379 & ~n1380;
  assign n1382 = \shift[1]  & n541;
  assign n1383 = \shift[1]  & n543;
  assign n1384 = ~n1382 & ~n1383;
  assign n1385 = n1381 & n1384;
  assign n1386 = n275 & ~n1385;
  assign n1387 = ~\shift[1]  & n536;
  assign n1388 = ~\shift[1]  & n538;
  assign n1389 = ~n1387 & ~n1388;
  assign n1390 = \shift[1]  & n553;
  assign n1391 = \shift[1]  & n555;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = n1389 & n1392;
  assign n1394 = n288 & ~n1393;
  assign n1395 = ~n1386 & ~n1394;
  assign n1396 = ~\shift[1]  & n573;
  assign n1397 = ~\shift[1]  & n575;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = \shift[1]  & n566;
  assign n1400 = \shift[1]  & n568;
  assign n1401 = ~n1399 & ~n1400;
  assign n1402 = n1398 & n1401;
  assign n1403 = n302 & ~n1402;
  assign n1404 = ~\shift[1]  & n548;
  assign n1405 = ~\shift[1]  & n550;
  assign n1406 = ~n1404 & ~n1405;
  assign n1407 = \shift[1]  & n578;
  assign n1408 = \shift[1]  & n580;
  assign n1409 = ~n1407 & ~n1408;
  assign n1410 = n1406 & n1409;
  assign n1411 = n315 & ~n1410;
  assign n1412 = ~n1403 & ~n1411;
  assign n1413 = n1395 & n1412;
  assign n1414 = n372 & ~n1413;
  assign n1415 = ~n1378 & ~n1414;
  assign n1416 = n1342 & n1415;
  assign n1417 = \shift[6]  & ~n1416;
  assign \result[2]  = n1269 | n1417;
  assign n1419 = \shift[1]  & n854;
  assign n1420 = ~\shift[1]  & n829;
  assign n1421 = ~n1419 & ~n1420;
  assign n1422 = \shift[1]  & n859;
  assign n1423 = ~\shift[1]  & n834;
  assign n1424 = ~n1422 & ~n1423;
  assign n1425 = n1421 & n1424;
  assign n1426 = n275 & ~n1425;
  assign n1427 = \shift[1]  & n866;
  assign n1428 = ~\shift[1]  & n856;
  assign n1429 = ~n1427 & ~n1428;
  assign n1430 = \shift[1]  & n871;
  assign n1431 = ~\shift[1]  & n861;
  assign n1432 = ~n1430 & ~n1431;
  assign n1433 = n1429 & n1432;
  assign n1434 = n288 & ~n1433;
  assign n1435 = ~n1426 & ~n1434;
  assign n1436 = \shift[1]  & n879;
  assign n1437 = ~\shift[1]  & n893;
  assign n1438 = ~n1436 & ~n1437;
  assign n1439 = \shift[1]  & n884;
  assign n1440 = ~\shift[1]  & n898;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = n1438 & n1441;
  assign n1443 = n302 & ~n1442;
  assign n1444 = \shift[1]  & n891;
  assign n1445 = ~\shift[1]  & n868;
  assign n1446 = ~n1444 & ~n1445;
  assign n1447 = \shift[1]  & n896;
  assign n1448 = ~\shift[1]  & n873;
  assign n1449 = ~n1447 & ~n1448;
  assign n1450 = n1446 & n1449;
  assign n1451 = n315 & ~n1450;
  assign n1452 = ~n1443 & ~n1451;
  assign n1453 = n1435 & n1452;
  assign n1454 = n479 & ~n1453;
  assign n1455 = \shift[1]  & n749;
  assign n1456 = ~\shift[1]  & n881;
  assign n1457 = ~n1455 & ~n1456;
  assign n1458 = \shift[1]  & n754;
  assign n1459 = ~\shift[1]  & n886;
  assign n1460 = ~n1458 & ~n1459;
  assign n1461 = n1457 & n1460;
  assign n1462 = n275 & ~n1461;
  assign n1463 = \shift[1]  & n761;
  assign n1464 = ~\shift[1]  & n751;
  assign n1465 = ~n1463 & ~n1464;
  assign n1466 = \shift[1]  & n766;
  assign n1467 = ~\shift[1]  & n756;
  assign n1468 = ~n1466 & ~n1467;
  assign n1469 = n1465 & n1468;
  assign n1470 = n288 & ~n1469;
  assign n1471 = ~n1462 & ~n1470;
  assign n1472 = \shift[1]  & n774;
  assign n1473 = ~\shift[1]  & n788;
  assign n1474 = ~n1472 & ~n1473;
  assign n1475 = \shift[1]  & n779;
  assign n1476 = ~\shift[1]  & n793;
  assign n1477 = ~n1475 & ~n1476;
  assign n1478 = n1474 & n1477;
  assign n1479 = n302 & ~n1478;
  assign n1480 = \shift[1]  & n786;
  assign n1481 = ~\shift[1]  & n763;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = \shift[1]  & n791;
  assign n1484 = ~\shift[1]  & n768;
  assign n1485 = ~n1483 & ~n1484;
  assign n1486 = n1482 & n1485;
  assign n1487 = n315 & ~n1486;
  assign n1488 = ~n1479 & ~n1487;
  assign n1489 = n1471 & n1488;
  assign n1490 = n372 & ~n1489;
  assign n1491 = ~n1454 & ~n1490;
  assign n1492 = \shift[1]  & n802;
  assign n1493 = ~\shift[1]  & n988;
  assign n1494 = ~n1492 & ~n1493;
  assign n1495 = \shift[1]  & n807;
  assign n1496 = ~\shift[1]  & n993;
  assign n1497 = ~n1495 & ~n1496;
  assign n1498 = n1494 & n1497;
  assign n1499 = n275 & ~n1498;
  assign n1500 = \shift[1]  & n814;
  assign n1501 = ~\shift[1]  & n804;
  assign n1502 = ~n1500 & ~n1501;
  assign n1503 = \shift[1]  & n819;
  assign n1504 = ~\shift[1]  & n809;
  assign n1505 = ~n1503 & ~n1504;
  assign n1506 = n1502 & n1505;
  assign n1507 = n288 & ~n1506;
  assign n1508 = ~n1499 & ~n1507;
  assign n1509 = \shift[1]  & n827;
  assign n1510 = ~\shift[1]  & n841;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = \shift[1]  & n832;
  assign n1513 = ~\shift[1]  & n846;
  assign n1514 = ~n1512 & ~n1513;
  assign n1515 = n1511 & n1514;
  assign n1516 = n302 & ~n1515;
  assign n1517 = \shift[1]  & n839;
  assign n1518 = ~\shift[1]  & n816;
  assign n1519 = ~n1517 & ~n1518;
  assign n1520 = \shift[1]  & n844;
  assign n1521 = ~\shift[1]  & n821;
  assign n1522 = ~n1520 & ~n1521;
  assign n1523 = n1519 & n1522;
  assign n1524 = n315 & ~n1523;
  assign n1525 = ~n1516 & ~n1524;
  assign n1526 = n1508 & n1525;
  assign n1527 = n426 & ~n1526;
  assign n1528 = \shift[1]  & n697;
  assign n1529 = ~\shift[1]  & n776;
  assign n1530 = ~n1528 & ~n1529;
  assign n1531 = \shift[1]  & n702;
  assign n1532 = ~\shift[1]  & n781;
  assign n1533 = ~n1531 & ~n1532;
  assign n1534 = n1530 & n1533;
  assign n1535 = n275 & ~n1534;
  assign n1536 = \shift[1]  & n709;
  assign n1537 = ~\shift[1]  & n699;
  assign n1538 = ~n1536 & ~n1537;
  assign n1539 = \shift[1]  & n714;
  assign n1540 = ~\shift[1]  & n704;
  assign n1541 = ~n1539 & ~n1540;
  assign n1542 = n1538 & n1541;
  assign n1543 = n288 & ~n1542;
  assign n1544 = ~n1535 & ~n1543;
  assign n1545 = \shift[1]  & n722;
  assign n1546 = ~\shift[1]  & n736;
  assign n1547 = ~n1545 & ~n1546;
  assign n1548 = \shift[1]  & n727;
  assign n1549 = ~\shift[1]  & n741;
  assign n1550 = ~n1548 & ~n1549;
  assign n1551 = n1547 & n1550;
  assign n1552 = n302 & ~n1551;
  assign n1553 = \shift[1]  & n734;
  assign n1554 = ~\shift[1]  & n711;
  assign n1555 = ~n1553 & ~n1554;
  assign n1556 = \shift[1]  & n739;
  assign n1557 = ~\shift[1]  & n716;
  assign n1558 = ~n1556 & ~n1557;
  assign n1559 = n1555 & n1558;
  assign n1560 = n315 & ~n1559;
  assign n1561 = ~n1552 & ~n1560;
  assign n1562 = n1544 & n1561;
  assign n1563 = n319 & ~n1562;
  assign n1564 = ~n1527 & ~n1563;
  assign n1565 = n1491 & n1564;
  assign n1566 = ~\shift[6]  & ~n1565;
  assign n1567 = \shift[1]  & n909;
  assign n1568 = ~\shift[1]  & n724;
  assign n1569 = ~n1567 & ~n1568;
  assign n1570 = \shift[1]  & n914;
  assign n1571 = ~\shift[1]  & n729;
  assign n1572 = ~n1570 & ~n1571;
  assign n1573 = n1569 & n1572;
  assign n1574 = n275 & ~n1573;
  assign n1575 = \shift[1]  & n921;
  assign n1576 = ~\shift[1]  & n911;
  assign n1577 = ~n1575 & ~n1576;
  assign n1578 = \shift[1]  & n926;
  assign n1579 = ~\shift[1]  & n916;
  assign n1580 = ~n1578 & ~n1579;
  assign n1581 = n1577 & n1580;
  assign n1582 = n288 & ~n1581;
  assign n1583 = ~n1574 & ~n1582;
  assign n1584 = \shift[1]  & n934;
  assign n1585 = ~\shift[1]  & n948;
  assign n1586 = ~n1584 & ~n1585;
  assign n1587 = \shift[1]  & n939;
  assign n1588 = ~\shift[1]  & n953;
  assign n1589 = ~n1587 & ~n1588;
  assign n1590 = n1586 & n1589;
  assign n1591 = n302 & ~n1590;
  assign n1592 = \shift[1]  & n946;
  assign n1593 = ~\shift[1]  & n923;
  assign n1594 = ~n1592 & ~n1593;
  assign n1595 = \shift[1]  & n951;
  assign n1596 = ~\shift[1]  & n928;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = n1594 & n1597;
  assign n1599 = n315 & ~n1598;
  assign n1600 = ~n1591 & ~n1599;
  assign n1601 = n1583 & n1600;
  assign n1602 = n426 & ~n1601;
  assign n1603 = \shift[1]  & n1014;
  assign n1604 = ~\shift[1]  & n936;
  assign n1605 = ~n1603 & ~n1604;
  assign n1606 = \shift[1]  & n1019;
  assign n1607 = ~\shift[1]  & n941;
  assign n1608 = ~n1606 & ~n1607;
  assign n1609 = n1605 & n1608;
  assign n1610 = n275 & ~n1609;
  assign n1611 = \shift[1]  & n1033;
  assign n1612 = \shift[1]  & n1031;
  assign n1613 = ~n1611 & ~n1612;
  assign n1614 = ~\shift[1]  & n1021;
  assign n1615 = ~\shift[1]  & n1016;
  assign n1616 = ~n1614 & ~n1615;
  assign n1617 = n1613 & n1616;
  assign n1618 = n288 & ~n1617;
  assign n1619 = ~n1610 & ~n1618;
  assign n1620 = \shift[1]  & n1039;
  assign n1621 = ~\shift[1]  & n1058;
  assign n1622 = ~n1620 & ~n1621;
  assign n1623 = \shift[1]  & n1044;
  assign n1624 = ~\shift[1]  & n1056;
  assign n1625 = ~n1623 & ~n1624;
  assign n1626 = n1622 & n1625;
  assign n1627 = n302 & ~n1626;
  assign n1628 = \shift[1]  & n1051;
  assign n1629 = ~\shift[1]  & n1026;
  assign n1630 = ~n1628 & ~n1629;
  assign n1631 = \shift[1]  & n1053;
  assign n1632 = ~\shift[1]  & n1028;
  assign n1633 = ~n1631 & ~n1632;
  assign n1634 = n1630 & n1633;
  assign n1635 = n315 & ~n1634;
  assign n1636 = ~n1627 & ~n1635;
  assign n1637 = n1619 & n1636;
  assign n1638 = n479 & ~n1637;
  assign n1639 = ~n1602 & ~n1638;
  assign n1640 = \shift[1]  & n961;
  assign n1641 = ~\shift[1]  & n1093;
  assign n1642 = ~n1640 & ~n1641;
  assign n1643 = \shift[1]  & n966;
  assign n1644 = ~\shift[1]  & n1098;
  assign n1645 = ~n1643 & ~n1644;
  assign n1646 = n1642 & n1645;
  assign n1647 = n275 & ~n1646;
  assign n1648 = \shift[1]  & n973;
  assign n1649 = ~\shift[1]  & n963;
  assign n1650 = ~n1648 & ~n1649;
  assign n1651 = \shift[1]  & n978;
  assign n1652 = ~\shift[1]  & n968;
  assign n1653 = ~n1651 & ~n1652;
  assign n1654 = n1650 & n1653;
  assign n1655 = n288 & ~n1654;
  assign n1656 = ~n1647 & ~n1655;
  assign n1657 = \shift[1]  & n986;
  assign n1658 = ~\shift[1]  & n1000;
  assign n1659 = ~n1657 & ~n1658;
  assign n1660 = \shift[1]  & n991;
  assign n1661 = ~\shift[1]  & n1005;
  assign n1662 = ~n1660 & ~n1661;
  assign n1663 = n1659 & n1662;
  assign n1664 = n302 & ~n1663;
  assign n1665 = \shift[1]  & n998;
  assign n1666 = ~\shift[1]  & n975;
  assign n1667 = ~n1665 & ~n1666;
  assign n1668 = \shift[1]  & n1003;
  assign n1669 = ~\shift[1]  & n980;
  assign n1670 = ~n1668 & ~n1669;
  assign n1671 = n1667 & n1670;
  assign n1672 = n315 & ~n1671;
  assign n1673 = ~n1664 & ~n1672;
  assign n1674 = n1656 & n1673;
  assign n1675 = n319 & ~n1674;
  assign n1676 = \shift[1]  & n1066;
  assign n1677 = ~\shift[1]  & n1041;
  assign n1678 = ~n1676 & ~n1677;
  assign n1679 = \shift[1]  & n1071;
  assign n1680 = ~\shift[1]  & n1046;
  assign n1681 = ~n1679 & ~n1680;
  assign n1682 = n1678 & n1681;
  assign n1683 = n275 & ~n1682;
  assign n1684 = \shift[1]  & n1078;
  assign n1685 = ~\shift[1]  & n1068;
  assign n1686 = ~n1684 & ~n1685;
  assign n1687 = \shift[1]  & n1083;
  assign n1688 = ~\shift[1]  & n1073;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = n1686 & n1689;
  assign n1691 = n288 & ~n1690;
  assign n1692 = ~n1683 & ~n1691;
  assign n1693 = \shift[1]  & n1091;
  assign n1694 = ~\shift[1]  & n1105;
  assign n1695 = ~n1693 & ~n1694;
  assign n1696 = \shift[1]  & n1096;
  assign n1697 = ~\shift[1]  & n1110;
  assign n1698 = ~n1696 & ~n1697;
  assign n1699 = n1695 & n1698;
  assign n1700 = n302 & ~n1699;
  assign n1701 = \shift[1]  & n1103;
  assign n1702 = ~\shift[1]  & n1080;
  assign n1703 = ~n1701 & ~n1702;
  assign n1704 = \shift[1]  & n1108;
  assign n1705 = ~\shift[1]  & n1085;
  assign n1706 = ~n1704 & ~n1705;
  assign n1707 = n1703 & n1706;
  assign n1708 = n315 & ~n1707;
  assign n1709 = ~n1700 & ~n1708;
  assign n1710 = n1692 & n1709;
  assign n1711 = n372 & ~n1710;
  assign n1712 = ~n1675 & ~n1711;
  assign n1713 = n1639 & n1712;
  assign n1714 = \shift[6]  & ~n1713;
  assign \result[3]  = n1566 | n1714;
  assign n1716 = n275 & ~n356;
  assign n1717 = ~n274 & n288;
  assign n1718 = ~n1716 & ~n1717;
  assign n1719 = n302 & ~n314;
  assign n1720 = ~n287 & n315;
  assign n1721 = ~n1719 & ~n1720;
  assign n1722 = n1718 & n1721;
  assign n1723 = n319 & ~n1722;
  assign n1724 = n275 & ~n463;
  assign n1725 = n288 & ~n331;
  assign n1726 = ~n1724 & ~n1725;
  assign n1727 = n302 & ~n368;
  assign n1728 = n315 & ~n343;
  assign n1729 = ~n1727 & ~n1728;
  assign n1730 = n1726 & n1729;
  assign n1731 = n372 & ~n1730;
  assign n1732 = ~n1723 & ~n1731;
  assign n1733 = n275 & ~n519;
  assign n1734 = n288 & ~n385;
  assign n1735 = ~n1733 & ~n1734;
  assign n1736 = n302 & ~n422;
  assign n1737 = n315 & ~n397;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = n1735 & n1738;
  assign n1740 = n426 & ~n1739;
  assign n1741 = n275 & ~n410;
  assign n1742 = n288 & ~n438;
  assign n1743 = ~n1741 & ~n1742;
  assign n1744 = n302 & ~n475;
  assign n1745 = n315 & ~n450;
  assign n1746 = ~n1744 & ~n1745;
  assign n1747 = n1743 & n1746;
  assign n1748 = n479 & ~n1747;
  assign n1749 = ~n1740 & ~n1748;
  assign n1750 = n1732 & n1749;
  assign n1751 = ~\shift[6]  & ~n1750;
  assign n1752 = n275 & ~n624;
  assign n1753 = n288 & ~n651;
  assign n1754 = ~n1752 & ~n1753;
  assign n1755 = n302 & ~n688;
  assign n1756 = n315 & ~n663;
  assign n1757 = ~n1755 & ~n1756;
  assign n1758 = n1754 & n1757;
  assign n1759 = n479 & ~n1758;
  assign n1760 = n275 & ~n301;
  assign n1761 = n288 & ~n599;
  assign n1762 = ~n1760 & ~n1761;
  assign n1763 = n302 & ~n636;
  assign n1764 = n315 & ~n611;
  assign n1765 = ~n1763 & ~n1764;
  assign n1766 = n1762 & n1765;
  assign n1767 = n426 & ~n1766;
  assign n1768 = ~n1759 & ~n1767;
  assign n1769 = n275 & ~n676;
  assign n1770 = n288 & ~n546;
  assign n1771 = ~n1769 & ~n1770;
  assign n1772 = n302 & ~n583;
  assign n1773 = n315 & ~n558;
  assign n1774 = ~n1772 & ~n1773;
  assign n1775 = n1771 & n1774;
  assign n1776 = n372 & ~n1775;
  assign n1777 = n275 & ~n571;
  assign n1778 = n288 & ~n494;
  assign n1779 = ~n1777 & ~n1778;
  assign n1780 = n302 & ~n531;
  assign n1781 = n315 & ~n506;
  assign n1782 = ~n1780 & ~n1781;
  assign n1783 = n1779 & n1782;
  assign n1784 = n319 & ~n1783;
  assign n1785 = ~n1776 & ~n1784;
  assign n1786 = n1768 & n1785;
  assign n1787 = \shift[6]  & ~n1786;
  assign \result[4]  = n1751 | n1787;
  assign n1789 = n275 & ~n784;
  assign n1790 = n288 & ~n707;
  assign n1791 = ~n1789 & ~n1790;
  assign n1792 = n302 & ~n744;
  assign n1793 = n315 & ~n719;
  assign n1794 = ~n1792 & ~n1793;
  assign n1795 = n1791 & n1794;
  assign n1796 = n319 & ~n1795;
  assign n1797 = n275 & ~n889;
  assign n1798 = n288 & ~n759;
  assign n1799 = ~n1797 & ~n1798;
  assign n1800 = n302 & ~n796;
  assign n1801 = n315 & ~n771;
  assign n1802 = ~n1800 & ~n1801;
  assign n1803 = n1799 & n1802;
  assign n1804 = n372 & ~n1803;
  assign n1805 = ~n1796 & ~n1804;
  assign n1806 = n275 & ~n996;
  assign n1807 = n288 & ~n812;
  assign n1808 = ~n1806 & ~n1807;
  assign n1809 = n302 & ~n849;
  assign n1810 = n315 & ~n824;
  assign n1811 = ~n1809 & ~n1810;
  assign n1812 = n1808 & n1811;
  assign n1813 = n426 & ~n1812;
  assign n1814 = n275 & ~n837;
  assign n1815 = n288 & ~n864;
  assign n1816 = ~n1814 & ~n1815;
  assign n1817 = n302 & ~n901;
  assign n1818 = n315 & ~n876;
  assign n1819 = ~n1817 & ~n1818;
  assign n1820 = n1816 & n1819;
  assign n1821 = n479 & ~n1820;
  assign n1822 = ~n1813 & ~n1821;
  assign n1823 = n1805 & n1822;
  assign n1824 = ~\shift[6]  & ~n1823;
  assign n1825 = n275 & ~n944;
  assign n1826 = n288 & ~n1024;
  assign n1827 = ~n1825 & ~n1826;
  assign n1828 = n302 & ~n1061;
  assign n1829 = n315 & ~n1036;
  assign n1830 = ~n1828 & ~n1829;
  assign n1831 = n1827 & n1830;
  assign n1832 = n479 & ~n1831;
  assign n1833 = n275 & ~n732;
  assign n1834 = n288 & ~n919;
  assign n1835 = ~n1833 & ~n1834;
  assign n1836 = n302 & ~n956;
  assign n1837 = n315 & ~n931;
  assign n1838 = ~n1836 & ~n1837;
  assign n1839 = n1835 & n1838;
  assign n1840 = n426 & ~n1839;
  assign n1841 = ~n1832 & ~n1840;
  assign n1842 = n275 & ~n1049;
  assign n1843 = n288 & ~n1076;
  assign n1844 = ~n1842 & ~n1843;
  assign n1845 = n302 & ~n1113;
  assign n1846 = n315 & ~n1088;
  assign n1847 = ~n1845 & ~n1846;
  assign n1848 = n1844 & n1847;
  assign n1849 = n372 & ~n1848;
  assign n1850 = n275 & ~n1101;
  assign n1851 = n288 & ~n971;
  assign n1852 = ~n1850 & ~n1851;
  assign n1853 = n302 & ~n1008;
  assign n1854 = n315 & ~n983;
  assign n1855 = ~n1853 & ~n1854;
  assign n1856 = n1852 & n1855;
  assign n1857 = n319 & ~n1856;
  assign n1858 = ~n1849 & ~n1857;
  assign n1859 = n1841 & n1858;
  assign n1860 = \shift[6]  & ~n1859;
  assign \result[5]  = n1824 | n1860;
  assign n1862 = n275 & ~n1181;
  assign n1863 = n288 & ~n1128;
  assign n1864 = ~n1862 & ~n1863;
  assign n1865 = n302 & ~n1153;
  assign n1866 = n315 & ~n1136;
  assign n1867 = ~n1865 & ~n1866;
  assign n1868 = n1864 & n1867;
  assign n1869 = n319 & ~n1868;
  assign n1870 = n275 & ~n1254;
  assign n1871 = n288 & ~n1164;
  assign n1872 = ~n1870 & ~n1871;
  assign n1873 = n302 & ~n1189;
  assign n1874 = n315 & ~n1172;
  assign n1875 = ~n1873 & ~n1874;
  assign n1876 = n1872 & n1875;
  assign n1877 = n372 & ~n1876;
  assign n1878 = ~n1869 & ~n1877;
  assign n1879 = n275 & ~n1329;
  assign n1880 = n288 & ~n1201;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = n302 & ~n1226;
  assign n1883 = n315 & ~n1209;
  assign n1884 = ~n1882 & ~n1883;
  assign n1885 = n1881 & n1884;
  assign n1886 = n426 & ~n1885;
  assign n1887 = n275 & ~n1218;
  assign n1888 = n288 & ~n1237;
  assign n1889 = ~n1887 & ~n1888;
  assign n1890 = n302 & ~n1262;
  assign n1891 = n315 & ~n1245;
  assign n1892 = ~n1890 & ~n1891;
  assign n1893 = n1889 & n1892;
  assign n1894 = n479 & ~n1893;
  assign n1895 = ~n1886 & ~n1894;
  assign n1896 = n1878 & n1895;
  assign n1897 = ~\shift[6]  & ~n1896;
  assign n1898 = n275 & ~n1293;
  assign n1899 = n288 & ~n1349;
  assign n1900 = ~n1898 & ~n1899;
  assign n1901 = n302 & ~n1374;
  assign n1902 = n315 & ~n1357;
  assign n1903 = ~n1901 & ~n1902;
  assign n1904 = n1900 & n1903;
  assign n1905 = n479 & ~n1904;
  assign n1906 = n275 & ~n1145;
  assign n1907 = n288 & ~n1276;
  assign n1908 = ~n1906 & ~n1907;
  assign n1909 = n302 & ~n1301;
  assign n1910 = n315 & ~n1284;
  assign n1911 = ~n1909 & ~n1910;
  assign n1912 = n1908 & n1911;
  assign n1913 = n426 & ~n1912;
  assign n1914 = ~n1905 & ~n1913;
  assign n1915 = n275 & ~n1366;
  assign n1916 = n288 & ~n1385;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = n302 & ~n1410;
  assign n1919 = n315 & ~n1393;
  assign n1920 = ~n1918 & ~n1919;
  assign n1921 = n1917 & n1920;
  assign n1922 = n372 & ~n1921;
  assign n1923 = n275 & ~n1402;
  assign n1924 = n288 & ~n1312;
  assign n1925 = ~n1923 & ~n1924;
  assign n1926 = n302 & ~n1337;
  assign n1927 = n315 & ~n1320;
  assign n1928 = ~n1926 & ~n1927;
  assign n1929 = n1925 & n1928;
  assign n1930 = n319 & ~n1929;
  assign n1931 = ~n1922 & ~n1930;
  assign n1932 = n1914 & n1931;
  assign n1933 = \shift[6]  & ~n1932;
  assign \result[6]  = n1897 | n1933;
  assign n1935 = n275 & ~n1478;
  assign n1936 = n288 & ~n1534;
  assign n1937 = ~n1935 & ~n1936;
  assign n1938 = n302 & ~n1559;
  assign n1939 = n315 & ~n1542;
  assign n1940 = ~n1938 & ~n1939;
  assign n1941 = n1937 & n1940;
  assign n1942 = n319 & ~n1941;
  assign n1943 = n275 & ~n1442;
  assign n1944 = n288 & ~n1461;
  assign n1945 = ~n1943 & ~n1944;
  assign n1946 = n302 & ~n1486;
  assign n1947 = n315 & ~n1469;
  assign n1948 = ~n1946 & ~n1947;
  assign n1949 = n1945 & n1948;
  assign n1950 = n372 & ~n1949;
  assign n1951 = ~n1942 & ~n1950;
  assign n1952 = n275 & ~n1663;
  assign n1953 = n288 & ~n1498;
  assign n1954 = ~n1952 & ~n1953;
  assign n1955 = n302 & ~n1523;
  assign n1956 = n315 & ~n1506;
  assign n1957 = ~n1955 & ~n1956;
  assign n1958 = n1954 & n1957;
  assign n1959 = n426 & ~n1958;
  assign n1960 = n275 & ~n1515;
  assign n1961 = n288 & ~n1425;
  assign n1962 = ~n1960 & ~n1961;
  assign n1963 = n302 & ~n1450;
  assign n1964 = n315 & ~n1433;
  assign n1965 = ~n1963 & ~n1964;
  assign n1966 = n1962 & n1965;
  assign n1967 = n479 & ~n1966;
  assign n1968 = ~n1959 & ~n1967;
  assign n1969 = n1951 & n1968;
  assign n1970 = ~\shift[6]  & ~n1969;
  assign n1971 = n288 & ~n1609;
  assign n1972 = n315 & ~n1617;
  assign n1973 = ~n1971 & ~n1972;
  assign n1974 = n302 & ~n1634;
  assign n1975 = n275 & ~n1590;
  assign n1976 = ~n1974 & ~n1975;
  assign n1977 = n1973 & n1976;
  assign n1978 = n479 & ~n1977;
  assign n1979 = n275 & ~n1551;
  assign n1980 = n288 & ~n1573;
  assign n1981 = ~n1979 & ~n1980;
  assign n1982 = n302 & ~n1598;
  assign n1983 = n315 & ~n1581;
  assign n1984 = ~n1982 & ~n1983;
  assign n1985 = n1981 & n1984;
  assign n1986 = n426 & ~n1985;
  assign n1987 = ~n1978 & ~n1986;
  assign n1988 = n275 & ~n1626;
  assign n1989 = n288 & ~n1682;
  assign n1990 = ~n1988 & ~n1989;
  assign n1991 = n302 & ~n1707;
  assign n1992 = n315 & ~n1690;
  assign n1993 = ~n1991 & ~n1992;
  assign n1994 = n1990 & n1993;
  assign n1995 = n372 & ~n1994;
  assign n1996 = n275 & ~n1699;
  assign n1997 = n288 & ~n1646;
  assign n1998 = ~n1996 & ~n1997;
  assign n1999 = n302 & ~n1671;
  assign n2000 = n315 & ~n1654;
  assign n2001 = ~n1999 & ~n2000;
  assign n2002 = n1998 & n2001;
  assign n2003 = n319 & ~n2002;
  assign n2004 = ~n1995 & ~n2003;
  assign n2005 = n1987 & n2004;
  assign n2006 = \shift[6]  & ~n2005;
  assign \result[7]  = n1970 | n2006;
  assign n2008 = n275 & ~n368;
  assign n2009 = n288 & ~n356;
  assign n2010 = ~n2008 & ~n2009;
  assign n2011 = ~n287 & n302;
  assign n2012 = ~n274 & n315;
  assign n2013 = ~n2011 & ~n2012;
  assign n2014 = n2010 & n2013;
  assign n2015 = n319 & ~n2014;
  assign n2016 = n275 & ~n475;
  assign n2017 = n288 & ~n463;
  assign n2018 = ~n2016 & ~n2017;
  assign n2019 = n302 & ~n343;
  assign n2020 = n315 & ~n331;
  assign n2021 = ~n2019 & ~n2020;
  assign n2022 = n2018 & n2021;
  assign n2023 = n372 & ~n2022;
  assign n2024 = ~n2015 & ~n2023;
  assign n2025 = n275 & ~n531;
  assign n2026 = n288 & ~n519;
  assign n2027 = ~n2025 & ~n2026;
  assign n2028 = n302 & ~n397;
  assign n2029 = n315 & ~n385;
  assign n2030 = ~n2028 & ~n2029;
  assign n2031 = n2027 & n2030;
  assign n2032 = n426 & ~n2031;
  assign n2033 = n275 & ~n422;
  assign n2034 = n288 & ~n410;
  assign n2035 = ~n2033 & ~n2034;
  assign n2036 = n302 & ~n450;
  assign n2037 = n315 & ~n438;
  assign n2038 = ~n2036 & ~n2037;
  assign n2039 = n2035 & n2038;
  assign n2040 = n479 & ~n2039;
  assign n2041 = ~n2032 & ~n2040;
  assign n2042 = n2024 & n2041;
  assign n2043 = ~\shift[6]  & ~n2042;
  assign n2044 = n275 & ~n636;
  assign n2045 = n288 & ~n624;
  assign n2046 = ~n2044 & ~n2045;
  assign n2047 = n302 & ~n663;
  assign n2048 = n315 & ~n651;
  assign n2049 = ~n2047 & ~n2048;
  assign n2050 = n2046 & n2049;
  assign n2051 = n479 & ~n2050;
  assign n2052 = n275 & ~n314;
  assign n2053 = n288 & ~n301;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055 = n302 & ~n611;
  assign n2056 = n315 & ~n599;
  assign n2057 = ~n2055 & ~n2056;
  assign n2058 = n2054 & n2057;
  assign n2059 = n426 & ~n2058;
  assign n2060 = ~n2051 & ~n2059;
  assign n2061 = n275 & ~n688;
  assign n2062 = n288 & ~n676;
  assign n2063 = ~n2061 & ~n2062;
  assign n2064 = n302 & ~n558;
  assign n2065 = n315 & ~n546;
  assign n2066 = ~n2064 & ~n2065;
  assign n2067 = n2063 & n2066;
  assign n2068 = n372 & ~n2067;
  assign n2069 = n275 & ~n583;
  assign n2070 = n288 & ~n571;
  assign n2071 = ~n2069 & ~n2070;
  assign n2072 = n302 & ~n506;
  assign n2073 = n315 & ~n494;
  assign n2074 = ~n2072 & ~n2073;
  assign n2075 = n2071 & n2074;
  assign n2076 = n319 & ~n2075;
  assign n2077 = ~n2068 & ~n2076;
  assign n2078 = n2060 & n2077;
  assign n2079 = \shift[6]  & ~n2078;
  assign \result[8]  = n2043 | n2079;
  assign n2081 = n275 & ~n796;
  assign n2082 = n288 & ~n784;
  assign n2083 = ~n2081 & ~n2082;
  assign n2084 = n302 & ~n719;
  assign n2085 = n315 & ~n707;
  assign n2086 = ~n2084 & ~n2085;
  assign n2087 = n2083 & n2086;
  assign n2088 = n319 & ~n2087;
  assign n2089 = n275 & ~n901;
  assign n2090 = n288 & ~n889;
  assign n2091 = ~n2089 & ~n2090;
  assign n2092 = n302 & ~n771;
  assign n2093 = n315 & ~n759;
  assign n2094 = ~n2092 & ~n2093;
  assign n2095 = n2091 & n2094;
  assign n2096 = n372 & ~n2095;
  assign n2097 = ~n2088 & ~n2096;
  assign n2098 = n275 & ~n1008;
  assign n2099 = n288 & ~n996;
  assign n2100 = ~n2098 & ~n2099;
  assign n2101 = n302 & ~n824;
  assign n2102 = n315 & ~n812;
  assign n2103 = ~n2101 & ~n2102;
  assign n2104 = n2100 & n2103;
  assign n2105 = n426 & ~n2104;
  assign n2106 = n275 & ~n849;
  assign n2107 = n288 & ~n837;
  assign n2108 = ~n2106 & ~n2107;
  assign n2109 = n302 & ~n876;
  assign n2110 = n315 & ~n864;
  assign n2111 = ~n2109 & ~n2110;
  assign n2112 = n2108 & n2111;
  assign n2113 = n479 & ~n2112;
  assign n2114 = ~n2105 & ~n2113;
  assign n2115 = n2097 & n2114;
  assign n2116 = ~\shift[6]  & ~n2115;
  assign n2117 = n275 & ~n956;
  assign n2118 = n288 & ~n944;
  assign n2119 = ~n2117 & ~n2118;
  assign n2120 = n302 & ~n1036;
  assign n2121 = n315 & ~n1024;
  assign n2122 = ~n2120 & ~n2121;
  assign n2123 = n2119 & n2122;
  assign n2124 = n479 & ~n2123;
  assign n2125 = n275 & ~n744;
  assign n2126 = n288 & ~n732;
  assign n2127 = ~n2125 & ~n2126;
  assign n2128 = n302 & ~n931;
  assign n2129 = n315 & ~n919;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = n2127 & n2130;
  assign n2132 = n426 & ~n2131;
  assign n2133 = ~n2124 & ~n2132;
  assign n2134 = n275 & ~n1061;
  assign n2135 = n288 & ~n1049;
  assign n2136 = ~n2134 & ~n2135;
  assign n2137 = n302 & ~n1088;
  assign n2138 = n315 & ~n1076;
  assign n2139 = ~n2137 & ~n2138;
  assign n2140 = n2136 & n2139;
  assign n2141 = n372 & ~n2140;
  assign n2142 = n275 & ~n1113;
  assign n2143 = n288 & ~n1101;
  assign n2144 = ~n2142 & ~n2143;
  assign n2145 = n302 & ~n983;
  assign n2146 = n315 & ~n971;
  assign n2147 = ~n2145 & ~n2146;
  assign n2148 = n2144 & n2147;
  assign n2149 = n319 & ~n2148;
  assign n2150 = ~n2141 & ~n2149;
  assign n2151 = n2133 & n2150;
  assign n2152 = \shift[6]  & ~n2151;
  assign \result[9]  = n2116 | n2152;
  assign n2154 = n275 & ~n1189;
  assign n2155 = n288 & ~n1181;
  assign n2156 = ~n2154 & ~n2155;
  assign n2157 = n302 & ~n1136;
  assign n2158 = n315 & ~n1128;
  assign n2159 = ~n2157 & ~n2158;
  assign n2160 = n2156 & n2159;
  assign n2161 = n319 & ~n2160;
  assign n2162 = n275 & ~n1262;
  assign n2163 = n288 & ~n1254;
  assign n2164 = ~n2162 & ~n2163;
  assign n2165 = n302 & ~n1172;
  assign n2166 = n315 & ~n1164;
  assign n2167 = ~n2165 & ~n2166;
  assign n2168 = n2164 & n2167;
  assign n2169 = n372 & ~n2168;
  assign n2170 = ~n2161 & ~n2169;
  assign n2171 = n275 & ~n1337;
  assign n2172 = n288 & ~n1329;
  assign n2173 = ~n2171 & ~n2172;
  assign n2174 = n302 & ~n1209;
  assign n2175 = n315 & ~n1201;
  assign n2176 = ~n2174 & ~n2175;
  assign n2177 = n2173 & n2176;
  assign n2178 = n426 & ~n2177;
  assign n2179 = n275 & ~n1226;
  assign n2180 = n288 & ~n1218;
  assign n2181 = ~n2179 & ~n2180;
  assign n2182 = n302 & ~n1245;
  assign n2183 = n315 & ~n1237;
  assign n2184 = ~n2182 & ~n2183;
  assign n2185 = n2181 & n2184;
  assign n2186 = n479 & ~n2185;
  assign n2187 = ~n2178 & ~n2186;
  assign n2188 = n2170 & n2187;
  assign n2189 = ~\shift[6]  & ~n2188;
  assign n2190 = n275 & ~n1301;
  assign n2191 = n288 & ~n1293;
  assign n2192 = ~n2190 & ~n2191;
  assign n2193 = n302 & ~n1357;
  assign n2194 = n315 & ~n1349;
  assign n2195 = ~n2193 & ~n2194;
  assign n2196 = n2192 & n2195;
  assign n2197 = n479 & ~n2196;
  assign n2198 = n275 & ~n1153;
  assign n2199 = n288 & ~n1145;
  assign n2200 = ~n2198 & ~n2199;
  assign n2201 = n302 & ~n1284;
  assign n2202 = n315 & ~n1276;
  assign n2203 = ~n2201 & ~n2202;
  assign n2204 = n2200 & n2203;
  assign n2205 = n426 & ~n2204;
  assign n2206 = ~n2197 & ~n2205;
  assign n2207 = n275 & ~n1374;
  assign n2208 = n288 & ~n1366;
  assign n2209 = ~n2207 & ~n2208;
  assign n2210 = n302 & ~n1393;
  assign n2211 = n315 & ~n1385;
  assign n2212 = ~n2210 & ~n2211;
  assign n2213 = n2209 & n2212;
  assign n2214 = n372 & ~n2213;
  assign n2215 = n275 & ~n1410;
  assign n2216 = n288 & ~n1402;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = n302 & ~n1320;
  assign n2219 = n315 & ~n1312;
  assign n2220 = ~n2218 & ~n2219;
  assign n2221 = n2217 & n2220;
  assign n2222 = n319 & ~n2221;
  assign n2223 = ~n2214 & ~n2222;
  assign n2224 = n2206 & n2223;
  assign n2225 = \shift[6]  & ~n2224;
  assign \result[10]  = n2189 | n2225;
  assign n2227 = n275 & ~n1486;
  assign n2228 = n288 & ~n1478;
  assign n2229 = ~n2227 & ~n2228;
  assign n2230 = n302 & ~n1542;
  assign n2231 = n315 & ~n1534;
  assign n2232 = ~n2230 & ~n2231;
  assign n2233 = n2229 & n2232;
  assign n2234 = n319 & ~n2233;
  assign n2235 = n275 & ~n1450;
  assign n2236 = n288 & ~n1442;
  assign n2237 = ~n2235 & ~n2236;
  assign n2238 = n302 & ~n1469;
  assign n2239 = n315 & ~n1461;
  assign n2240 = ~n2238 & ~n2239;
  assign n2241 = n2237 & n2240;
  assign n2242 = n372 & ~n2241;
  assign n2243 = ~n2234 & ~n2242;
  assign n2244 = n275 & ~n1671;
  assign n2245 = n288 & ~n1663;
  assign n2246 = ~n2244 & ~n2245;
  assign n2247 = n302 & ~n1506;
  assign n2248 = n315 & ~n1498;
  assign n2249 = ~n2247 & ~n2248;
  assign n2250 = n2246 & n2249;
  assign n2251 = n426 & ~n2250;
  assign n2252 = n275 & ~n1523;
  assign n2253 = n288 & ~n1515;
  assign n2254 = ~n2252 & ~n2253;
  assign n2255 = n302 & ~n1433;
  assign n2256 = n315 & ~n1425;
  assign n2257 = ~n2255 & ~n2256;
  assign n2258 = n2254 & n2257;
  assign n2259 = n479 & ~n2258;
  assign n2260 = ~n2251 & ~n2259;
  assign n2261 = n2243 & n2260;
  assign n2262 = ~\shift[6]  & ~n2261;
  assign n2263 = n275 & ~n1598;
  assign n2264 = n315 & ~n1609;
  assign n2265 = ~n2263 & ~n2264;
  assign n2266 = n302 & ~n1617;
  assign n2267 = n288 & ~n1590;
  assign n2268 = ~n2266 & ~n2267;
  assign n2269 = n2265 & n2268;
  assign n2270 = n479 & ~n2269;
  assign n2271 = n275 & ~n1559;
  assign n2272 = n288 & ~n1551;
  assign n2273 = ~n2271 & ~n2272;
  assign n2274 = n302 & ~n1581;
  assign n2275 = n315 & ~n1573;
  assign n2276 = ~n2274 & ~n2275;
  assign n2277 = n2273 & n2276;
  assign n2278 = n426 & ~n2277;
  assign n2279 = ~n2270 & ~n2278;
  assign n2280 = n275 & ~n1634;
  assign n2281 = n288 & ~n1626;
  assign n2282 = ~n2280 & ~n2281;
  assign n2283 = n302 & ~n1690;
  assign n2284 = n315 & ~n1682;
  assign n2285 = ~n2283 & ~n2284;
  assign n2286 = n2282 & n2285;
  assign n2287 = n372 & ~n2286;
  assign n2288 = n275 & ~n1707;
  assign n2289 = n288 & ~n1699;
  assign n2290 = ~n2288 & ~n2289;
  assign n2291 = n302 & ~n1654;
  assign n2292 = n315 & ~n1646;
  assign n2293 = ~n2291 & ~n2292;
  assign n2294 = n2290 & n2293;
  assign n2295 = n319 & ~n2294;
  assign n2296 = ~n2287 & ~n2295;
  assign n2297 = n2279 & n2296;
  assign n2298 = \shift[6]  & ~n2297;
  assign \result[11]  = n2262 | n2298;
  assign n2300 = n275 & ~n343;
  assign n2301 = n288 & ~n368;
  assign n2302 = ~n2300 & ~n2301;
  assign n2303 = ~n274 & n302;
  assign n2304 = n315 & ~n356;
  assign n2305 = ~n2303 & ~n2304;
  assign n2306 = n2302 & n2305;
  assign n2307 = n319 & ~n2306;
  assign n2308 = n275 & ~n450;
  assign n2309 = n288 & ~n475;
  assign n2310 = ~n2308 & ~n2309;
  assign n2311 = n302 & ~n331;
  assign n2312 = n315 & ~n463;
  assign n2313 = ~n2311 & ~n2312;
  assign n2314 = n2310 & n2313;
  assign n2315 = n372 & ~n2314;
  assign n2316 = ~n2307 & ~n2315;
  assign n2317 = n275 & ~n506;
  assign n2318 = n288 & ~n531;
  assign n2319 = ~n2317 & ~n2318;
  assign n2320 = n302 & ~n385;
  assign n2321 = n315 & ~n519;
  assign n2322 = ~n2320 & ~n2321;
  assign n2323 = n2319 & n2322;
  assign n2324 = n426 & ~n2323;
  assign n2325 = n275 & ~n397;
  assign n2326 = n288 & ~n422;
  assign n2327 = ~n2325 & ~n2326;
  assign n2328 = n302 & ~n438;
  assign n2329 = n315 & ~n410;
  assign n2330 = ~n2328 & ~n2329;
  assign n2331 = n2327 & n2330;
  assign n2332 = n479 & ~n2331;
  assign n2333 = ~n2324 & ~n2332;
  assign n2334 = n2316 & n2333;
  assign n2335 = ~\shift[6]  & ~n2334;
  assign n2336 = n275 & ~n611;
  assign n2337 = n288 & ~n636;
  assign n2338 = ~n2336 & ~n2337;
  assign n2339 = n302 & ~n651;
  assign n2340 = n315 & ~n624;
  assign n2341 = ~n2339 & ~n2340;
  assign n2342 = n2338 & n2341;
  assign n2343 = n479 & ~n2342;
  assign n2344 = n275 & ~n287;
  assign n2345 = n288 & ~n314;
  assign n2346 = ~n2344 & ~n2345;
  assign n2347 = n302 & ~n599;
  assign n2348 = ~n301 & n315;
  assign n2349 = ~n2347 & ~n2348;
  assign n2350 = n2346 & n2349;
  assign n2351 = n426 & ~n2350;
  assign n2352 = ~n2343 & ~n2351;
  assign n2353 = n275 & ~n663;
  assign n2354 = n288 & ~n688;
  assign n2355 = ~n2353 & ~n2354;
  assign n2356 = n302 & ~n546;
  assign n2357 = n315 & ~n676;
  assign n2358 = ~n2356 & ~n2357;
  assign n2359 = n2355 & n2358;
  assign n2360 = n372 & ~n2359;
  assign n2361 = n275 & ~n558;
  assign n2362 = n288 & ~n583;
  assign n2363 = ~n2361 & ~n2362;
  assign n2364 = n302 & ~n494;
  assign n2365 = n315 & ~n571;
  assign n2366 = ~n2364 & ~n2365;
  assign n2367 = n2363 & n2366;
  assign n2368 = n319 & ~n2367;
  assign n2369 = ~n2360 & ~n2368;
  assign n2370 = n2352 & n2369;
  assign n2371 = \shift[6]  & ~n2370;
  assign \result[12]  = n2335 | n2371;
  assign n2373 = n275 & ~n771;
  assign n2374 = n288 & ~n796;
  assign n2375 = ~n2373 & ~n2374;
  assign n2376 = n302 & ~n707;
  assign n2377 = n315 & ~n784;
  assign n2378 = ~n2376 & ~n2377;
  assign n2379 = n2375 & n2378;
  assign n2380 = n319 & ~n2379;
  assign n2381 = n275 & ~n876;
  assign n2382 = n288 & ~n901;
  assign n2383 = ~n2381 & ~n2382;
  assign n2384 = n302 & ~n759;
  assign n2385 = n315 & ~n889;
  assign n2386 = ~n2384 & ~n2385;
  assign n2387 = n2383 & n2386;
  assign n2388 = n372 & ~n2387;
  assign n2389 = ~n2380 & ~n2388;
  assign n2390 = n275 & ~n983;
  assign n2391 = n288 & ~n1008;
  assign n2392 = ~n2390 & ~n2391;
  assign n2393 = n302 & ~n812;
  assign n2394 = n315 & ~n996;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = n2392 & n2395;
  assign n2397 = n426 & ~n2396;
  assign n2398 = n275 & ~n824;
  assign n2399 = n288 & ~n849;
  assign n2400 = ~n2398 & ~n2399;
  assign n2401 = n302 & ~n864;
  assign n2402 = n315 & ~n837;
  assign n2403 = ~n2401 & ~n2402;
  assign n2404 = n2400 & n2403;
  assign n2405 = n479 & ~n2404;
  assign n2406 = ~n2397 & ~n2405;
  assign n2407 = n2389 & n2406;
  assign n2408 = ~\shift[6]  & ~n2407;
  assign n2409 = n275 & ~n931;
  assign n2410 = n288 & ~n956;
  assign n2411 = ~n2409 & ~n2410;
  assign n2412 = n302 & ~n1024;
  assign n2413 = n315 & ~n944;
  assign n2414 = ~n2412 & ~n2413;
  assign n2415 = n2411 & n2414;
  assign n2416 = n479 & ~n2415;
  assign n2417 = n275 & ~n719;
  assign n2418 = n288 & ~n744;
  assign n2419 = ~n2417 & ~n2418;
  assign n2420 = n302 & ~n919;
  assign n2421 = n315 & ~n732;
  assign n2422 = ~n2420 & ~n2421;
  assign n2423 = n2419 & n2422;
  assign n2424 = n426 & ~n2423;
  assign n2425 = ~n2416 & ~n2424;
  assign n2426 = n275 & ~n1036;
  assign n2427 = n288 & ~n1061;
  assign n2428 = ~n2426 & ~n2427;
  assign n2429 = n302 & ~n1076;
  assign n2430 = n315 & ~n1049;
  assign n2431 = ~n2429 & ~n2430;
  assign n2432 = n2428 & n2431;
  assign n2433 = n372 & ~n2432;
  assign n2434 = n275 & ~n1088;
  assign n2435 = n288 & ~n1113;
  assign n2436 = ~n2434 & ~n2435;
  assign n2437 = n302 & ~n971;
  assign n2438 = n315 & ~n1101;
  assign n2439 = ~n2437 & ~n2438;
  assign n2440 = n2436 & n2439;
  assign n2441 = n319 & ~n2440;
  assign n2442 = ~n2433 & ~n2441;
  assign n2443 = n2425 & n2442;
  assign n2444 = \shift[6]  & ~n2443;
  assign \result[13]  = n2408 | n2444;
  assign n2446 = n275 & ~n1172;
  assign n2447 = n288 & ~n1189;
  assign n2448 = ~n2446 & ~n2447;
  assign n2449 = n302 & ~n1128;
  assign n2450 = n315 & ~n1181;
  assign n2451 = ~n2449 & ~n2450;
  assign n2452 = n2448 & n2451;
  assign n2453 = n319 & ~n2452;
  assign n2454 = n275 & ~n1245;
  assign n2455 = n288 & ~n1262;
  assign n2456 = ~n2454 & ~n2455;
  assign n2457 = n302 & ~n1164;
  assign n2458 = n315 & ~n1254;
  assign n2459 = ~n2457 & ~n2458;
  assign n2460 = n2456 & n2459;
  assign n2461 = n372 & ~n2460;
  assign n2462 = ~n2453 & ~n2461;
  assign n2463 = n275 & ~n1320;
  assign n2464 = n288 & ~n1337;
  assign n2465 = ~n2463 & ~n2464;
  assign n2466 = n302 & ~n1201;
  assign n2467 = n315 & ~n1329;
  assign n2468 = ~n2466 & ~n2467;
  assign n2469 = n2465 & n2468;
  assign n2470 = n426 & ~n2469;
  assign n2471 = n275 & ~n1209;
  assign n2472 = n288 & ~n1226;
  assign n2473 = ~n2471 & ~n2472;
  assign n2474 = n302 & ~n1237;
  assign n2475 = n315 & ~n1218;
  assign n2476 = ~n2474 & ~n2475;
  assign n2477 = n2473 & n2476;
  assign n2478 = n479 & ~n2477;
  assign n2479 = ~n2470 & ~n2478;
  assign n2480 = n2462 & n2479;
  assign n2481 = ~\shift[6]  & ~n2480;
  assign n2482 = n275 & ~n1284;
  assign n2483 = n288 & ~n1301;
  assign n2484 = ~n2482 & ~n2483;
  assign n2485 = n302 & ~n1349;
  assign n2486 = n315 & ~n1293;
  assign n2487 = ~n2485 & ~n2486;
  assign n2488 = n2484 & n2487;
  assign n2489 = n479 & ~n2488;
  assign n2490 = n275 & ~n1136;
  assign n2491 = n288 & ~n1153;
  assign n2492 = ~n2490 & ~n2491;
  assign n2493 = n302 & ~n1276;
  assign n2494 = n315 & ~n1145;
  assign n2495 = ~n2493 & ~n2494;
  assign n2496 = n2492 & n2495;
  assign n2497 = n426 & ~n2496;
  assign n2498 = ~n2489 & ~n2497;
  assign n2499 = n275 & ~n1357;
  assign n2500 = n288 & ~n1374;
  assign n2501 = ~n2499 & ~n2500;
  assign n2502 = n302 & ~n1385;
  assign n2503 = n315 & ~n1366;
  assign n2504 = ~n2502 & ~n2503;
  assign n2505 = n2501 & n2504;
  assign n2506 = n372 & ~n2505;
  assign n2507 = n275 & ~n1393;
  assign n2508 = n288 & ~n1410;
  assign n2509 = ~n2507 & ~n2508;
  assign n2510 = n302 & ~n1312;
  assign n2511 = n315 & ~n1402;
  assign n2512 = ~n2510 & ~n2511;
  assign n2513 = n2509 & n2512;
  assign n2514 = n319 & ~n2513;
  assign n2515 = ~n2506 & ~n2514;
  assign n2516 = n2498 & n2515;
  assign n2517 = \shift[6]  & ~n2516;
  assign \result[14]  = n2481 | n2517;
  assign n2519 = n275 & ~n1469;
  assign n2520 = n288 & ~n1486;
  assign n2521 = ~n2519 & ~n2520;
  assign n2522 = n302 & ~n1534;
  assign n2523 = n315 & ~n1478;
  assign n2524 = ~n2522 & ~n2523;
  assign n2525 = n2521 & n2524;
  assign n2526 = n319 & ~n2525;
  assign n2527 = n275 & ~n1433;
  assign n2528 = n288 & ~n1450;
  assign n2529 = ~n2527 & ~n2528;
  assign n2530 = n302 & ~n1461;
  assign n2531 = n315 & ~n1442;
  assign n2532 = ~n2530 & ~n2531;
  assign n2533 = n2529 & n2532;
  assign n2534 = n372 & ~n2533;
  assign n2535 = ~n2526 & ~n2534;
  assign n2536 = n275 & ~n1654;
  assign n2537 = n288 & ~n1671;
  assign n2538 = ~n2536 & ~n2537;
  assign n2539 = n302 & ~n1498;
  assign n2540 = n315 & ~n1663;
  assign n2541 = ~n2539 & ~n2540;
  assign n2542 = n2538 & n2541;
  assign n2543 = n426 & ~n2542;
  assign n2544 = n275 & ~n1506;
  assign n2545 = n288 & ~n1523;
  assign n2546 = ~n2544 & ~n2545;
  assign n2547 = n302 & ~n1425;
  assign n2548 = n315 & ~n1515;
  assign n2549 = ~n2547 & ~n2548;
  assign n2550 = n2546 & n2549;
  assign n2551 = n479 & ~n2550;
  assign n2552 = ~n2543 & ~n2551;
  assign n2553 = n2535 & n2552;
  assign n2554 = ~\shift[6]  & ~n2553;
  assign n2555 = n275 & ~n1581;
  assign n2556 = n288 & ~n1598;
  assign n2557 = ~n2555 & ~n2556;
  assign n2558 = n302 & ~n1609;
  assign n2559 = n315 & ~n1590;
  assign n2560 = ~n2558 & ~n2559;
  assign n2561 = n2557 & n2560;
  assign n2562 = n479 & ~n2561;
  assign n2563 = n275 & ~n1542;
  assign n2564 = n288 & ~n1559;
  assign n2565 = ~n2563 & ~n2564;
  assign n2566 = n302 & ~n1573;
  assign n2567 = n315 & ~n1551;
  assign n2568 = ~n2566 & ~n2567;
  assign n2569 = n2565 & n2568;
  assign n2570 = n426 & ~n2569;
  assign n2571 = ~n2562 & ~n2570;
  assign n2572 = n275 & ~n1617;
  assign n2573 = n288 & ~n1634;
  assign n2574 = ~n2572 & ~n2573;
  assign n2575 = n302 & ~n1682;
  assign n2576 = n315 & ~n1626;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = n2574 & n2577;
  assign n2579 = n372 & ~n2578;
  assign n2580 = n275 & ~n1690;
  assign n2581 = n288 & ~n1707;
  assign n2582 = ~n2580 & ~n2581;
  assign n2583 = n302 & ~n1646;
  assign n2584 = n315 & ~n1699;
  assign n2585 = ~n2583 & ~n2584;
  assign n2586 = n2582 & n2585;
  assign n2587 = n319 & ~n2586;
  assign n2588 = ~n2579 & ~n2587;
  assign n2589 = n2571 & n2588;
  assign n2590 = \shift[6]  & ~n2589;
  assign \result[15]  = n2554 | n2590;
  assign n2592 = n319 & ~n371;
  assign n2593 = n372 & ~n478;
  assign n2594 = ~n2592 & ~n2593;
  assign n2595 = n426 & ~n534;
  assign n2596 = ~n425 & n479;
  assign n2597 = ~n2595 & ~n2596;
  assign n2598 = n2594 & n2597;
  assign n2599 = ~\shift[6]  & ~n2598;
  assign n2600 = ~n318 & n426;
  assign n2601 = n319 & ~n586;
  assign n2602 = ~n2600 & ~n2601;
  assign n2603 = n479 & ~n639;
  assign n2604 = n372 & ~n691;
  assign n2605 = ~n2603 & ~n2604;
  assign n2606 = n2602 & n2605;
  assign n2607 = \shift[6]  & ~n2606;
  assign \result[16]  = n2599 | n2607;
  assign n2609 = n319 & ~n799;
  assign n2610 = n372 & ~n904;
  assign n2611 = ~n2609 & ~n2610;
  assign n2612 = n426 & ~n1011;
  assign n2613 = n479 & ~n852;
  assign n2614 = ~n2612 & ~n2613;
  assign n2615 = n2611 & n2614;
  assign n2616 = ~\shift[6]  & ~n2615;
  assign n2617 = n479 & ~n959;
  assign n2618 = n426 & ~n747;
  assign n2619 = ~n2617 & ~n2618;
  assign n2620 = n372 & ~n1064;
  assign n2621 = n319 & ~n1116;
  assign n2622 = ~n2620 & ~n2621;
  assign n2623 = n2619 & n2622;
  assign n2624 = \shift[6]  & ~n2623;
  assign \result[17]  = n2616 | n2624;
  assign n2626 = n319 & ~n1192;
  assign n2627 = n372 & ~n1265;
  assign n2628 = ~n2626 & ~n2627;
  assign n2629 = n426 & ~n1340;
  assign n2630 = n479 & ~n1229;
  assign n2631 = ~n2629 & ~n2630;
  assign n2632 = n2628 & n2631;
  assign n2633 = ~\shift[6]  & ~n2632;
  assign n2634 = n479 & ~n1304;
  assign n2635 = n426 & ~n1156;
  assign n2636 = ~n2634 & ~n2635;
  assign n2637 = n372 & ~n1377;
  assign n2638 = n319 & ~n1413;
  assign n2639 = ~n2637 & ~n2638;
  assign n2640 = n2636 & n2639;
  assign n2641 = \shift[6]  & ~n2640;
  assign \result[18]  = n2633 | n2641;
  assign n2643 = n372 & ~n1453;
  assign n2644 = n319 & ~n1489;
  assign n2645 = ~n2643 & ~n2644;
  assign n2646 = n479 & ~n1526;
  assign n2647 = n426 & ~n1674;
  assign n2648 = ~n2646 & ~n2647;
  assign n2649 = n2645 & n2648;
  assign n2650 = ~\shift[6]  & ~n2649;
  assign n2651 = n479 & ~n1601;
  assign n2652 = n426 & ~n1562;
  assign n2653 = ~n2651 & ~n2652;
  assign n2654 = n319 & ~n1710;
  assign n2655 = n372 & ~n1637;
  assign n2656 = ~n2654 & ~n2655;
  assign n2657 = n2653 & n2656;
  assign n2658 = \shift[6]  & ~n2657;
  assign \result[19]  = n2650 | n2658;
  assign n2660 = n319 & ~n1730;
  assign n2661 = n372 & ~n1747;
  assign n2662 = ~n2660 & ~n2661;
  assign n2663 = n426 & ~n1783;
  assign n2664 = n479 & ~n1739;
  assign n2665 = ~n2663 & ~n2664;
  assign n2666 = n2662 & n2665;
  assign n2667 = ~\shift[6]  & ~n2666;
  assign n2668 = n426 & ~n1722;
  assign n2669 = n372 & ~n1758;
  assign n2670 = ~n2668 & ~n2669;
  assign n2671 = n319 & ~n1775;
  assign n2672 = n479 & ~n1766;
  assign n2673 = ~n2671 & ~n2672;
  assign n2674 = n2670 & n2673;
  assign n2675 = \shift[6]  & ~n2674;
  assign \result[20]  = n2667 | n2675;
  assign n2677 = n319 & ~n1803;
  assign n2678 = n372 & ~n1820;
  assign n2679 = ~n2677 & ~n2678;
  assign n2680 = n426 & ~n1856;
  assign n2681 = n479 & ~n1812;
  assign n2682 = ~n2680 & ~n2681;
  assign n2683 = n2679 & n2682;
  assign n2684 = ~\shift[6]  & ~n2683;
  assign n2685 = n426 & ~n1795;
  assign n2686 = n372 & ~n1831;
  assign n2687 = ~n2685 & ~n2686;
  assign n2688 = n319 & ~n1848;
  assign n2689 = n479 & ~n1839;
  assign n2690 = ~n2688 & ~n2689;
  assign n2691 = n2687 & n2690;
  assign n2692 = \shift[6]  & ~n2691;
  assign \result[21]  = n2684 | n2692;
  assign n2694 = n319 & ~n1876;
  assign n2695 = n372 & ~n1893;
  assign n2696 = ~n2694 & ~n2695;
  assign n2697 = n426 & ~n1929;
  assign n2698 = n479 & ~n1885;
  assign n2699 = ~n2697 & ~n2698;
  assign n2700 = n2696 & n2699;
  assign n2701 = ~\shift[6]  & ~n2700;
  assign n2702 = n426 & ~n1868;
  assign n2703 = n372 & ~n1904;
  assign n2704 = ~n2702 & ~n2703;
  assign n2705 = n319 & ~n1921;
  assign n2706 = n479 & ~n1912;
  assign n2707 = ~n2705 & ~n2706;
  assign n2708 = n2704 & n2707;
  assign n2709 = \shift[6]  & ~n2708;
  assign \result[22]  = n2701 | n2709;
  assign n2711 = n319 & ~n1949;
  assign n2712 = n426 & ~n2002;
  assign n2713 = ~n2711 & ~n2712;
  assign n2714 = n479 & ~n1958;
  assign n2715 = n372 & ~n1966;
  assign n2716 = ~n2714 & ~n2715;
  assign n2717 = n2713 & n2716;
  assign n2718 = ~\shift[6]  & ~n2717;
  assign n2719 = n372 & ~n1977;
  assign n2720 = n479 & ~n1985;
  assign n2721 = ~n2719 & ~n2720;
  assign n2722 = n319 & ~n1994;
  assign n2723 = n426 & ~n1941;
  assign n2724 = ~n2722 & ~n2723;
  assign n2725 = n2721 & n2724;
  assign n2726 = \shift[6]  & ~n2725;
  assign \result[23]  = n2718 | n2726;
  assign n2728 = n319 & ~n2022;
  assign n2729 = n426 & ~n2075;
  assign n2730 = ~n2728 & ~n2729;
  assign n2731 = n479 & ~n2031;
  assign n2732 = n372 & ~n2039;
  assign n2733 = ~n2731 & ~n2732;
  assign n2734 = n2730 & n2733;
  assign n2735 = ~\shift[6]  & ~n2734;
  assign n2736 = n372 & ~n2050;
  assign n2737 = n479 & ~n2058;
  assign n2738 = ~n2736 & ~n2737;
  assign n2739 = n319 & ~n2067;
  assign n2740 = n426 & ~n2014;
  assign n2741 = ~n2739 & ~n2740;
  assign n2742 = n2738 & n2741;
  assign n2743 = \shift[6]  & ~n2742;
  assign \result[24]  = n2735 | n2743;
  assign n2745 = n319 & ~n2095;
  assign n2746 = n426 & ~n2148;
  assign n2747 = ~n2745 & ~n2746;
  assign n2748 = n479 & ~n2104;
  assign n2749 = n372 & ~n2112;
  assign n2750 = ~n2748 & ~n2749;
  assign n2751 = n2747 & n2750;
  assign n2752 = ~\shift[6]  & ~n2751;
  assign n2753 = n372 & ~n2123;
  assign n2754 = n479 & ~n2131;
  assign n2755 = ~n2753 & ~n2754;
  assign n2756 = n319 & ~n2140;
  assign n2757 = n426 & ~n2087;
  assign n2758 = ~n2756 & ~n2757;
  assign n2759 = n2755 & n2758;
  assign n2760 = \shift[6]  & ~n2759;
  assign \result[25]  = n2752 | n2760;
  assign n2762 = n319 & ~n2168;
  assign n2763 = n372 & ~n2185;
  assign n2764 = ~n2762 & ~n2763;
  assign n2765 = n426 & ~n2221;
  assign n2766 = n479 & ~n2177;
  assign n2767 = ~n2765 & ~n2766;
  assign n2768 = n2764 & n2767;
  assign n2769 = ~\shift[6]  & ~n2768;
  assign n2770 = n372 & ~n2196;
  assign n2771 = n479 & ~n2204;
  assign n2772 = ~n2770 & ~n2771;
  assign n2773 = n319 & ~n2213;
  assign n2774 = n426 & ~n2160;
  assign n2775 = ~n2773 & ~n2774;
  assign n2776 = n2772 & n2775;
  assign n2777 = \shift[6]  & ~n2776;
  assign \result[26]  = n2769 | n2777;
  assign n2779 = n319 & ~n2241;
  assign n2780 = n372 & ~n2258;
  assign n2781 = ~n2779 & ~n2780;
  assign n2782 = n426 & ~n2294;
  assign n2783 = n479 & ~n2250;
  assign n2784 = ~n2782 & ~n2783;
  assign n2785 = n2781 & n2784;
  assign n2786 = ~\shift[6]  & ~n2785;
  assign n2787 = n372 & ~n2269;
  assign n2788 = n479 & ~n2277;
  assign n2789 = ~n2787 & ~n2788;
  assign n2790 = n319 & ~n2286;
  assign n2791 = n426 & ~n2233;
  assign n2792 = ~n2790 & ~n2791;
  assign n2793 = n2789 & n2792;
  assign n2794 = \shift[6]  & ~n2793;
  assign \result[27]  = n2786 | n2794;
  assign n2796 = n319 & ~n2314;
  assign n2797 = n372 & ~n2331;
  assign n2798 = ~n2796 & ~n2797;
  assign n2799 = n426 & ~n2367;
  assign n2800 = n479 & ~n2323;
  assign n2801 = ~n2799 & ~n2800;
  assign n2802 = n2798 & n2801;
  assign n2803 = ~\shift[6]  & ~n2802;
  assign n2804 = n372 & ~n2342;
  assign n2805 = n479 & ~n2350;
  assign n2806 = ~n2804 & ~n2805;
  assign n2807 = n319 & ~n2359;
  assign n2808 = n426 & ~n2306;
  assign n2809 = ~n2807 & ~n2808;
  assign n2810 = n2806 & n2809;
  assign n2811 = \shift[6]  & ~n2810;
  assign \result[28]  = n2803 | n2811;
  assign n2813 = n319 & ~n2387;
  assign n2814 = n372 & ~n2404;
  assign n2815 = ~n2813 & ~n2814;
  assign n2816 = n426 & ~n2440;
  assign n2817 = n479 & ~n2396;
  assign n2818 = ~n2816 & ~n2817;
  assign n2819 = n2815 & n2818;
  assign n2820 = ~\shift[6]  & ~n2819;
  assign n2821 = n372 & ~n2415;
  assign n2822 = n479 & ~n2423;
  assign n2823 = ~n2821 & ~n2822;
  assign n2824 = n319 & ~n2432;
  assign n2825 = n426 & ~n2379;
  assign n2826 = ~n2824 & ~n2825;
  assign n2827 = n2823 & n2826;
  assign n2828 = \shift[6]  & ~n2827;
  assign \result[29]  = n2820 | n2828;
  assign n2830 = n319 & ~n2460;
  assign n2831 = n372 & ~n2477;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = n426 & ~n2513;
  assign n2834 = n479 & ~n2469;
  assign n2835 = ~n2833 & ~n2834;
  assign n2836 = n2832 & n2835;
  assign n2837 = ~\shift[6]  & ~n2836;
  assign n2838 = n372 & ~n2488;
  assign n2839 = n479 & ~n2496;
  assign n2840 = ~n2838 & ~n2839;
  assign n2841 = n319 & ~n2505;
  assign n2842 = n426 & ~n2452;
  assign n2843 = ~n2841 & ~n2842;
  assign n2844 = n2840 & n2843;
  assign n2845 = \shift[6]  & ~n2844;
  assign \result[30]  = n2837 | n2845;
  assign n2847 = n319 & ~n2533;
  assign n2848 = n372 & ~n2550;
  assign n2849 = ~n2847 & ~n2848;
  assign n2850 = n426 & ~n2586;
  assign n2851 = n479 & ~n2542;
  assign n2852 = ~n2850 & ~n2851;
  assign n2853 = n2849 & n2852;
  assign n2854 = ~\shift[6]  & ~n2853;
  assign n2855 = n372 & ~n2561;
  assign n2856 = n479 & ~n2569;
  assign n2857 = ~n2855 & ~n2856;
  assign n2858 = n319 & ~n2578;
  assign n2859 = n426 & ~n2525;
  assign n2860 = ~n2858 & ~n2859;
  assign n2861 = n2857 & n2860;
  assign n2862 = \shift[6]  & ~n2861;
  assign \result[31]  = n2854 | n2862;
  assign n2864 = n319 & ~n478;
  assign n2865 = n372 & ~n425;
  assign n2866 = ~n2864 & ~n2865;
  assign n2867 = n426 & ~n586;
  assign n2868 = n479 & ~n534;
  assign n2869 = ~n2867 & ~n2868;
  assign n2870 = n2866 & n2869;
  assign n2871 = ~\shift[6]  & ~n2870;
  assign n2872 = ~n318 & n479;
  assign n2873 = ~n371 & n426;
  assign n2874 = ~n2872 & ~n2873;
  assign n2875 = n372 & ~n639;
  assign n2876 = n319 & ~n691;
  assign n2877 = ~n2875 & ~n2876;
  assign n2878 = n2874 & n2877;
  assign n2879 = \shift[6]  & ~n2878;
  assign \result[32]  = n2871 | n2879;
  assign n2881 = n319 & ~n904;
  assign n2882 = n372 & ~n852;
  assign n2883 = ~n2881 & ~n2882;
  assign n2884 = n426 & ~n1116;
  assign n2885 = n479 & ~n1011;
  assign n2886 = ~n2884 & ~n2885;
  assign n2887 = n2883 & n2886;
  assign n2888 = ~\shift[6]  & ~n2887;
  assign n2889 = n372 & ~n959;
  assign n2890 = n479 & ~n747;
  assign n2891 = ~n2889 & ~n2890;
  assign n2892 = n319 & ~n1064;
  assign n2893 = n426 & ~n799;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895 = n2891 & n2894;
  assign n2896 = \shift[6]  & ~n2895;
  assign \result[33]  = n2888 | n2896;
  assign n2898 = n319 & ~n1265;
  assign n2899 = n372 & ~n1229;
  assign n2900 = ~n2898 & ~n2899;
  assign n2901 = n426 & ~n1413;
  assign n2902 = n479 & ~n1340;
  assign n2903 = ~n2901 & ~n2902;
  assign n2904 = n2900 & n2903;
  assign n2905 = ~\shift[6]  & ~n2904;
  assign n2906 = n372 & ~n1304;
  assign n2907 = n479 & ~n1156;
  assign n2908 = ~n2906 & ~n2907;
  assign n2909 = n319 & ~n1377;
  assign n2910 = n426 & ~n1192;
  assign n2911 = ~n2909 & ~n2910;
  assign n2912 = n2908 & n2911;
  assign n2913 = \shift[6]  & ~n2912;
  assign \result[34]  = n2905 | n2913;
  assign n2915 = n319 & ~n1453;
  assign n2916 = n426 & ~n1710;
  assign n2917 = ~n2915 & ~n2916;
  assign n2918 = n372 & ~n1526;
  assign n2919 = n479 & ~n1674;
  assign n2920 = ~n2918 & ~n2919;
  assign n2921 = n2917 & n2920;
  assign n2922 = ~\shift[6]  & ~n2921;
  assign n2923 = n372 & ~n1601;
  assign n2924 = n426 & ~n1489;
  assign n2925 = ~n2923 & ~n2924;
  assign n2926 = n319 & ~n1637;
  assign n2927 = n479 & ~n1562;
  assign n2928 = ~n2926 & ~n2927;
  assign n2929 = n2925 & n2928;
  assign n2930 = \shift[6]  & ~n2929;
  assign \result[35]  = n2922 | n2930;
  assign n2932 = n319 & ~n1747;
  assign n2933 = n372 & ~n1739;
  assign n2934 = ~n2932 & ~n2933;
  assign n2935 = n426 & ~n1775;
  assign n2936 = n479 & ~n1783;
  assign n2937 = ~n2935 & ~n2936;
  assign n2938 = n2934 & n2937;
  assign n2939 = ~\shift[6]  & ~n2938;
  assign n2940 = n479 & ~n1722;
  assign n2941 = n426 & ~n1730;
  assign n2942 = ~n2940 & ~n2941;
  assign n2943 = n372 & ~n1766;
  assign n2944 = n319 & ~n1758;
  assign n2945 = ~n2943 & ~n2944;
  assign n2946 = n2942 & n2945;
  assign n2947 = \shift[6]  & ~n2946;
  assign \result[36]  = n2939 | n2947;
  assign n2949 = n319 & ~n1820;
  assign n2950 = n372 & ~n1812;
  assign n2951 = ~n2949 & ~n2950;
  assign n2952 = n426 & ~n1848;
  assign n2953 = n479 & ~n1856;
  assign n2954 = ~n2952 & ~n2953;
  assign n2955 = n2951 & n2954;
  assign n2956 = ~\shift[6]  & ~n2955;
  assign n2957 = n479 & ~n1795;
  assign n2958 = n426 & ~n1803;
  assign n2959 = ~n2957 & ~n2958;
  assign n2960 = n372 & ~n1839;
  assign n2961 = n319 & ~n1831;
  assign n2962 = ~n2960 & ~n2961;
  assign n2963 = n2959 & n2962;
  assign n2964 = \shift[6]  & ~n2963;
  assign \result[37]  = n2956 | n2964;
  assign n2966 = n319 & ~n1893;
  assign n2967 = n372 & ~n1885;
  assign n2968 = ~n2966 & ~n2967;
  assign n2969 = n426 & ~n1921;
  assign n2970 = n479 & ~n1929;
  assign n2971 = ~n2969 & ~n2970;
  assign n2972 = n2968 & n2971;
  assign n2973 = ~\shift[6]  & ~n2972;
  assign n2974 = n479 & ~n1868;
  assign n2975 = n426 & ~n1876;
  assign n2976 = ~n2974 & ~n2975;
  assign n2977 = n372 & ~n1912;
  assign n2978 = n319 & ~n1904;
  assign n2979 = ~n2977 & ~n2978;
  assign n2980 = n2976 & n2979;
  assign n2981 = \shift[6]  & ~n2980;
  assign \result[38]  = n2973 | n2981;
  assign n2983 = n479 & ~n2002;
  assign n2984 = n426 & ~n1994;
  assign n2985 = ~n2983 & ~n2984;
  assign n2986 = n372 & ~n1958;
  assign n2987 = n319 & ~n1966;
  assign n2988 = ~n2986 & ~n2987;
  assign n2989 = n2985 & n2988;
  assign n2990 = ~\shift[6]  & ~n2989;
  assign n2991 = n319 & ~n1977;
  assign n2992 = n372 & ~n1985;
  assign n2993 = ~n2991 & ~n2992;
  assign n2994 = n426 & ~n1949;
  assign n2995 = n479 & ~n1941;
  assign n2996 = ~n2994 & ~n2995;
  assign n2997 = n2993 & n2996;
  assign n2998 = \shift[6]  & ~n2997;
  assign \result[39]  = n2990 | n2998;
  assign n3000 = n479 & ~n2075;
  assign n3001 = n426 & ~n2067;
  assign n3002 = ~n3000 & ~n3001;
  assign n3003 = n372 & ~n2031;
  assign n3004 = n319 & ~n2039;
  assign n3005 = ~n3003 & ~n3004;
  assign n3006 = n3002 & n3005;
  assign n3007 = ~\shift[6]  & ~n3006;
  assign n3008 = n319 & ~n2050;
  assign n3009 = n372 & ~n2058;
  assign n3010 = ~n3008 & ~n3009;
  assign n3011 = n426 & ~n2022;
  assign n3012 = n479 & ~n2014;
  assign n3013 = ~n3011 & ~n3012;
  assign n3014 = n3010 & n3013;
  assign n3015 = \shift[6]  & ~n3014;
  assign \result[40]  = n3007 | n3015;
  assign n3017 = n479 & ~n2148;
  assign n3018 = n426 & ~n2140;
  assign n3019 = ~n3017 & ~n3018;
  assign n3020 = n372 & ~n2104;
  assign n3021 = n319 & ~n2112;
  assign n3022 = ~n3020 & ~n3021;
  assign n3023 = n3019 & n3022;
  assign n3024 = ~\shift[6]  & ~n3023;
  assign n3025 = n319 & ~n2123;
  assign n3026 = n372 & ~n2131;
  assign n3027 = ~n3025 & ~n3026;
  assign n3028 = n426 & ~n2095;
  assign n3029 = n479 & ~n2087;
  assign n3030 = ~n3028 & ~n3029;
  assign n3031 = n3027 & n3030;
  assign n3032 = \shift[6]  & ~n3031;
  assign \result[41]  = n3024 | n3032;
  assign n3034 = n319 & ~n2185;
  assign n3035 = n372 & ~n2177;
  assign n3036 = ~n3034 & ~n3035;
  assign n3037 = n426 & ~n2213;
  assign n3038 = n479 & ~n2221;
  assign n3039 = ~n3037 & ~n3038;
  assign n3040 = n3036 & n3039;
  assign n3041 = ~\shift[6]  & ~n3040;
  assign n3042 = n319 & ~n2196;
  assign n3043 = n372 & ~n2204;
  assign n3044 = ~n3042 & ~n3043;
  assign n3045 = n426 & ~n2168;
  assign n3046 = n479 & ~n2160;
  assign n3047 = ~n3045 & ~n3046;
  assign n3048 = n3044 & n3047;
  assign n3049 = \shift[6]  & ~n3048;
  assign \result[42]  = n3041 | n3049;
  assign n3051 = n319 & ~n2258;
  assign n3052 = n372 & ~n2250;
  assign n3053 = ~n3051 & ~n3052;
  assign n3054 = n426 & ~n2286;
  assign n3055 = n479 & ~n2294;
  assign n3056 = ~n3054 & ~n3055;
  assign n3057 = n3053 & n3056;
  assign n3058 = ~\shift[6]  & ~n3057;
  assign n3059 = n319 & ~n2269;
  assign n3060 = n372 & ~n2277;
  assign n3061 = ~n3059 & ~n3060;
  assign n3062 = n426 & ~n2241;
  assign n3063 = n479 & ~n2233;
  assign n3064 = ~n3062 & ~n3063;
  assign n3065 = n3061 & n3064;
  assign n3066 = \shift[6]  & ~n3065;
  assign \result[43]  = n3058 | n3066;
  assign n3068 = n319 & ~n2331;
  assign n3069 = n372 & ~n2323;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = n426 & ~n2359;
  assign n3072 = n479 & ~n2367;
  assign n3073 = ~n3071 & ~n3072;
  assign n3074 = n3070 & n3073;
  assign n3075 = ~\shift[6]  & ~n3074;
  assign n3076 = n319 & ~n2342;
  assign n3077 = n372 & ~n2350;
  assign n3078 = ~n3076 & ~n3077;
  assign n3079 = n426 & ~n2314;
  assign n3080 = n479 & ~n2306;
  assign n3081 = ~n3079 & ~n3080;
  assign n3082 = n3078 & n3081;
  assign n3083 = \shift[6]  & ~n3082;
  assign \result[44]  = n3075 | n3083;
  assign n3085 = n319 & ~n2404;
  assign n3086 = n372 & ~n2396;
  assign n3087 = ~n3085 & ~n3086;
  assign n3088 = n426 & ~n2432;
  assign n3089 = n479 & ~n2440;
  assign n3090 = ~n3088 & ~n3089;
  assign n3091 = n3087 & n3090;
  assign n3092 = ~\shift[6]  & ~n3091;
  assign n3093 = n319 & ~n2415;
  assign n3094 = n372 & ~n2423;
  assign n3095 = ~n3093 & ~n3094;
  assign n3096 = n426 & ~n2387;
  assign n3097 = n479 & ~n2379;
  assign n3098 = ~n3096 & ~n3097;
  assign n3099 = n3095 & n3098;
  assign n3100 = \shift[6]  & ~n3099;
  assign \result[45]  = n3092 | n3100;
  assign n3102 = n319 & ~n2477;
  assign n3103 = n372 & ~n2469;
  assign n3104 = ~n3102 & ~n3103;
  assign n3105 = n426 & ~n2505;
  assign n3106 = n479 & ~n2513;
  assign n3107 = ~n3105 & ~n3106;
  assign n3108 = n3104 & n3107;
  assign n3109 = ~\shift[6]  & ~n3108;
  assign n3110 = n319 & ~n2488;
  assign n3111 = n372 & ~n2496;
  assign n3112 = ~n3110 & ~n3111;
  assign n3113 = n426 & ~n2460;
  assign n3114 = n479 & ~n2452;
  assign n3115 = ~n3113 & ~n3114;
  assign n3116 = n3112 & n3115;
  assign n3117 = \shift[6]  & ~n3116;
  assign \result[46]  = n3109 | n3117;
  assign n3119 = n319 & ~n2550;
  assign n3120 = n372 & ~n2542;
  assign n3121 = ~n3119 & ~n3120;
  assign n3122 = n426 & ~n2578;
  assign n3123 = n479 & ~n2586;
  assign n3124 = ~n3122 & ~n3123;
  assign n3125 = n3121 & n3124;
  assign n3126 = ~\shift[6]  & ~n3125;
  assign n3127 = n319 & ~n2561;
  assign n3128 = n372 & ~n2569;
  assign n3129 = ~n3127 & ~n3128;
  assign n3130 = n426 & ~n2533;
  assign n3131 = n479 & ~n2525;
  assign n3132 = ~n3130 & ~n3131;
  assign n3133 = n3129 & n3132;
  assign n3134 = \shift[6]  & ~n3133;
  assign \result[47]  = n3126 | n3134;
  assign n3136 = n319 & ~n425;
  assign n3137 = n372 & ~n534;
  assign n3138 = ~n3136 & ~n3137;
  assign n3139 = n426 & ~n691;
  assign n3140 = n479 & ~n586;
  assign n3141 = ~n3139 & ~n3140;
  assign n3142 = n3138 & n3141;
  assign n3143 = ~\shift[6]  & ~n3142;
  assign n3144 = ~n318 & n372;
  assign n3145 = ~n371 & n479;
  assign n3146 = ~n3144 & ~n3145;
  assign n3147 = n319 & ~n639;
  assign n3148 = n426 & ~n478;
  assign n3149 = ~n3147 & ~n3148;
  assign n3150 = n3146 & n3149;
  assign n3151 = \shift[6]  & ~n3150;
  assign \result[48]  = n3143 | n3151;
  assign n3153 = n319 & ~n852;
  assign n3154 = n372 & ~n1011;
  assign n3155 = ~n3153 & ~n3154;
  assign n3156 = n426 & ~n1064;
  assign n3157 = n479 & ~n1116;
  assign n3158 = ~n3156 & ~n3157;
  assign n3159 = n3155 & n3158;
  assign n3160 = ~\shift[6]  & ~n3159;
  assign n3161 = n319 & ~n959;
  assign n3162 = n372 & ~n747;
  assign n3163 = ~n3161 & ~n3162;
  assign n3164 = n426 & ~n904;
  assign n3165 = n479 & ~n799;
  assign n3166 = ~n3164 & ~n3165;
  assign n3167 = n3163 & n3166;
  assign n3168 = \shift[6]  & ~n3167;
  assign \result[49]  = n3160 | n3168;
  assign n3170 = n319 & ~n1229;
  assign n3171 = n372 & ~n1340;
  assign n3172 = ~n3170 & ~n3171;
  assign n3173 = n426 & ~n1377;
  assign n3174 = n479 & ~n1413;
  assign n3175 = ~n3173 & ~n3174;
  assign n3176 = n3172 & n3175;
  assign n3177 = ~\shift[6]  & ~n3176;
  assign n3178 = n319 & ~n1304;
  assign n3179 = n372 & ~n1156;
  assign n3180 = ~n3178 & ~n3179;
  assign n3181 = n426 & ~n1265;
  assign n3182 = n479 & ~n1192;
  assign n3183 = ~n3181 & ~n3182;
  assign n3184 = n3180 & n3183;
  assign n3185 = \shift[6]  & ~n3184;
  assign \result[50]  = n3177 | n3185;
  assign n3187 = n426 & ~n1637;
  assign n3188 = n479 & ~n1710;
  assign n3189 = ~n3187 & ~n3188;
  assign n3190 = n319 & ~n1526;
  assign n3191 = n372 & ~n1674;
  assign n3192 = ~n3190 & ~n3191;
  assign n3193 = n3189 & n3192;
  assign n3194 = ~\shift[6]  & ~n3193;
  assign n3195 = n319 & ~n1601;
  assign n3196 = n426 & ~n1453;
  assign n3197 = ~n3195 & ~n3196;
  assign n3198 = n372 & ~n1562;
  assign n3199 = n479 & ~n1489;
  assign n3200 = ~n3198 & ~n3199;
  assign n3201 = n3197 & n3200;
  assign n3202 = \shift[6]  & ~n3201;
  assign \result[51]  = n3194 | n3202;
  assign n3204 = n426 & ~n1758;
  assign n3205 = n319 & ~n1739;
  assign n3206 = ~n3204 & ~n3205;
  assign n3207 = n479 & ~n1775;
  assign n3208 = n372 & ~n1783;
  assign n3209 = ~n3207 & ~n3208;
  assign n3210 = n3206 & n3209;
  assign n3211 = ~\shift[6]  & ~n3210;
  assign n3212 = n372 & ~n1722;
  assign n3213 = n479 & ~n1730;
  assign n3214 = ~n3212 & ~n3213;
  assign n3215 = n426 & ~n1747;
  assign n3216 = n319 & ~n1766;
  assign n3217 = ~n3215 & ~n3216;
  assign n3218 = n3214 & n3217;
  assign n3219 = \shift[6]  & ~n3218;
  assign \result[52]  = n3211 | n3219;
  assign n3221 = n426 & ~n1831;
  assign n3222 = n319 & ~n1812;
  assign n3223 = ~n3221 & ~n3222;
  assign n3224 = n479 & ~n1848;
  assign n3225 = n372 & ~n1856;
  assign n3226 = ~n3224 & ~n3225;
  assign n3227 = n3223 & n3226;
  assign n3228 = ~\shift[6]  & ~n3227;
  assign n3229 = n372 & ~n1795;
  assign n3230 = n479 & ~n1803;
  assign n3231 = ~n3229 & ~n3230;
  assign n3232 = n426 & ~n1820;
  assign n3233 = n319 & ~n1839;
  assign n3234 = ~n3232 & ~n3233;
  assign n3235 = n3231 & n3234;
  assign n3236 = \shift[6]  & ~n3235;
  assign \result[53]  = n3228 | n3236;
  assign n3238 = n426 & ~n1904;
  assign n3239 = n319 & ~n1885;
  assign n3240 = ~n3238 & ~n3239;
  assign n3241 = n479 & ~n1921;
  assign n3242 = n372 & ~n1929;
  assign n3243 = ~n3241 & ~n3242;
  assign n3244 = n3240 & n3243;
  assign n3245 = ~\shift[6]  & ~n3244;
  assign n3246 = n372 & ~n1868;
  assign n3247 = n479 & ~n1876;
  assign n3248 = ~n3246 & ~n3247;
  assign n3249 = n426 & ~n1893;
  assign n3250 = n319 & ~n1912;
  assign n3251 = ~n3249 & ~n3250;
  assign n3252 = n3248 & n3251;
  assign n3253 = \shift[6]  & ~n3252;
  assign \result[54]  = n3245 | n3253;
  assign n3255 = n426 & ~n1977;
  assign n3256 = n372 & ~n2002;
  assign n3257 = ~n3255 & ~n3256;
  assign n3258 = n319 & ~n1958;
  assign n3259 = n479 & ~n1994;
  assign n3260 = ~n3258 & ~n3259;
  assign n3261 = n3257 & n3260;
  assign n3262 = ~\shift[6]  & ~n3261;
  assign n3263 = n319 & ~n1985;
  assign n3264 = n372 & ~n1941;
  assign n3265 = ~n3263 & ~n3264;
  assign n3266 = n426 & ~n1966;
  assign n3267 = n479 & ~n1949;
  assign n3268 = ~n3266 & ~n3267;
  assign n3269 = n3265 & n3268;
  assign n3270 = \shift[6]  & ~n3269;
  assign \result[55]  = n3262 | n3270;
  assign n3272 = n426 & ~n2050;
  assign n3273 = n372 & ~n2075;
  assign n3274 = ~n3272 & ~n3273;
  assign n3275 = n319 & ~n2031;
  assign n3276 = n479 & ~n2067;
  assign n3277 = ~n3275 & ~n3276;
  assign n3278 = n3274 & n3277;
  assign n3279 = ~\shift[6]  & ~n3278;
  assign n3280 = n319 & ~n2058;
  assign n3281 = n372 & ~n2014;
  assign n3282 = ~n3280 & ~n3281;
  assign n3283 = n426 & ~n2039;
  assign n3284 = n479 & ~n2022;
  assign n3285 = ~n3283 & ~n3284;
  assign n3286 = n3282 & n3285;
  assign n3287 = \shift[6]  & ~n3286;
  assign \result[56]  = n3279 | n3287;
  assign n3289 = n426 & ~n2123;
  assign n3290 = n372 & ~n2148;
  assign n3291 = ~n3289 & ~n3290;
  assign n3292 = n319 & ~n2104;
  assign n3293 = n479 & ~n2140;
  assign n3294 = ~n3292 & ~n3293;
  assign n3295 = n3291 & n3294;
  assign n3296 = ~\shift[6]  & ~n3295;
  assign n3297 = n319 & ~n2131;
  assign n3298 = n372 & ~n2087;
  assign n3299 = ~n3297 & ~n3298;
  assign n3300 = n426 & ~n2112;
  assign n3301 = n479 & ~n2095;
  assign n3302 = ~n3300 & ~n3301;
  assign n3303 = n3299 & n3302;
  assign n3304 = \shift[6]  & ~n3303;
  assign \result[57]  = n3296 | n3304;
  assign n3306 = n426 & ~n2196;
  assign n3307 = n319 & ~n2177;
  assign n3308 = ~n3306 & ~n3307;
  assign n3309 = n479 & ~n2213;
  assign n3310 = n372 & ~n2221;
  assign n3311 = ~n3309 & ~n3310;
  assign n3312 = n3308 & n3311;
  assign n3313 = ~\shift[6]  & ~n3312;
  assign n3314 = n319 & ~n2204;
  assign n3315 = n372 & ~n2160;
  assign n3316 = ~n3314 & ~n3315;
  assign n3317 = n426 & ~n2185;
  assign n3318 = n479 & ~n2168;
  assign n3319 = ~n3317 & ~n3318;
  assign n3320 = n3316 & n3319;
  assign n3321 = \shift[6]  & ~n3320;
  assign \result[58]  = n3313 | n3321;
  assign n3323 = n426 & ~n2269;
  assign n3324 = n319 & ~n2250;
  assign n3325 = ~n3323 & ~n3324;
  assign n3326 = n479 & ~n2286;
  assign n3327 = n372 & ~n2294;
  assign n3328 = ~n3326 & ~n3327;
  assign n3329 = n3325 & n3328;
  assign n3330 = ~\shift[6]  & ~n3329;
  assign n3331 = n319 & ~n2277;
  assign n3332 = n372 & ~n2233;
  assign n3333 = ~n3331 & ~n3332;
  assign n3334 = n426 & ~n2258;
  assign n3335 = n479 & ~n2241;
  assign n3336 = ~n3334 & ~n3335;
  assign n3337 = n3333 & n3336;
  assign n3338 = \shift[6]  & ~n3337;
  assign \result[59]  = n3330 | n3338;
  assign n3340 = n426 & ~n2342;
  assign n3341 = n319 & ~n2323;
  assign n3342 = ~n3340 & ~n3341;
  assign n3343 = n479 & ~n2359;
  assign n3344 = n372 & ~n2367;
  assign n3345 = ~n3343 & ~n3344;
  assign n3346 = n3342 & n3345;
  assign n3347 = ~\shift[6]  & ~n3346;
  assign n3348 = n319 & ~n2350;
  assign n3349 = n372 & ~n2306;
  assign n3350 = ~n3348 & ~n3349;
  assign n3351 = n426 & ~n2331;
  assign n3352 = n479 & ~n2314;
  assign n3353 = ~n3351 & ~n3352;
  assign n3354 = n3350 & n3353;
  assign n3355 = \shift[6]  & ~n3354;
  assign \result[60]  = n3347 | n3355;
  assign n3357 = n426 & ~n2415;
  assign n3358 = n319 & ~n2396;
  assign n3359 = ~n3357 & ~n3358;
  assign n3360 = n479 & ~n2432;
  assign n3361 = n372 & ~n2440;
  assign n3362 = ~n3360 & ~n3361;
  assign n3363 = n3359 & n3362;
  assign n3364 = ~\shift[6]  & ~n3363;
  assign n3365 = n319 & ~n2423;
  assign n3366 = n372 & ~n2379;
  assign n3367 = ~n3365 & ~n3366;
  assign n3368 = n426 & ~n2404;
  assign n3369 = n479 & ~n2387;
  assign n3370 = ~n3368 & ~n3369;
  assign n3371 = n3367 & n3370;
  assign n3372 = \shift[6]  & ~n3371;
  assign \result[61]  = n3364 | n3372;
  assign n3374 = n426 & ~n2488;
  assign n3375 = n319 & ~n2469;
  assign n3376 = ~n3374 & ~n3375;
  assign n3377 = n479 & ~n2505;
  assign n3378 = n372 & ~n2513;
  assign n3379 = ~n3377 & ~n3378;
  assign n3380 = n3376 & n3379;
  assign n3381 = ~\shift[6]  & ~n3380;
  assign n3382 = n319 & ~n2496;
  assign n3383 = n372 & ~n2452;
  assign n3384 = ~n3382 & ~n3383;
  assign n3385 = n426 & ~n2477;
  assign n3386 = n479 & ~n2460;
  assign n3387 = ~n3385 & ~n3386;
  assign n3388 = n3384 & n3387;
  assign n3389 = \shift[6]  & ~n3388;
  assign \result[62]  = n3381 | n3389;
  assign n3391 = n426 & ~n2561;
  assign n3392 = n319 & ~n2542;
  assign n3393 = ~n3391 & ~n3392;
  assign n3394 = n479 & ~n2578;
  assign n3395 = n372 & ~n2586;
  assign n3396 = ~n3394 & ~n3395;
  assign n3397 = n3393 & n3396;
  assign n3398 = ~\shift[6]  & ~n3397;
  assign n3399 = n319 & ~n2569;
  assign n3400 = n372 & ~n2525;
  assign n3401 = ~n3399 & ~n3400;
  assign n3402 = n426 & ~n2550;
  assign n3403 = n479 & ~n2533;
  assign n3404 = ~n3402 & ~n3403;
  assign n3405 = n3401 & n3404;
  assign n3406 = \shift[6]  & ~n3405;
  assign \result[63]  = n3398 | n3406;
  assign n3408 = ~\shift[6]  & ~n694;
  assign n3409 = \shift[6]  & ~n482;
  assign \result[64]  = n3408 | n3409;
  assign n3411 = ~\shift[6]  & ~n1119;
  assign n3412 = \shift[6]  & ~n907;
  assign \result[65]  = n3411 | n3412;
  assign n3414 = ~\shift[6]  & ~n1416;
  assign n3415 = \shift[6]  & ~n1268;
  assign \result[66]  = n3414 | n3415;
  assign n3417 = ~\shift[6]  & ~n1713;
  assign n3418 = \shift[6]  & ~n1565;
  assign \result[67]  = n3417 | n3418;
  assign n3420 = ~\shift[6]  & ~n1786;
  assign n3421 = \shift[6]  & ~n1750;
  assign \result[68]  = n3420 | n3421;
  assign n3423 = ~\shift[6]  & ~n1859;
  assign n3424 = \shift[6]  & ~n1823;
  assign \result[69]  = n3423 | n3424;
  assign n3426 = ~\shift[6]  & ~n1932;
  assign n3427 = \shift[6]  & ~n1896;
  assign \result[70]  = n3426 | n3427;
  assign n3429 = ~\shift[6]  & ~n2005;
  assign n3430 = \shift[6]  & ~n1969;
  assign \result[71]  = n3429 | n3430;
  assign n3432 = ~\shift[6]  & ~n2078;
  assign n3433 = \shift[6]  & ~n2042;
  assign \result[72]  = n3432 | n3433;
  assign n3435 = ~\shift[6]  & ~n2151;
  assign n3436 = \shift[6]  & ~n2115;
  assign \result[73]  = n3435 | n3436;
  assign n3438 = ~\shift[6]  & ~n2224;
  assign n3439 = \shift[6]  & ~n2188;
  assign \result[74]  = n3438 | n3439;
  assign n3441 = ~\shift[6]  & ~n2297;
  assign n3442 = \shift[6]  & ~n2261;
  assign \result[75]  = n3441 | n3442;
  assign n3444 = ~\shift[6]  & ~n2370;
  assign n3445 = \shift[6]  & ~n2334;
  assign \result[76]  = n3444 | n3445;
  assign n3447 = ~\shift[6]  & ~n2443;
  assign n3448 = \shift[6]  & ~n2407;
  assign \result[77]  = n3447 | n3448;
  assign n3450 = ~\shift[6]  & ~n2516;
  assign n3451 = \shift[6]  & ~n2480;
  assign \result[78]  = n3450 | n3451;
  assign n3453 = ~\shift[6]  & ~n2589;
  assign n3454 = \shift[6]  & ~n2553;
  assign \result[79]  = n3453 | n3454;
  assign n3456 = ~\shift[6]  & ~n2606;
  assign n3457 = \shift[6]  & ~n2598;
  assign \result[80]  = n3456 | n3457;
  assign n3459 = ~\shift[6]  & ~n2623;
  assign n3460 = \shift[6]  & ~n2615;
  assign \result[81]  = n3459 | n3460;
  assign n3462 = ~\shift[6]  & ~n2640;
  assign n3463 = \shift[6]  & ~n2632;
  assign \result[82]  = n3462 | n3463;
  assign n3465 = ~\shift[6]  & ~n2657;
  assign n3466 = \shift[6]  & ~n2649;
  assign \result[83]  = n3465 | n3466;
  assign n3468 = ~\shift[6]  & ~n2674;
  assign n3469 = \shift[6]  & ~n2666;
  assign \result[84]  = n3468 | n3469;
  assign n3471 = ~\shift[6]  & ~n2691;
  assign n3472 = \shift[6]  & ~n2683;
  assign \result[85]  = n3471 | n3472;
  assign n3474 = ~\shift[6]  & ~n2708;
  assign n3475 = \shift[6]  & ~n2700;
  assign \result[86]  = n3474 | n3475;
  assign n3477 = ~\shift[6]  & ~n2725;
  assign n3478 = \shift[6]  & ~n2717;
  assign \result[87]  = n3477 | n3478;
  assign n3480 = ~\shift[6]  & ~n2742;
  assign n3481 = \shift[6]  & ~n2734;
  assign \result[88]  = n3480 | n3481;
  assign n3483 = ~\shift[6]  & ~n2759;
  assign n3484 = \shift[6]  & ~n2751;
  assign \result[89]  = n3483 | n3484;
  assign n3486 = ~\shift[6]  & ~n2776;
  assign n3487 = \shift[6]  & ~n2768;
  assign \result[90]  = n3486 | n3487;
  assign n3489 = ~\shift[6]  & ~n2793;
  assign n3490 = \shift[6]  & ~n2785;
  assign \result[91]  = n3489 | n3490;
  assign n3492 = ~\shift[6]  & ~n2810;
  assign n3493 = \shift[6]  & ~n2802;
  assign \result[92]  = n3492 | n3493;
  assign n3495 = ~\shift[6]  & ~n2827;
  assign n3496 = \shift[6]  & ~n2819;
  assign \result[93]  = n3495 | n3496;
  assign n3498 = ~\shift[6]  & ~n2844;
  assign n3499 = \shift[6]  & ~n2836;
  assign \result[94]  = n3498 | n3499;
  assign n3501 = ~\shift[6]  & ~n2861;
  assign n3502 = \shift[6]  & ~n2853;
  assign \result[95]  = n3501 | n3502;
  assign n3504 = ~\shift[6]  & ~n2878;
  assign n3505 = \shift[6]  & ~n2870;
  assign \result[96]  = n3504 | n3505;
  assign n3507 = ~\shift[6]  & ~n2895;
  assign n3508 = \shift[6]  & ~n2887;
  assign \result[97]  = n3507 | n3508;
  assign n3510 = ~\shift[6]  & ~n2912;
  assign n3511 = \shift[6]  & ~n2904;
  assign \result[98]  = n3510 | n3511;
  assign n3513 = ~\shift[6]  & ~n2929;
  assign n3514 = \shift[6]  & ~n2921;
  assign \result[99]  = n3513 | n3514;
  assign n3516 = ~\shift[6]  & ~n2946;
  assign n3517 = \shift[6]  & ~n2938;
  assign \result[100]  = n3516 | n3517;
  assign n3519 = ~\shift[6]  & ~n2963;
  assign n3520 = \shift[6]  & ~n2955;
  assign \result[101]  = n3519 | n3520;
  assign n3522 = ~\shift[6]  & ~n2980;
  assign n3523 = \shift[6]  & ~n2972;
  assign \result[102]  = n3522 | n3523;
  assign n3525 = ~\shift[6]  & ~n2997;
  assign n3526 = \shift[6]  & ~n2989;
  assign \result[103]  = n3525 | n3526;
  assign n3528 = ~\shift[6]  & ~n3014;
  assign n3529 = \shift[6]  & ~n3006;
  assign \result[104]  = n3528 | n3529;
  assign n3531 = ~\shift[6]  & ~n3031;
  assign n3532 = \shift[6]  & ~n3023;
  assign \result[105]  = n3531 | n3532;
  assign n3534 = ~\shift[6]  & ~n3048;
  assign n3535 = \shift[6]  & ~n3040;
  assign \result[106]  = n3534 | n3535;
  assign n3537 = ~\shift[6]  & ~n3065;
  assign n3538 = \shift[6]  & ~n3057;
  assign \result[107]  = n3537 | n3538;
  assign n3540 = ~\shift[6]  & ~n3082;
  assign n3541 = \shift[6]  & ~n3074;
  assign \result[108]  = n3540 | n3541;
  assign n3543 = ~\shift[6]  & ~n3099;
  assign n3544 = \shift[6]  & ~n3091;
  assign \result[109]  = n3543 | n3544;
  assign n3546 = ~\shift[6]  & ~n3116;
  assign n3547 = \shift[6]  & ~n3108;
  assign \result[110]  = n3546 | n3547;
  assign n3549 = ~\shift[6]  & ~n3133;
  assign n3550 = \shift[6]  & ~n3125;
  assign \result[111]  = n3549 | n3550;
  assign n3552 = ~\shift[6]  & ~n3150;
  assign n3553 = \shift[6]  & ~n3142;
  assign \result[112]  = n3552 | n3553;
  assign n3555 = ~\shift[6]  & ~n3167;
  assign n3556 = \shift[6]  & ~n3159;
  assign \result[113]  = n3555 | n3556;
  assign n3558 = ~\shift[6]  & ~n3184;
  assign n3559 = \shift[6]  & ~n3176;
  assign \result[114]  = n3558 | n3559;
  assign n3561 = ~\shift[6]  & ~n3201;
  assign n3562 = \shift[6]  & ~n3193;
  assign \result[115]  = n3561 | n3562;
  assign n3564 = ~\shift[6]  & ~n3218;
  assign n3565 = \shift[6]  & ~n3210;
  assign \result[116]  = n3564 | n3565;
  assign n3567 = ~\shift[6]  & ~n3235;
  assign n3568 = \shift[6]  & ~n3227;
  assign \result[117]  = n3567 | n3568;
  assign n3570 = ~\shift[6]  & ~n3252;
  assign n3571 = \shift[6]  & ~n3244;
  assign \result[118]  = n3570 | n3571;
  assign n3573 = ~\shift[6]  & ~n3269;
  assign n3574 = \shift[6]  & ~n3261;
  assign \result[119]  = n3573 | n3574;
  assign n3576 = ~\shift[6]  & ~n3286;
  assign n3577 = \shift[6]  & ~n3278;
  assign \result[120]  = n3576 | n3577;
  assign n3579 = ~\shift[6]  & ~n3303;
  assign n3580 = \shift[6]  & ~n3295;
  assign \result[121]  = n3579 | n3580;
  assign n3582 = ~\shift[6]  & ~n3320;
  assign n3583 = \shift[6]  & ~n3312;
  assign \result[122]  = n3582 | n3583;
  assign n3585 = ~\shift[6]  & ~n3337;
  assign n3586 = \shift[6]  & ~n3329;
  assign \result[123]  = n3585 | n3586;
  assign n3588 = ~\shift[6]  & ~n3354;
  assign n3589 = \shift[6]  & ~n3346;
  assign \result[124]  = n3588 | n3589;
  assign n3591 = ~\shift[6]  & ~n3371;
  assign n3592 = \shift[6]  & ~n3363;
  assign \result[125]  = n3591 | n3592;
  assign n3594 = ~\shift[6]  & ~n3388;
  assign n3595 = \shift[6]  & ~n3380;
  assign \result[126]  = n3594 | n3595;
  assign n3597 = ~\shift[6]  & ~n3405;
  assign n3598 = \shift[6]  & ~n3397;
  assign \result[127]  = n3597 | n3598;
endmodule


