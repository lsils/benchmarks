library ieee;
use ieee.std_logic_1164.all;

entity top is
port( in0,in1,in2,in3: in std_logic_vector(127 downto 0);
address: out std_logic_vector(1 downto 0);
result: out std_logic_vector(127 downto 0));
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864: std_logic;

begin

w0 <= in2(119) and not in3(119);
w1 <= not in2(119) and in3(119);
w2 <= not in2(118) and in3(118);
w3 <= not w1 and not w2;
w4 <= not in2(117) and in3(117);
w5 <= in2(116) and not in3(116);
w6 <= not w4 and w5;
w7 <= in2(117) and not in3(117);
w8 <= not w6 and not w7;
w9 <= w3 and not w8;
w10 <= not in3(118) and not w1;
w11 <= in2(118) and w10;
w12 <= not in2(112) and in3(112);
w13 <= not in2(115) and in3(115);
w14 <= not in2(114) and in3(114);
w15 <= not w13 and not w14;
w16 <= not in2(113) and in3(113);
w17 <= in2(111) and not in3(111);
w18 <= not in2(111) and in3(111);
w19 <= not in2(110) and in3(110);
w20 <= not w18 and not w19;
w21 <= not in2(109) and in3(109);
w22 <= in2(108) and not in3(108);
w23 <= not w21 and w22;
w24 <= in2(109) and not in3(109);
w25 <= not w23 and not w24;
w26 <= w20 and not w25;
w27 <= not in3(110) and not w18;
w28 <= in2(110) and w27;
w29 <= in2(103) and not in3(103);
w30 <= not in2(103) and in3(103);
w31 <= not in2(102) and in3(102);
w32 <= not w30 and not w31;
w33 <= not in2(101) and in3(101);
w34 <= in2(100) and not in3(100);
w35 <= not w33 and w34;
w36 <= in2(101) and not in3(101);
w37 <= not w35 and not w36;
w38 <= w32 and not w37;
w39 <= not in3(102) and not w30;
w40 <= in2(102) and w39;
w41 <= not in2(96) and in3(96);
w42 <= not in2(99) and in3(99);
w43 <= not in2(98) and in3(98);
w44 <= not w42 and not w43;
w45 <= not in2(97) and in3(97);
w46 <= in2(95) and not in3(95);
w47 <= not in2(95) and in3(95);
w48 <= not in2(94) and in3(94);
w49 <= not w47 and not w48;
w50 <= not in2(93) and in3(93);
w51 <= in2(92) and not in3(92);
w52 <= not w50 and w51;
w53 <= in2(93) and not in3(93);
w54 <= not w52 and not w53;
w55 <= w49 and not w54;
w56 <= not in3(94) and not w47;
w57 <= in2(94) and w56;
w58 <= in2(87) and not in3(87);
w59 <= not in2(87) and in3(87);
w60 <= not in2(86) and in3(86);
w61 <= not w59 and not w60;
w62 <= not in2(85) and in3(85);
w63 <= in2(84) and not in3(84);
w64 <= not w62 and w63;
w65 <= in2(85) and not in3(85);
w66 <= not w64 and not w65;
w67 <= w61 and not w66;
w68 <= not in3(86) and not w59;
w69 <= in2(86) and w68;
w70 <= not in2(80) and in3(80);
w71 <= not in2(83) and in3(83);
w72 <= not in2(82) and in3(82);
w73 <= not w71 and not w72;
w74 <= not in2(81) and in3(81);
w75 <= in2(79) and not in3(79);
w76 <= not in2(79) and in3(79);
w77 <= not in2(78) and in3(78);
w78 <= not w76 and not w77;
w79 <= not in2(77) and in3(77);
w80 <= in2(76) and not in3(76);
w81 <= not w79 and w80;
w82 <= in2(77) and not in3(77);
w83 <= not w81 and not w82;
w84 <= w78 and not w83;
w85 <= not in3(78) and not w76;
w86 <= in2(78) and w85;
w87 <= in2(71) and not in3(71);
w88 <= not in2(71) and in3(71);
w89 <= not in2(70) and in3(70);
w90 <= not w88 and not w89;
w91 <= not in2(69) and in3(69);
w92 <= in2(68) and not in3(68);
w93 <= not w91 and w92;
w94 <= in2(69) and not in3(69);
w95 <= not w93 and not w94;
w96 <= w90 and not w95;
w97 <= not in3(70) and not w88;
w98 <= in2(70) and w97;
w99 <= not in2(67) and in3(67);
w100 <= not in2(66) and in3(66);
w101 <= not w99 and not w100;
w102 <= not in2(65) and in3(65);
w103 <= in2(63) and not in3(63);
w104 <= not in2(63) and in3(63);
w105 <= not in2(62) and in3(62);
w106 <= not w104 and not w105;
w107 <= not in2(60) and in3(60);
w108 <= not in2(61) and in3(61);
w109 <= not w107 and not w108;
w110 <= w106 and w109;
w111 <= in2(59) and not in3(59);
w112 <= not in2(59) and in3(59);
w113 <= not in2(58) and in3(58);
w114 <= not w112 and not w113;
w115 <= not in2(57) and in3(57);
w116 <= in2(56) and not in3(56);
w117 <= not w115 and w116;
w118 <= in2(57) and not in3(57);
w119 <= not w117 and not w118;
w120 <= in2(58) and not in3(58);
w121 <= w119 and not w120;
w122 <= w114 and not w121;
w123 <= not w111 and not w122;
w124 <= w110 and not w123;
w125 <= in2(60) and not in3(60);
w126 <= not w108 and w125;
w127 <= in2(61) and not in3(61);
w128 <= not w126 and not w127;
w129 <= w106 and not w128;
w130 <= not in3(62) and not w104;
w131 <= in2(62) and w130;
w132 <= in2(47) and not in3(47);
w133 <= not in2(47) and in3(47);
w134 <= not in2(46) and in3(46);
w135 <= not w133 and not w134;
w136 <= not in2(44) and in3(44);
w137 <= not in2(45) and in3(45);
w138 <= not w136 and not w137;
w139 <= w135 and w138;
w140 <= in2(43) and not in3(43);
w141 <= not in2(43) and in3(43);
w142 <= not in2(42) and in3(42);
w143 <= not w141 and not w142;
w144 <= not in2(41) and in3(41);
w145 <= in2(40) and not in3(40);
w146 <= not w144 and w145;
w147 <= in2(41) and not in3(41);
w148 <= not w146 and not w147;
w149 <= in2(42) and not in3(42);
w150 <= w148 and not w149;
w151 <= w143 and not w150;
w152 <= not w140 and not w151;
w153 <= w139 and not w152;
w154 <= in2(44) and not in3(44);
w155 <= not w137 and w154;
w156 <= in2(45) and not in3(45);
w157 <= not w155 and not w156;
w158 <= w135 and not w157;
w159 <= not in3(46) and not w133;
w160 <= in2(46) and w159;
w161 <= not in2(32) and in3(32);
w162 <= not in2(31) and in3(31);
w163 <= not in2(30) and in3(30);
w164 <= not in2(29) and in3(29);
w165 <= not in2(28) and in3(28);
w166 <= not in2(27) and in3(27);
w167 <= not in2(26) and in3(26);
w168 <= not in2(23) and in3(23);
w169 <= not in2(22) and in3(22);
w170 <= not in2(21) and in3(21);
w171 <= not in2(20) and in3(20);
w172 <= not in2(19) and in3(19);
w173 <= not in2(18) and in3(18);
w174 <= not in2(15) and in3(15);
w175 <= not in2(14) and in3(14);
w176 <= not in2(13) and in3(13);
w177 <= not in2(12) and in3(12);
w178 <= not in2(11) and in3(11);
w179 <= not in2(10) and in3(10);
w180 <= not in2(7) and in3(7);
w181 <= not in2(6) and in3(6);
w182 <= not in2(3) and in3(3);
w183 <= in2(0) and not in3(0);
w184 <= in2(1) and w183;
w185 <= in3(1) and not w184;
w186 <= not in2(2) and in3(2);
w187 <= not in2(1) and not w183;
w188 <= not w186 and not w187;
w189 <= not w185 and w188;
w190 <= in2(2) and not in3(2);
w191 <= not w189 and not w190;
w192 <= not w182 and not w191;
w193 <= in2(3) and not in3(3);
w194 <= not w192 and not w193;
w195 <= not in2(4) and w194;
w196 <= not in3(4) and not w195;
w197 <= in2(4) and not w194;
w198 <= not w196 and not w197;
w199 <= not in2(5) and w198;
w200 <= not in3(5) and not w199;
w201 <= in2(5) and not w198;
w202 <= not w200 and not w201;
w203 <= not w181 and not w202;
w204 <= in2(6) and not in3(6);
w205 <= not w203 and not w204;
w206 <= not w180 and not w205;
w207 <= in2(7) and not in3(7);
w208 <= not w206 and not w207;
w209 <= not in2(8) and w208;
w210 <= not in3(8) and not w209;
w211 <= in2(8) and not w208;
w212 <= not w210 and not w211;
w213 <= not in2(9) and w212;
w214 <= not in3(9) and not w213;
w215 <= in2(9) and not w212;
w216 <= not w214 and not w215;
w217 <= not w179 and not w216;
w218 <= in2(10) and not in3(10);
w219 <= not w217 and not w218;
w220 <= not w178 and not w219;
w221 <= in2(11) and not in3(11);
w222 <= not w220 and not w221;
w223 <= not w177 and not w222;
w224 <= in2(12) and not in3(12);
w225 <= not w223 and not w224;
w226 <= not w176 and not w225;
w227 <= in2(13) and not in3(13);
w228 <= not w226 and not w227;
w229 <= not w175 and not w228;
w230 <= in2(14) and not in3(14);
w231 <= not w229 and not w230;
w232 <= not w174 and not w231;
w233 <= in2(15) and not in3(15);
w234 <= not w232 and not w233;
w235 <= not in2(16) and w234;
w236 <= not in3(16) and not w235;
w237 <= in2(16) and not w234;
w238 <= not w236 and not w237;
w239 <= not in2(17) and w238;
w240 <= not in3(17) and not w239;
w241 <= in2(17) and not w238;
w242 <= not w240 and not w241;
w243 <= not w173 and not w242;
w244 <= in2(18) and not in3(18);
w245 <= not w243 and not w244;
w246 <= not w172 and not w245;
w247 <= in2(19) and not in3(19);
w248 <= not w246 and not w247;
w249 <= not w171 and not w248;
w250 <= in2(20) and not in3(20);
w251 <= not w249 and not w250;
w252 <= not w170 and not w251;
w253 <= in2(21) and not in3(21);
w254 <= not w252 and not w253;
w255 <= not w169 and not w254;
w256 <= in2(22) and not in3(22);
w257 <= not w255 and not w256;
w258 <= not w168 and not w257;
w259 <= in2(23) and not in3(23);
w260 <= not w258 and not w259;
w261 <= not in2(24) and w260;
w262 <= not in3(24) and not w261;
w263 <= in2(24) and not w260;
w264 <= not w262 and not w263;
w265 <= not in2(25) and w264;
w266 <= not in3(25) and not w265;
w267 <= in2(25) and not w264;
w268 <= not w266 and not w267;
w269 <= not w167 and not w268;
w270 <= in2(26) and not in3(26);
w271 <= not w269 and not w270;
w272 <= not w166 and not w271;
w273 <= in2(27) and not in3(27);
w274 <= not w272 and not w273;
w275 <= not w165 and not w274;
w276 <= in2(28) and not in3(28);
w277 <= not w275 and not w276;
w278 <= not w164 and not w277;
w279 <= in2(29) and not in3(29);
w280 <= not w278 and not w279;
w281 <= not w163 and not w280;
w282 <= in2(30) and not in3(30);
w283 <= not w281 and not w282;
w284 <= not w162 and not w283;
w285 <= in2(31) and not in3(31);
w286 <= not w284 and not w285;
w287 <= not in2(39) and in3(39);
w288 <= not in2(38) and in3(38);
w289 <= not w287 and not w288;
w290 <= not in2(36) and in3(36);
w291 <= not in2(37) and in3(37);
w292 <= not w290 and not w291;
w293 <= w289 and w292;
w294 <= not in2(33) and in3(33);
w295 <= not in2(35) and in3(35);
w296 <= not in2(34) and in3(34);
w297 <= not w295 and not w296;
w298 <= not w294 and w297;
w299 <= w293 and w298;
w300 <= not w286 and w299;
w301 <= not w161 and w300;
w302 <= in2(39) and not in3(39);
w303 <= in2(36) and not in3(36);
w304 <= not w291 and w303;
w305 <= in2(37) and not in3(37);
w306 <= not w304 and not w305;
w307 <= w289 and not w306;
w308 <= not in3(38) and not w287;
w309 <= in2(38) and w308;
w310 <= in2(35) and not in3(35);
w311 <= not in3(32) and not w294;
w312 <= in2(32) and w311;
w313 <= in2(33) and not in3(33);
w314 <= not w312 and not w313;
w315 <= in2(34) and not in3(34);
w316 <= w314 and not w315;
w317 <= w297 and not w316;
w318 <= not w310 and not w317;
w319 <= w293 and not w318;
w320 <= not w309 and not w319;
w321 <= not w307 and w320;
w322 <= not w302 and w321;
w323 <= not w301 and w322;
w324 <= not in2(40) and in3(40);
w325 <= not w144 and not w324;
w326 <= w143 and w325;
w327 <= w139 and w326;
w328 <= not w323 and w327;
w329 <= not w160 and not w328;
w330 <= not w158 and w329;
w331 <= not w153 and w330;
w332 <= not w132 and w331;
w333 <= not in2(48) and in3(48);
w334 <= not in2(55) and in3(55);
w335 <= not in2(54) and in3(54);
w336 <= not w334 and not w335;
w337 <= not in2(53) and in3(53);
w338 <= not in2(52) and in3(52);
w339 <= not w337 and not w338;
w340 <= w336 and w339;
w341 <= not in2(49) and in3(49);
w342 <= not in2(51) and in3(51);
w343 <= not in2(50) and in3(50);
w344 <= not w342 and not w343;
w345 <= not w341 and w344;
w346 <= w340 and w345;
w347 <= not w333 and w346;
w348 <= not w332 and w347;
w349 <= in2(55) and not in3(55);
w350 <= in2(51) and not in3(51);
w351 <= not in3(48) and not w341;
w352 <= in2(48) and w351;
w353 <= in2(49) and not in3(49);
w354 <= not w352 and not w353;
w355 <= in2(50) and not in3(50);
w356 <= w354 and not w355;
w357 <= w344 and not w356;
w358 <= not w350 and not w357;
w359 <= w340 and not w358;
w360 <= in2(52) and not in3(52);
w361 <= not w337 and w360;
w362 <= in2(53) and not in3(53);
w363 <= not w361 and not w362;
w364 <= in2(54) and not in3(54);
w365 <= w363 and not w364;
w366 <= w336 and not w365;
w367 <= not w359 and not w366;
w368 <= not w349 and w367;
w369 <= not w348 and w368;
w370 <= not in2(56) and in3(56);
w371 <= not w115 and not w370;
w372 <= w110 and w371;
w373 <= w114 and w372;
w374 <= not w369 and w373;
w375 <= not w131 and not w374;
w376 <= not w129 and w375;
w377 <= not w124 and w376;
w378 <= not w103 and w377;
w379 <= not in2(64) and in3(64);
w380 <= not w378 and not w379;
w381 <= not w102 and w380;
w382 <= w101 and w381;
w383 <= in2(67) and not in3(67);
w384 <= in2(64) and not in3(64);
w385 <= not w102 and w384;
w386 <= in2(65) and not in3(65);
w387 <= not w385 and not w386;
w388 <= in2(66) and not in3(66);
w389 <= w387 and not w388;
w390 <= w101 and not w389;
w391 <= not w383 and not w390;
w392 <= not w382 and w391;
w393 <= not in2(68) and in3(68);
w394 <= not w91 and not w393;
w395 <= w90 and w394;
w396 <= not w392 and w395;
w397 <= not w98 and not w396;
w398 <= not w96 and w397;
w399 <= not w87 and w398;
w400 <= not in2(75) and in3(75);
w401 <= not in2(74) and in3(74);
w402 <= not w400 and not w401;
w403 <= not in2(73) and in3(73);
w404 <= not in2(72) and in3(72);
w405 <= not w403 and not w404;
w406 <= w402 and w405;
w407 <= not w399 and w406;
w408 <= in2(75) and not in3(75);
w409 <= in2(72) and not in3(72);
w410 <= not w403 and w409;
w411 <= in2(73) and not in3(73);
w412 <= not w410 and not w411;
w413 <= in2(74) and not in3(74);
w414 <= w412 and not w413;
w415 <= w402 and not w414;
w416 <= not w408 and not w415;
w417 <= not w407 and w416;
w418 <= not in2(76) and in3(76);
w419 <= not w79 and not w418;
w420 <= w78 and w419;
w421 <= not w417 and w420;
w422 <= not w86 and not w421;
w423 <= not w84 and w422;
w424 <= not w75 and w423;
w425 <= not w74 and not w424;
w426 <= w73 and w425;
w427 <= not w70 and w426;
w428 <= in2(83) and not in3(83);
w429 <= not in3(80) and not w74;
w430 <= in2(80) and w429;
w431 <= in2(81) and not in3(81);
w432 <= not w430 and not w431;
w433 <= in2(82) and not in3(82);
w434 <= w432 and not w433;
w435 <= w73 and not w434;
w436 <= not w428 and not w435;
w437 <= not w427 and w436;
w438 <= not in2(84) and in3(84);
w439 <= not w62 and not w438;
w440 <= w61 and w439;
w441 <= not w437 and w440;
w442 <= not w69 and not w441;
w443 <= not w67 and w442;
w444 <= not w58 and w443;
w445 <= not in2(91) and in3(91);
w446 <= not in2(90) and in3(90);
w447 <= not w445 and not w446;
w448 <= not in2(89) and in3(89);
w449 <= not in2(88) and in3(88);
w450 <= not w448 and not w449;
w451 <= w447 and w450;
w452 <= not w444 and w451;
w453 <= in2(91) and not in3(91);
w454 <= in2(88) and not in3(88);
w455 <= not w448 and w454;
w456 <= in2(89) and not in3(89);
w457 <= not w455 and not w456;
w458 <= in2(90) and not in3(90);
w459 <= w457 and not w458;
w460 <= w447 and not w459;
w461 <= not w453 and not w460;
w462 <= not w452 and w461;
w463 <= not in2(92) and in3(92);
w464 <= not w50 and not w463;
w465 <= w49 and w464;
w466 <= not w462 and w465;
w467 <= not w57 and not w466;
w468 <= not w55 and w467;
w469 <= not w46 and w468;
w470 <= not w45 and not w469;
w471 <= w44 and w470;
w472 <= not w41 and w471;
w473 <= in2(99) and not in3(99);
w474 <= not in3(96) and not w45;
w475 <= in2(96) and w474;
w476 <= in2(97) and not in3(97);
w477 <= not w475 and not w476;
w478 <= in2(98) and not in3(98);
w479 <= w477 and not w478;
w480 <= w44 and not w479;
w481 <= not w473 and not w480;
w482 <= not w472 and w481;
w483 <= not in2(100) and in3(100);
w484 <= not w33 and not w483;
w485 <= w32 and w484;
w486 <= not w482 and w485;
w487 <= not w40 and not w486;
w488 <= not w38 and w487;
w489 <= not w29 and w488;
w490 <= not in2(107) and in3(107);
w491 <= not in2(106) and in3(106);
w492 <= not w490 and not w491;
w493 <= not in2(105) and in3(105);
w494 <= not in2(104) and in3(104);
w495 <= not w493 and not w494;
w496 <= w492 and w495;
w497 <= not w489 and w496;
w498 <= in2(107) and not in3(107);
w499 <= in2(104) and not in3(104);
w500 <= not w493 and w499;
w501 <= in2(105) and not in3(105);
w502 <= not w500 and not w501;
w503 <= in2(106) and not in3(106);
w504 <= w502 and not w503;
w505 <= w492 and not w504;
w506 <= not w498 and not w505;
w507 <= not w497 and w506;
w508 <= not in2(108) and in3(108);
w509 <= not w21 and not w508;
w510 <= w20 and w509;
w511 <= not w507 and w510;
w512 <= not w28 and not w511;
w513 <= not w26 and w512;
w514 <= not w17 and w513;
w515 <= not w16 and not w514;
w516 <= w15 and w515;
w517 <= not w12 and w516;
w518 <= in2(115) and not in3(115);
w519 <= not in3(112) and not w16;
w520 <= in2(112) and w519;
w521 <= in2(113) and not in3(113);
w522 <= not w520 and not w521;
w523 <= in2(114) and not in3(114);
w524 <= w522 and not w523;
w525 <= w15 and not w524;
w526 <= not w518 and not w525;
w527 <= not w517 and w526;
w528 <= not in2(116) and in3(116);
w529 <= not w4 and not w528;
w530 <= w3 and w529;
w531 <= not w527 and w530;
w532 <= not w11 and not w531;
w533 <= not w9 and w532;
w534 <= not w0 and w533;
w535 <= not in2(123) and in3(123);
w536 <= not in2(122) and in3(122);
w537 <= not w535 and not w536;
w538 <= not in2(121) and in3(121);
w539 <= not in2(120) and in3(120);
w540 <= not w538 and not w539;
w541 <= w537 and w540;
w542 <= not w534 and w541;
w543 <= in2(123) and not in3(123);
w544 <= in2(120) and not in3(120);
w545 <= not w538 and w544;
w546 <= in2(121) and not in3(121);
w547 <= not w545 and not w546;
w548 <= in2(122) and not in3(122);
w549 <= w547 and not w548;
w550 <= w537 and not w549;
w551 <= not w543 and not w550;
w552 <= not w542 and w551;
w553 <= not in2(124) and in3(124);
w554 <= in2(127) and not in3(127);
w555 <= not in2(126) and in3(126);
w556 <= not in2(125) and in3(125);
w557 <= not w555 and not w556;
w558 <= not w554 and w557;
w559 <= not w553 and w558;
w560 <= not w552 and w559;
w561 <= in2(124) and not in3(124);
w562 <= in2(125) and not in3(125);
w563 <= not w561 and not w562;
w564 <= w557 and not w563;
w565 <= in2(126) and not in3(126);
w566 <= not w564 and not w565;
w567 <= not w554 and not w566;
w568 <= not w560 and not w567;
w569 <= not in3(127) and w568;
w570 <= in2(127) and not w569;
w571 <= in0(119) and not in1(119);
w572 <= not in0(119) and in1(119);
w573 <= not in0(118) and in1(118);
w574 <= not w572 and not w573;
w575 <= not in0(117) and in1(117);
w576 <= in0(116) and not in1(116);
w577 <= not w575 and w576;
w578 <= in0(117) and not in1(117);
w579 <= not w577 and not w578;
w580 <= w574 and not w579;
w581 <= not in1(118) and not w572;
w582 <= in0(118) and w581;
w583 <= not in0(112) and in1(112);
w584 <= not in0(115) and in1(115);
w585 <= not in0(114) and in1(114);
w586 <= not w584 and not w585;
w587 <= not in0(113) and in1(113);
w588 <= in0(111) and not in1(111);
w589 <= not in0(111) and in1(111);
w590 <= not in0(110) and in1(110);
w591 <= not w589 and not w590;
w592 <= not in0(109) and in1(109);
w593 <= in0(108) and not in1(108);
w594 <= not w592 and w593;
w595 <= in0(109) and not in1(109);
w596 <= not w594 and not w595;
w597 <= w591 and not w596;
w598 <= not in1(110) and not w589;
w599 <= in0(110) and w598;
w600 <= in0(103) and not in1(103);
w601 <= not in0(103) and in1(103);
w602 <= not in0(102) and in1(102);
w603 <= not w601 and not w602;
w604 <= not in0(101) and in1(101);
w605 <= in0(100) and not in1(100);
w606 <= not w604 and w605;
w607 <= in0(101) and not in1(101);
w608 <= not w606 and not w607;
w609 <= w603 and not w608;
w610 <= not in1(102) and not w601;
w611 <= in0(102) and w610;
w612 <= not in0(96) and in1(96);
w613 <= not in0(99) and in1(99);
w614 <= not in0(98) and in1(98);
w615 <= not w613 and not w614;
w616 <= not in0(97) and in1(97);
w617 <= in0(95) and not in1(95);
w618 <= not in0(95) and in1(95);
w619 <= not in0(94) and in1(94);
w620 <= not w618 and not w619;
w621 <= not in0(93) and in1(93);
w622 <= in0(92) and not in1(92);
w623 <= not w621 and w622;
w624 <= in0(93) and not in1(93);
w625 <= not w623 and not w624;
w626 <= w620 and not w625;
w627 <= not in1(94) and not w618;
w628 <= in0(94) and w627;
w629 <= in0(87) and not in1(87);
w630 <= not in0(87) and in1(87);
w631 <= not in0(86) and in1(86);
w632 <= not w630 and not w631;
w633 <= not in0(85) and in1(85);
w634 <= in0(84) and not in1(84);
w635 <= not w633 and w634;
w636 <= in0(85) and not in1(85);
w637 <= not w635 and not w636;
w638 <= w632 and not w637;
w639 <= not in1(86) and not w630;
w640 <= in0(86) and w639;
w641 <= not in0(80) and in1(80);
w642 <= not in0(83) and in1(83);
w643 <= not in0(82) and in1(82);
w644 <= not w642 and not w643;
w645 <= not in0(81) and in1(81);
w646 <= in0(79) and not in1(79);
w647 <= not in0(79) and in1(79);
w648 <= not in0(78) and in1(78);
w649 <= not w647 and not w648;
w650 <= not in0(77) and in1(77);
w651 <= in0(76) and not in1(76);
w652 <= not w650 and w651;
w653 <= in0(77) and not in1(77);
w654 <= not w652 and not w653;
w655 <= w649 and not w654;
w656 <= not in1(78) and not w647;
w657 <= in0(78) and w656;
w658 <= in0(71) and not in1(71);
w659 <= not in0(71) and in1(71);
w660 <= not in0(70) and in1(70);
w661 <= not w659 and not w660;
w662 <= not in0(69) and in1(69);
w663 <= in0(68) and not in1(68);
w664 <= not w662 and w663;
w665 <= in0(69) and not in1(69);
w666 <= not w664 and not w665;
w667 <= w661 and not w666;
w668 <= not in1(70) and not w659;
w669 <= in0(70) and w668;
w670 <= not in0(67) and in1(67);
w671 <= not in0(66) and in1(66);
w672 <= not w670 and not w671;
w673 <= not in0(65) and in1(65);
w674 <= in0(63) and not in1(63);
w675 <= not in0(63) and in1(63);
w676 <= not in0(62) and in1(62);
w677 <= not w675 and not w676;
w678 <= not in0(60) and in1(60);
w679 <= not in0(61) and in1(61);
w680 <= not w678 and not w679;
w681 <= w677 and w680;
w682 <= in0(59) and not in1(59);
w683 <= not in0(59) and in1(59);
w684 <= not in0(58) and in1(58);
w685 <= not w683 and not w684;
w686 <= not in0(57) and in1(57);
w687 <= in0(56) and not in1(56);
w688 <= not w686 and w687;
w689 <= in0(57) and not in1(57);
w690 <= not w688 and not w689;
w691 <= in0(58) and not in1(58);
w692 <= w690 and not w691;
w693 <= w685 and not w692;
w694 <= not w682 and not w693;
w695 <= w681 and not w694;
w696 <= in0(60) and not in1(60);
w697 <= not w679 and w696;
w698 <= in0(61) and not in1(61);
w699 <= not w697 and not w698;
w700 <= w677 and not w699;
w701 <= not in1(62) and not w675;
w702 <= in0(62) and w701;
w703 <= in0(47) and not in1(47);
w704 <= not in0(47) and in1(47);
w705 <= not in0(46) and in1(46);
w706 <= not w704 and not w705;
w707 <= not in0(44) and in1(44);
w708 <= not in0(45) and in1(45);
w709 <= not w707 and not w708;
w710 <= w706 and w709;
w711 <= in0(43) and not in1(43);
w712 <= not in0(43) and in1(43);
w713 <= not in0(42) and in1(42);
w714 <= not w712 and not w713;
w715 <= not in0(41) and in1(41);
w716 <= in0(40) and not in1(40);
w717 <= not w715 and w716;
w718 <= in0(41) and not in1(41);
w719 <= not w717 and not w718;
w720 <= in0(42) and not in1(42);
w721 <= w719 and not w720;
w722 <= w714 and not w721;
w723 <= not w711 and not w722;
w724 <= w710 and not w723;
w725 <= in0(44) and not in1(44);
w726 <= not w708 and w725;
w727 <= in0(45) and not in1(45);
w728 <= not w726 and not w727;
w729 <= w706 and not w728;
w730 <= not in1(46) and not w704;
w731 <= in0(46) and w730;
w732 <= not in0(32) and in1(32);
w733 <= not in0(31) and in1(31);
w734 <= not in0(30) and in1(30);
w735 <= not in0(29) and in1(29);
w736 <= not in0(28) and in1(28);
w737 <= not in0(27) and in1(27);
w738 <= not in0(26) and in1(26);
w739 <= not in0(23) and in1(23);
w740 <= not in0(22) and in1(22);
w741 <= not in0(21) and in1(21);
w742 <= not in0(20) and in1(20);
w743 <= not in0(19) and in1(19);
w744 <= not in0(18) and in1(18);
w745 <= not in0(15) and in1(15);
w746 <= not in0(14) and in1(14);
w747 <= not in0(13) and in1(13);
w748 <= not in0(12) and in1(12);
w749 <= not in0(11) and in1(11);
w750 <= not in0(10) and in1(10);
w751 <= not in0(7) and in1(7);
w752 <= not in0(6) and in1(6);
w753 <= not in0(3) and in1(3);
w754 <= in0(0) and not in1(0);
w755 <= in0(1) and not in1(1);
w756 <= not w754 and not w755;
w757 <= not in0(2) and in1(2);
w758 <= not in0(1) and in1(1);
w759 <= not w757 and not w758;
w760 <= not w756 and w759;
w761 <= in0(2) and not in1(2);
w762 <= not w760 and not w761;
w763 <= not w753 and not w762;
w764 <= in0(3) and not in1(3);
w765 <= not w763 and not w764;
w766 <= not in0(4) and w765;
w767 <= not in1(4) and not w766;
w768 <= in0(4) and not w765;
w769 <= not w767 and not w768;
w770 <= not in0(5) and w769;
w771 <= not in1(5) and not w770;
w772 <= in0(5) and not w769;
w773 <= not w771 and not w772;
w774 <= not w752 and not w773;
w775 <= in0(6) and not in1(6);
w776 <= not w774 and not w775;
w777 <= not w751 and not w776;
w778 <= in0(7) and not in1(7);
w779 <= not w777 and not w778;
w780 <= not in0(8) and w779;
w781 <= not in1(8) and not w780;
w782 <= in0(8) and not w779;
w783 <= not w781 and not w782;
w784 <= not in0(9) and w783;
w785 <= not in1(9) and not w784;
w786 <= in0(9) and not w783;
w787 <= not w785 and not w786;
w788 <= not w750 and not w787;
w789 <= in0(10) and not in1(10);
w790 <= not w788 and not w789;
w791 <= not w749 and not w790;
w792 <= in0(11) and not in1(11);
w793 <= not w791 and not w792;
w794 <= not w748 and not w793;
w795 <= in0(12) and not in1(12);
w796 <= not w794 and not w795;
w797 <= not w747 and not w796;
w798 <= in0(13) and not in1(13);
w799 <= not w797 and not w798;
w800 <= not w746 and not w799;
w801 <= in0(14) and not in1(14);
w802 <= not w800 and not w801;
w803 <= not w745 and not w802;
w804 <= in0(15) and not in1(15);
w805 <= not w803 and not w804;
w806 <= not in0(16) and w805;
w807 <= not in1(16) and not w806;
w808 <= in0(16) and not w805;
w809 <= not w807 and not w808;
w810 <= not in0(17) and w809;
w811 <= not in1(17) and not w810;
w812 <= in0(17) and not w809;
w813 <= not w811 and not w812;
w814 <= not w744 and not w813;
w815 <= in0(18) and not in1(18);
w816 <= not w814 and not w815;
w817 <= not w743 and not w816;
w818 <= in0(19) and not in1(19);
w819 <= not w817 and not w818;
w820 <= not w742 and not w819;
w821 <= in0(20) and not in1(20);
w822 <= not w820 and not w821;
w823 <= not w741 and not w822;
w824 <= in0(21) and not in1(21);
w825 <= not w823 and not w824;
w826 <= not w740 and not w825;
w827 <= in0(22) and not in1(22);
w828 <= not w826 and not w827;
w829 <= not w739 and not w828;
w830 <= in0(23) and not in1(23);
w831 <= not w829 and not w830;
w832 <= not in0(24) and w831;
w833 <= not in1(24) and not w832;
w834 <= in0(24) and not w831;
w835 <= not w833 and not w834;
w836 <= not in0(25) and w835;
w837 <= not in1(25) and not w836;
w838 <= in0(25) and not w835;
w839 <= not w837 and not w838;
w840 <= not w738 and not w839;
w841 <= in0(26) and not in1(26);
w842 <= not w840 and not w841;
w843 <= not w737 and not w842;
w844 <= in0(27) and not in1(27);
w845 <= not w843 and not w844;
w846 <= not w736 and not w845;
w847 <= in0(28) and not in1(28);
w848 <= not w846 and not w847;
w849 <= not w735 and not w848;
w850 <= in0(29) and not in1(29);
w851 <= not w849 and not w850;
w852 <= not w734 and not w851;
w853 <= in0(30) and not in1(30);
w854 <= not w852 and not w853;
w855 <= not w733 and not w854;
w856 <= in0(31) and not in1(31);
w857 <= not w855 and not w856;
w858 <= not in0(39) and in1(39);
w859 <= not in0(38) and in1(38);
w860 <= not w858 and not w859;
w861 <= not in0(36) and in1(36);
w862 <= not in0(37) and in1(37);
w863 <= not w861 and not w862;
w864 <= w860 and w863;
w865 <= not in0(33) and in1(33);
w866 <= not in0(35) and in1(35);
w867 <= not in0(34) and in1(34);
w868 <= not w866 and not w867;
w869 <= not w865 and w868;
w870 <= w864 and w869;
w871 <= not w857 and w870;
w872 <= not w732 and w871;
w873 <= in0(39) and not in1(39);
w874 <= in0(36) and not in1(36);
w875 <= not w862 and w874;
w876 <= in0(37) and not in1(37);
w877 <= not w875 and not w876;
w878 <= w860 and not w877;
w879 <= not in1(38) and not w858;
w880 <= in0(38) and w879;
w881 <= in0(35) and not in1(35);
w882 <= not in1(32) and not w865;
w883 <= in0(32) and w882;
w884 <= in0(33) and not in1(33);
w885 <= not w883 and not w884;
w886 <= in0(34) and not in1(34);
w887 <= w885 and not w886;
w888 <= w868 and not w887;
w889 <= not w881 and not w888;
w890 <= w864 and not w889;
w891 <= not w880 and not w890;
w892 <= not w878 and w891;
w893 <= not w873 and w892;
w894 <= not w872 and w893;
w895 <= not in0(40) and in1(40);
w896 <= not w715 and not w895;
w897 <= w714 and w896;
w898 <= w710 and w897;
w899 <= not w894 and w898;
w900 <= not w731 and not w899;
w901 <= not w729 and w900;
w902 <= not w724 and w901;
w903 <= not w703 and w902;
w904 <= not in0(48) and in1(48);
w905 <= not in0(55) and in1(55);
w906 <= not in0(54) and in1(54);
w907 <= not w905 and not w906;
w908 <= not in0(53) and in1(53);
w909 <= not in0(52) and in1(52);
w910 <= not w908 and not w909;
w911 <= w907 and w910;
w912 <= not in0(49) and in1(49);
w913 <= not in0(51) and in1(51);
w914 <= not in0(50) and in1(50);
w915 <= not w913 and not w914;
w916 <= not w912 and w915;
w917 <= w911 and w916;
w918 <= not w904 and w917;
w919 <= not w903 and w918;
w920 <= in0(55) and not in1(55);
w921 <= in0(51) and not in1(51);
w922 <= not in1(48) and not w912;
w923 <= in0(48) and w922;
w924 <= in0(49) and not in1(49);
w925 <= not w923 and not w924;
w926 <= in0(50) and not in1(50);
w927 <= w925 and not w926;
w928 <= w915 and not w927;
w929 <= not w921 and not w928;
w930 <= w911 and not w929;
w931 <= in0(52) and not in1(52);
w932 <= not w908 and w931;
w933 <= in0(53) and not in1(53);
w934 <= not w932 and not w933;
w935 <= in0(54) and not in1(54);
w936 <= w934 and not w935;
w937 <= w907 and not w936;
w938 <= not w930 and not w937;
w939 <= not w920 and w938;
w940 <= not w919 and w939;
w941 <= not in0(56) and in1(56);
w942 <= not w686 and not w941;
w943 <= w681 and w942;
w944 <= w685 and w943;
w945 <= not w940 and w944;
w946 <= not w702 and not w945;
w947 <= not w700 and w946;
w948 <= not w695 and w947;
w949 <= not w674 and w948;
w950 <= not in0(64) and in1(64);
w951 <= not w949 and not w950;
w952 <= not w673 and w951;
w953 <= w672 and w952;
w954 <= in0(67) and not in1(67);
w955 <= in0(64) and not in1(64);
w956 <= not w673 and w955;
w957 <= in0(65) and not in1(65);
w958 <= not w956 and not w957;
w959 <= in0(66) and not in1(66);
w960 <= w958 and not w959;
w961 <= w672 and not w960;
w962 <= not w954 and not w961;
w963 <= not w953 and w962;
w964 <= not in0(68) and in1(68);
w965 <= not w662 and not w964;
w966 <= w661 and w965;
w967 <= not w963 and w966;
w968 <= not w669 and not w967;
w969 <= not w667 and w968;
w970 <= not w658 and w969;
w971 <= not in0(75) and in1(75);
w972 <= not in0(74) and in1(74);
w973 <= not w971 and not w972;
w974 <= not in0(73) and in1(73);
w975 <= not in0(72) and in1(72);
w976 <= not w974 and not w975;
w977 <= w973 and w976;
w978 <= not w970 and w977;
w979 <= in0(75) and not in1(75);
w980 <= in0(72) and not in1(72);
w981 <= not w974 and w980;
w982 <= in0(73) and not in1(73);
w983 <= not w981 and not w982;
w984 <= in0(74) and not in1(74);
w985 <= w983 and not w984;
w986 <= w973 and not w985;
w987 <= not w979 and not w986;
w988 <= not w978 and w987;
w989 <= not in0(76) and in1(76);
w990 <= not w650 and not w989;
w991 <= w649 and w990;
w992 <= not w988 and w991;
w993 <= not w657 and not w992;
w994 <= not w655 and w993;
w995 <= not w646 and w994;
w996 <= not w645 and not w995;
w997 <= w644 and w996;
w998 <= not w641 and w997;
w999 <= in0(83) and not in1(83);
w1000 <= not in1(80) and not w645;
w1001 <= in0(80) and w1000;
w1002 <= in0(81) and not in1(81);
w1003 <= not w1001 and not w1002;
w1004 <= in0(82) and not in1(82);
w1005 <= w1003 and not w1004;
w1006 <= w644 and not w1005;
w1007 <= not w999 and not w1006;
w1008 <= not w998 and w1007;
w1009 <= not in0(84) and in1(84);
w1010 <= not w633 and not w1009;
w1011 <= w632 and w1010;
w1012 <= not w1008 and w1011;
w1013 <= not w640 and not w1012;
w1014 <= not w638 and w1013;
w1015 <= not w629 and w1014;
w1016 <= not in0(91) and in1(91);
w1017 <= not in0(90) and in1(90);
w1018 <= not w1016 and not w1017;
w1019 <= not in0(89) and in1(89);
w1020 <= not in0(88) and in1(88);
w1021 <= not w1019 and not w1020;
w1022 <= w1018 and w1021;
w1023 <= not w1015 and w1022;
w1024 <= in0(91) and not in1(91);
w1025 <= in0(88) and not in1(88);
w1026 <= not w1019 and w1025;
w1027 <= in0(89) and not in1(89);
w1028 <= not w1026 and not w1027;
w1029 <= in0(90) and not in1(90);
w1030 <= w1028 and not w1029;
w1031 <= w1018 and not w1030;
w1032 <= not w1024 and not w1031;
w1033 <= not w1023 and w1032;
w1034 <= not in0(92) and in1(92);
w1035 <= not w621 and not w1034;
w1036 <= w620 and w1035;
w1037 <= not w1033 and w1036;
w1038 <= not w628 and not w1037;
w1039 <= not w626 and w1038;
w1040 <= not w617 and w1039;
w1041 <= not w616 and not w1040;
w1042 <= w615 and w1041;
w1043 <= not w612 and w1042;
w1044 <= in0(99) and not in1(99);
w1045 <= not in1(96) and not w616;
w1046 <= in0(96) and w1045;
w1047 <= in0(97) and not in1(97);
w1048 <= not w1046 and not w1047;
w1049 <= in0(98) and not in1(98);
w1050 <= w1048 and not w1049;
w1051 <= w615 and not w1050;
w1052 <= not w1044 and not w1051;
w1053 <= not w1043 and w1052;
w1054 <= not in0(100) and in1(100);
w1055 <= not w604 and not w1054;
w1056 <= w603 and w1055;
w1057 <= not w1053 and w1056;
w1058 <= not w611 and not w1057;
w1059 <= not w609 and w1058;
w1060 <= not w600 and w1059;
w1061 <= not in0(107) and in1(107);
w1062 <= not in0(106) and in1(106);
w1063 <= not w1061 and not w1062;
w1064 <= not in0(105) and in1(105);
w1065 <= not in0(104) and in1(104);
w1066 <= not w1064 and not w1065;
w1067 <= w1063 and w1066;
w1068 <= not w1060 and w1067;
w1069 <= in0(107) and not in1(107);
w1070 <= in0(104) and not in1(104);
w1071 <= not w1064 and w1070;
w1072 <= in0(105) and not in1(105);
w1073 <= not w1071 and not w1072;
w1074 <= in0(106) and not in1(106);
w1075 <= w1073 and not w1074;
w1076 <= w1063 and not w1075;
w1077 <= not w1069 and not w1076;
w1078 <= not w1068 and w1077;
w1079 <= not in0(108) and in1(108);
w1080 <= not w592 and not w1079;
w1081 <= w591 and w1080;
w1082 <= not w1078 and w1081;
w1083 <= not w599 and not w1082;
w1084 <= not w597 and w1083;
w1085 <= not w588 and w1084;
w1086 <= not w587 and not w1085;
w1087 <= w586 and w1086;
w1088 <= not w583 and w1087;
w1089 <= in0(115) and not in1(115);
w1090 <= not in1(112) and not w587;
w1091 <= in0(112) and w1090;
w1092 <= in0(113) and not in1(113);
w1093 <= not w1091 and not w1092;
w1094 <= in0(114) and not in1(114);
w1095 <= w1093 and not w1094;
w1096 <= w586 and not w1095;
w1097 <= not w1089 and not w1096;
w1098 <= not w1088 and w1097;
w1099 <= not in0(116) and in1(116);
w1100 <= not w575 and not w1099;
w1101 <= w574 and w1100;
w1102 <= not w1098 and w1101;
w1103 <= not w582 and not w1102;
w1104 <= not w580 and w1103;
w1105 <= not w571 and w1104;
w1106 <= not in0(123) and in1(123);
w1107 <= not in0(122) and in1(122);
w1108 <= not w1106 and not w1107;
w1109 <= not in0(121) and in1(121);
w1110 <= not in0(120) and in1(120);
w1111 <= not w1109 and not w1110;
w1112 <= w1108 and w1111;
w1113 <= not w1105 and w1112;
w1114 <= in0(123) and not in1(123);
w1115 <= in0(120) and not in1(120);
w1116 <= not w1109 and w1115;
w1117 <= in0(121) and not in1(121);
w1118 <= not w1116 and not w1117;
w1119 <= in0(122) and not in1(122);
w1120 <= w1118 and not w1119;
w1121 <= w1108 and not w1120;
w1122 <= not w1114 and not w1121;
w1123 <= not w1113 and w1122;
w1124 <= not in0(124) and in1(124);
w1125 <= in0(127) and not in1(127);
w1126 <= not in0(126) and in1(126);
w1127 <= not in0(125) and in1(125);
w1128 <= not w1126 and not w1127;
w1129 <= not w1125 and w1128;
w1130 <= not w1124 and w1129;
w1131 <= not w1123 and w1130;
w1132 <= in0(124) and not in1(124);
w1133 <= in0(125) and not in1(125);
w1134 <= not w1132 and not w1133;
w1135 <= w1128 and not w1134;
w1136 <= in0(126) and not in1(126);
w1137 <= not w1135 and not w1136;
w1138 <= not w1125 and not w1137;
w1139 <= not w1131 and not w1138;
w1140 <= not in1(127) and w1139;
w1141 <= in0(127) and not w1140;
w1142 <= w570 and not w1141;
w1143 <= not in0(127) and in1(127);
w1144 <= w1139 and not w1143;
w1145 <= in1(119) and w1144;
w1146 <= in0(119) and not w1144;
w1147 <= not w1145 and not w1146;
w1148 <= not in2(127) and in3(127);
w1149 <= w568 and not w1148;
w1150 <= in3(119) and w1149;
w1151 <= in2(119) and not w1149;
w1152 <= not w1150 and not w1151;
w1153 <= not w1147 and w1152;
w1154 <= w1147 and not w1152;
w1155 <= in3(118) and w1149;
w1156 <= in2(118) and not w1149;
w1157 <= not w1155 and not w1156;
w1158 <= in1(118) and w1144;
w1159 <= in0(118) and not w1144;
w1160 <= not w1158 and not w1159;
w1161 <= not w1157 and w1160;
w1162 <= not w1154 and not w1161;
w1163 <= in1(116) and w1144;
w1164 <= in0(116) and not w1144;
w1165 <= not w1163 and not w1164;
w1166 <= in1(117) and w1144;
w1167 <= in0(117) and not w1144;
w1168 <= not w1166 and not w1167;
w1169 <= in3(117) and w1149;
w1170 <= in2(117) and not w1149;
w1171 <= not w1169 and not w1170;
w1172 <= w1168 and not w1171;
w1173 <= in3(116) and w1149;
w1174 <= in2(116) and not w1149;
w1175 <= not w1173 and not w1174;
w1176 <= not w1172 and w1175;
w1177 <= not w1165 and w1176;
w1178 <= not w1168 and w1171;
w1179 <= not w1177 and not w1178;
w1180 <= w1162 and not w1179;
w1181 <= w1157 and not w1160;
w1182 <= not w1154 and w1181;
w1183 <= in3(112) and w1149;
w1184 <= in2(112) and not w1149;
w1185 <= not w1183 and not w1184;
w1186 <= in1(112) and w1144;
w1187 <= in0(112) and not w1144;
w1188 <= not w1186 and not w1187;
w1189 <= not w1185 and w1188;
w1190 <= in1(115) and w1144;
w1191 <= in0(115) and not w1144;
w1192 <= not w1190 and not w1191;
w1193 <= in3(115) and w1149;
w1194 <= in2(115) and not w1149;
w1195 <= not w1193 and not w1194;
w1196 <= w1192 and not w1195;
w1197 <= in3(114) and w1149;
w1198 <= in2(114) and not w1149;
w1199 <= not w1197 and not w1198;
w1200 <= in1(114) and w1144;
w1201 <= in0(114) and not w1144;
w1202 <= not w1200 and not w1201;
w1203 <= not w1199 and w1202;
w1204 <= not w1196 and not w1203;
w1205 <= in1(113) and w1144;
w1206 <= in0(113) and not w1144;
w1207 <= not w1205 and not w1206;
w1208 <= in3(113) and w1149;
w1209 <= in2(113) and not w1149;
w1210 <= not w1208 and not w1209;
w1211 <= w1207 and not w1210;
w1212 <= in1(111) and w1144;
w1213 <= in0(111) and not w1144;
w1214 <= not w1212 and not w1213;
w1215 <= in3(111) and w1149;
w1216 <= in2(111) and not w1149;
w1217 <= not w1215 and not w1216;
w1218 <= not w1214 and w1217;
w1219 <= w1214 and not w1217;
w1220 <= in3(110) and w1149;
w1221 <= in2(110) and not w1149;
w1222 <= not w1220 and not w1221;
w1223 <= in1(110) and w1144;
w1224 <= in0(110) and not w1144;
w1225 <= not w1223 and not w1224;
w1226 <= not w1222 and w1225;
w1227 <= not w1219 and not w1226;
w1228 <= in1(109) and w1144;
w1229 <= in0(109) and not w1144;
w1230 <= not w1228 and not w1229;
w1231 <= in3(109) and w1149;
w1232 <= in2(109) and not w1149;
w1233 <= not w1231 and not w1232;
w1234 <= w1230 and not w1233;
w1235 <= in1(108) and w1144;
w1236 <= in0(108) and not w1144;
w1237 <= not w1235 and not w1236;
w1238 <= in3(108) and w1149;
w1239 <= in2(108) and not w1149;
w1240 <= not w1238 and not w1239;
w1241 <= not w1237 and w1240;
w1242 <= not w1234 and w1241;
w1243 <= not w1230 and w1233;
w1244 <= not w1242 and not w1243;
w1245 <= w1227 and not w1244;
w1246 <= w1222 and not w1225;
w1247 <= not w1219 and w1246;
w1248 <= in1(103) and w1144;
w1249 <= in0(103) and not w1144;
w1250 <= not w1248 and not w1249;
w1251 <= in3(103) and w1149;
w1252 <= in2(103) and not w1149;
w1253 <= not w1251 and not w1252;
w1254 <= not w1250 and w1253;
w1255 <= w1250 and not w1253;
w1256 <= in3(102) and w1149;
w1257 <= in2(102) and not w1149;
w1258 <= not w1256 and not w1257;
w1259 <= in1(102) and w1144;
w1260 <= in0(102) and not w1144;
w1261 <= not w1259 and not w1260;
w1262 <= not w1258 and w1261;
w1263 <= not w1255 and not w1262;
w1264 <= in1(101) and w1144;
w1265 <= in0(101) and not w1144;
w1266 <= not w1264 and not w1265;
w1267 <= in3(101) and w1149;
w1268 <= in2(101) and not w1149;
w1269 <= not w1267 and not w1268;
w1270 <= w1266 and not w1269;
w1271 <= in1(100) and w1144;
w1272 <= in0(100) and not w1144;
w1273 <= not w1271 and not w1272;
w1274 <= in3(100) and w1149;
w1275 <= in2(100) and not w1149;
w1276 <= not w1274 and not w1275;
w1277 <= not w1273 and w1276;
w1278 <= not w1270 and w1277;
w1279 <= not w1266 and w1269;
w1280 <= not w1278 and not w1279;
w1281 <= w1263 and not w1280;
w1282 <= w1258 and not w1261;
w1283 <= not w1255 and w1282;
w1284 <= in3(96) and w1149;
w1285 <= in2(96) and not w1149;
w1286 <= not w1284 and not w1285;
w1287 <= in1(96) and w1144;
w1288 <= in0(96) and not w1144;
w1289 <= not w1287 and not w1288;
w1290 <= not w1286 and w1289;
w1291 <= in1(99) and w1144;
w1292 <= in0(99) and not w1144;
w1293 <= not w1291 and not w1292;
w1294 <= in3(99) and w1149;
w1295 <= in2(99) and not w1149;
w1296 <= not w1294 and not w1295;
w1297 <= w1293 and not w1296;
w1298 <= in3(98) and w1149;
w1299 <= in2(98) and not w1149;
w1300 <= not w1298 and not w1299;
w1301 <= in1(98) and w1144;
w1302 <= in0(98) and not w1144;
w1303 <= not w1301 and not w1302;
w1304 <= not w1300 and w1303;
w1305 <= not w1297 and not w1304;
w1306 <= in1(97) and w1144;
w1307 <= in0(97) and not w1144;
w1308 <= not w1306 and not w1307;
w1309 <= in3(97) and w1149;
w1310 <= in2(97) and not w1149;
w1311 <= not w1309 and not w1310;
w1312 <= w1308 and not w1311;
w1313 <= in1(95) and w1144;
w1314 <= in0(95) and not w1144;
w1315 <= not w1313 and not w1314;
w1316 <= in3(95) and w1149;
w1317 <= in2(95) and not w1149;
w1318 <= not w1316 and not w1317;
w1319 <= not w1315 and w1318;
w1320 <= w1315 and not w1318;
w1321 <= in3(94) and w1149;
w1322 <= in2(94) and not w1149;
w1323 <= not w1321 and not w1322;
w1324 <= in1(94) and w1144;
w1325 <= in0(94) and not w1144;
w1326 <= not w1324 and not w1325;
w1327 <= not w1323 and w1326;
w1328 <= not w1320 and not w1327;
w1329 <= in1(93) and w1144;
w1330 <= in0(93) and not w1144;
w1331 <= not w1329 and not w1330;
w1332 <= in3(93) and w1149;
w1333 <= in2(93) and not w1149;
w1334 <= not w1332 and not w1333;
w1335 <= w1331 and not w1334;
w1336 <= in1(92) and w1144;
w1337 <= in0(92) and not w1144;
w1338 <= not w1336 and not w1337;
w1339 <= in3(92) and w1149;
w1340 <= in2(92) and not w1149;
w1341 <= not w1339 and not w1340;
w1342 <= not w1338 and w1341;
w1343 <= not w1335 and w1342;
w1344 <= not w1331 and w1334;
w1345 <= not w1343 and not w1344;
w1346 <= w1328 and not w1345;
w1347 <= w1323 and not w1326;
w1348 <= not w1320 and w1347;
w1349 <= in1(87) and w1144;
w1350 <= in0(87) and not w1144;
w1351 <= not w1349 and not w1350;
w1352 <= in3(87) and w1149;
w1353 <= in2(87) and not w1149;
w1354 <= not w1352 and not w1353;
w1355 <= not w1351 and w1354;
w1356 <= w1351 and not w1354;
w1357 <= in3(86) and w1149;
w1358 <= in2(86) and not w1149;
w1359 <= not w1357 and not w1358;
w1360 <= in1(86) and w1144;
w1361 <= in0(86) and not w1144;
w1362 <= not w1360 and not w1361;
w1363 <= not w1359 and w1362;
w1364 <= not w1356 and not w1363;
w1365 <= in1(85) and w1144;
w1366 <= in0(85) and not w1144;
w1367 <= not w1365 and not w1366;
w1368 <= in3(85) and w1149;
w1369 <= in2(85) and not w1149;
w1370 <= not w1368 and not w1369;
w1371 <= w1367 and not w1370;
w1372 <= in1(84) and w1144;
w1373 <= in0(84) and not w1144;
w1374 <= not w1372 and not w1373;
w1375 <= in3(84) and w1149;
w1376 <= in2(84) and not w1149;
w1377 <= not w1375 and not w1376;
w1378 <= not w1374 and w1377;
w1379 <= not w1371 and w1378;
w1380 <= not w1367 and w1370;
w1381 <= not w1379 and not w1380;
w1382 <= w1364 and not w1381;
w1383 <= w1359 and not w1362;
w1384 <= not w1356 and w1383;
w1385 <= in3(80) and w1149;
w1386 <= in2(80) and not w1149;
w1387 <= not w1385 and not w1386;
w1388 <= in1(80) and w1144;
w1389 <= in0(80) and not w1144;
w1390 <= not w1388 and not w1389;
w1391 <= not w1387 and w1390;
w1392 <= in1(83) and w1144;
w1393 <= in0(83) and not w1144;
w1394 <= not w1392 and not w1393;
w1395 <= in3(83) and w1149;
w1396 <= in2(83) and not w1149;
w1397 <= not w1395 and not w1396;
w1398 <= w1394 and not w1397;
w1399 <= in3(82) and w1149;
w1400 <= in2(82) and not w1149;
w1401 <= not w1399 and not w1400;
w1402 <= in1(82) and w1144;
w1403 <= in0(82) and not w1144;
w1404 <= not w1402 and not w1403;
w1405 <= not w1401 and w1404;
w1406 <= not w1398 and not w1405;
w1407 <= in1(81) and w1144;
w1408 <= in0(81) and not w1144;
w1409 <= not w1407 and not w1408;
w1410 <= in3(81) and w1149;
w1411 <= in2(81) and not w1149;
w1412 <= not w1410 and not w1411;
w1413 <= w1409 and not w1412;
w1414 <= in1(79) and w1144;
w1415 <= in0(79) and not w1144;
w1416 <= not w1414 and not w1415;
w1417 <= in3(79) and w1149;
w1418 <= in2(79) and not w1149;
w1419 <= not w1417 and not w1418;
w1420 <= not w1416 and w1419;
w1421 <= w1416 and not w1419;
w1422 <= in3(78) and w1149;
w1423 <= in2(78) and not w1149;
w1424 <= not w1422 and not w1423;
w1425 <= in1(78) and w1144;
w1426 <= in0(78) and not w1144;
w1427 <= not w1425 and not w1426;
w1428 <= not w1424 and w1427;
w1429 <= not w1421 and not w1428;
w1430 <= in1(77) and w1144;
w1431 <= in0(77) and not w1144;
w1432 <= not w1430 and not w1431;
w1433 <= in3(77) and w1149;
w1434 <= in2(77) and not w1149;
w1435 <= not w1433 and not w1434;
w1436 <= w1432 and not w1435;
w1437 <= in1(76) and w1144;
w1438 <= in0(76) and not w1144;
w1439 <= not w1437 and not w1438;
w1440 <= in3(76) and w1149;
w1441 <= in2(76) and not w1149;
w1442 <= not w1440 and not w1441;
w1443 <= not w1439 and w1442;
w1444 <= not w1436 and w1443;
w1445 <= not w1432 and w1435;
w1446 <= not w1444 and not w1445;
w1447 <= w1429 and not w1446;
w1448 <= w1424 and not w1427;
w1449 <= not w1421 and w1448;
w1450 <= in1(71) and w1144;
w1451 <= in0(71) and not w1144;
w1452 <= not w1450 and not w1451;
w1453 <= in3(71) and w1149;
w1454 <= in2(71) and not w1149;
w1455 <= not w1453 and not w1454;
w1456 <= not w1452 and w1455;
w1457 <= w1452 and not w1455;
w1458 <= in3(70) and w1149;
w1459 <= in2(70) and not w1149;
w1460 <= not w1458 and not w1459;
w1461 <= in1(70) and w1144;
w1462 <= in0(70) and not w1144;
w1463 <= not w1461 and not w1462;
w1464 <= not w1460 and w1463;
w1465 <= not w1457 and not w1464;
w1466 <= in1(69) and w1144;
w1467 <= in0(69) and not w1144;
w1468 <= not w1466 and not w1467;
w1469 <= in3(69) and w1149;
w1470 <= in2(69) and not w1149;
w1471 <= not w1469 and not w1470;
w1472 <= w1468 and not w1471;
w1473 <= in1(68) and w1144;
w1474 <= in0(68) and not w1144;
w1475 <= not w1473 and not w1474;
w1476 <= in3(68) and w1149;
w1477 <= in2(68) and not w1149;
w1478 <= not w1476 and not w1477;
w1479 <= not w1475 and w1478;
w1480 <= not w1472 and w1479;
w1481 <= not w1468 and w1471;
w1482 <= not w1480 and not w1481;
w1483 <= w1465 and not w1482;
w1484 <= w1460 and not w1463;
w1485 <= not w1457 and w1484;
w1486 <= in1(67) and w1144;
w1487 <= in0(67) and not w1144;
w1488 <= not w1486 and not w1487;
w1489 <= in3(67) and w1149;
w1490 <= in2(67) and not w1149;
w1491 <= not w1489 and not w1490;
w1492 <= w1488 and not w1491;
w1493 <= in3(66) and w1149;
w1494 <= in2(66) and not w1149;
w1495 <= not w1493 and not w1494;
w1496 <= in1(66) and w1144;
w1497 <= in0(66) and not w1144;
w1498 <= not w1496 and not w1497;
w1499 <= not w1495 and w1498;
w1500 <= not w1492 and not w1499;
w1501 <= in3(64) and w1149;
w1502 <= in2(64) and not w1149;
w1503 <= not w1501 and not w1502;
w1504 <= in1(64) and w1144;
w1505 <= in0(64) and not w1144;
w1506 <= not w1504 and not w1505;
w1507 <= not w1503 and w1506;
w1508 <= in1(65) and w1144;
w1509 <= in0(65) and not w1144;
w1510 <= not w1508 and not w1509;
w1511 <= in3(65) and w1149;
w1512 <= in2(65) and not w1149;
w1513 <= not w1511 and not w1512;
w1514 <= w1510 and not w1513;
w1515 <= in1(63) and w1144;
w1516 <= in0(63) and not w1144;
w1517 <= not w1515 and not w1516;
w1518 <= in3(63) and w1149;
w1519 <= in2(63) and not w1149;
w1520 <= not w1518 and not w1519;
w1521 <= not w1517 and w1520;
w1522 <= w1517 and not w1520;
w1523 <= in3(62) and w1149;
w1524 <= in2(62) and not w1149;
w1525 <= not w1523 and not w1524;
w1526 <= in1(62) and w1144;
w1527 <= in0(62) and not w1144;
w1528 <= not w1526 and not w1527;
w1529 <= not w1525 and w1528;
w1530 <= not w1522 and not w1529;
w1531 <= in1(60) and w1144;
w1532 <= in0(60) and not w1144;
w1533 <= not w1531 and not w1532;
w1534 <= in3(60) and w1149;
w1535 <= in2(60) and not w1149;
w1536 <= not w1534 and not w1535;
w1537 <= w1533 and not w1536;
w1538 <= in1(61) and w1144;
w1539 <= in0(61) and not w1144;
w1540 <= not w1538 and not w1539;
w1541 <= in3(61) and w1149;
w1542 <= in2(61) and not w1149;
w1543 <= not w1541 and not w1542;
w1544 <= w1540 and not w1543;
w1545 <= not w1537 and not w1544;
w1546 <= w1530 and w1545;
w1547 <= in1(59) and w1144;
w1548 <= in0(59) and not w1144;
w1549 <= not w1547 and not w1548;
w1550 <= in3(59) and w1149;
w1551 <= in2(59) and not w1149;
w1552 <= not w1550 and not w1551;
w1553 <= not w1549 and w1552;
w1554 <= w1549 and not w1552;
w1555 <= in1(58) and w1144;
w1556 <= in0(58) and not w1144;
w1557 <= not w1555 and not w1556;
w1558 <= in3(58) and w1149;
w1559 <= in2(58) and not w1149;
w1560 <= not w1558 and not w1559;
w1561 <= w1557 and not w1560;
w1562 <= not w1554 and not w1561;
w1563 <= in1(57) and w1144;
w1564 <= in0(57) and not w1144;
w1565 <= not w1563 and not w1564;
w1566 <= in3(57) and w1149;
w1567 <= in2(57) and not w1149;
w1568 <= not w1566 and not w1567;
w1569 <= w1565 and not w1568;
w1570 <= in1(56) and w1144;
w1571 <= in0(56) and not w1144;
w1572 <= not w1570 and not w1571;
w1573 <= in3(56) and w1149;
w1574 <= in2(56) and not w1149;
w1575 <= not w1573 and not w1574;
w1576 <= not w1572 and w1575;
w1577 <= not w1569 and w1576;
w1578 <= not w1565 and w1568;
w1579 <= not w1577 and not w1578;
w1580 <= not w1557 and w1560;
w1581 <= w1579 and not w1580;
w1582 <= w1562 and not w1581;
w1583 <= not w1553 and not w1582;
w1584 <= w1546 and not w1583;
w1585 <= not w1533 and w1536;
w1586 <= not w1544 and w1585;
w1587 <= not w1540 and w1543;
w1588 <= not w1586 and not w1587;
w1589 <= w1530 and not w1588;
w1590 <= w1525 and not w1528;
w1591 <= not w1522 and w1590;
w1592 <= in1(47) and w1144;
w1593 <= in0(47) and not w1144;
w1594 <= not w1592 and not w1593;
w1595 <= in3(47) and w1149;
w1596 <= in2(47) and not w1149;
w1597 <= not w1595 and not w1596;
w1598 <= not w1594 and w1597;
w1599 <= w1594 and not w1597;
w1600 <= in3(46) and w1149;
w1601 <= in2(46) and not w1149;
w1602 <= not w1600 and not w1601;
w1603 <= in1(46) and w1144;
w1604 <= in0(46) and not w1144;
w1605 <= not w1603 and not w1604;
w1606 <= not w1602 and w1605;
w1607 <= not w1599 and not w1606;
w1608 <= in1(44) and w1144;
w1609 <= in0(44) and not w1144;
w1610 <= not w1608 and not w1609;
w1611 <= in3(44) and w1149;
w1612 <= in2(44) and not w1149;
w1613 <= not w1611 and not w1612;
w1614 <= w1610 and not w1613;
w1615 <= in1(45) and w1144;
w1616 <= in0(45) and not w1144;
w1617 <= not w1615 and not w1616;
w1618 <= in3(45) and w1149;
w1619 <= in2(45) and not w1149;
w1620 <= not w1618 and not w1619;
w1621 <= w1617 and not w1620;
w1622 <= not w1614 and not w1621;
w1623 <= w1607 and w1622;
w1624 <= in1(43) and w1144;
w1625 <= in0(43) and not w1144;
w1626 <= not w1624 and not w1625;
w1627 <= in3(43) and w1149;
w1628 <= in2(43) and not w1149;
w1629 <= not w1627 and not w1628;
w1630 <= not w1626 and w1629;
w1631 <= w1626 and not w1629;
w1632 <= in1(42) and w1144;
w1633 <= in0(42) and not w1144;
w1634 <= not w1632 and not w1633;
w1635 <= in3(42) and w1149;
w1636 <= in2(42) and not w1149;
w1637 <= not w1635 and not w1636;
w1638 <= w1634 and not w1637;
w1639 <= not w1631 and not w1638;
w1640 <= in1(41) and w1144;
w1641 <= in0(41) and not w1144;
w1642 <= not w1640 and not w1641;
w1643 <= in3(41) and w1149;
w1644 <= in2(41) and not w1149;
w1645 <= not w1643 and not w1644;
w1646 <= w1642 and not w1645;
w1647 <= in1(40) and w1144;
w1648 <= in0(40) and not w1144;
w1649 <= not w1647 and not w1648;
w1650 <= in3(40) and w1149;
w1651 <= in2(40) and not w1149;
w1652 <= not w1650 and not w1651;
w1653 <= not w1649 and w1652;
w1654 <= not w1646 and w1653;
w1655 <= not w1642 and w1645;
w1656 <= not w1654 and not w1655;
w1657 <= not w1634 and w1637;
w1658 <= w1656 and not w1657;
w1659 <= w1639 and not w1658;
w1660 <= not w1630 and not w1659;
w1661 <= w1623 and not w1660;
w1662 <= not w1610 and w1613;
w1663 <= not w1621 and w1662;
w1664 <= not w1617 and w1620;
w1665 <= not w1663 and not w1664;
w1666 <= w1607 and not w1665;
w1667 <= w1602 and not w1605;
w1668 <= not w1599 and w1667;
w1669 <= in3(32) and w1149;
w1670 <= in2(32) and not w1149;
w1671 <= not w1669 and not w1670;
w1672 <= in1(32) and w1144;
w1673 <= in0(32) and not w1144;
w1674 <= not w1672 and not w1673;
w1675 <= not w1671 and w1674;
w1676 <= in1(31) and w1144;
w1677 <= in0(31) and not w1144;
w1678 <= not w1676 and not w1677;
w1679 <= in3(31) and w1149;
w1680 <= in2(31) and not w1149;
w1681 <= not w1679 and not w1680;
w1682 <= w1678 and not w1681;
w1683 <= in1(30) and w1144;
w1684 <= in0(30) and not w1144;
w1685 <= not w1683 and not w1684;
w1686 <= in3(30) and w1149;
w1687 <= in2(30) and not w1149;
w1688 <= not w1686 and not w1687;
w1689 <= w1685 and not w1688;
w1690 <= in1(29) and w1144;
w1691 <= in0(29) and not w1144;
w1692 <= not w1690 and not w1691;
w1693 <= in3(29) and w1149;
w1694 <= in2(29) and not w1149;
w1695 <= not w1693 and not w1694;
w1696 <= w1692 and not w1695;
w1697 <= in1(28) and w1144;
w1698 <= in0(28) and not w1144;
w1699 <= not w1697 and not w1698;
w1700 <= in3(28) and w1149;
w1701 <= in2(28) and not w1149;
w1702 <= not w1700 and not w1701;
w1703 <= w1699 and not w1702;
w1704 <= in1(27) and w1144;
w1705 <= in0(27) and not w1144;
w1706 <= not w1704 and not w1705;
w1707 <= in3(27) and w1149;
w1708 <= in2(27) and not w1149;
w1709 <= not w1707 and not w1708;
w1710 <= w1706 and not w1709;
w1711 <= in1(26) and w1144;
w1712 <= in0(26) and not w1144;
w1713 <= not w1711 and not w1712;
w1714 <= in3(26) and w1149;
w1715 <= in2(26) and not w1149;
w1716 <= not w1714 and not w1715;
w1717 <= w1713 and not w1716;
w1718 <= in3(25) and w1149;
w1719 <= in2(25) and not w1149;
w1720 <= not w1718 and not w1719;
w1721 <= in3(24) and w1149;
w1722 <= in2(24) and not w1149;
w1723 <= not w1721 and not w1722;
w1724 <= in1(23) and w1144;
w1725 <= in0(23) and not w1144;
w1726 <= not w1724 and not w1725;
w1727 <= in3(23) and w1149;
w1728 <= in2(23) and not w1149;
w1729 <= not w1727 and not w1728;
w1730 <= w1726 and not w1729;
w1731 <= in1(22) and w1144;
w1732 <= in0(22) and not w1144;
w1733 <= not w1731 and not w1732;
w1734 <= in3(22) and w1149;
w1735 <= in2(22) and not w1149;
w1736 <= not w1734 and not w1735;
w1737 <= w1733 and not w1736;
w1738 <= in1(21) and w1144;
w1739 <= in0(21) and not w1144;
w1740 <= not w1738 and not w1739;
w1741 <= in3(21) and w1149;
w1742 <= in2(21) and not w1149;
w1743 <= not w1741 and not w1742;
w1744 <= w1740 and not w1743;
w1745 <= in1(20) and w1144;
w1746 <= in0(20) and not w1144;
w1747 <= not w1745 and not w1746;
w1748 <= in3(20) and w1149;
w1749 <= in2(20) and not w1149;
w1750 <= not w1748 and not w1749;
w1751 <= w1747 and not w1750;
w1752 <= in1(19) and w1144;
w1753 <= in0(19) and not w1144;
w1754 <= not w1752 and not w1753;
w1755 <= in3(19) and w1149;
w1756 <= in2(19) and not w1149;
w1757 <= not w1755 and not w1756;
w1758 <= w1754 and not w1757;
w1759 <= in1(18) and w1144;
w1760 <= in0(18) and not w1144;
w1761 <= not w1759 and not w1760;
w1762 <= in3(18) and w1149;
w1763 <= in2(18) and not w1149;
w1764 <= not w1762 and not w1763;
w1765 <= w1761 and not w1764;
w1766 <= in3(17) and w1149;
w1767 <= in2(17) and not w1149;
w1768 <= not w1766 and not w1767;
w1769 <= in3(16) and w1149;
w1770 <= in2(16) and not w1149;
w1771 <= not w1769 and not w1770;
w1772 <= in1(15) and w1144;
w1773 <= in0(15) and not w1144;
w1774 <= not w1772 and not w1773;
w1775 <= in3(15) and w1149;
w1776 <= in2(15) and not w1149;
w1777 <= not w1775 and not w1776;
w1778 <= w1774 and not w1777;
w1779 <= in1(14) and w1144;
w1780 <= in0(14) and not w1144;
w1781 <= not w1779 and not w1780;
w1782 <= in3(14) and w1149;
w1783 <= in2(14) and not w1149;
w1784 <= not w1782 and not w1783;
w1785 <= w1781 and not w1784;
w1786 <= in1(13) and w1144;
w1787 <= in0(13) and not w1144;
w1788 <= not w1786 and not w1787;
w1789 <= in3(13) and w1149;
w1790 <= in2(13) and not w1149;
w1791 <= not w1789 and not w1790;
w1792 <= w1788 and not w1791;
w1793 <= in1(12) and w1144;
w1794 <= in0(12) and not w1144;
w1795 <= not w1793 and not w1794;
w1796 <= in3(12) and w1149;
w1797 <= in2(12) and not w1149;
w1798 <= not w1796 and not w1797;
w1799 <= w1795 and not w1798;
w1800 <= in1(11) and w1144;
w1801 <= in0(11) and not w1144;
w1802 <= not w1800 and not w1801;
w1803 <= in3(11) and w1149;
w1804 <= in2(11) and not w1149;
w1805 <= not w1803 and not w1804;
w1806 <= w1802 and not w1805;
w1807 <= in1(10) and w1144;
w1808 <= in0(10) and not w1144;
w1809 <= not w1807 and not w1808;
w1810 <= in3(10) and w1149;
w1811 <= in2(10) and not w1149;
w1812 <= not w1810 and not w1811;
w1813 <= w1809 and not w1812;
w1814 <= in3(9) and w1149;
w1815 <= in2(9) and not w1149;
w1816 <= not w1814 and not w1815;
w1817 <= in3(8) and w1149;
w1818 <= in2(8) and not w1149;
w1819 <= not w1817 and not w1818;
w1820 <= in1(7) and w1144;
w1821 <= in0(7) and not w1144;
w1822 <= not w1820 and not w1821;
w1823 <= in3(7) and w1149;
w1824 <= in2(7) and not w1149;
w1825 <= not w1823 and not w1824;
w1826 <= w1822 and not w1825;
w1827 <= in3(6) and w1149;
w1828 <= in2(6) and not w1149;
w1829 <= not w1827 and not w1828;
w1830 <= in1(6) and w1144;
w1831 <= in0(6) and not w1144;
w1832 <= not w1830 and not w1831;
w1833 <= in3(5) and w1149;
w1834 <= in2(5) and not w1149;
w1835 <= not w1833 and not w1834;
w1836 <= in1(5) and w1144;
w1837 <= in0(5) and not w1144;
w1838 <= not w1836 and not w1837;
w1839 <= in3(4) and w1149;
w1840 <= in2(4) and not w1149;
w1841 <= not w1839 and not w1840;
w1842 <= in1(4) and w1144;
w1843 <= in0(4) and not w1144;
w1844 <= not w1842 and not w1843;
w1845 <= in1(3) and w1144;
w1846 <= in0(3) and not w1144;
w1847 <= not w1845 and not w1846;
w1848 <= in3(3) and w1149;
w1849 <= in2(3) and not w1149;
w1850 <= not w1848 and not w1849;
w1851 <= w1847 and not w1850;
w1852 <= in3(1) and w1149;
w1853 <= in2(1) and not w1149;
w1854 <= not w1852 and not w1853;
w1855 <= in1(0) and w1144;
w1856 <= in0(0) and not w1144;
w1857 <= not w1855 and not w1856;
w1858 <= in3(0) and w1149;
w1859 <= in2(0) and not w1149;
w1860 <= not w1858 and not w1859;
w1861 <= not w1857 and w1860;
w1862 <= w1854 and w1861;
w1863 <= in1(1) and w1144;
w1864 <= in0(1) and not w1144;
w1865 <= not w1863 and not w1864;
w1866 <= not w1862 and w1865;
w1867 <= in1(2) and w1144;
w1868 <= in0(2) and not w1144;
w1869 <= not w1867 and not w1868;
w1870 <= in3(2) and w1149;
w1871 <= in2(2) and not w1149;
w1872 <= not w1870 and not w1871;
w1873 <= w1869 and not w1872;
w1874 <= not w1854 and not w1861;
w1875 <= not w1873 and not w1874;
w1876 <= not w1866 and w1875;
w1877 <= not w1869 and w1872;
w1878 <= not w1876 and not w1877;
w1879 <= not w1851 and not w1878;
w1880 <= not w1847 and w1850;
w1881 <= not w1879 and not w1880;
w1882 <= w1844 and w1881;
w1883 <= w1841 and not w1882;
w1884 <= not w1844 and not w1881;
w1885 <= not w1883 and not w1884;
w1886 <= w1838 and w1885;
w1887 <= w1835 and not w1886;
w1888 <= not w1838 and not w1885;
w1889 <= not w1887 and not w1888;
w1890 <= w1832 and w1889;
w1891 <= w1829 and not w1890;
w1892 <= not w1832 and not w1889;
w1893 <= not w1891 and not w1892;
w1894 <= not w1826 and not w1893;
w1895 <= not w1822 and w1825;
w1896 <= not w1894 and not w1895;
w1897 <= in1(8) and w1144;
w1898 <= in0(8) and not w1144;
w1899 <= not w1897 and not w1898;
w1900 <= w1896 and w1899;
w1901 <= w1819 and not w1900;
w1902 <= not w1896 and not w1899;
w1903 <= not w1901 and not w1902;
w1904 <= in1(9) and w1144;
w1905 <= in0(9) and not w1144;
w1906 <= not w1904 and not w1905;
w1907 <= w1903 and w1906;
w1908 <= w1816 and not w1907;
w1909 <= not w1903 and not w1906;
w1910 <= not w1908 and not w1909;
w1911 <= not w1813 and not w1910;
w1912 <= not w1809 and w1812;
w1913 <= not w1911 and not w1912;
w1914 <= not w1806 and not w1913;
w1915 <= not w1802 and w1805;
w1916 <= not w1914 and not w1915;
w1917 <= not w1799 and not w1916;
w1918 <= not w1795 and w1798;
w1919 <= not w1917 and not w1918;
w1920 <= not w1792 and not w1919;
w1921 <= not w1788 and w1791;
w1922 <= not w1920 and not w1921;
w1923 <= not w1785 and not w1922;
w1924 <= not w1781 and w1784;
w1925 <= not w1923 and not w1924;
w1926 <= not w1778 and not w1925;
w1927 <= not w1774 and w1777;
w1928 <= not w1926 and not w1927;
w1929 <= in1(16) and w1144;
w1930 <= in0(16) and not w1144;
w1931 <= not w1929 and not w1930;
w1932 <= w1928 and w1931;
w1933 <= w1771 and not w1932;
w1934 <= not w1928 and not w1931;
w1935 <= not w1933 and not w1934;
w1936 <= in1(17) and w1144;
w1937 <= in0(17) and not w1144;
w1938 <= not w1936 and not w1937;
w1939 <= w1935 and w1938;
w1940 <= w1768 and not w1939;
w1941 <= not w1935 and not w1938;
w1942 <= not w1940 and not w1941;
w1943 <= not w1765 and not w1942;
w1944 <= not w1761 and w1764;
w1945 <= not w1943 and not w1944;
w1946 <= not w1758 and not w1945;
w1947 <= not w1754 and w1757;
w1948 <= not w1946 and not w1947;
w1949 <= not w1751 and not w1948;
w1950 <= not w1747 and w1750;
w1951 <= not w1949 and not w1950;
w1952 <= not w1744 and not w1951;
w1953 <= not w1740 and w1743;
w1954 <= not w1952 and not w1953;
w1955 <= not w1737 and not w1954;
w1956 <= not w1733 and w1736;
w1957 <= not w1955 and not w1956;
w1958 <= not w1730 and not w1957;
w1959 <= not w1726 and w1729;
w1960 <= not w1958 and not w1959;
w1961 <= in1(24) and w1144;
w1962 <= in0(24) and not w1144;
w1963 <= not w1961 and not w1962;
w1964 <= w1960 and w1963;
w1965 <= w1723 and not w1964;
w1966 <= not w1960 and not w1963;
w1967 <= not w1965 and not w1966;
w1968 <= in1(25) and w1144;
w1969 <= in0(25) and not w1144;
w1970 <= not w1968 and not w1969;
w1971 <= w1967 and w1970;
w1972 <= w1720 and not w1971;
w1973 <= not w1967 and not w1970;
w1974 <= not w1972 and not w1973;
w1975 <= not w1717 and not w1974;
w1976 <= not w1713 and w1716;
w1977 <= not w1975 and not w1976;
w1978 <= not w1710 and not w1977;
w1979 <= not w1706 and w1709;
w1980 <= not w1978 and not w1979;
w1981 <= not w1703 and not w1980;
w1982 <= not w1699 and w1702;
w1983 <= not w1981 and not w1982;
w1984 <= not w1696 and not w1983;
w1985 <= not w1692 and w1695;
w1986 <= not w1984 and not w1985;
w1987 <= not w1689 and not w1986;
w1988 <= not w1685 and w1688;
w1989 <= not w1987 and not w1988;
w1990 <= not w1682 and not w1989;
w1991 <= not w1678 and w1681;
w1992 <= not w1990 and not w1991;
w1993 <= in1(39) and w1144;
w1994 <= in0(39) and not w1144;
w1995 <= not w1993 and not w1994;
w1996 <= in3(39) and w1149;
w1997 <= in2(39) and not w1149;
w1998 <= not w1996 and not w1997;
w1999 <= w1995 and not w1998;
w2000 <= in3(38) and w1149;
w2001 <= in2(38) and not w1149;
w2002 <= not w2000 and not w2001;
w2003 <= in1(38) and w1144;
w2004 <= in0(38) and not w1144;
w2005 <= not w2003 and not w2004;
w2006 <= not w2002 and w2005;
w2007 <= not w1999 and not w2006;
w2008 <= in1(36) and w1144;
w2009 <= in0(36) and not w1144;
w2010 <= not w2008 and not w2009;
w2011 <= in3(36) and w1149;
w2012 <= in2(36) and not w1149;
w2013 <= not w2011 and not w2012;
w2014 <= w2010 and not w2013;
w2015 <= in1(37) and w1144;
w2016 <= in0(37) and not w1144;
w2017 <= not w2015 and not w2016;
w2018 <= in3(37) and w1149;
w2019 <= in2(37) and not w1149;
w2020 <= not w2018 and not w2019;
w2021 <= w2017 and not w2020;
w2022 <= not w2014 and not w2021;
w2023 <= w2007 and w2022;
w2024 <= in1(33) and w1144;
w2025 <= in0(33) and not w1144;
w2026 <= not w2024 and not w2025;
w2027 <= in3(33) and w1149;
w2028 <= in2(33) and not w1149;
w2029 <= not w2027 and not w2028;
w2030 <= w2026 and not w2029;
w2031 <= in1(35) and w1144;
w2032 <= in0(35) and not w1144;
w2033 <= not w2031 and not w2032;
w2034 <= in3(35) and w1149;
w2035 <= in2(35) and not w1149;
w2036 <= not w2034 and not w2035;
w2037 <= w2033 and not w2036;
w2038 <= in3(34) and w1149;
w2039 <= in2(34) and not w1149;
w2040 <= not w2038 and not w2039;
w2041 <= in1(34) and w1144;
w2042 <= in0(34) and not w1144;
w2043 <= not w2041 and not w2042;
w2044 <= not w2040 and w2043;
w2045 <= not w2037 and not w2044;
w2046 <= not w2030 and w2045;
w2047 <= w2023 and w2046;
w2048 <= not w1992 and w2047;
w2049 <= not w1675 and w2048;
w2050 <= not w1995 and w1998;
w2051 <= not w2010 and w2013;
w2052 <= not w2021 and w2051;
w2053 <= not w2017 and w2020;
w2054 <= not w2052 and not w2053;
w2055 <= w2007 and not w2054;
w2056 <= not w1999 and w2002;
w2057 <= not w2005 and w2056;
w2058 <= not w2033 and w2036;
w2059 <= not w2037 and w2040;
w2060 <= not w2043 and w2059;
w2061 <= w1671 and not w1674;
w2062 <= not w2026 and w2029;
w2063 <= not w2061 and not w2062;
w2064 <= w2046 and not w2063;
w2065 <= not w2060 and not w2064;
w2066 <= not w2058 and w2065;
w2067 <= w2023 and not w2066;
w2068 <= not w2057 and not w2067;
w2069 <= not w2055 and w2068;
w2070 <= not w2050 and w2069;
w2071 <= not w2049 and w2070;
w2072 <= w1649 and not w1652;
w2073 <= not w1646 and not w2072;
w2074 <= w1639 and w2073;
w2075 <= w1623 and w2074;
w2076 <= not w2071 and w2075;
w2077 <= not w1668 and not w2076;
w2078 <= not w1666 and w2077;
w2079 <= not w1661 and w2078;
w2080 <= not w1598 and w2079;
w2081 <= in3(48) and w1149;
w2082 <= in2(48) and not w1149;
w2083 <= not w2081 and not w2082;
w2084 <= in1(48) and w1144;
w2085 <= in0(48) and not w1144;
w2086 <= not w2084 and not w2085;
w2087 <= not w2083 and w2086;
w2088 <= in1(55) and w1144;
w2089 <= in0(55) and not w1144;
w2090 <= not w2088 and not w2089;
w2091 <= in3(55) and w1149;
w2092 <= in2(55) and not w1149;
w2093 <= not w2091 and not w2092;
w2094 <= w2090 and not w2093;
w2095 <= in3(54) and w1149;
w2096 <= in2(54) and not w1149;
w2097 <= not w2095 and not w2096;
w2098 <= in1(54) and w1144;
w2099 <= in0(54) and not w1144;
w2100 <= not w2098 and not w2099;
w2101 <= not w2097 and w2100;
w2102 <= not w2094 and not w2101;
w2103 <= in1(53) and w1144;
w2104 <= in0(53) and not w1144;
w2105 <= not w2103 and not w2104;
w2106 <= in3(53) and w1149;
w2107 <= in2(53) and not w1149;
w2108 <= not w2106 and not w2107;
w2109 <= w2105 and not w2108;
w2110 <= in3(52) and w1149;
w2111 <= in2(52) and not w1149;
w2112 <= not w2110 and not w2111;
w2113 <= in1(52) and w1144;
w2114 <= in0(52) and not w1144;
w2115 <= not w2113 and not w2114;
w2116 <= not w2112 and w2115;
w2117 <= not w2109 and not w2116;
w2118 <= w2102 and w2117;
w2119 <= in1(49) and w1144;
w2120 <= in0(49) and not w1144;
w2121 <= not w2119 and not w2120;
w2122 <= in3(49) and w1149;
w2123 <= in2(49) and not w1149;
w2124 <= not w2122 and not w2123;
w2125 <= w2121 and not w2124;
w2126 <= in1(51) and w1144;
w2127 <= in0(51) and not w1144;
w2128 <= not w2126 and not w2127;
w2129 <= in3(51) and w1149;
w2130 <= in2(51) and not w1149;
w2131 <= not w2129 and not w2130;
w2132 <= w2128 and not w2131;
w2133 <= in3(50) and w1149;
w2134 <= in2(50) and not w1149;
w2135 <= not w2133 and not w2134;
w2136 <= in1(50) and w1144;
w2137 <= in0(50) and not w1144;
w2138 <= not w2136 and not w2137;
w2139 <= not w2135 and w2138;
w2140 <= not w2132 and not w2139;
w2141 <= not w2125 and w2140;
w2142 <= w2118 and w2141;
w2143 <= not w2087 and w2142;
w2144 <= not w2080 and w2143;
w2145 <= not w2090 and w2093;
w2146 <= not w2128 and w2131;
w2147 <= not w2132 and w2135;
w2148 <= not w2138 and w2147;
w2149 <= w2083 and not w2086;
w2150 <= not w2121 and w2124;
w2151 <= not w2149 and not w2150;
w2152 <= w2141 and not w2151;
w2153 <= not w2148 and not w2152;
w2154 <= not w2146 and w2153;
w2155 <= w2118 and not w2154;
w2156 <= w2112 and not w2115;
w2157 <= not w2109 and w2156;
w2158 <= not w2105 and w2108;
w2159 <= not w2157 and not w2158;
w2160 <= w2097 and not w2100;
w2161 <= w2159 and not w2160;
w2162 <= w2102 and not w2161;
w2163 <= not w2155 and not w2162;
w2164 <= not w2145 and w2163;
w2165 <= not w2144 and w2164;
w2166 <= w1572 and not w1575;
w2167 <= not w1569 and not w2166;
w2168 <= w1546 and w2167;
w2169 <= w1562 and w2168;
w2170 <= not w2165 and w2169;
w2171 <= not w1591 and not w2170;
w2172 <= not w1589 and w2171;
w2173 <= not w1584 and w2172;
w2174 <= not w1521 and w2173;
w2175 <= not w1514 and not w2174;
w2176 <= not w1507 and w2175;
w2177 <= w1500 and w2176;
w2178 <= not w1488 and w1491;
w2179 <= w1503 and not w1514;
w2180 <= not w1506 and w2179;
w2181 <= not w1510 and w1513;
w2182 <= not w2180 and not w2181;
w2183 <= w1495 and not w1498;
w2184 <= w2182 and not w2183;
w2185 <= w1500 and not w2184;
w2186 <= not w2178 and not w2185;
w2187 <= not w2177 and w2186;
w2188 <= w1475 and not w1478;
w2189 <= not w1472 and not w2188;
w2190 <= w1465 and w2189;
w2191 <= not w2187 and w2190;
w2192 <= not w1485 and not w2191;
w2193 <= not w1483 and w2192;
w2194 <= not w1456 and w2193;
w2195 <= in1(75) and w1144;
w2196 <= in0(75) and not w1144;
w2197 <= not w2195 and not w2196;
w2198 <= in3(75) and w1149;
w2199 <= in2(75) and not w1149;
w2200 <= not w2198 and not w2199;
w2201 <= w2197 and not w2200;
w2202 <= in3(74) and w1149;
w2203 <= in2(74) and not w1149;
w2204 <= not w2202 and not w2203;
w2205 <= in1(74) and w1144;
w2206 <= in0(74) and not w1144;
w2207 <= not w2205 and not w2206;
w2208 <= not w2204 and w2207;
w2209 <= not w2201 and not w2208;
w2210 <= in1(73) and w1144;
w2211 <= in0(73) and not w1144;
w2212 <= not w2210 and not w2211;
w2213 <= in3(73) and w1149;
w2214 <= in2(73) and not w1149;
w2215 <= not w2213 and not w2214;
w2216 <= w2212 and not w2215;
w2217 <= in3(72) and w1149;
w2218 <= in2(72) and not w1149;
w2219 <= not w2217 and not w2218;
w2220 <= in1(72) and w1144;
w2221 <= in0(72) and not w1144;
w2222 <= not w2220 and not w2221;
w2223 <= not w2219 and w2222;
w2224 <= not w2216 and not w2223;
w2225 <= w2209 and w2224;
w2226 <= not w2194 and w2225;
w2227 <= not w2197 and w2200;
w2228 <= w2219 and not w2222;
w2229 <= not w2216 and w2228;
w2230 <= not w2212 and w2215;
w2231 <= not w2229 and not w2230;
w2232 <= w2204 and not w2207;
w2233 <= w2231 and not w2232;
w2234 <= w2209 and not w2233;
w2235 <= not w2227 and not w2234;
w2236 <= not w2226 and w2235;
w2237 <= w1439 and not w1442;
w2238 <= not w1436 and not w2237;
w2239 <= w1429 and w2238;
w2240 <= not w2236 and w2239;
w2241 <= not w1449 and not w2240;
w2242 <= not w1447 and w2241;
w2243 <= not w1420 and w2242;
w2244 <= not w1413 and not w2243;
w2245 <= w1406 and w2244;
w2246 <= not w1391 and w2245;
w2247 <= not w1394 and w1397;
w2248 <= w1387 and not w1413;
w2249 <= not w1390 and w2248;
w2250 <= not w1409 and w1412;
w2251 <= not w2249 and not w2250;
w2252 <= w1401 and not w1404;
w2253 <= w2251 and not w2252;
w2254 <= w1406 and not w2253;
w2255 <= not w2247 and not w2254;
w2256 <= not w2246 and w2255;
w2257 <= w1374 and not w1377;
w2258 <= not w1371 and not w2257;
w2259 <= w1364 and w2258;
w2260 <= not w2256 and w2259;
w2261 <= not w1384 and not w2260;
w2262 <= not w1382 and w2261;
w2263 <= not w1355 and w2262;
w2264 <= in1(91) and w1144;
w2265 <= in0(91) and not w1144;
w2266 <= not w2264 and not w2265;
w2267 <= in3(91) and w1149;
w2268 <= in2(91) and not w1149;
w2269 <= not w2267 and not w2268;
w2270 <= w2266 and not w2269;
w2271 <= in3(90) and w1149;
w2272 <= in2(90) and not w1149;
w2273 <= not w2271 and not w2272;
w2274 <= in1(90) and w1144;
w2275 <= in0(90) and not w1144;
w2276 <= not w2274 and not w2275;
w2277 <= not w2273 and w2276;
w2278 <= not w2270 and not w2277;
w2279 <= in1(89) and w1144;
w2280 <= in0(89) and not w1144;
w2281 <= not w2279 and not w2280;
w2282 <= in3(89) and w1149;
w2283 <= in2(89) and not w1149;
w2284 <= not w2282 and not w2283;
w2285 <= w2281 and not w2284;
w2286 <= in3(88) and w1149;
w2287 <= in2(88) and not w1149;
w2288 <= not w2286 and not w2287;
w2289 <= in1(88) and w1144;
w2290 <= in0(88) and not w1144;
w2291 <= not w2289 and not w2290;
w2292 <= not w2288 and w2291;
w2293 <= not w2285 and not w2292;
w2294 <= w2278 and w2293;
w2295 <= not w2263 and w2294;
w2296 <= not w2266 and w2269;
w2297 <= w2288 and not w2291;
w2298 <= not w2285 and w2297;
w2299 <= not w2281 and w2284;
w2300 <= not w2298 and not w2299;
w2301 <= w2273 and not w2276;
w2302 <= w2300 and not w2301;
w2303 <= w2278 and not w2302;
w2304 <= not w2296 and not w2303;
w2305 <= not w2295 and w2304;
w2306 <= w1338 and not w1341;
w2307 <= not w1335 and not w2306;
w2308 <= w1328 and w2307;
w2309 <= not w2305 and w2308;
w2310 <= not w1348 and not w2309;
w2311 <= not w1346 and w2310;
w2312 <= not w1319 and w2311;
w2313 <= not w1312 and not w2312;
w2314 <= w1305 and w2313;
w2315 <= not w1290 and w2314;
w2316 <= not w1293 and w1296;
w2317 <= w1286 and not w1312;
w2318 <= not w1289 and w2317;
w2319 <= not w1308 and w1311;
w2320 <= not w2318 and not w2319;
w2321 <= w1300 and not w1303;
w2322 <= w2320 and not w2321;
w2323 <= w1305 and not w2322;
w2324 <= not w2316 and not w2323;
w2325 <= not w2315 and w2324;
w2326 <= w1273 and not w1276;
w2327 <= not w1270 and not w2326;
w2328 <= w1263 and w2327;
w2329 <= not w2325 and w2328;
w2330 <= not w1283 and not w2329;
w2331 <= not w1281 and w2330;
w2332 <= not w1254 and w2331;
w2333 <= in1(107) and w1144;
w2334 <= in0(107) and not w1144;
w2335 <= not w2333 and not w2334;
w2336 <= in3(107) and w1149;
w2337 <= in2(107) and not w1149;
w2338 <= not w2336 and not w2337;
w2339 <= w2335 and not w2338;
w2340 <= in3(106) and w1149;
w2341 <= in2(106) and not w1149;
w2342 <= not w2340 and not w2341;
w2343 <= in1(106) and w1144;
w2344 <= in0(106) and not w1144;
w2345 <= not w2343 and not w2344;
w2346 <= not w2342 and w2345;
w2347 <= not w2339 and not w2346;
w2348 <= in1(105) and w1144;
w2349 <= in0(105) and not w1144;
w2350 <= not w2348 and not w2349;
w2351 <= in3(105) and w1149;
w2352 <= in2(105) and not w1149;
w2353 <= not w2351 and not w2352;
w2354 <= w2350 and not w2353;
w2355 <= in3(104) and w1149;
w2356 <= in2(104) and not w1149;
w2357 <= not w2355 and not w2356;
w2358 <= in1(104) and w1144;
w2359 <= in0(104) and not w1144;
w2360 <= not w2358 and not w2359;
w2361 <= not w2357 and w2360;
w2362 <= not w2354 and not w2361;
w2363 <= w2347 and w2362;
w2364 <= not w2332 and w2363;
w2365 <= not w2335 and w2338;
w2366 <= w2357 and not w2360;
w2367 <= not w2354 and w2366;
w2368 <= not w2350 and w2353;
w2369 <= not w2367 and not w2368;
w2370 <= w2342 and not w2345;
w2371 <= w2369 and not w2370;
w2372 <= w2347 and not w2371;
w2373 <= not w2365 and not w2372;
w2374 <= not w2364 and w2373;
w2375 <= w1237 and not w1240;
w2376 <= not w1234 and not w2375;
w2377 <= w1227 and w2376;
w2378 <= not w2374 and w2377;
w2379 <= not w1247 and not w2378;
w2380 <= not w1245 and w2379;
w2381 <= not w1218 and w2380;
w2382 <= not w1211 and not w2381;
w2383 <= w1204 and w2382;
w2384 <= not w1189 and w2383;
w2385 <= not w1192 and w1195;
w2386 <= w1185 and not w1211;
w2387 <= not w1188 and w2386;
w2388 <= not w1207 and w1210;
w2389 <= not w2387 and not w2388;
w2390 <= w1199 and not w1202;
w2391 <= w2389 and not w2390;
w2392 <= w1204 and not w2391;
w2393 <= not w2385 and not w2392;
w2394 <= not w2384 and w2393;
w2395 <= w1165 and not w1175;
w2396 <= not w1172 and not w2395;
w2397 <= w1162 and w2396;
w2398 <= not w2394 and w2397;
w2399 <= not w1182 and not w2398;
w2400 <= not w1180 and w2399;
w2401 <= not w1153 and w2400;
w2402 <= in1(123) and w1144;
w2403 <= in0(123) and not w1144;
w2404 <= not w2402 and not w2403;
w2405 <= in3(123) and w1149;
w2406 <= in2(123) and not w1149;
w2407 <= not w2405 and not w2406;
w2408 <= w2404 and not w2407;
w2409 <= in3(122) and w1149;
w2410 <= in2(122) and not w1149;
w2411 <= not w2409 and not w2410;
w2412 <= in1(122) and w1144;
w2413 <= in0(122) and not w1144;
w2414 <= not w2412 and not w2413;
w2415 <= not w2411 and w2414;
w2416 <= not w2408 and not w2415;
w2417 <= in1(121) and w1144;
w2418 <= in0(121) and not w1144;
w2419 <= not w2417 and not w2418;
w2420 <= in3(121) and w1149;
w2421 <= in2(121) and not w1149;
w2422 <= not w2420 and not w2421;
w2423 <= w2419 and not w2422;
w2424 <= in3(120) and w1149;
w2425 <= in2(120) and not w1149;
w2426 <= not w2424 and not w2425;
w2427 <= in1(120) and w1144;
w2428 <= in0(120) and not w1144;
w2429 <= not w2427 and not w2428;
w2430 <= not w2426 and w2429;
w2431 <= not w2423 and not w2430;
w2432 <= w2416 and w2431;
w2433 <= not w2401 and w2432;
w2434 <= not w2404 and w2407;
w2435 <= not w2423 and w2426;
w2436 <= not w2429 and w2435;
w2437 <= not w2419 and w2422;
w2438 <= not w2436 and not w2437;
w2439 <= w2411 and not w2414;
w2440 <= w2438 and not w2439;
w2441 <= w2416 and not w2440;
w2442 <= not w2434 and not w2441;
w2443 <= not w2433 and w2442;
w2444 <= in1(124) and w1144;
w2445 <= in0(124) and not w1144;
w2446 <= not w2444 and not w2445;
w2447 <= in3(124) and w1149;
w2448 <= in2(124) and not w1149;
w2449 <= not w2447 and not w2448;
w2450 <= w2446 and not w2449;
w2451 <= not w570 and w1141;
w2452 <= in1(126) and w1144;
w2453 <= in0(126) and not w1144;
w2454 <= not w2452 and not w2453;
w2455 <= in3(126) and w1149;
w2456 <= in2(126) and not w1149;
w2457 <= not w2455 and not w2456;
w2458 <= w2454 and not w2457;
w2459 <= in1(125) and w1144;
w2460 <= in0(125) and not w1144;
w2461 <= not w2459 and not w2460;
w2462 <= in3(125) and w1149;
w2463 <= in2(125) and not w1149;
w2464 <= not w2462 and not w2463;
w2465 <= w2461 and not w2464;
w2466 <= not w2458 and not w2465;
w2467 <= not w2451 and w2466;
w2468 <= not w2450 and w2467;
w2469 <= not w2443 and w2468;
w2470 <= not w2446 and w2449;
w2471 <= not w2461 and w2464;
w2472 <= not w2470 and not w2471;
w2473 <= w2466 and not w2472;
w2474 <= not w2454 and w2457;
w2475 <= not w2473 and not w2474;
w2476 <= not w2451 and not w2475;
w2477 <= not w2469 and not w2476;
w2478 <= not w1142 and w2477;
w2479 <= not w1860 and w2478;
w2480 <= not w1857 and not w2478;
w2481 <= not w2479 and not w2480;
w2482 <= not w1854 and w2478;
w2483 <= not w1865 and not w2478;
w2484 <= not w2482 and not w2483;
w2485 <= not w1872 and w2478;
w2486 <= not w1869 and not w2478;
w2487 <= not w2485 and not w2486;
w2488 <= not w1850 and w2478;
w2489 <= not w1847 and not w2478;
w2490 <= not w2488 and not w2489;
w2491 <= not w1841 and w2478;
w2492 <= not w1844 and not w2478;
w2493 <= not w2491 and not w2492;
w2494 <= not w1835 and w2478;
w2495 <= not w1838 and not w2478;
w2496 <= not w2494 and not w2495;
w2497 <= not w1829 and w2478;
w2498 <= not w1832 and not w2478;
w2499 <= not w2497 and not w2498;
w2500 <= not w1825 and w2478;
w2501 <= not w1822 and not w2478;
w2502 <= not w2500 and not w2501;
w2503 <= not w1819 and w2478;
w2504 <= not w1899 and not w2478;
w2505 <= not w2503 and not w2504;
w2506 <= not w1816 and w2478;
w2507 <= not w1906 and not w2478;
w2508 <= not w2506 and not w2507;
w2509 <= not w1812 and w2478;
w2510 <= not w1809 and not w2478;
w2511 <= not w2509 and not w2510;
w2512 <= not w1805 and w2478;
w2513 <= not w1802 and not w2478;
w2514 <= not w2512 and not w2513;
w2515 <= not w1798 and w2478;
w2516 <= not w1795 and not w2478;
w2517 <= not w2515 and not w2516;
w2518 <= not w1791 and w2478;
w2519 <= not w1788 and not w2478;
w2520 <= not w2518 and not w2519;
w2521 <= not w1784 and w2478;
w2522 <= not w1781 and not w2478;
w2523 <= not w2521 and not w2522;
w2524 <= not w1777 and w2478;
w2525 <= not w1774 and not w2478;
w2526 <= not w2524 and not w2525;
w2527 <= not w1771 and w2478;
w2528 <= not w1931 and not w2478;
w2529 <= not w2527 and not w2528;
w2530 <= not w1768 and w2478;
w2531 <= not w1938 and not w2478;
w2532 <= not w2530 and not w2531;
w2533 <= not w1764 and w2478;
w2534 <= not w1761 and not w2478;
w2535 <= not w2533 and not w2534;
w2536 <= not w1757 and w2478;
w2537 <= not w1754 and not w2478;
w2538 <= not w2536 and not w2537;
w2539 <= not w1750 and w2478;
w2540 <= not w1747 and not w2478;
w2541 <= not w2539 and not w2540;
w2542 <= not w1743 and w2478;
w2543 <= not w1740 and not w2478;
w2544 <= not w2542 and not w2543;
w2545 <= not w1736 and w2478;
w2546 <= not w1733 and not w2478;
w2547 <= not w2545 and not w2546;
w2548 <= not w1729 and w2478;
w2549 <= not w1726 and not w2478;
w2550 <= not w2548 and not w2549;
w2551 <= not w1723 and w2478;
w2552 <= not w1963 and not w2478;
w2553 <= not w2551 and not w2552;
w2554 <= not w1720 and w2478;
w2555 <= not w1970 and not w2478;
w2556 <= not w2554 and not w2555;
w2557 <= not w1716 and w2478;
w2558 <= not w1713 and not w2478;
w2559 <= not w2557 and not w2558;
w2560 <= not w1709 and w2478;
w2561 <= not w1706 and not w2478;
w2562 <= not w2560 and not w2561;
w2563 <= not w1702 and w2478;
w2564 <= not w1699 and not w2478;
w2565 <= not w2563 and not w2564;
w2566 <= not w1695 and w2478;
w2567 <= not w1692 and not w2478;
w2568 <= not w2566 and not w2567;
w2569 <= not w1688 and w2478;
w2570 <= not w1685 and not w2478;
w2571 <= not w2569 and not w2570;
w2572 <= not w1681 and w2478;
w2573 <= not w1678 and not w2478;
w2574 <= not w2572 and not w2573;
w2575 <= not w1671 and w2478;
w2576 <= not w1674 and not w2478;
w2577 <= not w2575 and not w2576;
w2578 <= not w2029 and w2478;
w2579 <= not w2026 and not w2478;
w2580 <= not w2578 and not w2579;
w2581 <= not w2040 and w2478;
w2582 <= not w2043 and not w2478;
w2583 <= not w2581 and not w2582;
w2584 <= not w2036 and w2478;
w2585 <= not w2033 and not w2478;
w2586 <= not w2584 and not w2585;
w2587 <= not w2013 and w2478;
w2588 <= not w2010 and not w2478;
w2589 <= not w2587 and not w2588;
w2590 <= not w2020 and w2478;
w2591 <= not w2017 and not w2478;
w2592 <= not w2590 and not w2591;
w2593 <= not w2002 and w2478;
w2594 <= not w2005 and not w2478;
w2595 <= not w2593 and not w2594;
w2596 <= not w1998 and w2478;
w2597 <= not w1995 and not w2478;
w2598 <= not w2596 and not w2597;
w2599 <= not w1652 and w2478;
w2600 <= not w1649 and not w2478;
w2601 <= not w2599 and not w2600;
w2602 <= not w1645 and w2478;
w2603 <= not w1642 and not w2478;
w2604 <= not w2602 and not w2603;
w2605 <= not w1637 and w2478;
w2606 <= not w1634 and not w2478;
w2607 <= not w2605 and not w2606;
w2608 <= not w1629 and w2478;
w2609 <= not w1626 and not w2478;
w2610 <= not w2608 and not w2609;
w2611 <= not w1613 and w2478;
w2612 <= not w1610 and not w2478;
w2613 <= not w2611 and not w2612;
w2614 <= not w1620 and w2478;
w2615 <= not w1617 and not w2478;
w2616 <= not w2614 and not w2615;
w2617 <= not w1602 and w2478;
w2618 <= not w1605 and not w2478;
w2619 <= not w2617 and not w2618;
w2620 <= not w1597 and w2478;
w2621 <= not w1594 and not w2478;
w2622 <= not w2620 and not w2621;
w2623 <= not w2083 and w2478;
w2624 <= not w2086 and not w2478;
w2625 <= not w2623 and not w2624;
w2626 <= not w2124 and w2478;
w2627 <= not w2121 and not w2478;
w2628 <= not w2626 and not w2627;
w2629 <= not w2135 and w2478;
w2630 <= not w2138 and not w2478;
w2631 <= not w2629 and not w2630;
w2632 <= not w2131 and w2478;
w2633 <= not w2128 and not w2478;
w2634 <= not w2632 and not w2633;
w2635 <= not w2112 and w2478;
w2636 <= not w2115 and not w2478;
w2637 <= not w2635 and not w2636;
w2638 <= not w2108 and w2478;
w2639 <= not w2105 and not w2478;
w2640 <= not w2638 and not w2639;
w2641 <= not w2097 and w2478;
w2642 <= not w2100 and not w2478;
w2643 <= not w2641 and not w2642;
w2644 <= not w2093 and w2478;
w2645 <= not w2090 and not w2478;
w2646 <= not w2644 and not w2645;
w2647 <= not w1575 and w2478;
w2648 <= not w1572 and not w2478;
w2649 <= not w2647 and not w2648;
w2650 <= not w1568 and w2478;
w2651 <= not w1565 and not w2478;
w2652 <= not w2650 and not w2651;
w2653 <= not w1560 and w2478;
w2654 <= not w1557 and not w2478;
w2655 <= not w2653 and not w2654;
w2656 <= not w1552 and w2478;
w2657 <= not w1549 and not w2478;
w2658 <= not w2656 and not w2657;
w2659 <= not w1536 and w2478;
w2660 <= not w1533 and not w2478;
w2661 <= not w2659 and not w2660;
w2662 <= not w1543 and w2478;
w2663 <= not w1540 and not w2478;
w2664 <= not w2662 and not w2663;
w2665 <= not w1525 and w2478;
w2666 <= not w1528 and not w2478;
w2667 <= not w2665 and not w2666;
w2668 <= not w1520 and w2478;
w2669 <= not w1517 and not w2478;
w2670 <= not w2668 and not w2669;
w2671 <= not w1503 and w2478;
w2672 <= not w1506 and not w2478;
w2673 <= not w2671 and not w2672;
w2674 <= not w1513 and w2478;
w2675 <= not w1510 and not w2478;
w2676 <= not w2674 and not w2675;
w2677 <= not w1495 and w2478;
w2678 <= not w1498 and not w2478;
w2679 <= not w2677 and not w2678;
w2680 <= not w1491 and w2478;
w2681 <= not w1488 and not w2478;
w2682 <= not w2680 and not w2681;
w2683 <= not w1478 and w2478;
w2684 <= not w1475 and not w2478;
w2685 <= not w2683 and not w2684;
w2686 <= not w1471 and w2478;
w2687 <= not w1468 and not w2478;
w2688 <= not w2686 and not w2687;
w2689 <= not w1460 and w2478;
w2690 <= not w1463 and not w2478;
w2691 <= not w2689 and not w2690;
w2692 <= not w1455 and w2478;
w2693 <= not w1452 and not w2478;
w2694 <= not w2692 and not w2693;
w2695 <= not w2219 and w2478;
w2696 <= not w2222 and not w2478;
w2697 <= not w2695 and not w2696;
w2698 <= not w2215 and w2478;
w2699 <= not w2212 and not w2478;
w2700 <= not w2698 and not w2699;
w2701 <= not w2204 and w2478;
w2702 <= not w2207 and not w2478;
w2703 <= not w2701 and not w2702;
w2704 <= not w2200 and w2478;
w2705 <= not w2197 and not w2478;
w2706 <= not w2704 and not w2705;
w2707 <= not w1442 and w2478;
w2708 <= not w1439 and not w2478;
w2709 <= not w2707 and not w2708;
w2710 <= not w1435 and w2478;
w2711 <= not w1432 and not w2478;
w2712 <= not w2710 and not w2711;
w2713 <= not w1424 and w2478;
w2714 <= not w1427 and not w2478;
w2715 <= not w2713 and not w2714;
w2716 <= not w1419 and w2478;
w2717 <= not w1416 and not w2478;
w2718 <= not w2716 and not w2717;
w2719 <= not w1387 and w2478;
w2720 <= not w1390 and not w2478;
w2721 <= not w2719 and not w2720;
w2722 <= not w1412 and w2478;
w2723 <= not w1409 and not w2478;
w2724 <= not w2722 and not w2723;
w2725 <= not w1401 and w2478;
w2726 <= not w1404 and not w2478;
w2727 <= not w2725 and not w2726;
w2728 <= not w1397 and w2478;
w2729 <= not w1394 and not w2478;
w2730 <= not w2728 and not w2729;
w2731 <= not w1377 and w2478;
w2732 <= not w1374 and not w2478;
w2733 <= not w2731 and not w2732;
w2734 <= not w1370 and w2478;
w2735 <= not w1367 and not w2478;
w2736 <= not w2734 and not w2735;
w2737 <= not w1359 and w2478;
w2738 <= not w1362 and not w2478;
w2739 <= not w2737 and not w2738;
w2740 <= not w1354 and w2478;
w2741 <= not w1351 and not w2478;
w2742 <= not w2740 and not w2741;
w2743 <= not w2288 and w2478;
w2744 <= not w2291 and not w2478;
w2745 <= not w2743 and not w2744;
w2746 <= not w2284 and w2478;
w2747 <= not w2281 and not w2478;
w2748 <= not w2746 and not w2747;
w2749 <= not w2273 and w2478;
w2750 <= not w2276 and not w2478;
w2751 <= not w2749 and not w2750;
w2752 <= not w2269 and w2478;
w2753 <= not w2266 and not w2478;
w2754 <= not w2752 and not w2753;
w2755 <= not w1341 and w2478;
w2756 <= not w1338 and not w2478;
w2757 <= not w2755 and not w2756;
w2758 <= not w1334 and w2478;
w2759 <= not w1331 and not w2478;
w2760 <= not w2758 and not w2759;
w2761 <= not w1323 and w2478;
w2762 <= not w1326 and not w2478;
w2763 <= not w2761 and not w2762;
w2764 <= not w1318 and w2478;
w2765 <= not w1315 and not w2478;
w2766 <= not w2764 and not w2765;
w2767 <= not w1286 and w2478;
w2768 <= not w1289 and not w2478;
w2769 <= not w2767 and not w2768;
w2770 <= not w1311 and w2478;
w2771 <= not w1308 and not w2478;
w2772 <= not w2770 and not w2771;
w2773 <= not w1300 and w2478;
w2774 <= not w1303 and not w2478;
w2775 <= not w2773 and not w2774;
w2776 <= not w1296 and w2478;
w2777 <= not w1293 and not w2478;
w2778 <= not w2776 and not w2777;
w2779 <= not w1276 and w2478;
w2780 <= not w1273 and not w2478;
w2781 <= not w2779 and not w2780;
w2782 <= not w1269 and w2478;
w2783 <= not w1266 and not w2478;
w2784 <= not w2782 and not w2783;
w2785 <= not w1258 and w2478;
w2786 <= not w1261 and not w2478;
w2787 <= not w2785 and not w2786;
w2788 <= not w1253 and w2478;
w2789 <= not w1250 and not w2478;
w2790 <= not w2788 and not w2789;
w2791 <= not w2357 and w2478;
w2792 <= not w2360 and not w2478;
w2793 <= not w2791 and not w2792;
w2794 <= not w2353 and w2478;
w2795 <= not w2350 and not w2478;
w2796 <= not w2794 and not w2795;
w2797 <= not w2342 and w2478;
w2798 <= not w2345 and not w2478;
w2799 <= not w2797 and not w2798;
w2800 <= not w2338 and w2478;
w2801 <= not w2335 and not w2478;
w2802 <= not w2800 and not w2801;
w2803 <= not w1240 and w2478;
w2804 <= not w1237 and not w2478;
w2805 <= not w2803 and not w2804;
w2806 <= not w1233 and w2478;
w2807 <= not w1230 and not w2478;
w2808 <= not w2806 and not w2807;
w2809 <= not w1222 and w2478;
w2810 <= not w1225 and not w2478;
w2811 <= not w2809 and not w2810;
w2812 <= not w1217 and w2478;
w2813 <= not w1214 and not w2478;
w2814 <= not w2812 and not w2813;
w2815 <= not w1185 and w2478;
w2816 <= not w1188 and not w2478;
w2817 <= not w2815 and not w2816;
w2818 <= not w1210 and w2478;
w2819 <= not w1207 and not w2478;
w2820 <= not w2818 and not w2819;
w2821 <= not w1199 and w2478;
w2822 <= not w1202 and not w2478;
w2823 <= not w2821 and not w2822;
w2824 <= not w1195 and w2478;
w2825 <= not w1192 and not w2478;
w2826 <= not w2824 and not w2825;
w2827 <= not w1175 and w2478;
w2828 <= not w1165 and not w2478;
w2829 <= not w2827 and not w2828;
w2830 <= not w1171 and w2478;
w2831 <= not w1168 and not w2478;
w2832 <= not w2830 and not w2831;
w2833 <= not w1157 and w2478;
w2834 <= not w1160 and not w2478;
w2835 <= not w2833 and not w2834;
w2836 <= not w1152 and w2478;
w2837 <= not w1147 and not w2478;
w2838 <= not w2836 and not w2837;
w2839 <= not w2426 and w2478;
w2840 <= not w2429 and not w2478;
w2841 <= not w2839 and not w2840;
w2842 <= not w2422 and w2478;
w2843 <= not w2419 and not w2478;
w2844 <= not w2842 and not w2843;
w2845 <= not w2411 and w2478;
w2846 <= not w2414 and not w2478;
w2847 <= not w2845 and not w2846;
w2848 <= not w2407 and w2478;
w2849 <= not w2404 and not w2478;
w2850 <= not w2848 and not w2849;
w2851 <= not w2449 and w2478;
w2852 <= not w2446 and not w2478;
w2853 <= not w2851 and not w2852;
w2854 <= not w2464 and w2478;
w2855 <= not w2461 and not w2478;
w2856 <= not w2854 and not w2855;
w2857 <= not w2457 and w2478;
w2858 <= not w2454 and not w2478;
w2859 <= not w2857 and not w2858;
w2860 <= not w570 and w2477;
w2861 <= w1141 and not w2860;
w2862 <= w1149 and w2478;
w2863 <= w1144 and not w2478;
w2864 <= not w2862 and not w2863;
one <= '1';
result(0) <= not w2481;-- level 287
result(1) <= not w2484;-- level 287
result(2) <= not w2487;-- level 287
result(3) <= not w2490;-- level 287
result(4) <= not w2493;-- level 287
result(5) <= not w2496;-- level 287
result(6) <= not w2499;-- level 287
result(7) <= not w2502;-- level 287
result(8) <= not w2505;-- level 287
result(9) <= not w2508;-- level 287
result(10) <= not w2511;-- level 287
result(11) <= not w2514;-- level 287
result(12) <= not w2517;-- level 287
result(13) <= not w2520;-- level 287
result(14) <= not w2523;-- level 287
result(15) <= not w2526;-- level 287
result(16) <= not w2529;-- level 287
result(17) <= not w2532;-- level 287
result(18) <= not w2535;-- level 287
result(19) <= not w2538;-- level 287
result(20) <= not w2541;-- level 287
result(21) <= not w2544;-- level 287
result(22) <= not w2547;-- level 287
result(23) <= not w2550;-- level 287
result(24) <= not w2553;-- level 287
result(25) <= not w2556;-- level 287
result(26) <= not w2559;-- level 287
result(27) <= not w2562;-- level 287
result(28) <= not w2565;-- level 287
result(29) <= not w2568;-- level 287
result(30) <= not w2571;-- level 287
result(31) <= not w2574;-- level 287
result(32) <= not w2577;-- level 287
result(33) <= not w2580;-- level 287
result(34) <= not w2583;-- level 287
result(35) <= not w2586;-- level 287
result(36) <= not w2589;-- level 287
result(37) <= not w2592;-- level 287
result(38) <= not w2595;-- level 287
result(39) <= not w2598;-- level 287
result(40) <= not w2601;-- level 287
result(41) <= not w2604;-- level 287
result(42) <= not w2607;-- level 287
result(43) <= not w2610;-- level 287
result(44) <= not w2613;-- level 287
result(45) <= not w2616;-- level 287
result(46) <= not w2619;-- level 287
result(47) <= not w2622;-- level 287
result(48) <= not w2625;-- level 287
result(49) <= not w2628;-- level 287
result(50) <= not w2631;-- level 287
result(51) <= not w2634;-- level 287
result(52) <= not w2637;-- level 287
result(53) <= not w2640;-- level 287
result(54) <= not w2643;-- level 287
result(55) <= not w2646;-- level 287
result(56) <= not w2649;-- level 287
result(57) <= not w2652;-- level 287
result(58) <= not w2655;-- level 287
result(59) <= not w2658;-- level 287
result(60) <= not w2661;-- level 287
result(61) <= not w2664;-- level 287
result(62) <= not w2667;-- level 287
result(63) <= not w2670;-- level 287
result(64) <= not w2673;-- level 287
result(65) <= not w2676;-- level 287
result(66) <= not w2679;-- level 287
result(67) <= not w2682;-- level 287
result(68) <= not w2685;-- level 287
result(69) <= not w2688;-- level 287
result(70) <= not w2691;-- level 287
result(71) <= not w2694;-- level 287
result(72) <= not w2697;-- level 287
result(73) <= not w2700;-- level 287
result(74) <= not w2703;-- level 287
result(75) <= not w2706;-- level 287
result(76) <= not w2709;-- level 287
result(77) <= not w2712;-- level 287
result(78) <= not w2715;-- level 287
result(79) <= not w2718;-- level 287
result(80) <= not w2721;-- level 287
result(81) <= not w2724;-- level 287
result(82) <= not w2727;-- level 287
result(83) <= not w2730;-- level 287
result(84) <= not w2733;-- level 287
result(85) <= not w2736;-- level 287
result(86) <= not w2739;-- level 287
result(87) <= not w2742;-- level 287
result(88) <= not w2745;-- level 287
result(89) <= not w2748;-- level 287
result(90) <= not w2751;-- level 287
result(91) <= not w2754;-- level 287
result(92) <= not w2757;-- level 287
result(93) <= not w2760;-- level 287
result(94) <= not w2763;-- level 287
result(95) <= not w2766;-- level 287
result(96) <= not w2769;-- level 287
result(97) <= not w2772;-- level 287
result(98) <= not w2775;-- level 287
result(99) <= not w2778;-- level 287
result(100) <= not w2781;-- level 287
result(101) <= not w2784;-- level 287
result(102) <= not w2787;-- level 287
result(103) <= not w2790;-- level 287
result(104) <= not w2793;-- level 287
result(105) <= not w2796;-- level 287
result(106) <= not w2799;-- level 287
result(107) <= not w2802;-- level 287
result(108) <= not w2805;-- level 287
result(109) <= not w2808;-- level 287
result(110) <= not w2811;-- level 287
result(111) <= not w2814;-- level 287
result(112) <= not w2817;-- level 287
result(113) <= not w2820;-- level 287
result(114) <= not w2823;-- level 287
result(115) <= not w2826;-- level 287
result(116) <= not w2829;-- level 287
result(117) <= not w2832;-- level 287
result(118) <= not w2835;-- level 287
result(119) <= not w2838;-- level 287
result(120) <= not w2841;-- level 287
result(121) <= not w2844;-- level 287
result(122) <= not w2847;-- level 287
result(123) <= not w2850;-- level 287
result(124) <= not w2853;-- level 287
result(125) <= not w2856;-- level 287
result(126) <= not w2859;-- level 287
result(127) <= w2861;-- level 286
address(0) <= not w2864;-- level 287
address(1) <= w2478;-- level 285
end Behavioral;
