library ieee;
use ieee.std_logic_1164.all;

entity top is
	port( A: in std_logic_vector(1000 downto 0); 
maj: out std_logic);
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757: std_logic;

begin

w0 <= A(718) and A(719);
w1 <= A(718) and not A(719);
w2 <= not A(718) and A(719);
w3 <= not w1 and not w2;
w4 <= A(720) and not w3;
w5 <= not w0 and not w4;
w6 <= A(715) and A(716);
w7 <= A(715) and not A(716);
w8 <= not A(715) and A(716);
w9 <= not w7 and not w8;
w10 <= A(717) and not w9;
w11 <= not w6 and not w10;
w12 <= w5 and not w11;
w13 <= not w5 and w11;
w14 <= A(717) and not w7;
w15 <= not w8 and w14;
w16 <= not A(717) and not w9;
w17 <= not w15 and not w16;
w18 <= A(720) and not w1;
w19 <= not w2 and w18;
w20 <= not A(720) and not w3;
w21 <= not w19 and not w20;
w22 <= not w17 and not w21;
w23 <= not w13 and w22;
w24 <= not w12 and w23;
w25 <= not w12 and not w13;
w26 <= not w22 and not w25;
w27 <= not w24 and not w26;
w28 <= not w17 and w21;
w29 <= w17 and not w21;
w30 <= not w28 and not w29;
w31 <= w22 and not w25;
w32 <= not w5 and not w11;
w33 <= not w31 and not w32;
w34 <= not w30 and not w33;
w35 <= not w27 and not w34;
w36 <= not w27 and not w33;
w37 <= A(724) and A(725);
w38 <= A(724) and not A(725);
w39 <= not A(724) and A(725);
w40 <= not w38 and not w39;
w41 <= A(726) and not w40;
w42 <= not w37 and not w41;
w43 <= A(721) and A(722);
w44 <= A(721) and not A(722);
w45 <= not A(721) and A(722);
w46 <= not w44 and not w45;
w47 <= A(723) and not w46;
w48 <= not w43 and not w47;
w49 <= not w42 and w48;
w50 <= w42 and not w48;
w51 <= not w49 and not w50;
w52 <= A(723) and not w44;
w53 <= not w45 and w52;
w54 <= not A(723) and not w46;
w55 <= not w53 and not w54;
w56 <= A(726) and not w38;
w57 <= not w39 and w56;
w58 <= not A(726) and not w40;
w59 <= not w57 and not w58;
w60 <= not w55 and not w59;
w61 <= not w51 and w60;
w62 <= not w42 and not w48;
w63 <= not w61 and not w62;
w64 <= not w49 and w60;
w65 <= not w50 and w64;
w66 <= not w51 and not w60;
w67 <= not w65 and not w66;
w68 <= not w63 and not w67;
w69 <= not w55 and w59;
w70 <= w55 and not w59;
w71 <= not w69 and not w70;
w72 <= not w30 and not w71;
w73 <= not w68 and w72;
w74 <= not w36 and w73;
w75 <= not w63 and not w71;
w76 <= not w67 and not w75;
w77 <= not w74 and not w76;
w78 <= not w67 and w72;
w79 <= not w68 and w78;
w80 <= not w36 and not w75;
w81 <= w79 and w80;
w82 <= not w77 and not w81;
w83 <= w35 and not w82;
w84 <= not w74 and w76;
w85 <= w74 and not w76;
w86 <= not w84 and not w85;
w87 <= not w35 and not w86;
w88 <= not w68 and not w71;
w89 <= not w30 and not w36;
w90 <= not w88 and w89;
w91 <= w88 and not w89;
w92 <= not w90 and not w91;
w93 <= not A(709) and A(710);
w94 <= A(709) and not A(710);
w95 <= A(711) and not w94;
w96 <= not w93 and w95;
w97 <= not w93 and not w94;
w98 <= not A(711) and not w97;
w99 <= not w96 and not w98;
w100 <= not A(712) and A(713);
w101 <= A(712) and not A(713);
w102 <= A(714) and not w101;
w103 <= not w100 and w102;
w104 <= not w100 and not w101;
w105 <= not A(714) and not w104;
w106 <= not w103 and not w105;
w107 <= not w99 and w106;
w108 <= w99 and not w106;
w109 <= not w107 and not w108;
w110 <= A(712) and A(713);
w111 <= A(714) and not w104;
w112 <= not w110 and not w111;
w113 <= A(709) and A(710);
w114 <= A(711) and not w97;
w115 <= not w113 and not w114;
w116 <= not w112 and w115;
w117 <= w112 and not w115;
w118 <= not w116 and not w117;
w119 <= not w99 and not w106;
w120 <= not w118 and w119;
w121 <= not w112 and not w115;
w122 <= not w120 and not w121;
w123 <= not w116 and w119;
w124 <= not w117 and w123;
w125 <= not w118 and not w119;
w126 <= not w124 and not w125;
w127 <= not w122 and not w126;
w128 <= not w109 and not w127;
w129 <= not A(703) and A(704);
w130 <= A(703) and not A(704);
w131 <= A(705) and not w130;
w132 <= not w129 and w131;
w133 <= not w129 and not w130;
w134 <= not A(705) and not w133;
w135 <= not w132 and not w134;
w136 <= not A(706) and A(707);
w137 <= A(706) and not A(707);
w138 <= A(708) and not w137;
w139 <= not w136 and w138;
w140 <= not w136 and not w137;
w141 <= not A(708) and not w140;
w142 <= not w139 and not w141;
w143 <= not w135 and w142;
w144 <= w135 and not w142;
w145 <= not w143 and not w144;
w146 <= A(706) and A(707);
w147 <= A(708) and not w140;
w148 <= not w146 and not w147;
w149 <= A(703) and A(704);
w150 <= A(705) and not w133;
w151 <= not w149 and not w150;
w152 <= not w148 and w151;
w153 <= w148 and not w151;
w154 <= not w152 and not w153;
w155 <= not w135 and not w142;
w156 <= not w154 and w155;
w157 <= not w148 and not w151;
w158 <= not w156 and not w157;
w159 <= not w152 and w155;
w160 <= not w153 and w159;
w161 <= not w154 and not w155;
w162 <= not w160 and not w161;
w163 <= not w158 and not w162;
w164 <= not w145 and not w163;
w165 <= not w128 and w164;
w166 <= w128 and not w164;
w167 <= not w165 and not w166;
w168 <= not w92 and not w167;
w169 <= not w87 and w168;
w170 <= not w83 and w169;
w171 <= not w83 and not w87;
w172 <= not w168 and not w171;
w173 <= not w170 and not w172;
w174 <= not w145 and not w158;
w175 <= not w162 and not w174;
w176 <= not w109 and not w145;
w177 <= not w127 and w176;
w178 <= not w163 and w177;
w179 <= not w109 and not w122;
w180 <= not w126 and not w179;
w181 <= not w178 and w180;
w182 <= w178 and not w180;
w183 <= not w181 and not w182;
w184 <= not w175 and not w183;
w185 <= not w178 and not w180;
w186 <= not w126 and w176;
w187 <= not w127 and w186;
w188 <= not w163 and not w179;
w189 <= w187 and w188;
w190 <= not w185 and not w189;
w191 <= w175 and not w190;
w192 <= not w184 and not w191;
w193 <= not w173 and w192;
w194 <= not w87 and not w168;
w195 <= not w83 and w194;
w196 <= w168 and not w171;
w197 <= not w195 and not w196;
w198 <= not w192 and not w197;
w199 <= not w193 and not w198;
w200 <= A(730) and A(731);
w201 <= A(730) and not A(731);
w202 <= not A(730) and A(731);
w203 <= not w201 and not w202;
w204 <= A(732) and not w203;
w205 <= not w200 and not w204;
w206 <= A(727) and A(728);
w207 <= A(727) and not A(728);
w208 <= not A(727) and A(728);
w209 <= not w207 and not w208;
w210 <= A(729) and not w209;
w211 <= not w206 and not w210;
w212 <= w205 and not w211;
w213 <= not w205 and w211;
w214 <= A(729) and not w207;
w215 <= not w208 and w214;
w216 <= not A(729) and not w209;
w217 <= not w215 and not w216;
w218 <= A(732) and not w201;
w219 <= not w202 and w218;
w220 <= not A(732) and not w203;
w221 <= not w219 and not w220;
w222 <= not w217 and not w221;
w223 <= not w213 and w222;
w224 <= not w212 and w223;
w225 <= not w212 and not w213;
w226 <= not w222 and not w225;
w227 <= not w224 and not w226;
w228 <= not w217 and w221;
w229 <= w217 and not w221;
w230 <= not w228 and not w229;
w231 <= w222 and not w225;
w232 <= not w205 and not w211;
w233 <= not w231 and not w232;
w234 <= not w230 and not w233;
w235 <= not w227 and not w234;
w236 <= not w227 and not w233;
w237 <= A(736) and A(737);
w238 <= A(736) and not A(737);
w239 <= not A(736) and A(737);
w240 <= not w238 and not w239;
w241 <= A(738) and not w240;
w242 <= not w237 and not w241;
w243 <= A(733) and A(734);
w244 <= A(733) and not A(734);
w245 <= not A(733) and A(734);
w246 <= not w244 and not w245;
w247 <= A(735) and not w246;
w248 <= not w243 and not w247;
w249 <= not w242 and w248;
w250 <= w242 and not w248;
w251 <= not w249 and not w250;
w252 <= A(735) and not w244;
w253 <= not w245 and w252;
w254 <= not A(735) and not w246;
w255 <= not w253 and not w254;
w256 <= A(738) and not w238;
w257 <= not w239 and w256;
w258 <= not A(738) and not w240;
w259 <= not w257 and not w258;
w260 <= not w255 and not w259;
w261 <= not w251 and w260;
w262 <= not w242 and not w248;
w263 <= not w261 and not w262;
w264 <= not w249 and w260;
w265 <= not w250 and w264;
w266 <= not w251 and not w260;
w267 <= not w265 and not w266;
w268 <= not w263 and not w267;
w269 <= not w255 and w259;
w270 <= w255 and not w259;
w271 <= not w269 and not w270;
w272 <= not w230 and not w271;
w273 <= not w268 and w272;
w274 <= not w236 and w273;
w275 <= not w263 and not w271;
w276 <= not w267 and not w275;
w277 <= not w274 and w276;
w278 <= w274 and not w276;
w279 <= not w277 and not w278;
w280 <= not w235 and not w279;
w281 <= not w274 and not w276;
w282 <= not w267 and w272;
w283 <= not w268 and w282;
w284 <= not w236 and not w275;
w285 <= w283 and w284;
w286 <= not w281 and not w285;
w287 <= w235 and not w286;
w288 <= not w280 and not w287;
w289 <= A(742) and A(743);
w290 <= A(742) and not A(743);
w291 <= not A(742) and A(743);
w292 <= not w290 and not w291;
w293 <= A(744) and not w292;
w294 <= not w289 and not w293;
w295 <= A(739) and A(740);
w296 <= A(739) and not A(740);
w297 <= not A(739) and A(740);
w298 <= not w296 and not w297;
w299 <= A(741) and not w298;
w300 <= not w295 and not w299;
w301 <= w294 and not w300;
w302 <= not w294 and w300;
w303 <= A(741) and not w296;
w304 <= not w297 and w303;
w305 <= not A(741) and not w298;
w306 <= not w304 and not w305;
w307 <= A(744) and not w290;
w308 <= not w291 and w307;
w309 <= not A(744) and not w292;
w310 <= not w308 and not w309;
w311 <= not w306 and not w310;
w312 <= not w302 and w311;
w313 <= not w301 and w312;
w314 <= not w301 and not w302;
w315 <= not w311 and not w314;
w316 <= not w313 and not w315;
w317 <= not w306 and w310;
w318 <= w306 and not w310;
w319 <= not w317 and not w318;
w320 <= w311 and not w314;
w321 <= not w294 and not w300;
w322 <= not w320 and not w321;
w323 <= not w319 and not w322;
w324 <= not w316 and not w323;
w325 <= not w316 and not w322;
w326 <= A(748) and A(749);
w327 <= A(748) and not A(749);
w328 <= not A(748) and A(749);
w329 <= not w327 and not w328;
w330 <= A(750) and not w329;
w331 <= not w326 and not w330;
w332 <= A(745) and A(746);
w333 <= A(745) and not A(746);
w334 <= not A(745) and A(746);
w335 <= not w333 and not w334;
w336 <= A(747) and not w335;
w337 <= not w332 and not w336;
w338 <= not w331 and w337;
w339 <= w331 and not w337;
w340 <= not w338 and not w339;
w341 <= A(747) and not w333;
w342 <= not w334 and w341;
w343 <= not A(747) and not w335;
w344 <= not w342 and not w343;
w345 <= A(750) and not w327;
w346 <= not w328 and w345;
w347 <= not A(750) and not w329;
w348 <= not w346 and not w347;
w349 <= not w344 and not w348;
w350 <= not w340 and w349;
w351 <= not w331 and not w337;
w352 <= not w350 and not w351;
w353 <= not w338 and w349;
w354 <= not w339 and w353;
w355 <= not w340 and not w349;
w356 <= not w354 and not w355;
w357 <= not w352 and not w356;
w358 <= not w344 and w348;
w359 <= w344 and not w348;
w360 <= not w358 and not w359;
w361 <= not w319 and not w360;
w362 <= not w357 and w361;
w363 <= not w325 and w362;
w364 <= not w352 and not w360;
w365 <= not w356 and not w364;
w366 <= not w363 and not w365;
w367 <= not w356 and w361;
w368 <= not w357 and w367;
w369 <= not w325 and not w364;
w370 <= w368 and w369;
w371 <= not w366 and not w370;
w372 <= w324 and not w371;
w373 <= not w363 and w365;
w374 <= w363 and not w365;
w375 <= not w373 and not w374;
w376 <= not w324 and not w375;
w377 <= not w357 and not w360;
w378 <= not w319 and not w325;
w379 <= not w377 and w378;
w380 <= w377 and not w378;
w381 <= not w379 and not w380;
w382 <= not w268 and not w271;
w383 <= not w230 and not w236;
w384 <= not w382 and w383;
w385 <= w382 and not w383;
w386 <= not w384 and not w385;
w387 <= not w381 and not w386;
w388 <= not w376 and not w387;
w389 <= not w372 and w388;
w390 <= not w372 and not w376;
w391 <= w387 and not w390;
w392 <= not w389 and not w391;
w393 <= not w288 and not w392;
w394 <= not w376 and w387;
w395 <= not w372 and w394;
w396 <= not w387 and not w390;
w397 <= not w395 and not w396;
w398 <= w288 and not w397;
w399 <= not w381 and w386;
w400 <= w381 and not w386;
w401 <= not w399 and not w400;
w402 <= not w92 and w167;
w403 <= w92 and not w167;
w404 <= not w402 and not w403;
w405 <= not w401 and not w404;
w406 <= not w398 and not w405;
w407 <= not w393 and w406;
w408 <= not w393 and not w398;
w409 <= w405 and not w408;
w410 <= not w407 and not w409;
w411 <= not w199 and not w410;
w412 <= not w398 and w405;
w413 <= not w393 and w412;
w414 <= not w405 and not w408;
w415 <= not w413 and not w414;
w416 <= w199 and not w415;
w417 <= not w401 and w404;
w418 <= w401 and not w404;
w419 <= not w417 and not w418;
w420 <= not A(697) and A(698);
w421 <= A(697) and not A(698);
w422 <= A(699) and not w421;
w423 <= not w420 and w422;
w424 <= not w420 and not w421;
w425 <= not A(699) and not w424;
w426 <= not w423 and not w425;
w427 <= not A(700) and A(701);
w428 <= A(700) and not A(701);
w429 <= A(702) and not w428;
w430 <= not w427 and w429;
w431 <= not w427 and not w428;
w432 <= not A(702) and not w431;
w433 <= not w430 and not w432;
w434 <= not w426 and w433;
w435 <= w426 and not w433;
w436 <= not w434 and not w435;
w437 <= A(700) and A(701);
w438 <= A(702) and not w431;
w439 <= not w437 and not w438;
w440 <= A(697) and A(698);
w441 <= A(699) and not w424;
w442 <= not w440 and not w441;
w443 <= not w439 and w442;
w444 <= w439 and not w442;
w445 <= not w443 and not w444;
w446 <= not w426 and not w433;
w447 <= not w445 and w446;
w448 <= not w439 and not w442;
w449 <= not w447 and not w448;
w450 <= not w443 and w446;
w451 <= not w444 and w450;
w452 <= not w445 and not w446;
w453 <= not w451 and not w452;
w454 <= not w449 and not w453;
w455 <= not w436 and not w454;
w456 <= not A(691) and A(692);
w457 <= A(691) and not A(692);
w458 <= A(693) and not w457;
w459 <= not w456 and w458;
w460 <= not w456 and not w457;
w461 <= not A(693) and not w460;
w462 <= not w459 and not w461;
w463 <= not A(694) and A(695);
w464 <= A(694) and not A(695);
w465 <= A(696) and not w464;
w466 <= not w463 and w465;
w467 <= not w463 and not w464;
w468 <= not A(696) and not w467;
w469 <= not w466 and not w468;
w470 <= not w462 and w469;
w471 <= w462 and not w469;
w472 <= not w470 and not w471;
w473 <= A(694) and A(695);
w474 <= A(696) and not w467;
w475 <= not w473 and not w474;
w476 <= A(691) and A(692);
w477 <= A(693) and not w460;
w478 <= not w476 and not w477;
w479 <= not w475 and w478;
w480 <= w475 and not w478;
w481 <= not w479 and not w480;
w482 <= not w462 and not w469;
w483 <= not w481 and w482;
w484 <= not w475 and not w478;
w485 <= not w483 and not w484;
w486 <= not w479 and w482;
w487 <= not w480 and w486;
w488 <= not w481 and not w482;
w489 <= not w487 and not w488;
w490 <= not w485 and not w489;
w491 <= not w472 and not w490;
w492 <= not w455 and w491;
w493 <= w455 and not w491;
w494 <= not w492 and not w493;
w495 <= not A(685) and A(686);
w496 <= A(685) and not A(686);
w497 <= A(687) and not w496;
w498 <= not w495 and w497;
w499 <= not w495 and not w496;
w500 <= not A(687) and not w499;
w501 <= not w498 and not w500;
w502 <= not A(688) and A(689);
w503 <= A(688) and not A(689);
w504 <= A(690) and not w503;
w505 <= not w502 and w504;
w506 <= not w502 and not w503;
w507 <= not A(690) and not w506;
w508 <= not w505 and not w507;
w509 <= not w501 and w508;
w510 <= w501 and not w508;
w511 <= not w509 and not w510;
w512 <= A(688) and A(689);
w513 <= A(690) and not w506;
w514 <= not w512 and not w513;
w515 <= A(685) and A(686);
w516 <= A(687) and not w499;
w517 <= not w515 and not w516;
w518 <= not w514 and w517;
w519 <= w514 and not w517;
w520 <= not w518 and not w519;
w521 <= not w501 and not w508;
w522 <= not w520 and w521;
w523 <= not w514 and not w517;
w524 <= not w522 and not w523;
w525 <= not w518 and w521;
w526 <= not w519 and w525;
w527 <= not w520 and not w521;
w528 <= not w526 and not w527;
w529 <= not w524 and not w528;
w530 <= not w511 and not w529;
w531 <= not A(679) and A(680);
w532 <= A(679) and not A(680);
w533 <= A(681) and not w532;
w534 <= not w531 and w533;
w535 <= not w531 and not w532;
w536 <= not A(681) and not w535;
w537 <= not w534 and not w536;
w538 <= not A(682) and A(683);
w539 <= A(682) and not A(683);
w540 <= A(684) and not w539;
w541 <= not w538 and w540;
w542 <= not w538 and not w539;
w543 <= not A(684) and not w542;
w544 <= not w541 and not w543;
w545 <= not w537 and w544;
w546 <= w537 and not w544;
w547 <= not w545 and not w546;
w548 <= A(682) and A(683);
w549 <= A(684) and not w542;
w550 <= not w548 and not w549;
w551 <= A(679) and A(680);
w552 <= A(681) and not w535;
w553 <= not w551 and not w552;
w554 <= not w550 and w553;
w555 <= w550 and not w553;
w556 <= not w554 and not w555;
w557 <= not w537 and not w544;
w558 <= not w556 and w557;
w559 <= not w550 and not w553;
w560 <= not w558 and not w559;
w561 <= not w554 and w557;
w562 <= not w555 and w561;
w563 <= not w556 and not w557;
w564 <= not w562 and not w563;
w565 <= not w560 and not w564;
w566 <= not w547 and not w565;
w567 <= not w530 and w566;
w568 <= w530 and not w566;
w569 <= not w567 and not w568;
w570 <= not w494 and w569;
w571 <= w494 and not w569;
w572 <= not w570 and not w571;
w573 <= not A(673) and A(674);
w574 <= A(673) and not A(674);
w575 <= A(675) and not w574;
w576 <= not w573 and w575;
w577 <= not w573 and not w574;
w578 <= not A(675) and not w577;
w579 <= not w576 and not w578;
w580 <= not A(676) and A(677);
w581 <= A(676) and not A(677);
w582 <= A(678) and not w581;
w583 <= not w580 and w582;
w584 <= not w580 and not w581;
w585 <= not A(678) and not w584;
w586 <= not w583 and not w585;
w587 <= not w579 and w586;
w588 <= w579 and not w586;
w589 <= not w587 and not w588;
w590 <= A(676) and A(677);
w591 <= A(678) and not w584;
w592 <= not w590 and not w591;
w593 <= A(673) and A(674);
w594 <= A(675) and not w577;
w595 <= not w593 and not w594;
w596 <= not w592 and w595;
w597 <= w592 and not w595;
w598 <= not w596 and not w597;
w599 <= not w579 and not w586;
w600 <= not w598 and w599;
w601 <= not w592 and not w595;
w602 <= not w600 and not w601;
w603 <= not w596 and w599;
w604 <= not w597 and w603;
w605 <= not w598 and not w599;
w606 <= not w604 and not w605;
w607 <= not w602 and not w606;
w608 <= not w589 and not w607;
w609 <= not A(667) and A(668);
w610 <= A(667) and not A(668);
w611 <= A(669) and not w610;
w612 <= not w609 and w611;
w613 <= not w609 and not w610;
w614 <= not A(669) and not w613;
w615 <= not w612 and not w614;
w616 <= not A(670) and A(671);
w617 <= A(670) and not A(671);
w618 <= A(672) and not w617;
w619 <= not w616 and w618;
w620 <= not w616 and not w617;
w621 <= not A(672) and not w620;
w622 <= not w619 and not w621;
w623 <= not w615 and w622;
w624 <= w615 and not w622;
w625 <= not w623 and not w624;
w626 <= A(670) and A(671);
w627 <= A(672) and not w620;
w628 <= not w626 and not w627;
w629 <= A(667) and A(668);
w630 <= A(669) and not w613;
w631 <= not w629 and not w630;
w632 <= not w628 and w631;
w633 <= w628 and not w631;
w634 <= not w632 and not w633;
w635 <= not w615 and not w622;
w636 <= not w634 and w635;
w637 <= not w628 and not w631;
w638 <= not w636 and not w637;
w639 <= not w632 and w635;
w640 <= not w633 and w639;
w641 <= not w634 and not w635;
w642 <= not w640 and not w641;
w643 <= not w638 and not w642;
w644 <= not w625 and not w643;
w645 <= not w608 and w644;
w646 <= w608 and not w644;
w647 <= not w645 and not w646;
w648 <= not A(661) and A(662);
w649 <= A(661) and not A(662);
w650 <= A(663) and not w649;
w651 <= not w648 and w650;
w652 <= not w648 and not w649;
w653 <= not A(663) and not w652;
w654 <= not w651 and not w653;
w655 <= not A(664) and A(665);
w656 <= A(664) and not A(665);
w657 <= A(666) and not w656;
w658 <= not w655 and w657;
w659 <= not w655 and not w656;
w660 <= not A(666) and not w659;
w661 <= not w658 and not w660;
w662 <= not w654 and w661;
w663 <= w654 and not w661;
w664 <= not w662 and not w663;
w665 <= A(664) and A(665);
w666 <= A(666) and not w659;
w667 <= not w665 and not w666;
w668 <= A(661) and A(662);
w669 <= A(663) and not w652;
w670 <= not w668 and not w669;
w671 <= not w667 and w670;
w672 <= w667 and not w670;
w673 <= not w671 and not w672;
w674 <= not w654 and not w661;
w675 <= not w673 and w674;
w676 <= not w667 and not w670;
w677 <= not w675 and not w676;
w678 <= not w671 and w674;
w679 <= not w672 and w678;
w680 <= not w673 and not w674;
w681 <= not w679 and not w680;
w682 <= not w677 and not w681;
w683 <= not w664 and not w682;
w684 <= not A(655) and A(656);
w685 <= A(655) and not A(656);
w686 <= A(657) and not w685;
w687 <= not w684 and w686;
w688 <= not w684 and not w685;
w689 <= not A(657) and not w688;
w690 <= not w687 and not w689;
w691 <= not A(658) and A(659);
w692 <= A(658) and not A(659);
w693 <= A(660) and not w692;
w694 <= not w691 and w693;
w695 <= not w691 and not w692;
w696 <= not A(660) and not w695;
w697 <= not w694 and not w696;
w698 <= not w690 and w697;
w699 <= w690 and not w697;
w700 <= not w698 and not w699;
w701 <= A(658) and A(659);
w702 <= A(660) and not w695;
w703 <= not w701 and not w702;
w704 <= A(655) and A(656);
w705 <= A(657) and not w688;
w706 <= not w704 and not w705;
w707 <= not w703 and w706;
w708 <= w703 and not w706;
w709 <= not w707 and not w708;
w710 <= not w690 and not w697;
w711 <= not w709 and w710;
w712 <= not w703 and not w706;
w713 <= not w711 and not w712;
w714 <= not w707 and w710;
w715 <= not w708 and w714;
w716 <= not w709 and not w710;
w717 <= not w715 and not w716;
w718 <= not w713 and not w717;
w719 <= not w700 and not w718;
w720 <= not w683 and w719;
w721 <= w683 and not w719;
w722 <= not w720 and not w721;
w723 <= not w647 and w722;
w724 <= w647 and not w722;
w725 <= not w723 and not w724;
w726 <= not w572 and w725;
w727 <= w572 and not w725;
w728 <= not w726 and not w727;
w729 <= not w419 and not w728;
w730 <= not w416 and w729;
w731 <= not w411 and w730;
w732 <= not w411 and not w416;
w733 <= not w729 and not w732;
w734 <= not w731 and not w733;
w735 <= not w547 and not w560;
w736 <= not w564 and not w735;
w737 <= not w511 and not w547;
w738 <= not w529 and w737;
w739 <= not w565 and w738;
w740 <= not w511 and not w524;
w741 <= not w528 and not w740;
w742 <= not w739 and w741;
w743 <= w739 and not w741;
w744 <= not w742 and not w743;
w745 <= not w736 and not w744;
w746 <= not w739 and not w741;
w747 <= not w528 and w737;
w748 <= not w529 and w747;
w749 <= not w565 and not w740;
w750 <= w748 and w749;
w751 <= not w746 and not w750;
w752 <= w736 and not w751;
w753 <= not w745 and not w752;
w754 <= not w472 and not w485;
w755 <= not w489 and not w754;
w756 <= not w436 and not w472;
w757 <= not w454 and w756;
w758 <= not w490 and w757;
w759 <= not w436 and not w449;
w760 <= not w453 and not w759;
w761 <= not w758 and not w760;
w762 <= not w453 and w756;
w763 <= not w454 and w762;
w764 <= not w490 and not w759;
w765 <= w763 and w764;
w766 <= not w761 and not w765;
w767 <= w755 and not w766;
w768 <= not w758 and w760;
w769 <= w758 and not w760;
w770 <= not w768 and not w769;
w771 <= not w755 and not w770;
w772 <= not w494 and not w569;
w773 <= not w771 and not w772;
w774 <= not w767 and w773;
w775 <= not w767 and not w771;
w776 <= w772 and not w775;
w777 <= not w774 and not w776;
w778 <= not w753 and not w777;
w779 <= not w771 and w772;
w780 <= not w767 and w779;
w781 <= not w772 and not w775;
w782 <= not w780 and not w781;
w783 <= w753 and not w782;
w784 <= not w572 and not w725;
w785 <= not w783 and w784;
w786 <= not w778 and w785;
w787 <= not w778 and not w783;
w788 <= not w784 and not w787;
w789 <= not w786 and not w788;
w790 <= not w625 and not w638;
w791 <= not w642 and not w790;
w792 <= not w589 and not w625;
w793 <= not w607 and w792;
w794 <= not w643 and w793;
w795 <= not w589 and not w602;
w796 <= not w606 and not w795;
w797 <= not w794 and not w796;
w798 <= not w606 and w792;
w799 <= not w607 and w798;
w800 <= not w643 and not w795;
w801 <= w799 and w800;
w802 <= not w797 and not w801;
w803 <= w791 and not w802;
w804 <= not w794 and w796;
w805 <= w794 and not w796;
w806 <= not w804 and not w805;
w807 <= not w791 and not w806;
w808 <= not w647 and not w722;
w809 <= not w807 and w808;
w810 <= not w803 and w809;
w811 <= not w803 and not w807;
w812 <= not w808 and not w811;
w813 <= not w810 and not w812;
w814 <= not w700 and not w713;
w815 <= not w717 and not w814;
w816 <= not w664 and not w700;
w817 <= not w682 and w816;
w818 <= not w718 and w817;
w819 <= not w664 and not w677;
w820 <= not w681 and not w819;
w821 <= not w818 and w820;
w822 <= w818 and not w820;
w823 <= not w821 and not w822;
w824 <= not w815 and not w823;
w825 <= not w818 and not w820;
w826 <= not w681 and w816;
w827 <= not w682 and w826;
w828 <= not w718 and not w819;
w829 <= w827 and w828;
w830 <= not w825 and not w829;
w831 <= w815 and not w830;
w832 <= not w824 and not w831;
w833 <= not w813 and w832;
w834 <= not w807 and not w808;
w835 <= not w803 and w834;
w836 <= w808 and not w811;
w837 <= not w835 and not w836;
w838 <= not w832 and not w837;
w839 <= not w833 and not w838;
w840 <= not w789 and w839;
w841 <= not w783 and not w784;
w842 <= not w778 and w841;
w843 <= w784 and not w787;
w844 <= not w842 and not w843;
w845 <= not w839 and not w844;
w846 <= not w840 and not w845;
w847 <= not w734 and w846;
w848 <= not w416 and not w729;
w849 <= not w411 and w848;
w850 <= w729 and not w732;
w851 <= not w849 and not w850;
w852 <= not w846 and not w851;
w853 <= not w847 and not w852;
w854 <= A(778) and A(779);
w855 <= A(778) and not A(779);
w856 <= not A(778) and A(779);
w857 <= not w855 and not w856;
w858 <= A(780) and not w857;
w859 <= not w854 and not w858;
w860 <= A(775) and A(776);
w861 <= A(775) and not A(776);
w862 <= not A(775) and A(776);
w863 <= not w861 and not w862;
w864 <= A(777) and not w863;
w865 <= not w860 and not w864;
w866 <= w859 and not w865;
w867 <= not w859 and w865;
w868 <= A(777) and not w861;
w869 <= not w862 and w868;
w870 <= not A(777) and not w863;
w871 <= not w869 and not w870;
w872 <= A(780) and not w855;
w873 <= not w856 and w872;
w874 <= not A(780) and not w857;
w875 <= not w873 and not w874;
w876 <= not w871 and not w875;
w877 <= not w867 and w876;
w878 <= not w866 and w877;
w879 <= not w866 and not w867;
w880 <= not w876 and not w879;
w881 <= not w878 and not w880;
w882 <= not w871 and w875;
w883 <= w871 and not w875;
w884 <= not w882 and not w883;
w885 <= w876 and not w879;
w886 <= not w859 and not w865;
w887 <= not w885 and not w886;
w888 <= not w884 and not w887;
w889 <= not w881 and not w888;
w890 <= not w881 and not w887;
w891 <= A(784) and A(785);
w892 <= A(784) and not A(785);
w893 <= not A(784) and A(785);
w894 <= not w892 and not w893;
w895 <= A(786) and not w894;
w896 <= not w891 and not w895;
w897 <= A(781) and A(782);
w898 <= A(781) and not A(782);
w899 <= not A(781) and A(782);
w900 <= not w898 and not w899;
w901 <= A(783) and not w900;
w902 <= not w897 and not w901;
w903 <= not w896 and w902;
w904 <= w896 and not w902;
w905 <= not w903 and not w904;
w906 <= A(783) and not w898;
w907 <= not w899 and w906;
w908 <= not A(783) and not w900;
w909 <= not w907 and not w908;
w910 <= A(786) and not w892;
w911 <= not w893 and w910;
w912 <= not A(786) and not w894;
w913 <= not w911 and not w912;
w914 <= not w909 and not w913;
w915 <= not w905 and w914;
w916 <= not w896 and not w902;
w917 <= not w915 and not w916;
w918 <= not w903 and w914;
w919 <= not w904 and w918;
w920 <= not w905 and not w914;
w921 <= not w919 and not w920;
w922 <= not w917 and not w921;
w923 <= not w909 and w913;
w924 <= w909 and not w913;
w925 <= not w923 and not w924;
w926 <= not w884 and not w925;
w927 <= not w922 and w926;
w928 <= not w890 and w927;
w929 <= not w917 and not w925;
w930 <= not w921 and not w929;
w931 <= not w928 and w930;
w932 <= w928 and not w930;
w933 <= not w931 and not w932;
w934 <= not w889 and not w933;
w935 <= not w928 and not w930;
w936 <= not w921 and w926;
w937 <= not w922 and w936;
w938 <= not w890 and not w929;
w939 <= w937 and w938;
w940 <= not w935 and not w939;
w941 <= w889 and not w940;
w942 <= not w934 and not w941;
w943 <= A(790) and A(791);
w944 <= A(790) and not A(791);
w945 <= not A(790) and A(791);
w946 <= not w944 and not w945;
w947 <= A(792) and not w946;
w948 <= not w943 and not w947;
w949 <= A(787) and A(788);
w950 <= A(787) and not A(788);
w951 <= not A(787) and A(788);
w952 <= not w950 and not w951;
w953 <= A(789) and not w952;
w954 <= not w949 and not w953;
w955 <= w948 and not w954;
w956 <= not w948 and w954;
w957 <= A(789) and not w950;
w958 <= not w951 and w957;
w959 <= not A(789) and not w952;
w960 <= not w958 and not w959;
w961 <= A(792) and not w944;
w962 <= not w945 and w961;
w963 <= not A(792) and not w946;
w964 <= not w962 and not w963;
w965 <= not w960 and not w964;
w966 <= not w956 and w965;
w967 <= not w955 and w966;
w968 <= not w955 and not w956;
w969 <= not w965 and not w968;
w970 <= not w967 and not w969;
w971 <= not w960 and w964;
w972 <= w960 and not w964;
w973 <= not w971 and not w972;
w974 <= w965 and not w968;
w975 <= not w948 and not w954;
w976 <= not w974 and not w975;
w977 <= not w973 and not w976;
w978 <= not w970 and not w977;
w979 <= not w970 and not w976;
w980 <= A(796) and A(797);
w981 <= A(796) and not A(797);
w982 <= not A(796) and A(797);
w983 <= not w981 and not w982;
w984 <= A(798) and not w983;
w985 <= not w980 and not w984;
w986 <= A(793) and A(794);
w987 <= A(793) and not A(794);
w988 <= not A(793) and A(794);
w989 <= not w987 and not w988;
w990 <= A(795) and not w989;
w991 <= not w986 and not w990;
w992 <= not w985 and w991;
w993 <= w985 and not w991;
w994 <= not w992 and not w993;
w995 <= A(795) and not w987;
w996 <= not w988 and w995;
w997 <= not A(795) and not w989;
w998 <= not w996 and not w997;
w999 <= A(798) and not w981;
w1000 <= not w982 and w999;
w1001 <= not A(798) and not w983;
w1002 <= not w1000 and not w1001;
w1003 <= not w998 and not w1002;
w1004 <= not w994 and w1003;
w1005 <= not w985 and not w991;
w1006 <= not w1004 and not w1005;
w1007 <= not w992 and w1003;
w1008 <= not w993 and w1007;
w1009 <= not w994 and not w1003;
w1010 <= not w1008 and not w1009;
w1011 <= not w1006 and not w1010;
w1012 <= not w998 and w1002;
w1013 <= w998 and not w1002;
w1014 <= not w1012 and not w1013;
w1015 <= not w973 and not w1014;
w1016 <= not w1011 and w1015;
w1017 <= not w979 and w1016;
w1018 <= not w1006 and not w1014;
w1019 <= not w1010 and not w1018;
w1020 <= not w1017 and not w1019;
w1021 <= not w1010 and w1015;
w1022 <= not w1011 and w1021;
w1023 <= not w979 and not w1018;
w1024 <= w1022 and w1023;
w1025 <= not w1020 and not w1024;
w1026 <= w978 and not w1025;
w1027 <= not w1017 and w1019;
w1028 <= w1017 and not w1019;
w1029 <= not w1027 and not w1028;
w1030 <= not w978 and not w1029;
w1031 <= not w1011 and not w1014;
w1032 <= not w973 and not w979;
w1033 <= not w1031 and w1032;
w1034 <= w1031 and not w1032;
w1035 <= not w1033 and not w1034;
w1036 <= not w922 and not w925;
w1037 <= not w884 and not w890;
w1038 <= not w1036 and w1037;
w1039 <= w1036 and not w1037;
w1040 <= not w1038 and not w1039;
w1041 <= not w1035 and not w1040;
w1042 <= not w1030 and not w1041;
w1043 <= not w1026 and w1042;
w1044 <= not w1026 and not w1030;
w1045 <= w1041 and not w1044;
w1046 <= not w1043 and not w1045;
w1047 <= not w942 and not w1046;
w1048 <= not w1030 and w1041;
w1049 <= not w1026 and w1048;
w1050 <= not w1041 and not w1044;
w1051 <= not w1049 and not w1050;
w1052 <= w942 and not w1051;
w1053 <= not w1035 and w1040;
w1054 <= w1035 and not w1040;
w1055 <= not w1053 and not w1054;
w1056 <= not A(769) and A(770);
w1057 <= A(769) and not A(770);
w1058 <= A(771) and not w1057;
w1059 <= not w1056 and w1058;
w1060 <= not w1056 and not w1057;
w1061 <= not A(771) and not w1060;
w1062 <= not w1059 and not w1061;
w1063 <= not A(772) and A(773);
w1064 <= A(772) and not A(773);
w1065 <= A(774) and not w1064;
w1066 <= not w1063 and w1065;
w1067 <= not w1063 and not w1064;
w1068 <= not A(774) and not w1067;
w1069 <= not w1066 and not w1068;
w1070 <= not w1062 and w1069;
w1071 <= w1062 and not w1069;
w1072 <= not w1070 and not w1071;
w1073 <= A(772) and A(773);
w1074 <= A(774) and not w1067;
w1075 <= not w1073 and not w1074;
w1076 <= A(769) and A(770);
w1077 <= A(771) and not w1060;
w1078 <= not w1076 and not w1077;
w1079 <= not w1075 and w1078;
w1080 <= w1075 and not w1078;
w1081 <= not w1079 and not w1080;
w1082 <= not w1062 and not w1069;
w1083 <= not w1081 and w1082;
w1084 <= not w1075 and not w1078;
w1085 <= not w1083 and not w1084;
w1086 <= not w1079 and w1082;
w1087 <= not w1080 and w1086;
w1088 <= not w1081 and not w1082;
w1089 <= not w1087 and not w1088;
w1090 <= not w1085 and not w1089;
w1091 <= not w1072 and not w1090;
w1092 <= not A(763) and A(764);
w1093 <= A(763) and not A(764);
w1094 <= A(765) and not w1093;
w1095 <= not w1092 and w1094;
w1096 <= not w1092 and not w1093;
w1097 <= not A(765) and not w1096;
w1098 <= not w1095 and not w1097;
w1099 <= not A(766) and A(767);
w1100 <= A(766) and not A(767);
w1101 <= A(768) and not w1100;
w1102 <= not w1099 and w1101;
w1103 <= not w1099 and not w1100;
w1104 <= not A(768) and not w1103;
w1105 <= not w1102 and not w1104;
w1106 <= not w1098 and w1105;
w1107 <= w1098 and not w1105;
w1108 <= not w1106 and not w1107;
w1109 <= A(766) and A(767);
w1110 <= A(768) and not w1103;
w1111 <= not w1109 and not w1110;
w1112 <= A(763) and A(764);
w1113 <= A(765) and not w1096;
w1114 <= not w1112 and not w1113;
w1115 <= not w1111 and w1114;
w1116 <= w1111 and not w1114;
w1117 <= not w1115 and not w1116;
w1118 <= not w1098 and not w1105;
w1119 <= not w1117 and w1118;
w1120 <= not w1111 and not w1114;
w1121 <= not w1119 and not w1120;
w1122 <= not w1115 and w1118;
w1123 <= not w1116 and w1122;
w1124 <= not w1117 and not w1118;
w1125 <= not w1123 and not w1124;
w1126 <= not w1121 and not w1125;
w1127 <= not w1108 and not w1126;
w1128 <= not w1091 and w1127;
w1129 <= w1091 and not w1127;
w1130 <= not w1128 and not w1129;
w1131 <= not A(757) and A(758);
w1132 <= A(757) and not A(758);
w1133 <= A(759) and not w1132;
w1134 <= not w1131 and w1133;
w1135 <= not w1131 and not w1132;
w1136 <= not A(759) and not w1135;
w1137 <= not w1134 and not w1136;
w1138 <= not A(760) and A(761);
w1139 <= A(760) and not A(761);
w1140 <= A(762) and not w1139;
w1141 <= not w1138 and w1140;
w1142 <= not w1138 and not w1139;
w1143 <= not A(762) and not w1142;
w1144 <= not w1141 and not w1143;
w1145 <= not w1137 and w1144;
w1146 <= w1137 and not w1144;
w1147 <= not w1145 and not w1146;
w1148 <= A(760) and A(761);
w1149 <= A(762) and not w1142;
w1150 <= not w1148 and not w1149;
w1151 <= A(757) and A(758);
w1152 <= A(759) and not w1135;
w1153 <= not w1151 and not w1152;
w1154 <= not w1150 and w1153;
w1155 <= w1150 and not w1153;
w1156 <= not w1154 and not w1155;
w1157 <= not w1137 and not w1144;
w1158 <= not w1156 and w1157;
w1159 <= not w1150 and not w1153;
w1160 <= not w1158 and not w1159;
w1161 <= not w1154 and w1157;
w1162 <= not w1155 and w1161;
w1163 <= not w1156 and not w1157;
w1164 <= not w1162 and not w1163;
w1165 <= not w1160 and not w1164;
w1166 <= not w1147 and not w1165;
w1167 <= not A(751) and A(752);
w1168 <= A(751) and not A(752);
w1169 <= A(753) and not w1168;
w1170 <= not w1167 and w1169;
w1171 <= not w1167 and not w1168;
w1172 <= not A(753) and not w1171;
w1173 <= not w1170 and not w1172;
w1174 <= not A(754) and A(755);
w1175 <= A(754) and not A(755);
w1176 <= A(756) and not w1175;
w1177 <= not w1174 and w1176;
w1178 <= not w1174 and not w1175;
w1179 <= not A(756) and not w1178;
w1180 <= not w1177 and not w1179;
w1181 <= not w1173 and w1180;
w1182 <= w1173 and not w1180;
w1183 <= not w1181 and not w1182;
w1184 <= A(754) and A(755);
w1185 <= A(756) and not w1178;
w1186 <= not w1184 and not w1185;
w1187 <= A(751) and A(752);
w1188 <= A(753) and not w1171;
w1189 <= not w1187 and not w1188;
w1190 <= not w1186 and w1189;
w1191 <= w1186 and not w1189;
w1192 <= not w1190 and not w1191;
w1193 <= not w1173 and not w1180;
w1194 <= not w1192 and w1193;
w1195 <= not w1186 and not w1189;
w1196 <= not w1194 and not w1195;
w1197 <= not w1190 and w1193;
w1198 <= not w1191 and w1197;
w1199 <= not w1192 and not w1193;
w1200 <= not w1198 and not w1199;
w1201 <= not w1196 and not w1200;
w1202 <= not w1183 and not w1201;
w1203 <= not w1166 and w1202;
w1204 <= w1166 and not w1202;
w1205 <= not w1203 and not w1204;
w1206 <= not w1130 and w1205;
w1207 <= w1130 and not w1205;
w1208 <= not w1206 and not w1207;
w1209 <= not w1055 and not w1208;
w1210 <= not w1052 and w1209;
w1211 <= not w1047 and w1210;
w1212 <= not w1047 and not w1052;
w1213 <= not w1209 and not w1212;
w1214 <= not w1211 and not w1213;
w1215 <= not w1108 and not w1121;
w1216 <= not w1125 and not w1215;
w1217 <= not w1072 and not w1108;
w1218 <= not w1090 and w1217;
w1219 <= not w1126 and w1218;
w1220 <= not w1072 and not w1085;
w1221 <= not w1089 and not w1220;
w1222 <= not w1219 and not w1221;
w1223 <= not w1089 and w1217;
w1224 <= not w1090 and w1223;
w1225 <= not w1126 and not w1220;
w1226 <= w1224 and w1225;
w1227 <= not w1222 and not w1226;
w1228 <= w1216 and not w1227;
w1229 <= not w1219 and w1221;
w1230 <= w1219 and not w1221;
w1231 <= not w1229 and not w1230;
w1232 <= not w1216 and not w1231;
w1233 <= not w1130 and not w1205;
w1234 <= not w1232 and w1233;
w1235 <= not w1228 and w1234;
w1236 <= not w1228 and not w1232;
w1237 <= not w1233 and not w1236;
w1238 <= not w1235 and not w1237;
w1239 <= not w1183 and not w1196;
w1240 <= not w1200 and not w1239;
w1241 <= not w1147 and not w1183;
w1242 <= not w1165 and w1241;
w1243 <= not w1201 and w1242;
w1244 <= not w1147 and not w1160;
w1245 <= not w1164 and not w1244;
w1246 <= not w1243 and w1245;
w1247 <= w1243 and not w1245;
w1248 <= not w1246 and not w1247;
w1249 <= not w1240 and not w1248;
w1250 <= not w1243 and not w1245;
w1251 <= not w1164 and w1241;
w1252 <= not w1165 and w1251;
w1253 <= not w1201 and not w1244;
w1254 <= w1252 and w1253;
w1255 <= not w1250 and not w1254;
w1256 <= w1240 and not w1255;
w1257 <= not w1249 and not w1256;
w1258 <= not w1238 and w1257;
w1259 <= not w1232 and not w1233;
w1260 <= not w1228 and w1259;
w1261 <= w1233 and not w1236;
w1262 <= not w1260 and not w1261;
w1263 <= not w1257 and not w1262;
w1264 <= not w1258 and not w1263;
w1265 <= not w1214 and w1264;
w1266 <= not w1052 and not w1209;
w1267 <= not w1047 and w1266;
w1268 <= w1209 and not w1212;
w1269 <= not w1267 and not w1268;
w1270 <= not w1264 and not w1269;
w1271 <= not w1265 and not w1270;
w1272 <= A(814) and A(815);
w1273 <= A(814) and not A(815);
w1274 <= not A(814) and A(815);
w1275 <= not w1273 and not w1274;
w1276 <= A(816) and not w1275;
w1277 <= not w1272 and not w1276;
w1278 <= A(811) and A(812);
w1279 <= A(811) and not A(812);
w1280 <= not A(811) and A(812);
w1281 <= not w1279 and not w1280;
w1282 <= A(813) and not w1281;
w1283 <= not w1278 and not w1282;
w1284 <= w1277 and not w1283;
w1285 <= not w1277 and w1283;
w1286 <= A(813) and not w1279;
w1287 <= not w1280 and w1286;
w1288 <= not A(813) and not w1281;
w1289 <= not w1287 and not w1288;
w1290 <= A(816) and not w1273;
w1291 <= not w1274 and w1290;
w1292 <= not A(816) and not w1275;
w1293 <= not w1291 and not w1292;
w1294 <= not w1289 and not w1293;
w1295 <= not w1285 and w1294;
w1296 <= not w1284 and w1295;
w1297 <= not w1284 and not w1285;
w1298 <= not w1294 and not w1297;
w1299 <= not w1296 and not w1298;
w1300 <= not w1289 and w1293;
w1301 <= w1289 and not w1293;
w1302 <= not w1300 and not w1301;
w1303 <= w1294 and not w1297;
w1304 <= not w1277 and not w1283;
w1305 <= not w1303 and not w1304;
w1306 <= not w1302 and not w1305;
w1307 <= not w1299 and not w1306;
w1308 <= not w1299 and not w1305;
w1309 <= A(820) and A(821);
w1310 <= A(820) and not A(821);
w1311 <= not A(820) and A(821);
w1312 <= not w1310 and not w1311;
w1313 <= A(822) and not w1312;
w1314 <= not w1309 and not w1313;
w1315 <= A(817) and A(818);
w1316 <= A(817) and not A(818);
w1317 <= not A(817) and A(818);
w1318 <= not w1316 and not w1317;
w1319 <= A(819) and not w1318;
w1320 <= not w1315 and not w1319;
w1321 <= not w1314 and w1320;
w1322 <= w1314 and not w1320;
w1323 <= not w1321 and not w1322;
w1324 <= A(819) and not w1316;
w1325 <= not w1317 and w1324;
w1326 <= not A(819) and not w1318;
w1327 <= not w1325 and not w1326;
w1328 <= A(822) and not w1310;
w1329 <= not w1311 and w1328;
w1330 <= not A(822) and not w1312;
w1331 <= not w1329 and not w1330;
w1332 <= not w1327 and not w1331;
w1333 <= not w1323 and w1332;
w1334 <= not w1314 and not w1320;
w1335 <= not w1333 and not w1334;
w1336 <= not w1321 and w1332;
w1337 <= not w1322 and w1336;
w1338 <= not w1323 and not w1332;
w1339 <= not w1337 and not w1338;
w1340 <= not w1335 and not w1339;
w1341 <= not w1327 and w1331;
w1342 <= w1327 and not w1331;
w1343 <= not w1341 and not w1342;
w1344 <= not w1302 and not w1343;
w1345 <= not w1340 and w1344;
w1346 <= not w1308 and w1345;
w1347 <= not w1335 and not w1343;
w1348 <= not w1339 and not w1347;
w1349 <= not w1346 and not w1348;
w1350 <= not w1339 and w1344;
w1351 <= not w1340 and w1350;
w1352 <= not w1308 and not w1347;
w1353 <= w1351 and w1352;
w1354 <= not w1349 and not w1353;
w1355 <= w1307 and not w1354;
w1356 <= not w1346 and w1348;
w1357 <= w1346 and not w1348;
w1358 <= not w1356 and not w1357;
w1359 <= not w1307 and not w1358;
w1360 <= not w1340 and not w1343;
w1361 <= not w1302 and not w1308;
w1362 <= not w1360 and w1361;
w1363 <= w1360 and not w1361;
w1364 <= not w1362 and not w1363;
w1365 <= not A(805) and A(806);
w1366 <= A(805) and not A(806);
w1367 <= A(807) and not w1366;
w1368 <= not w1365 and w1367;
w1369 <= not w1365 and not w1366;
w1370 <= not A(807) and not w1369;
w1371 <= not w1368 and not w1370;
w1372 <= not A(808) and A(809);
w1373 <= A(808) and not A(809);
w1374 <= A(810) and not w1373;
w1375 <= not w1372 and w1374;
w1376 <= not w1372 and not w1373;
w1377 <= not A(810) and not w1376;
w1378 <= not w1375 and not w1377;
w1379 <= not w1371 and w1378;
w1380 <= w1371 and not w1378;
w1381 <= not w1379 and not w1380;
w1382 <= A(808) and A(809);
w1383 <= A(810) and not w1376;
w1384 <= not w1382 and not w1383;
w1385 <= A(805) and A(806);
w1386 <= A(807) and not w1369;
w1387 <= not w1385 and not w1386;
w1388 <= not w1384 and w1387;
w1389 <= w1384 and not w1387;
w1390 <= not w1388 and not w1389;
w1391 <= not w1371 and not w1378;
w1392 <= not w1390 and w1391;
w1393 <= not w1384 and not w1387;
w1394 <= not w1392 and not w1393;
w1395 <= not w1388 and w1391;
w1396 <= not w1389 and w1395;
w1397 <= not w1390 and not w1391;
w1398 <= not w1396 and not w1397;
w1399 <= not w1394 and not w1398;
w1400 <= not w1381 and not w1399;
w1401 <= not A(799) and A(800);
w1402 <= A(799) and not A(800);
w1403 <= A(801) and not w1402;
w1404 <= not w1401 and w1403;
w1405 <= not w1401 and not w1402;
w1406 <= not A(801) and not w1405;
w1407 <= not w1404 and not w1406;
w1408 <= not A(802) and A(803);
w1409 <= A(802) and not A(803);
w1410 <= A(804) and not w1409;
w1411 <= not w1408 and w1410;
w1412 <= not w1408 and not w1409;
w1413 <= not A(804) and not w1412;
w1414 <= not w1411 and not w1413;
w1415 <= not w1407 and w1414;
w1416 <= w1407 and not w1414;
w1417 <= not w1415 and not w1416;
w1418 <= A(802) and A(803);
w1419 <= A(804) and not w1412;
w1420 <= not w1418 and not w1419;
w1421 <= A(799) and A(800);
w1422 <= A(801) and not w1405;
w1423 <= not w1421 and not w1422;
w1424 <= not w1420 and w1423;
w1425 <= w1420 and not w1423;
w1426 <= not w1424 and not w1425;
w1427 <= not w1407 and not w1414;
w1428 <= not w1426 and w1427;
w1429 <= not w1420 and not w1423;
w1430 <= not w1428 and not w1429;
w1431 <= not w1424 and w1427;
w1432 <= not w1425 and w1431;
w1433 <= not w1426 and not w1427;
w1434 <= not w1432 and not w1433;
w1435 <= not w1430 and not w1434;
w1436 <= not w1417 and not w1435;
w1437 <= not w1400 and w1436;
w1438 <= w1400 and not w1436;
w1439 <= not w1437 and not w1438;
w1440 <= not w1364 and not w1439;
w1441 <= not w1359 and w1440;
w1442 <= not w1355 and w1441;
w1443 <= not w1355 and not w1359;
w1444 <= not w1440 and not w1443;
w1445 <= not w1442 and not w1444;
w1446 <= not w1417 and not w1430;
w1447 <= not w1434 and not w1446;
w1448 <= not w1381 and not w1417;
w1449 <= not w1399 and w1448;
w1450 <= not w1435 and w1449;
w1451 <= not w1381 and not w1394;
w1452 <= not w1398 and not w1451;
w1453 <= not w1450 and w1452;
w1454 <= w1450 and not w1452;
w1455 <= not w1453 and not w1454;
w1456 <= not w1447 and not w1455;
w1457 <= not w1450 and not w1452;
w1458 <= not w1398 and w1448;
w1459 <= not w1399 and w1458;
w1460 <= not w1435 and not w1451;
w1461 <= w1459 and w1460;
w1462 <= not w1457 and not w1461;
w1463 <= w1447 and not w1462;
w1464 <= not w1456 and not w1463;
w1465 <= not w1445 and w1464;
w1466 <= not w1359 and not w1440;
w1467 <= not w1355 and w1466;
w1468 <= w1440 and not w1443;
w1469 <= not w1467 and not w1468;
w1470 <= not w1464 and not w1469;
w1471 <= not w1465 and not w1470;
w1472 <= A(826) and A(827);
w1473 <= A(826) and not A(827);
w1474 <= not A(826) and A(827);
w1475 <= not w1473 and not w1474;
w1476 <= A(828) and not w1475;
w1477 <= not w1472 and not w1476;
w1478 <= A(823) and A(824);
w1479 <= A(823) and not A(824);
w1480 <= not A(823) and A(824);
w1481 <= not w1479 and not w1480;
w1482 <= A(825) and not w1481;
w1483 <= not w1478 and not w1482;
w1484 <= w1477 and not w1483;
w1485 <= not w1477 and w1483;
w1486 <= A(825) and not w1479;
w1487 <= not w1480 and w1486;
w1488 <= not A(825) and not w1481;
w1489 <= not w1487 and not w1488;
w1490 <= A(828) and not w1473;
w1491 <= not w1474 and w1490;
w1492 <= not A(828) and not w1475;
w1493 <= not w1491 and not w1492;
w1494 <= not w1489 and not w1493;
w1495 <= not w1485 and w1494;
w1496 <= not w1484 and w1495;
w1497 <= not w1484 and not w1485;
w1498 <= not w1494 and not w1497;
w1499 <= not w1496 and not w1498;
w1500 <= not w1489 and w1493;
w1501 <= w1489 and not w1493;
w1502 <= not w1500 and not w1501;
w1503 <= w1494 and not w1497;
w1504 <= not w1477 and not w1483;
w1505 <= not w1503 and not w1504;
w1506 <= not w1502 and not w1505;
w1507 <= not w1499 and not w1506;
w1508 <= not w1499 and not w1505;
w1509 <= A(832) and A(833);
w1510 <= A(832) and not A(833);
w1511 <= not A(832) and A(833);
w1512 <= not w1510 and not w1511;
w1513 <= A(834) and not w1512;
w1514 <= not w1509 and not w1513;
w1515 <= A(829) and A(830);
w1516 <= A(829) and not A(830);
w1517 <= not A(829) and A(830);
w1518 <= not w1516 and not w1517;
w1519 <= A(831) and not w1518;
w1520 <= not w1515 and not w1519;
w1521 <= not w1514 and w1520;
w1522 <= w1514 and not w1520;
w1523 <= not w1521 and not w1522;
w1524 <= A(831) and not w1516;
w1525 <= not w1517 and w1524;
w1526 <= not A(831) and not w1518;
w1527 <= not w1525 and not w1526;
w1528 <= A(834) and not w1510;
w1529 <= not w1511 and w1528;
w1530 <= not A(834) and not w1512;
w1531 <= not w1529 and not w1530;
w1532 <= not w1527 and not w1531;
w1533 <= not w1523 and w1532;
w1534 <= not w1514 and not w1520;
w1535 <= not w1533 and not w1534;
w1536 <= not w1521 and w1532;
w1537 <= not w1522 and w1536;
w1538 <= not w1523 and not w1532;
w1539 <= not w1537 and not w1538;
w1540 <= not w1535 and not w1539;
w1541 <= not w1527 and w1531;
w1542 <= w1527 and not w1531;
w1543 <= not w1541 and not w1542;
w1544 <= not w1502 and not w1543;
w1545 <= not w1540 and w1544;
w1546 <= not w1508 and w1545;
w1547 <= not w1535 and not w1543;
w1548 <= not w1539 and not w1547;
w1549 <= not w1546 and w1548;
w1550 <= w1546 and not w1548;
w1551 <= not w1549 and not w1550;
w1552 <= not w1507 and not w1551;
w1553 <= not w1546 and not w1548;
w1554 <= not w1539 and w1544;
w1555 <= not w1540 and w1554;
w1556 <= not w1508 and not w1547;
w1557 <= w1555 and w1556;
w1558 <= not w1553 and not w1557;
w1559 <= w1507 and not w1558;
w1560 <= not w1552 and not w1559;
w1561 <= A(838) and A(839);
w1562 <= A(838) and not A(839);
w1563 <= not A(838) and A(839);
w1564 <= not w1562 and not w1563;
w1565 <= A(840) and not w1564;
w1566 <= not w1561 and not w1565;
w1567 <= A(835) and A(836);
w1568 <= A(835) and not A(836);
w1569 <= not A(835) and A(836);
w1570 <= not w1568 and not w1569;
w1571 <= A(837) and not w1570;
w1572 <= not w1567 and not w1571;
w1573 <= w1566 and not w1572;
w1574 <= not w1566 and w1572;
w1575 <= A(837) and not w1568;
w1576 <= not w1569 and w1575;
w1577 <= not A(837) and not w1570;
w1578 <= not w1576 and not w1577;
w1579 <= A(840) and not w1562;
w1580 <= not w1563 and w1579;
w1581 <= not A(840) and not w1564;
w1582 <= not w1580 and not w1581;
w1583 <= not w1578 and not w1582;
w1584 <= not w1574 and w1583;
w1585 <= not w1573 and w1584;
w1586 <= not w1573 and not w1574;
w1587 <= not w1583 and not w1586;
w1588 <= not w1585 and not w1587;
w1589 <= not w1578 and w1582;
w1590 <= w1578 and not w1582;
w1591 <= not w1589 and not w1590;
w1592 <= w1583 and not w1586;
w1593 <= not w1566 and not w1572;
w1594 <= not w1592 and not w1593;
w1595 <= not w1591 and not w1594;
w1596 <= not w1588 and not w1595;
w1597 <= not w1588 and not w1594;
w1598 <= A(844) and A(845);
w1599 <= A(844) and not A(845);
w1600 <= not A(844) and A(845);
w1601 <= not w1599 and not w1600;
w1602 <= A(846) and not w1601;
w1603 <= not w1598 and not w1602;
w1604 <= A(841) and A(842);
w1605 <= A(841) and not A(842);
w1606 <= not A(841) and A(842);
w1607 <= not w1605 and not w1606;
w1608 <= A(843) and not w1607;
w1609 <= not w1604 and not w1608;
w1610 <= not w1603 and w1609;
w1611 <= w1603 and not w1609;
w1612 <= not w1610 and not w1611;
w1613 <= A(843) and not w1605;
w1614 <= not w1606 and w1613;
w1615 <= not A(843) and not w1607;
w1616 <= not w1614 and not w1615;
w1617 <= A(846) and not w1599;
w1618 <= not w1600 and w1617;
w1619 <= not A(846) and not w1601;
w1620 <= not w1618 and not w1619;
w1621 <= not w1616 and not w1620;
w1622 <= not w1612 and w1621;
w1623 <= not w1603 and not w1609;
w1624 <= not w1622 and not w1623;
w1625 <= not w1610 and w1621;
w1626 <= not w1611 and w1625;
w1627 <= not w1612 and not w1621;
w1628 <= not w1626 and not w1627;
w1629 <= not w1624 and not w1628;
w1630 <= not w1616 and w1620;
w1631 <= w1616 and not w1620;
w1632 <= not w1630 and not w1631;
w1633 <= not w1591 and not w1632;
w1634 <= not w1629 and w1633;
w1635 <= not w1597 and w1634;
w1636 <= not w1624 and not w1632;
w1637 <= not w1628 and not w1636;
w1638 <= not w1635 and not w1637;
w1639 <= not w1628 and w1633;
w1640 <= not w1629 and w1639;
w1641 <= not w1597 and not w1636;
w1642 <= w1640 and w1641;
w1643 <= not w1638 and not w1642;
w1644 <= w1596 and not w1643;
w1645 <= not w1635 and w1637;
w1646 <= w1635 and not w1637;
w1647 <= not w1645 and not w1646;
w1648 <= not w1596 and not w1647;
w1649 <= not w1629 and not w1632;
w1650 <= not w1591 and not w1597;
w1651 <= not w1649 and w1650;
w1652 <= w1649 and not w1650;
w1653 <= not w1651 and not w1652;
w1654 <= not w1540 and not w1543;
w1655 <= not w1502 and not w1508;
w1656 <= not w1654 and w1655;
w1657 <= w1654 and not w1655;
w1658 <= not w1656 and not w1657;
w1659 <= not w1653 and not w1658;
w1660 <= not w1648 and not w1659;
w1661 <= not w1644 and w1660;
w1662 <= not w1644 and not w1648;
w1663 <= w1659 and not w1662;
w1664 <= not w1661 and not w1663;
w1665 <= not w1560 and not w1664;
w1666 <= not w1648 and w1659;
w1667 <= not w1644 and w1666;
w1668 <= not w1659 and not w1662;
w1669 <= not w1667 and not w1668;
w1670 <= w1560 and not w1669;
w1671 <= not w1653 and w1658;
w1672 <= w1653 and not w1658;
w1673 <= not w1671 and not w1672;
w1674 <= not w1364 and w1439;
w1675 <= w1364 and not w1439;
w1676 <= not w1674 and not w1675;
w1677 <= not w1673 and not w1676;
w1678 <= not w1670 and not w1677;
w1679 <= not w1665 and w1678;
w1680 <= not w1665 and not w1670;
w1681 <= w1677 and not w1680;
w1682 <= not w1679 and not w1681;
w1683 <= not w1471 and not w1682;
w1684 <= not w1670 and w1677;
w1685 <= not w1665 and w1684;
w1686 <= not w1677 and not w1680;
w1687 <= not w1685 and not w1686;
w1688 <= w1471 and not w1687;
w1689 <= not w1673 and w1676;
w1690 <= w1673 and not w1676;
w1691 <= not w1689 and not w1690;
w1692 <= not w1055 and w1208;
w1693 <= w1055 and not w1208;
w1694 <= not w1692 and not w1693;
w1695 <= not w1691 and not w1694;
w1696 <= not w1688 and not w1695;
w1697 <= not w1683 and w1696;
w1698 <= not w1683 and not w1688;
w1699 <= w1695 and not w1698;
w1700 <= not w1697 and not w1699;
w1701 <= not w1271 and not w1700;
w1702 <= not w1688 and w1695;
w1703 <= not w1683 and w1702;
w1704 <= not w1695 and not w1698;
w1705 <= not w1703 and not w1704;
w1706 <= w1271 and not w1705;
w1707 <= not w1691 and w1694;
w1708 <= w1691 and not w1694;
w1709 <= not w1707 and not w1708;
w1710 <= not w419 and w728;
w1711 <= w419 and not w728;
w1712 <= not w1710 and not w1711;
w1713 <= not w1709 and not w1712;
w1714 <= not w1706 and not w1713;
w1715 <= not w1701 and w1714;
w1716 <= not w1701 and not w1706;
w1717 <= w1713 and not w1716;
w1718 <= not w1715 and not w1717;
w1719 <= not w853 and not w1718;
w1720 <= not w1706 and w1713;
w1721 <= not w1701 and w1720;
w1722 <= not w1713 and not w1716;
w1723 <= not w1721 and not w1722;
w1724 <= w853 and not w1723;
w1725 <= not A(469) and A(470);
w1726 <= A(469) and not A(470);
w1727 <= A(471) and not w1726;
w1728 <= not w1725 and w1727;
w1729 <= not w1725 and not w1726;
w1730 <= not A(471) and not w1729;
w1731 <= not w1728 and not w1730;
w1732 <= not A(472) and A(473);
w1733 <= A(472) and not A(473);
w1734 <= A(474) and not w1733;
w1735 <= not w1732 and w1734;
w1736 <= not w1732 and not w1733;
w1737 <= not A(474) and not w1736;
w1738 <= not w1735 and not w1737;
w1739 <= not w1731 and w1738;
w1740 <= w1731 and not w1738;
w1741 <= not w1739 and not w1740;
w1742 <= A(472) and A(473);
w1743 <= A(474) and not w1736;
w1744 <= not w1742 and not w1743;
w1745 <= A(469) and A(470);
w1746 <= A(471) and not w1729;
w1747 <= not w1745 and not w1746;
w1748 <= not w1744 and w1747;
w1749 <= w1744 and not w1747;
w1750 <= not w1748 and not w1749;
w1751 <= not w1731 and not w1738;
w1752 <= not w1750 and w1751;
w1753 <= not w1744 and not w1747;
w1754 <= not w1752 and not w1753;
w1755 <= not w1748 and w1751;
w1756 <= not w1749 and w1755;
w1757 <= not w1750 and not w1751;
w1758 <= not w1756 and not w1757;
w1759 <= not w1754 and not w1758;
w1760 <= not w1741 and not w1759;
w1761 <= not A(466) and A(467);
w1762 <= A(466) and not A(467);
w1763 <= A(468) and not w1762;
w1764 <= not w1761 and w1763;
w1765 <= not w1761 and not w1762;
w1766 <= not A(468) and not w1765;
w1767 <= not w1764 and not w1766;
w1768 <= not A(463) and A(464);
w1769 <= A(463) and not A(464);
w1770 <= A(465) and not w1769;
w1771 <= not w1768 and w1770;
w1772 <= not w1768 and not w1769;
w1773 <= not A(465) and not w1772;
w1774 <= not w1771 and not w1773;
w1775 <= not w1767 and w1774;
w1776 <= w1767 and not w1774;
w1777 <= not w1775 and not w1776;
w1778 <= A(466) and A(467);
w1779 <= A(468) and not w1765;
w1780 <= not w1778 and not w1779;
w1781 <= A(463) and A(464);
w1782 <= A(465) and not w1772;
w1783 <= not w1781 and not w1782;
w1784 <= w1780 and not w1783;
w1785 <= not w1780 and w1783;
w1786 <= not w1767 and not w1774;
w1787 <= not w1785 and w1786;
w1788 <= not w1784 and w1787;
w1789 <= not w1784 and not w1785;
w1790 <= not w1786 and not w1789;
w1791 <= not w1788 and not w1790;
w1792 <= w1786 and not w1789;
w1793 <= not w1780 and not w1783;
w1794 <= not w1792 and not w1793;
w1795 <= not w1791 and not w1794;
w1796 <= not w1777 and not w1795;
w1797 <= not w1760 and w1796;
w1798 <= w1760 and not w1796;
w1799 <= not w1797 and not w1798;
w1800 <= not A(481) and A(482);
w1801 <= A(481) and not A(482);
w1802 <= A(483) and not w1801;
w1803 <= not w1800 and w1802;
w1804 <= not w1800 and not w1801;
w1805 <= not A(483) and not w1804;
w1806 <= not w1803 and not w1805;
w1807 <= not A(484) and A(485);
w1808 <= A(484) and not A(485);
w1809 <= A(486) and not w1808;
w1810 <= not w1807 and w1809;
w1811 <= not w1807 and not w1808;
w1812 <= not A(486) and not w1811;
w1813 <= not w1810 and not w1812;
w1814 <= not w1806 and w1813;
w1815 <= w1806 and not w1813;
w1816 <= not w1814 and not w1815;
w1817 <= A(484) and A(485);
w1818 <= A(486) and not w1811;
w1819 <= not w1817 and not w1818;
w1820 <= A(481) and A(482);
w1821 <= A(483) and not w1804;
w1822 <= not w1820 and not w1821;
w1823 <= not w1819 and w1822;
w1824 <= w1819 and not w1822;
w1825 <= not w1823 and not w1824;
w1826 <= not w1806 and not w1813;
w1827 <= not w1825 and w1826;
w1828 <= not w1819 and not w1822;
w1829 <= not w1827 and not w1828;
w1830 <= not w1823 and w1826;
w1831 <= not w1824 and w1830;
w1832 <= not w1825 and not w1826;
w1833 <= not w1831 and not w1832;
w1834 <= not w1829 and not w1833;
w1835 <= not w1816 and not w1834;
w1836 <= not A(475) and A(476);
w1837 <= A(475) and not A(476);
w1838 <= A(477) and not w1837;
w1839 <= not w1836 and w1838;
w1840 <= not w1836 and not w1837;
w1841 <= not A(477) and not w1840;
w1842 <= not w1839 and not w1841;
w1843 <= not A(478) and A(479);
w1844 <= A(478) and not A(479);
w1845 <= A(480) and not w1844;
w1846 <= not w1843 and w1845;
w1847 <= not w1843 and not w1844;
w1848 <= not A(480) and not w1847;
w1849 <= not w1846 and not w1848;
w1850 <= not w1842 and w1849;
w1851 <= w1842 and not w1849;
w1852 <= not w1850 and not w1851;
w1853 <= A(478) and A(479);
w1854 <= A(480) and not w1847;
w1855 <= not w1853 and not w1854;
w1856 <= A(475) and A(476);
w1857 <= A(477) and not w1840;
w1858 <= not w1856 and not w1857;
w1859 <= not w1855 and w1858;
w1860 <= w1855 and not w1858;
w1861 <= not w1859 and not w1860;
w1862 <= not w1842 and not w1849;
w1863 <= not w1861 and w1862;
w1864 <= not w1855 and not w1858;
w1865 <= not w1863 and not w1864;
w1866 <= not w1859 and w1862;
w1867 <= not w1860 and w1866;
w1868 <= not w1861 and not w1862;
w1869 <= not w1867 and not w1868;
w1870 <= not w1865 and not w1869;
w1871 <= not w1852 and not w1870;
w1872 <= not w1835 and w1871;
w1873 <= w1835 and not w1871;
w1874 <= not w1872 and not w1873;
w1875 <= not w1799 and w1874;
w1876 <= w1799 and not w1874;
w1877 <= not w1875 and not w1876;
w1878 <= not A(505) and A(506);
w1879 <= A(505) and not A(506);
w1880 <= A(507) and not w1879;
w1881 <= not w1878 and w1880;
w1882 <= not w1878 and not w1879;
w1883 <= not A(507) and not w1882;
w1884 <= not w1881 and not w1883;
w1885 <= not A(508) and A(509);
w1886 <= A(508) and not A(509);
w1887 <= A(510) and not w1886;
w1888 <= not w1885 and w1887;
w1889 <= not w1885 and not w1886;
w1890 <= not A(510) and not w1889;
w1891 <= not w1888 and not w1890;
w1892 <= not w1884 and w1891;
w1893 <= w1884 and not w1891;
w1894 <= not w1892 and not w1893;
w1895 <= A(508) and A(509);
w1896 <= A(510) and not w1889;
w1897 <= not w1895 and not w1896;
w1898 <= A(505) and A(506);
w1899 <= A(507) and not w1882;
w1900 <= not w1898 and not w1899;
w1901 <= not w1897 and w1900;
w1902 <= w1897 and not w1900;
w1903 <= not w1901 and not w1902;
w1904 <= not w1884 and not w1891;
w1905 <= not w1903 and w1904;
w1906 <= not w1897 and not w1900;
w1907 <= not w1905 and not w1906;
w1908 <= not w1901 and w1904;
w1909 <= not w1902 and w1908;
w1910 <= not w1903 and not w1904;
w1911 <= not w1909 and not w1910;
w1912 <= not w1907 and not w1911;
w1913 <= not w1894 and not w1912;
w1914 <= not A(499) and A(500);
w1915 <= A(499) and not A(500);
w1916 <= A(501) and not w1915;
w1917 <= not w1914 and w1916;
w1918 <= not w1914 and not w1915;
w1919 <= not A(501) and not w1918;
w1920 <= not w1917 and not w1919;
w1921 <= not A(502) and A(503);
w1922 <= A(502) and not A(503);
w1923 <= A(504) and not w1922;
w1924 <= not w1921 and w1923;
w1925 <= not w1921 and not w1922;
w1926 <= not A(504) and not w1925;
w1927 <= not w1924 and not w1926;
w1928 <= not w1920 and w1927;
w1929 <= w1920 and not w1927;
w1930 <= not w1928 and not w1929;
w1931 <= A(502) and A(503);
w1932 <= A(504) and not w1925;
w1933 <= not w1931 and not w1932;
w1934 <= A(499) and A(500);
w1935 <= A(501) and not w1918;
w1936 <= not w1934 and not w1935;
w1937 <= not w1933 and w1936;
w1938 <= w1933 and not w1936;
w1939 <= not w1937 and not w1938;
w1940 <= not w1920 and not w1927;
w1941 <= not w1939 and w1940;
w1942 <= not w1933 and not w1936;
w1943 <= not w1941 and not w1942;
w1944 <= not w1937 and w1940;
w1945 <= not w1938 and w1944;
w1946 <= not w1939 and not w1940;
w1947 <= not w1945 and not w1946;
w1948 <= not w1943 and not w1947;
w1949 <= not w1930 and not w1948;
w1950 <= not w1913 and w1949;
w1951 <= w1913 and not w1949;
w1952 <= not w1950 and not w1951;
w1953 <= not A(493) and A(494);
w1954 <= A(493) and not A(494);
w1955 <= A(495) and not w1954;
w1956 <= not w1953 and w1955;
w1957 <= not w1953 and not w1954;
w1958 <= not A(495) and not w1957;
w1959 <= not w1956 and not w1958;
w1960 <= not A(496) and A(497);
w1961 <= A(496) and not A(497);
w1962 <= A(498) and not w1961;
w1963 <= not w1960 and w1962;
w1964 <= not w1960 and not w1961;
w1965 <= not A(498) and not w1964;
w1966 <= not w1963 and not w1965;
w1967 <= not w1959 and w1966;
w1968 <= w1959 and not w1966;
w1969 <= not w1967 and not w1968;
w1970 <= A(496) and A(497);
w1971 <= A(498) and not w1964;
w1972 <= not w1970 and not w1971;
w1973 <= A(493) and A(494);
w1974 <= A(495) and not w1957;
w1975 <= not w1973 and not w1974;
w1976 <= not w1972 and w1975;
w1977 <= w1972 and not w1975;
w1978 <= not w1976 and not w1977;
w1979 <= not w1959 and not w1966;
w1980 <= not w1978 and w1979;
w1981 <= not w1972 and not w1975;
w1982 <= not w1980 and not w1981;
w1983 <= not w1976 and w1979;
w1984 <= not w1977 and w1983;
w1985 <= not w1978 and not w1979;
w1986 <= not w1984 and not w1985;
w1987 <= not w1982 and not w1986;
w1988 <= not w1969 and not w1987;
w1989 <= not A(487) and A(488);
w1990 <= A(487) and not A(488);
w1991 <= A(489) and not w1990;
w1992 <= not w1989 and w1991;
w1993 <= not w1989 and not w1990;
w1994 <= not A(489) and not w1993;
w1995 <= not w1992 and not w1994;
w1996 <= not A(490) and A(491);
w1997 <= A(490) and not A(491);
w1998 <= A(492) and not w1997;
w1999 <= not w1996 and w1998;
w2000 <= not w1996 and not w1997;
w2001 <= not A(492) and not w2000;
w2002 <= not w1999 and not w2001;
w2003 <= not w1995 and w2002;
w2004 <= w1995 and not w2002;
w2005 <= not w2003 and not w2004;
w2006 <= A(490) and A(491);
w2007 <= A(492) and not w2000;
w2008 <= not w2006 and not w2007;
w2009 <= A(487) and A(488);
w2010 <= A(489) and not w1993;
w2011 <= not w2009 and not w2010;
w2012 <= not w2008 and w2011;
w2013 <= w2008 and not w2011;
w2014 <= not w2012 and not w2013;
w2015 <= not w1995 and not w2002;
w2016 <= not w2014 and w2015;
w2017 <= not w2008 and not w2011;
w2018 <= not w2016 and not w2017;
w2019 <= not w2012 and w2015;
w2020 <= not w2013 and w2019;
w2021 <= not w2014 and not w2015;
w2022 <= not w2020 and not w2021;
w2023 <= not w2018 and not w2022;
w2024 <= not w2005 and not w2023;
w2025 <= not w1988 and w2024;
w2026 <= w1988 and not w2024;
w2027 <= not w2025 and not w2026;
w2028 <= not w1952 and w2027;
w2029 <= w1952 and not w2027;
w2030 <= not w2028 and not w2029;
w2031 <= not w1877 and w2030;
w2032 <= w1877 and not w2030;
w2033 <= not w2031 and not w2032;
w2034 <= not A(553) and A(554);
w2035 <= A(553) and not A(554);
w2036 <= A(555) and not w2035;
w2037 <= not w2034 and w2036;
w2038 <= not w2034 and not w2035;
w2039 <= not A(555) and not w2038;
w2040 <= not w2037 and not w2039;
w2041 <= not A(556) and A(557);
w2042 <= A(556) and not A(557);
w2043 <= A(558) and not w2042;
w2044 <= not w2041 and w2043;
w2045 <= not w2041 and not w2042;
w2046 <= not A(558) and not w2045;
w2047 <= not w2044 and not w2046;
w2048 <= not w2040 and w2047;
w2049 <= w2040 and not w2047;
w2050 <= not w2048 and not w2049;
w2051 <= A(556) and A(557);
w2052 <= A(558) and not w2045;
w2053 <= not w2051 and not w2052;
w2054 <= A(553) and A(554);
w2055 <= A(555) and not w2038;
w2056 <= not w2054 and not w2055;
w2057 <= not w2053 and w2056;
w2058 <= w2053 and not w2056;
w2059 <= not w2057 and not w2058;
w2060 <= not w2040 and not w2047;
w2061 <= not w2059 and w2060;
w2062 <= not w2053 and not w2056;
w2063 <= not w2061 and not w2062;
w2064 <= not w2057 and w2060;
w2065 <= not w2058 and w2064;
w2066 <= not w2059 and not w2060;
w2067 <= not w2065 and not w2066;
w2068 <= not w2063 and not w2067;
w2069 <= not w2050 and not w2068;
w2070 <= not A(547) and A(548);
w2071 <= A(547) and not A(548);
w2072 <= A(549) and not w2071;
w2073 <= not w2070 and w2072;
w2074 <= not w2070 and not w2071;
w2075 <= not A(549) and not w2074;
w2076 <= not w2073 and not w2075;
w2077 <= not A(550) and A(551);
w2078 <= A(550) and not A(551);
w2079 <= A(552) and not w2078;
w2080 <= not w2077 and w2079;
w2081 <= not w2077 and not w2078;
w2082 <= not A(552) and not w2081;
w2083 <= not w2080 and not w2082;
w2084 <= not w2076 and w2083;
w2085 <= w2076 and not w2083;
w2086 <= not w2084 and not w2085;
w2087 <= A(550) and A(551);
w2088 <= A(552) and not w2081;
w2089 <= not w2087 and not w2088;
w2090 <= A(547) and A(548);
w2091 <= A(549) and not w2074;
w2092 <= not w2090 and not w2091;
w2093 <= not w2089 and w2092;
w2094 <= w2089 and not w2092;
w2095 <= not w2093 and not w2094;
w2096 <= not w2076 and not w2083;
w2097 <= not w2095 and w2096;
w2098 <= not w2089 and not w2092;
w2099 <= not w2097 and not w2098;
w2100 <= not w2093 and w2096;
w2101 <= not w2094 and w2100;
w2102 <= not w2095 and not w2096;
w2103 <= not w2101 and not w2102;
w2104 <= not w2099 and not w2103;
w2105 <= not w2086 and not w2104;
w2106 <= not w2069 and w2105;
w2107 <= w2069 and not w2105;
w2108 <= not w2106 and not w2107;
w2109 <= not A(541) and A(542);
w2110 <= A(541) and not A(542);
w2111 <= A(543) and not w2110;
w2112 <= not w2109 and w2111;
w2113 <= not w2109 and not w2110;
w2114 <= not A(543) and not w2113;
w2115 <= not w2112 and not w2114;
w2116 <= not A(544) and A(545);
w2117 <= A(544) and not A(545);
w2118 <= A(546) and not w2117;
w2119 <= not w2116 and w2118;
w2120 <= not w2116 and not w2117;
w2121 <= not A(546) and not w2120;
w2122 <= not w2119 and not w2121;
w2123 <= not w2115 and w2122;
w2124 <= w2115 and not w2122;
w2125 <= not w2123 and not w2124;
w2126 <= A(544) and A(545);
w2127 <= A(546) and not w2120;
w2128 <= not w2126 and not w2127;
w2129 <= A(541) and A(542);
w2130 <= A(543) and not w2113;
w2131 <= not w2129 and not w2130;
w2132 <= not w2128 and w2131;
w2133 <= w2128 and not w2131;
w2134 <= not w2132 and not w2133;
w2135 <= not w2115 and not w2122;
w2136 <= not w2134 and w2135;
w2137 <= not w2128 and not w2131;
w2138 <= not w2136 and not w2137;
w2139 <= not w2132 and w2135;
w2140 <= not w2133 and w2139;
w2141 <= not w2134 and not w2135;
w2142 <= not w2140 and not w2141;
w2143 <= not w2138 and not w2142;
w2144 <= not w2125 and not w2143;
w2145 <= not A(535) and A(536);
w2146 <= A(535) and not A(536);
w2147 <= A(537) and not w2146;
w2148 <= not w2145 and w2147;
w2149 <= not w2145 and not w2146;
w2150 <= not A(537) and not w2149;
w2151 <= not w2148 and not w2150;
w2152 <= not A(538) and A(539);
w2153 <= A(538) and not A(539);
w2154 <= A(540) and not w2153;
w2155 <= not w2152 and w2154;
w2156 <= not w2152 and not w2153;
w2157 <= not A(540) and not w2156;
w2158 <= not w2155 and not w2157;
w2159 <= not w2151 and w2158;
w2160 <= w2151 and not w2158;
w2161 <= not w2159 and not w2160;
w2162 <= A(538) and A(539);
w2163 <= A(540) and not w2156;
w2164 <= not w2162 and not w2163;
w2165 <= A(535) and A(536);
w2166 <= A(537) and not w2149;
w2167 <= not w2165 and not w2166;
w2168 <= not w2164 and w2167;
w2169 <= w2164 and not w2167;
w2170 <= not w2168 and not w2169;
w2171 <= not w2151 and not w2158;
w2172 <= not w2170 and w2171;
w2173 <= not w2164 and not w2167;
w2174 <= not w2172 and not w2173;
w2175 <= not w2168 and w2171;
w2176 <= not w2169 and w2175;
w2177 <= not w2170 and not w2171;
w2178 <= not w2176 and not w2177;
w2179 <= not w2174 and not w2178;
w2180 <= not w2161 and not w2179;
w2181 <= not w2144 and w2180;
w2182 <= w2144 and not w2180;
w2183 <= not w2181 and not w2182;
w2184 <= not w2108 and w2183;
w2185 <= w2108 and not w2183;
w2186 <= not w2184 and not w2185;
w2187 <= not A(529) and A(530);
w2188 <= A(529) and not A(530);
w2189 <= A(531) and not w2188;
w2190 <= not w2187 and w2189;
w2191 <= not w2187 and not w2188;
w2192 <= not A(531) and not w2191;
w2193 <= not w2190 and not w2192;
w2194 <= not A(532) and A(533);
w2195 <= A(532) and not A(533);
w2196 <= A(534) and not w2195;
w2197 <= not w2194 and w2196;
w2198 <= not w2194 and not w2195;
w2199 <= not A(534) and not w2198;
w2200 <= not w2197 and not w2199;
w2201 <= not w2193 and w2200;
w2202 <= w2193 and not w2200;
w2203 <= not w2201 and not w2202;
w2204 <= A(532) and A(533);
w2205 <= A(534) and not w2198;
w2206 <= not w2204 and not w2205;
w2207 <= A(529) and A(530);
w2208 <= A(531) and not w2191;
w2209 <= not w2207 and not w2208;
w2210 <= not w2206 and w2209;
w2211 <= w2206 and not w2209;
w2212 <= not w2210 and not w2211;
w2213 <= not w2193 and not w2200;
w2214 <= not w2212 and w2213;
w2215 <= not w2206 and not w2209;
w2216 <= not w2214 and not w2215;
w2217 <= not w2210 and w2213;
w2218 <= not w2211 and w2217;
w2219 <= not w2212 and not w2213;
w2220 <= not w2218 and not w2219;
w2221 <= not w2216 and not w2220;
w2222 <= not w2203 and not w2221;
w2223 <= not A(523) and A(524);
w2224 <= A(523) and not A(524);
w2225 <= A(525) and not w2224;
w2226 <= not w2223 and w2225;
w2227 <= not w2223 and not w2224;
w2228 <= not A(525) and not w2227;
w2229 <= not w2226 and not w2228;
w2230 <= not A(526) and A(527);
w2231 <= A(526) and not A(527);
w2232 <= A(528) and not w2231;
w2233 <= not w2230 and w2232;
w2234 <= not w2230 and not w2231;
w2235 <= not A(528) and not w2234;
w2236 <= not w2233 and not w2235;
w2237 <= not w2229 and w2236;
w2238 <= w2229 and not w2236;
w2239 <= not w2237 and not w2238;
w2240 <= A(526) and A(527);
w2241 <= A(528) and not w2234;
w2242 <= not w2240 and not w2241;
w2243 <= A(523) and A(524);
w2244 <= A(525) and not w2227;
w2245 <= not w2243 and not w2244;
w2246 <= not w2242 and w2245;
w2247 <= w2242 and not w2245;
w2248 <= not w2246 and not w2247;
w2249 <= not w2229 and not w2236;
w2250 <= not w2248 and w2249;
w2251 <= not w2242 and not w2245;
w2252 <= not w2250 and not w2251;
w2253 <= not w2246 and w2249;
w2254 <= not w2247 and w2253;
w2255 <= not w2248 and not w2249;
w2256 <= not w2254 and not w2255;
w2257 <= not w2252 and not w2256;
w2258 <= not w2239 and not w2257;
w2259 <= not w2222 and w2258;
w2260 <= w2222 and not w2258;
w2261 <= not w2259 and not w2260;
w2262 <= not A(517) and A(518);
w2263 <= A(517) and not A(518);
w2264 <= A(519) and not w2263;
w2265 <= not w2262 and w2264;
w2266 <= not w2262 and not w2263;
w2267 <= not A(519) and not w2266;
w2268 <= not w2265 and not w2267;
w2269 <= not A(520) and A(521);
w2270 <= A(520) and not A(521);
w2271 <= A(522) and not w2270;
w2272 <= not w2269 and w2271;
w2273 <= not w2269 and not w2270;
w2274 <= not A(522) and not w2273;
w2275 <= not w2272 and not w2274;
w2276 <= not w2268 and w2275;
w2277 <= w2268 and not w2275;
w2278 <= not w2276 and not w2277;
w2279 <= A(520) and A(521);
w2280 <= A(522) and not w2273;
w2281 <= not w2279 and not w2280;
w2282 <= A(517) and A(518);
w2283 <= A(519) and not w2266;
w2284 <= not w2282 and not w2283;
w2285 <= not w2281 and w2284;
w2286 <= w2281 and not w2284;
w2287 <= not w2285 and not w2286;
w2288 <= not w2268 and not w2275;
w2289 <= not w2287 and w2288;
w2290 <= not w2281 and not w2284;
w2291 <= not w2289 and not w2290;
w2292 <= not w2285 and w2288;
w2293 <= not w2286 and w2292;
w2294 <= not w2287 and not w2288;
w2295 <= not w2293 and not w2294;
w2296 <= not w2291 and not w2295;
w2297 <= not w2278 and not w2296;
w2298 <= not A(511) and A(512);
w2299 <= A(511) and not A(512);
w2300 <= A(513) and not w2299;
w2301 <= not w2298 and w2300;
w2302 <= not w2298 and not w2299;
w2303 <= not A(513) and not w2302;
w2304 <= not w2301 and not w2303;
w2305 <= not A(514) and A(515);
w2306 <= A(514) and not A(515);
w2307 <= A(516) and not w2306;
w2308 <= not w2305 and w2307;
w2309 <= not w2305 and not w2306;
w2310 <= not A(516) and not w2309;
w2311 <= not w2308 and not w2310;
w2312 <= not w2304 and w2311;
w2313 <= w2304 and not w2311;
w2314 <= not w2312 and not w2313;
w2315 <= A(514) and A(515);
w2316 <= A(516) and not w2309;
w2317 <= not w2315 and not w2316;
w2318 <= A(511) and A(512);
w2319 <= A(513) and not w2302;
w2320 <= not w2318 and not w2319;
w2321 <= not w2317 and w2320;
w2322 <= w2317 and not w2320;
w2323 <= not w2321 and not w2322;
w2324 <= not w2304 and not w2311;
w2325 <= not w2323 and w2324;
w2326 <= not w2317 and not w2320;
w2327 <= not w2325 and not w2326;
w2328 <= not w2321 and w2324;
w2329 <= not w2322 and w2328;
w2330 <= not w2323 and not w2324;
w2331 <= not w2329 and not w2330;
w2332 <= not w2327 and not w2331;
w2333 <= not w2314 and not w2332;
w2334 <= not w2297 and w2333;
w2335 <= w2297 and not w2333;
w2336 <= not w2334 and not w2335;
w2337 <= not w2261 and w2336;
w2338 <= w2261 and not w2336;
w2339 <= not w2337 and not w2338;
w2340 <= not w2186 and w2339;
w2341 <= w2186 and not w2339;
w2342 <= not w2340 and not w2341;
w2343 <= not w2033 and w2342;
w2344 <= w2033 and not w2342;
w2345 <= not w2343 and not w2344;
w2346 <= not A(649) and A(650);
w2347 <= A(649) and not A(650);
w2348 <= A(651) and not w2347;
w2349 <= not w2346 and w2348;
w2350 <= not w2346 and not w2347;
w2351 <= not A(651) and not w2350;
w2352 <= not w2349 and not w2351;
w2353 <= not A(652) and A(653);
w2354 <= A(652) and not A(653);
w2355 <= A(654) and not w2354;
w2356 <= not w2353 and w2355;
w2357 <= not w2353 and not w2354;
w2358 <= not A(654) and not w2357;
w2359 <= not w2356 and not w2358;
w2360 <= not w2352 and w2359;
w2361 <= w2352 and not w2359;
w2362 <= not w2360 and not w2361;
w2363 <= A(652) and A(653);
w2364 <= A(654) and not w2357;
w2365 <= not w2363 and not w2364;
w2366 <= A(649) and A(650);
w2367 <= A(651) and not w2350;
w2368 <= not w2366 and not w2367;
w2369 <= not w2365 and w2368;
w2370 <= w2365 and not w2368;
w2371 <= not w2369 and not w2370;
w2372 <= not w2352 and not w2359;
w2373 <= not w2371 and w2372;
w2374 <= not w2365 and not w2368;
w2375 <= not w2373 and not w2374;
w2376 <= not w2369 and w2372;
w2377 <= not w2370 and w2376;
w2378 <= not w2371 and not w2372;
w2379 <= not w2377 and not w2378;
w2380 <= not w2375 and not w2379;
w2381 <= not w2362 and not w2380;
w2382 <= not A(643) and A(644);
w2383 <= A(643) and not A(644);
w2384 <= A(645) and not w2383;
w2385 <= not w2382 and w2384;
w2386 <= not w2382 and not w2383;
w2387 <= not A(645) and not w2386;
w2388 <= not w2385 and not w2387;
w2389 <= not A(646) and A(647);
w2390 <= A(646) and not A(647);
w2391 <= A(648) and not w2390;
w2392 <= not w2389 and w2391;
w2393 <= not w2389 and not w2390;
w2394 <= not A(648) and not w2393;
w2395 <= not w2392 and not w2394;
w2396 <= not w2388 and w2395;
w2397 <= w2388 and not w2395;
w2398 <= not w2396 and not w2397;
w2399 <= A(646) and A(647);
w2400 <= A(648) and not w2393;
w2401 <= not w2399 and not w2400;
w2402 <= A(643) and A(644);
w2403 <= A(645) and not w2386;
w2404 <= not w2402 and not w2403;
w2405 <= not w2401 and w2404;
w2406 <= w2401 and not w2404;
w2407 <= not w2405 and not w2406;
w2408 <= not w2388 and not w2395;
w2409 <= not w2407 and w2408;
w2410 <= not w2401 and not w2404;
w2411 <= not w2409 and not w2410;
w2412 <= not w2405 and w2408;
w2413 <= not w2406 and w2412;
w2414 <= not w2407 and not w2408;
w2415 <= not w2413 and not w2414;
w2416 <= not w2411 and not w2415;
w2417 <= not w2398 and not w2416;
w2418 <= not w2381 and w2417;
w2419 <= w2381 and not w2417;
w2420 <= not w2418 and not w2419;
w2421 <= not A(637) and A(638);
w2422 <= A(637) and not A(638);
w2423 <= A(639) and not w2422;
w2424 <= not w2421 and w2423;
w2425 <= not w2421 and not w2422;
w2426 <= not A(639) and not w2425;
w2427 <= not w2424 and not w2426;
w2428 <= not A(640) and A(641);
w2429 <= A(640) and not A(641);
w2430 <= A(642) and not w2429;
w2431 <= not w2428 and w2430;
w2432 <= not w2428 and not w2429;
w2433 <= not A(642) and not w2432;
w2434 <= not w2431 and not w2433;
w2435 <= not w2427 and w2434;
w2436 <= w2427 and not w2434;
w2437 <= not w2435 and not w2436;
w2438 <= A(640) and A(641);
w2439 <= A(642) and not w2432;
w2440 <= not w2438 and not w2439;
w2441 <= A(637) and A(638);
w2442 <= A(639) and not w2425;
w2443 <= not w2441 and not w2442;
w2444 <= not w2440 and w2443;
w2445 <= w2440 and not w2443;
w2446 <= not w2444 and not w2445;
w2447 <= not w2427 and not w2434;
w2448 <= not w2446 and w2447;
w2449 <= not w2440 and not w2443;
w2450 <= not w2448 and not w2449;
w2451 <= not w2444 and w2447;
w2452 <= not w2445 and w2451;
w2453 <= not w2446 and not w2447;
w2454 <= not w2452 and not w2453;
w2455 <= not w2450 and not w2454;
w2456 <= not w2437 and not w2455;
w2457 <= not A(631) and A(632);
w2458 <= A(631) and not A(632);
w2459 <= A(633) and not w2458;
w2460 <= not w2457 and w2459;
w2461 <= not w2457 and not w2458;
w2462 <= not A(633) and not w2461;
w2463 <= not w2460 and not w2462;
w2464 <= not A(634) and A(635);
w2465 <= A(634) and not A(635);
w2466 <= A(636) and not w2465;
w2467 <= not w2464 and w2466;
w2468 <= not w2464 and not w2465;
w2469 <= not A(636) and not w2468;
w2470 <= not w2467 and not w2469;
w2471 <= not w2463 and w2470;
w2472 <= w2463 and not w2470;
w2473 <= not w2471 and not w2472;
w2474 <= A(634) and A(635);
w2475 <= A(636) and not w2468;
w2476 <= not w2474 and not w2475;
w2477 <= A(631) and A(632);
w2478 <= A(633) and not w2461;
w2479 <= not w2477 and not w2478;
w2480 <= not w2476 and w2479;
w2481 <= w2476 and not w2479;
w2482 <= not w2480 and not w2481;
w2483 <= not w2463 and not w2470;
w2484 <= not w2482 and w2483;
w2485 <= not w2476 and not w2479;
w2486 <= not w2484 and not w2485;
w2487 <= not w2480 and w2483;
w2488 <= not w2481 and w2487;
w2489 <= not w2482 and not w2483;
w2490 <= not w2488 and not w2489;
w2491 <= not w2486 and not w2490;
w2492 <= not w2473 and not w2491;
w2493 <= not w2456 and w2492;
w2494 <= w2456 and not w2492;
w2495 <= not w2493 and not w2494;
w2496 <= not w2420 and w2495;
w2497 <= w2420 and not w2495;
w2498 <= not w2496 and not w2497;
w2499 <= not A(625) and A(626);
w2500 <= A(625) and not A(626);
w2501 <= A(627) and not w2500;
w2502 <= not w2499 and w2501;
w2503 <= not w2499 and not w2500;
w2504 <= not A(627) and not w2503;
w2505 <= not w2502 and not w2504;
w2506 <= not A(628) and A(629);
w2507 <= A(628) and not A(629);
w2508 <= A(630) and not w2507;
w2509 <= not w2506 and w2508;
w2510 <= not w2506 and not w2507;
w2511 <= not A(630) and not w2510;
w2512 <= not w2509 and not w2511;
w2513 <= not w2505 and w2512;
w2514 <= w2505 and not w2512;
w2515 <= not w2513 and not w2514;
w2516 <= A(628) and A(629);
w2517 <= A(630) and not w2510;
w2518 <= not w2516 and not w2517;
w2519 <= A(625) and A(626);
w2520 <= A(627) and not w2503;
w2521 <= not w2519 and not w2520;
w2522 <= not w2518 and w2521;
w2523 <= w2518 and not w2521;
w2524 <= not w2522 and not w2523;
w2525 <= not w2505 and not w2512;
w2526 <= not w2524 and w2525;
w2527 <= not w2518 and not w2521;
w2528 <= not w2526 and not w2527;
w2529 <= not w2522 and w2525;
w2530 <= not w2523 and w2529;
w2531 <= not w2524 and not w2525;
w2532 <= not w2530 and not w2531;
w2533 <= not w2528 and not w2532;
w2534 <= not w2515 and not w2533;
w2535 <= not A(619) and A(620);
w2536 <= A(619) and not A(620);
w2537 <= A(621) and not w2536;
w2538 <= not w2535 and w2537;
w2539 <= not w2535 and not w2536;
w2540 <= not A(621) and not w2539;
w2541 <= not w2538 and not w2540;
w2542 <= not A(622) and A(623);
w2543 <= A(622) and not A(623);
w2544 <= A(624) and not w2543;
w2545 <= not w2542 and w2544;
w2546 <= not w2542 and not w2543;
w2547 <= not A(624) and not w2546;
w2548 <= not w2545 and not w2547;
w2549 <= not w2541 and w2548;
w2550 <= w2541 and not w2548;
w2551 <= not w2549 and not w2550;
w2552 <= A(622) and A(623);
w2553 <= A(624) and not w2546;
w2554 <= not w2552 and not w2553;
w2555 <= A(619) and A(620);
w2556 <= A(621) and not w2539;
w2557 <= not w2555 and not w2556;
w2558 <= not w2554 and w2557;
w2559 <= w2554 and not w2557;
w2560 <= not w2558 and not w2559;
w2561 <= not w2541 and not w2548;
w2562 <= not w2560 and w2561;
w2563 <= not w2554 and not w2557;
w2564 <= not w2562 and not w2563;
w2565 <= not w2558 and w2561;
w2566 <= not w2559 and w2565;
w2567 <= not w2560 and not w2561;
w2568 <= not w2566 and not w2567;
w2569 <= not w2564 and not w2568;
w2570 <= not w2551 and not w2569;
w2571 <= not w2534 and w2570;
w2572 <= w2534 and not w2570;
w2573 <= not w2571 and not w2572;
w2574 <= not A(613) and A(614);
w2575 <= A(613) and not A(614);
w2576 <= A(615) and not w2575;
w2577 <= not w2574 and w2576;
w2578 <= not w2574 and not w2575;
w2579 <= not A(615) and not w2578;
w2580 <= not w2577 and not w2579;
w2581 <= not A(616) and A(617);
w2582 <= A(616) and not A(617);
w2583 <= A(618) and not w2582;
w2584 <= not w2581 and w2583;
w2585 <= not w2581 and not w2582;
w2586 <= not A(618) and not w2585;
w2587 <= not w2584 and not w2586;
w2588 <= not w2580 and w2587;
w2589 <= w2580 and not w2587;
w2590 <= not w2588 and not w2589;
w2591 <= A(616) and A(617);
w2592 <= A(618) and not w2585;
w2593 <= not w2591 and not w2592;
w2594 <= A(613) and A(614);
w2595 <= A(615) and not w2578;
w2596 <= not w2594 and not w2595;
w2597 <= not w2593 and w2596;
w2598 <= w2593 and not w2596;
w2599 <= not w2597 and not w2598;
w2600 <= not w2580 and not w2587;
w2601 <= not w2599 and w2600;
w2602 <= not w2593 and not w2596;
w2603 <= not w2601 and not w2602;
w2604 <= not w2597 and w2600;
w2605 <= not w2598 and w2604;
w2606 <= not w2599 and not w2600;
w2607 <= not w2605 and not w2606;
w2608 <= not w2603 and not w2607;
w2609 <= not w2590 and not w2608;
w2610 <= not A(607) and A(608);
w2611 <= A(607) and not A(608);
w2612 <= A(609) and not w2611;
w2613 <= not w2610 and w2612;
w2614 <= not w2610 and not w2611;
w2615 <= not A(609) and not w2614;
w2616 <= not w2613 and not w2615;
w2617 <= not A(610) and A(611);
w2618 <= A(610) and not A(611);
w2619 <= A(612) and not w2618;
w2620 <= not w2617 and w2619;
w2621 <= not w2617 and not w2618;
w2622 <= not A(612) and not w2621;
w2623 <= not w2620 and not w2622;
w2624 <= not w2616 and w2623;
w2625 <= w2616 and not w2623;
w2626 <= not w2624 and not w2625;
w2627 <= A(610) and A(611);
w2628 <= A(612) and not w2621;
w2629 <= not w2627 and not w2628;
w2630 <= A(607) and A(608);
w2631 <= A(609) and not w2614;
w2632 <= not w2630 and not w2631;
w2633 <= not w2629 and w2632;
w2634 <= w2629 and not w2632;
w2635 <= not w2633 and not w2634;
w2636 <= not w2616 and not w2623;
w2637 <= not w2635 and w2636;
w2638 <= not w2629 and not w2632;
w2639 <= not w2637 and not w2638;
w2640 <= not w2633 and w2636;
w2641 <= not w2634 and w2640;
w2642 <= not w2635 and not w2636;
w2643 <= not w2641 and not w2642;
w2644 <= not w2639 and not w2643;
w2645 <= not w2626 and not w2644;
w2646 <= not w2609 and w2645;
w2647 <= w2609 and not w2645;
w2648 <= not w2646 and not w2647;
w2649 <= not w2573 and w2648;
w2650 <= w2573 and not w2648;
w2651 <= not w2649 and not w2650;
w2652 <= not w2498 and w2651;
w2653 <= w2498 and not w2651;
w2654 <= not w2652 and not w2653;
w2655 <= not A(601) and A(602);
w2656 <= A(601) and not A(602);
w2657 <= A(603) and not w2656;
w2658 <= not w2655 and w2657;
w2659 <= not w2655 and not w2656;
w2660 <= not A(603) and not w2659;
w2661 <= not w2658 and not w2660;
w2662 <= not A(604) and A(605);
w2663 <= A(604) and not A(605);
w2664 <= A(606) and not w2663;
w2665 <= not w2662 and w2664;
w2666 <= not w2662 and not w2663;
w2667 <= not A(606) and not w2666;
w2668 <= not w2665 and not w2667;
w2669 <= not w2661 and w2668;
w2670 <= w2661 and not w2668;
w2671 <= not w2669 and not w2670;
w2672 <= A(604) and A(605);
w2673 <= A(606) and not w2666;
w2674 <= not w2672 and not w2673;
w2675 <= A(601) and A(602);
w2676 <= A(603) and not w2659;
w2677 <= not w2675 and not w2676;
w2678 <= not w2674 and w2677;
w2679 <= w2674 and not w2677;
w2680 <= not w2678 and not w2679;
w2681 <= not w2661 and not w2668;
w2682 <= not w2680 and w2681;
w2683 <= not w2674 and not w2677;
w2684 <= not w2682 and not w2683;
w2685 <= not w2678 and w2681;
w2686 <= not w2679 and w2685;
w2687 <= not w2680 and not w2681;
w2688 <= not w2686 and not w2687;
w2689 <= not w2684 and not w2688;
w2690 <= not w2671 and not w2689;
w2691 <= not A(595) and A(596);
w2692 <= A(595) and not A(596);
w2693 <= A(597) and not w2692;
w2694 <= not w2691 and w2693;
w2695 <= not w2691 and not w2692;
w2696 <= not A(597) and not w2695;
w2697 <= not w2694 and not w2696;
w2698 <= not A(598) and A(599);
w2699 <= A(598) and not A(599);
w2700 <= A(600) and not w2699;
w2701 <= not w2698 and w2700;
w2702 <= not w2698 and not w2699;
w2703 <= not A(600) and not w2702;
w2704 <= not w2701 and not w2703;
w2705 <= not w2697 and w2704;
w2706 <= w2697 and not w2704;
w2707 <= not w2705 and not w2706;
w2708 <= A(598) and A(599);
w2709 <= A(600) and not w2702;
w2710 <= not w2708 and not w2709;
w2711 <= A(595) and A(596);
w2712 <= A(597) and not w2695;
w2713 <= not w2711 and not w2712;
w2714 <= not w2710 and w2713;
w2715 <= w2710 and not w2713;
w2716 <= not w2714 and not w2715;
w2717 <= not w2697 and not w2704;
w2718 <= not w2716 and w2717;
w2719 <= not w2710 and not w2713;
w2720 <= not w2718 and not w2719;
w2721 <= not w2714 and w2717;
w2722 <= not w2715 and w2721;
w2723 <= not w2716 and not w2717;
w2724 <= not w2722 and not w2723;
w2725 <= not w2720 and not w2724;
w2726 <= not w2707 and not w2725;
w2727 <= not w2690 and w2726;
w2728 <= w2690 and not w2726;
w2729 <= not w2727 and not w2728;
w2730 <= not A(589) and A(590);
w2731 <= A(589) and not A(590);
w2732 <= A(591) and not w2731;
w2733 <= not w2730 and w2732;
w2734 <= not w2730 and not w2731;
w2735 <= not A(591) and not w2734;
w2736 <= not w2733 and not w2735;
w2737 <= not A(592) and A(593);
w2738 <= A(592) and not A(593);
w2739 <= A(594) and not w2738;
w2740 <= not w2737 and w2739;
w2741 <= not w2737 and not w2738;
w2742 <= not A(594) and not w2741;
w2743 <= not w2740 and not w2742;
w2744 <= not w2736 and w2743;
w2745 <= w2736 and not w2743;
w2746 <= not w2744 and not w2745;
w2747 <= A(592) and A(593);
w2748 <= A(594) and not w2741;
w2749 <= not w2747 and not w2748;
w2750 <= A(589) and A(590);
w2751 <= A(591) and not w2734;
w2752 <= not w2750 and not w2751;
w2753 <= not w2749 and w2752;
w2754 <= w2749 and not w2752;
w2755 <= not w2753 and not w2754;
w2756 <= not w2736 and not w2743;
w2757 <= not w2755 and w2756;
w2758 <= not w2749 and not w2752;
w2759 <= not w2757 and not w2758;
w2760 <= not w2753 and w2756;
w2761 <= not w2754 and w2760;
w2762 <= not w2755 and not w2756;
w2763 <= not w2761 and not w2762;
w2764 <= not w2759 and not w2763;
w2765 <= not w2746 and not w2764;
w2766 <= not A(583) and A(584);
w2767 <= A(583) and not A(584);
w2768 <= A(585) and not w2767;
w2769 <= not w2766 and w2768;
w2770 <= not w2766 and not w2767;
w2771 <= not A(585) and not w2770;
w2772 <= not w2769 and not w2771;
w2773 <= not A(586) and A(587);
w2774 <= A(586) and not A(587);
w2775 <= A(588) and not w2774;
w2776 <= not w2773 and w2775;
w2777 <= not w2773 and not w2774;
w2778 <= not A(588) and not w2777;
w2779 <= not w2776 and not w2778;
w2780 <= not w2772 and w2779;
w2781 <= w2772 and not w2779;
w2782 <= not w2780 and not w2781;
w2783 <= A(586) and A(587);
w2784 <= A(588) and not w2777;
w2785 <= not w2783 and not w2784;
w2786 <= A(583) and A(584);
w2787 <= A(585) and not w2770;
w2788 <= not w2786 and not w2787;
w2789 <= not w2785 and w2788;
w2790 <= w2785 and not w2788;
w2791 <= not w2789 and not w2790;
w2792 <= not w2772 and not w2779;
w2793 <= not w2791 and w2792;
w2794 <= not w2785 and not w2788;
w2795 <= not w2793 and not w2794;
w2796 <= not w2789 and w2792;
w2797 <= not w2790 and w2796;
w2798 <= not w2791 and not w2792;
w2799 <= not w2797 and not w2798;
w2800 <= not w2795 and not w2799;
w2801 <= not w2782 and not w2800;
w2802 <= not w2765 and w2801;
w2803 <= w2765 and not w2801;
w2804 <= not w2802 and not w2803;
w2805 <= not w2729 and w2804;
w2806 <= w2729 and not w2804;
w2807 <= not w2805 and not w2806;
w2808 <= not A(577) and A(578);
w2809 <= A(577) and not A(578);
w2810 <= A(579) and not w2809;
w2811 <= not w2808 and w2810;
w2812 <= not w2808 and not w2809;
w2813 <= not A(579) and not w2812;
w2814 <= not w2811 and not w2813;
w2815 <= not A(580) and A(581);
w2816 <= A(580) and not A(581);
w2817 <= A(582) and not w2816;
w2818 <= not w2815 and w2817;
w2819 <= not w2815 and not w2816;
w2820 <= not A(582) and not w2819;
w2821 <= not w2818 and not w2820;
w2822 <= not w2814 and w2821;
w2823 <= w2814 and not w2821;
w2824 <= not w2822 and not w2823;
w2825 <= A(580) and A(581);
w2826 <= A(582) and not w2819;
w2827 <= not w2825 and not w2826;
w2828 <= A(577) and A(578);
w2829 <= A(579) and not w2812;
w2830 <= not w2828 and not w2829;
w2831 <= not w2827 and w2830;
w2832 <= w2827 and not w2830;
w2833 <= not w2831 and not w2832;
w2834 <= not w2814 and not w2821;
w2835 <= not w2833 and w2834;
w2836 <= not w2827 and not w2830;
w2837 <= not w2835 and not w2836;
w2838 <= not w2831 and w2834;
w2839 <= not w2832 and w2838;
w2840 <= not w2833 and not w2834;
w2841 <= not w2839 and not w2840;
w2842 <= not w2837 and not w2841;
w2843 <= not w2824 and not w2842;
w2844 <= not A(571) and A(572);
w2845 <= A(571) and not A(572);
w2846 <= A(573) and not w2845;
w2847 <= not w2844 and w2846;
w2848 <= not w2844 and not w2845;
w2849 <= not A(573) and not w2848;
w2850 <= not w2847 and not w2849;
w2851 <= not A(574) and A(575);
w2852 <= A(574) and not A(575);
w2853 <= A(576) and not w2852;
w2854 <= not w2851 and w2853;
w2855 <= not w2851 and not w2852;
w2856 <= not A(576) and not w2855;
w2857 <= not w2854 and not w2856;
w2858 <= not w2850 and w2857;
w2859 <= w2850 and not w2857;
w2860 <= not w2858 and not w2859;
w2861 <= A(574) and A(575);
w2862 <= A(576) and not w2855;
w2863 <= not w2861 and not w2862;
w2864 <= A(571) and A(572);
w2865 <= A(573) and not w2848;
w2866 <= not w2864 and not w2865;
w2867 <= not w2863 and w2866;
w2868 <= w2863 and not w2866;
w2869 <= not w2867 and not w2868;
w2870 <= not w2850 and not w2857;
w2871 <= not w2869 and w2870;
w2872 <= not w2863 and not w2866;
w2873 <= not w2871 and not w2872;
w2874 <= not w2867 and w2870;
w2875 <= not w2868 and w2874;
w2876 <= not w2869 and not w2870;
w2877 <= not w2875 and not w2876;
w2878 <= not w2873 and not w2877;
w2879 <= not w2860 and not w2878;
w2880 <= not w2843 and w2879;
w2881 <= w2843 and not w2879;
w2882 <= not w2880 and not w2881;
w2883 <= not A(565) and A(566);
w2884 <= A(565) and not A(566);
w2885 <= A(567) and not w2884;
w2886 <= not w2883 and w2885;
w2887 <= not w2883 and not w2884;
w2888 <= not A(567) and not w2887;
w2889 <= not w2886 and not w2888;
w2890 <= not A(568) and A(569);
w2891 <= A(568) and not A(569);
w2892 <= A(570) and not w2891;
w2893 <= not w2890 and w2892;
w2894 <= not w2890 and not w2891;
w2895 <= not A(570) and not w2894;
w2896 <= not w2893 and not w2895;
w2897 <= not w2889 and w2896;
w2898 <= w2889 and not w2896;
w2899 <= not w2897 and not w2898;
w2900 <= A(568) and A(569);
w2901 <= A(570) and not w2894;
w2902 <= not w2900 and not w2901;
w2903 <= A(565) and A(566);
w2904 <= A(567) and not w2887;
w2905 <= not w2903 and not w2904;
w2906 <= not w2902 and w2905;
w2907 <= w2902 and not w2905;
w2908 <= not w2906 and not w2907;
w2909 <= not w2889 and not w2896;
w2910 <= not w2908 and w2909;
w2911 <= not w2902 and not w2905;
w2912 <= not w2910 and not w2911;
w2913 <= not w2906 and w2909;
w2914 <= not w2907 and w2913;
w2915 <= not w2908 and not w2909;
w2916 <= not w2914 and not w2915;
w2917 <= not w2912 and not w2916;
w2918 <= not w2899 and not w2917;
w2919 <= not A(559) and A(560);
w2920 <= A(559) and not A(560);
w2921 <= A(561) and not w2920;
w2922 <= not w2919 and w2921;
w2923 <= not w2919 and not w2920;
w2924 <= not A(561) and not w2923;
w2925 <= not w2922 and not w2924;
w2926 <= not A(562) and A(563);
w2927 <= A(562) and not A(563);
w2928 <= A(564) and not w2927;
w2929 <= not w2926 and w2928;
w2930 <= not w2926 and not w2927;
w2931 <= not A(564) and not w2930;
w2932 <= not w2929 and not w2931;
w2933 <= not w2925 and w2932;
w2934 <= w2925 and not w2932;
w2935 <= not w2933 and not w2934;
w2936 <= A(562) and A(563);
w2937 <= A(564) and not w2930;
w2938 <= not w2936 and not w2937;
w2939 <= A(559) and A(560);
w2940 <= A(561) and not w2923;
w2941 <= not w2939 and not w2940;
w2942 <= not w2938 and w2941;
w2943 <= w2938 and not w2941;
w2944 <= not w2942 and not w2943;
w2945 <= not w2925 and not w2932;
w2946 <= not w2944 and w2945;
w2947 <= not w2938 and not w2941;
w2948 <= not w2946 and not w2947;
w2949 <= not w2942 and w2945;
w2950 <= not w2943 and w2949;
w2951 <= not w2944 and not w2945;
w2952 <= not w2950 and not w2951;
w2953 <= not w2948 and not w2952;
w2954 <= not w2935 and not w2953;
w2955 <= not w2918 and w2954;
w2956 <= w2918 and not w2954;
w2957 <= not w2955 and not w2956;
w2958 <= not w2882 and w2957;
w2959 <= w2882 and not w2957;
w2960 <= not w2958 and not w2959;
w2961 <= not w2807 and w2960;
w2962 <= w2807 and not w2960;
w2963 <= not w2961 and not w2962;
w2964 <= not w2654 and w2963;
w2965 <= w2654 and not w2963;
w2966 <= not w2964 and not w2965;
w2967 <= not w2345 and w2966;
w2968 <= w2345 and not w2966;
w2969 <= not w2967 and not w2968;
w2970 <= not w1709 and w1712;
w2971 <= w1709 and not w1712;
w2972 <= not w2970 and not w2971;
w2973 <= not w2969 and not w2972;
w2974 <= not w1724 and w2973;
w2975 <= not w1719 and w2974;
w2976 <= not w1719 and not w1724;
w2977 <= not w2973 and not w2976;
w2978 <= not w2975 and not w2977;
w2979 <= not w2782 and not w2795;
w2980 <= not w2799 and not w2979;
w2981 <= not w2746 and not w2782;
w2982 <= not w2764 and w2981;
w2983 <= not w2800 and w2982;
w2984 <= not w2746 and not w2759;
w2985 <= not w2763 and not w2984;
w2986 <= not w2983 and w2985;
w2987 <= w2983 and not w2985;
w2988 <= not w2986 and not w2987;
w2989 <= not w2980 and not w2988;
w2990 <= not w2983 and not w2985;
w2991 <= not w2763 and w2981;
w2992 <= not w2764 and w2991;
w2993 <= not w2800 and not w2984;
w2994 <= w2992 and w2993;
w2995 <= not w2990 and not w2994;
w2996 <= w2980 and not w2995;
w2997 <= not w2989 and not w2996;
w2998 <= not w2707 and not w2720;
w2999 <= not w2724 and not w2998;
w3000 <= not w2671 and not w2707;
w3001 <= not w2689 and w3000;
w3002 <= not w2725 and w3001;
w3003 <= not w2671 and not w2684;
w3004 <= not w2688 and not w3003;
w3005 <= not w3002 and not w3004;
w3006 <= not w2688 and w3000;
w3007 <= not w2689 and w3006;
w3008 <= not w2725 and not w3003;
w3009 <= w3007 and w3008;
w3010 <= not w3005 and not w3009;
w3011 <= w2999 and not w3010;
w3012 <= not w3002 and w3004;
w3013 <= w3002 and not w3004;
w3014 <= not w3012 and not w3013;
w3015 <= not w2999 and not w3014;
w3016 <= not w2729 and not w2804;
w3017 <= not w3015 and not w3016;
w3018 <= not w3011 and w3017;
w3019 <= not w3011 and not w3015;
w3020 <= w3016 and not w3019;
w3021 <= not w3018 and not w3020;
w3022 <= not w2997 and not w3021;
w3023 <= not w3015 and w3016;
w3024 <= not w3011 and w3023;
w3025 <= not w3016 and not w3019;
w3026 <= not w3024 and not w3025;
w3027 <= w2997 and not w3026;
w3028 <= not w2807 and not w2960;
w3029 <= not w3027 and w3028;
w3030 <= not w3022 and w3029;
w3031 <= not w3022 and not w3027;
w3032 <= not w3028 and not w3031;
w3033 <= not w3030 and not w3032;
w3034 <= not w2860 and not w2873;
w3035 <= not w2877 and not w3034;
w3036 <= not w2824 and not w2860;
w3037 <= not w2842 and w3036;
w3038 <= not w2878 and w3037;
w3039 <= not w2824 and not w2837;
w3040 <= not w2841 and not w3039;
w3041 <= not w3038 and not w3040;
w3042 <= not w2841 and w3036;
w3043 <= not w2842 and w3042;
w3044 <= not w2878 and not w3039;
w3045 <= w3043 and w3044;
w3046 <= not w3041 and not w3045;
w3047 <= w3035 and not w3046;
w3048 <= not w3038 and w3040;
w3049 <= w3038 and not w3040;
w3050 <= not w3048 and not w3049;
w3051 <= not w3035 and not w3050;
w3052 <= not w2882 and not w2957;
w3053 <= not w3051 and w3052;
w3054 <= not w3047 and w3053;
w3055 <= not w3047 and not w3051;
w3056 <= not w3052 and not w3055;
w3057 <= not w3054 and not w3056;
w3058 <= not w2935 and not w2948;
w3059 <= not w2952 and not w3058;
w3060 <= not w2899 and not w2935;
w3061 <= not w2917 and w3060;
w3062 <= not w2953 and w3061;
w3063 <= not w2899 and not w2912;
w3064 <= not w2916 and not w3063;
w3065 <= not w3062 and w3064;
w3066 <= w3062 and not w3064;
w3067 <= not w3065 and not w3066;
w3068 <= not w3059 and not w3067;
w3069 <= not w3062 and not w3064;
w3070 <= not w2916 and w3060;
w3071 <= not w2917 and w3070;
w3072 <= not w2953 and not w3063;
w3073 <= w3071 and w3072;
w3074 <= not w3069 and not w3073;
w3075 <= w3059 and not w3074;
w3076 <= not w3068 and not w3075;
w3077 <= not w3057 and w3076;
w3078 <= not w3051 and not w3052;
w3079 <= not w3047 and w3078;
w3080 <= w3052 and not w3055;
w3081 <= not w3079 and not w3080;
w3082 <= not w3076 and not w3081;
w3083 <= not w3077 and not w3082;
w3084 <= not w3033 and w3083;
w3085 <= not w3027 and not w3028;
w3086 <= not w3022 and w3085;
w3087 <= w3028 and not w3031;
w3088 <= not w3086 and not w3087;
w3089 <= not w3083 and not w3088;
w3090 <= not w3084 and not w3089;
w3091 <= not w2551 and not w2564;
w3092 <= not w2568 and not w3091;
w3093 <= not w2515 and not w2551;
w3094 <= not w2533 and w3093;
w3095 <= not w2569 and w3094;
w3096 <= not w2515 and not w2528;
w3097 <= not w2532 and not w3096;
w3098 <= not w3095 and not w3097;
w3099 <= not w2532 and w3093;
w3100 <= not w2533 and w3099;
w3101 <= not w2569 and not w3096;
w3102 <= w3100 and w3101;
w3103 <= not w3098 and not w3102;
w3104 <= w3092 and not w3103;
w3105 <= not w3095 and w3097;
w3106 <= w3095 and not w3097;
w3107 <= not w3105 and not w3106;
w3108 <= not w3092 and not w3107;
w3109 <= not w2573 and not w2648;
w3110 <= not w3108 and w3109;
w3111 <= not w3104 and w3110;
w3112 <= not w3104 and not w3108;
w3113 <= not w3109 and not w3112;
w3114 <= not w3111 and not w3113;
w3115 <= not w2626 and not w2639;
w3116 <= not w2643 and not w3115;
w3117 <= not w2590 and not w2626;
w3118 <= not w2608 and w3117;
w3119 <= not w2644 and w3118;
w3120 <= not w2590 and not w2603;
w3121 <= not w2607 and not w3120;
w3122 <= not w3119 and w3121;
w3123 <= w3119 and not w3121;
w3124 <= not w3122 and not w3123;
w3125 <= not w3116 and not w3124;
w3126 <= not w3119 and not w3121;
w3127 <= not w2607 and w3117;
w3128 <= not w2608 and w3127;
w3129 <= not w2644 and not w3120;
w3130 <= w3128 and w3129;
w3131 <= not w3126 and not w3130;
w3132 <= w3116 and not w3131;
w3133 <= not w3125 and not w3132;
w3134 <= not w3114 and w3133;
w3135 <= not w3108 and not w3109;
w3136 <= not w3104 and w3135;
w3137 <= w3109 and not w3112;
w3138 <= not w3136 and not w3137;
w3139 <= not w3133 and not w3138;
w3140 <= not w3134 and not w3139;
w3141 <= not w2473 and not w2486;
w3142 <= not w2490 and not w3141;
w3143 <= not w2437 and not w2473;
w3144 <= not w2455 and w3143;
w3145 <= not w2491 and w3144;
w3146 <= not w2437 and not w2450;
w3147 <= not w2454 and not w3146;
w3148 <= not w3145 and w3147;
w3149 <= w3145 and not w3147;
w3150 <= not w3148 and not w3149;
w3151 <= not w3142 and not w3150;
w3152 <= not w3145 and not w3147;
w3153 <= not w2454 and w3143;
w3154 <= not w2455 and w3153;
w3155 <= not w2491 and not w3146;
w3156 <= w3154 and w3155;
w3157 <= not w3152 and not w3156;
w3158 <= w3142 and not w3157;
w3159 <= not w3151 and not w3158;
w3160 <= not w2398 and not w2411;
w3161 <= not w2415 and not w3160;
w3162 <= not w2362 and not w2398;
w3163 <= not w2380 and w3162;
w3164 <= not w2416 and w3163;
w3165 <= not w2362 and not w2375;
w3166 <= not w2379 and not w3165;
w3167 <= not w3164 and not w3166;
w3168 <= not w2379 and w3162;
w3169 <= not w2380 and w3168;
w3170 <= not w2416 and not w3165;
w3171 <= w3169 and w3170;
w3172 <= not w3167 and not w3171;
w3173 <= w3161 and not w3172;
w3174 <= not w3164 and w3166;
w3175 <= w3164 and not w3166;
w3176 <= not w3174 and not w3175;
w3177 <= not w3161 and not w3176;
w3178 <= not w2420 and not w2495;
w3179 <= not w3177 and not w3178;
w3180 <= not w3173 and w3179;
w3181 <= not w3173 and not w3177;
w3182 <= w3178 and not w3181;
w3183 <= not w3180 and not w3182;
w3184 <= not w3159 and not w3183;
w3185 <= not w3177 and w3178;
w3186 <= not w3173 and w3185;
w3187 <= not w3178 and not w3181;
w3188 <= not w3186 and not w3187;
w3189 <= w3159 and not w3188;
w3190 <= not w2498 and not w2651;
w3191 <= not w3189 and not w3190;
w3192 <= not w3184 and w3191;
w3193 <= not w3184 and not w3189;
w3194 <= w3190 and not w3193;
w3195 <= not w3192 and not w3194;
w3196 <= not w3140 and not w3195;
w3197 <= not w3189 and w3190;
w3198 <= not w3184 and w3197;
w3199 <= not w3190 and not w3193;
w3200 <= not w3198 and not w3199;
w3201 <= w3140 and not w3200;
w3202 <= not w2654 and not w2963;
w3203 <= not w3201 and not w3202;
w3204 <= not w3196 and w3203;
w3205 <= not w3196 and not w3201;
w3206 <= w3202 and not w3205;
w3207 <= not w3204 and not w3206;
w3208 <= not w3090 and not w3207;
w3209 <= not w3201 and w3202;
w3210 <= not w3196 and w3209;
w3211 <= not w3202 and not w3205;
w3212 <= not w3210 and not w3211;
w3213 <= w3090 and not w3212;
w3214 <= not w2345 and not w2966;
w3215 <= not w3213 and w3214;
w3216 <= not w3208 and w3215;
w3217 <= not w3208 and not w3213;
w3218 <= not w3214 and not w3217;
w3219 <= not w3216 and not w3218;
w3220 <= not w2239 and not w2252;
w3221 <= not w2256 and not w3220;
w3222 <= not w2203 and not w2239;
w3223 <= not w2221 and w3222;
w3224 <= not w2257 and w3223;
w3225 <= not w2203 and not w2216;
w3226 <= not w2220 and not w3225;
w3227 <= not w3224 and not w3226;
w3228 <= not w2220 and w3222;
w3229 <= not w2221 and w3228;
w3230 <= not w2257 and not w3225;
w3231 <= w3229 and w3230;
w3232 <= not w3227 and not w3231;
w3233 <= w3221 and not w3232;
w3234 <= not w3224 and w3226;
w3235 <= w3224 and not w3226;
w3236 <= not w3234 and not w3235;
w3237 <= not w3221 and not w3236;
w3238 <= not w2261 and not w2336;
w3239 <= not w3237 and w3238;
w3240 <= not w3233 and w3239;
w3241 <= not w3233 and not w3237;
w3242 <= not w3238 and not w3241;
w3243 <= not w3240 and not w3242;
w3244 <= not w2314 and not w2327;
w3245 <= not w2331 and not w3244;
w3246 <= not w2278 and not w2314;
w3247 <= not w2296 and w3246;
w3248 <= not w2332 and w3247;
w3249 <= not w2278 and not w2291;
w3250 <= not w2295 and not w3249;
w3251 <= not w3248 and w3250;
w3252 <= w3248 and not w3250;
w3253 <= not w3251 and not w3252;
w3254 <= not w3245 and not w3253;
w3255 <= not w3248 and not w3250;
w3256 <= not w2295 and w3246;
w3257 <= not w2296 and w3256;
w3258 <= not w2332 and not w3249;
w3259 <= w3257 and w3258;
w3260 <= not w3255 and not w3259;
w3261 <= w3245 and not w3260;
w3262 <= not w3254 and not w3261;
w3263 <= not w3243 and w3262;
w3264 <= not w3237 and not w3238;
w3265 <= not w3233 and w3264;
w3266 <= w3238 and not w3241;
w3267 <= not w3265 and not w3266;
w3268 <= not w3262 and not w3267;
w3269 <= not w3263 and not w3268;
w3270 <= not w2161 and not w2174;
w3271 <= not w2178 and not w3270;
w3272 <= not w2125 and not w2161;
w3273 <= not w2143 and w3272;
w3274 <= not w2179 and w3273;
w3275 <= not w2125 and not w2138;
w3276 <= not w2142 and not w3275;
w3277 <= not w3274 and w3276;
w3278 <= w3274 and not w3276;
w3279 <= not w3277 and not w3278;
w3280 <= not w3271 and not w3279;
w3281 <= not w3274 and not w3276;
w3282 <= not w2142 and w3272;
w3283 <= not w2143 and w3282;
w3284 <= not w2179 and not w3275;
w3285 <= w3283 and w3284;
w3286 <= not w3281 and not w3285;
w3287 <= w3271 and not w3286;
w3288 <= not w3280 and not w3287;
w3289 <= not w2086 and not w2099;
w3290 <= not w2103 and not w3289;
w3291 <= not w2050 and not w2086;
w3292 <= not w2068 and w3291;
w3293 <= not w2104 and w3292;
w3294 <= not w2050 and not w2063;
w3295 <= not w2067 and not w3294;
w3296 <= not w3293 and not w3295;
w3297 <= not w2067 and w3291;
w3298 <= not w2068 and w3297;
w3299 <= not w2104 and not w3294;
w3300 <= w3298 and w3299;
w3301 <= not w3296 and not w3300;
w3302 <= w3290 and not w3301;
w3303 <= not w3293 and w3295;
w3304 <= w3293 and not w3295;
w3305 <= not w3303 and not w3304;
w3306 <= not w3290 and not w3305;
w3307 <= not w2108 and not w2183;
w3308 <= not w3306 and not w3307;
w3309 <= not w3302 and w3308;
w3310 <= not w3302 and not w3306;
w3311 <= w3307 and not w3310;
w3312 <= not w3309 and not w3311;
w3313 <= not w3288 and not w3312;
w3314 <= not w3306 and w3307;
w3315 <= not w3302 and w3314;
w3316 <= not w3307 and not w3310;
w3317 <= not w3315 and not w3316;
w3318 <= w3288 and not w3317;
w3319 <= not w2186 and not w2339;
w3320 <= not w3318 and not w3319;
w3321 <= not w3313 and w3320;
w3322 <= not w3313 and not w3318;
w3323 <= w3319 and not w3322;
w3324 <= not w3321 and not w3323;
w3325 <= not w3269 and not w3324;
w3326 <= not w3318 and w3319;
w3327 <= not w3313 and w3326;
w3328 <= not w3319 and not w3322;
w3329 <= not w3327 and not w3328;
w3330 <= w3269 and not w3329;
w3331 <= not w2033 and not w2342;
w3332 <= not w3330 and w3331;
w3333 <= not w3325 and w3332;
w3334 <= not w3325 and not w3330;
w3335 <= not w3331 and not w3334;
w3336 <= not w3333 and not w3335;
w3337 <= not w2005 and not w2018;
w3338 <= not w2022 and not w3337;
w3339 <= not w1969 and not w2005;
w3340 <= not w1987 and w3339;
w3341 <= not w2023 and w3340;
w3342 <= not w1969 and not w1982;
w3343 <= not w1986 and not w3342;
w3344 <= not w3341 and w3343;
w3345 <= w3341 and not w3343;
w3346 <= not w3344 and not w3345;
w3347 <= not w3338 and not w3346;
w3348 <= not w3341 and not w3343;
w3349 <= not w1986 and w3339;
w3350 <= not w1987 and w3349;
w3351 <= not w2023 and not w3342;
w3352 <= w3350 and w3351;
w3353 <= not w3348 and not w3352;
w3354 <= w3338 and not w3353;
w3355 <= not w3347 and not w3354;
w3356 <= not w1930 and not w1943;
w3357 <= not w1947 and not w3356;
w3358 <= not w1894 and not w1930;
w3359 <= not w1912 and w3358;
w3360 <= not w1948 and w3359;
w3361 <= not w1894 and not w1907;
w3362 <= not w1911 and not w3361;
w3363 <= not w3360 and not w3362;
w3364 <= not w1911 and w3358;
w3365 <= not w1912 and w3364;
w3366 <= not w1948 and not w3361;
w3367 <= w3365 and w3366;
w3368 <= not w3363 and not w3367;
w3369 <= w3357 and not w3368;
w3370 <= not w3360 and w3362;
w3371 <= w3360 and not w3362;
w3372 <= not w3370 and not w3371;
w3373 <= not w3357 and not w3372;
w3374 <= not w1952 and not w2027;
w3375 <= not w3373 and not w3374;
w3376 <= not w3369 and w3375;
w3377 <= not w3369 and not w3373;
w3378 <= w3374 and not w3377;
w3379 <= not w3376 and not w3378;
w3380 <= not w3355 and not w3379;
w3381 <= not w3373 and w3374;
w3382 <= not w3369 and w3381;
w3383 <= not w3374 and not w3377;
w3384 <= not w3382 and not w3383;
w3385 <= w3355 and not w3384;
w3386 <= not w1877 and not w2030;
w3387 <= not w3385 and w3386;
w3388 <= not w3380 and w3387;
w3389 <= not w3380 and not w3385;
w3390 <= not w3386 and not w3389;
w3391 <= not w3388 and not w3390;
w3392 <= not w1852 and not w1865;
w3393 <= not w1869 and not w3392;
w3394 <= not w1816 and not w1852;
w3395 <= not w1834 and w3394;
w3396 <= not w1870 and w3395;
w3397 <= not w1816 and not w1829;
w3398 <= not w1833 and not w3397;
w3399 <= not w3396 and not w3398;
w3400 <= not w1833 and w3394;
w3401 <= not w1834 and w3400;
w3402 <= not w1870 and not w3397;
w3403 <= w3401 and w3402;
w3404 <= not w3399 and not w3403;
w3405 <= w3393 and not w3404;
w3406 <= not w3396 and w3398;
w3407 <= w3396 and not w3398;
w3408 <= not w3406 and not w3407;
w3409 <= not w3393 and not w3408;
w3410 <= not w1799 and not w1874;
w3411 <= not w3409 and w3410;
w3412 <= not w3405 and w3411;
w3413 <= not w3405 and not w3409;
w3414 <= not w3410 and not w3413;
w3415 <= not w3412 and not w3414;
w3416 <= not w1777 and not w1794;
w3417 <= not w1791 and not w3416;
w3418 <= not w1741 and not w1777;
w3419 <= not w1759 and w3418;
w3420 <= not w1795 and w3419;
w3421 <= not w1741 and not w1754;
w3422 <= not w1758 and not w3421;
w3423 <= not w3420 and w3422;
w3424 <= w3420 and not w3422;
w3425 <= not w3423 and not w3424;
w3426 <= not w3417 and not w3425;
w3427 <= not w3420 and not w3422;
w3428 <= not w1758 and w3418;
w3429 <= not w1759 and w3428;
w3430 <= not w1795 and not w3421;
w3431 <= w3429 and w3430;
w3432 <= not w3427 and not w3431;
w3433 <= w3417 and not w3432;
w3434 <= not w3426 and not w3433;
w3435 <= not w3415 and w3434;
w3436 <= not w3409 and not w3410;
w3437 <= not w3405 and w3436;
w3438 <= w3410 and not w3413;
w3439 <= not w3437 and not w3438;
w3440 <= not w3434 and not w3439;
w3441 <= not w3435 and not w3440;
w3442 <= not w3391 and w3441;
w3443 <= not w3385 and not w3386;
w3444 <= not w3380 and w3443;
w3445 <= w3386 and not w3389;
w3446 <= not w3444 and not w3445;
w3447 <= not w3441 and not w3446;
w3448 <= not w3442 and not w3447;
w3449 <= not w3336 and w3448;
w3450 <= not w3330 and not w3331;
w3451 <= not w3325 and w3450;
w3452 <= w3331 and not w3334;
w3453 <= not w3451 and not w3452;
w3454 <= not w3448 and not w3453;
w3455 <= not w3449 and not w3454;
w3456 <= not w3219 and w3455;
w3457 <= not w3213 and not w3214;
w3458 <= not w3208 and w3457;
w3459 <= w3214 and not w3217;
w3460 <= not w3458 and not w3459;
w3461 <= not w3455 and not w3460;
w3462 <= not w3456 and not w3461;
w3463 <= not w2978 and w3462;
w3464 <= not w1724 and not w2973;
w3465 <= not w1719 and w3464;
w3466 <= w2973 and not w2976;
w3467 <= not w3465 and not w3466;
w3468 <= not w3462 and not w3467;
w3469 <= not w3463 and not w3468;
w3470 <= A(970) and A(971);
w3471 <= A(970) and not A(971);
w3472 <= not A(970) and A(971);
w3473 <= not w3471 and not w3472;
w3474 <= A(972) and not w3473;
w3475 <= not w3470 and not w3474;
w3476 <= A(967) and A(968);
w3477 <= A(967) and not A(968);
w3478 <= not A(967) and A(968);
w3479 <= not w3477 and not w3478;
w3480 <= A(969) and not w3479;
w3481 <= not w3476 and not w3480;
w3482 <= w3475 and not w3481;
w3483 <= not w3475 and w3481;
w3484 <= A(969) and not w3477;
w3485 <= not w3478 and w3484;
w3486 <= not A(969) and not w3479;
w3487 <= not w3485 and not w3486;
w3488 <= A(972) and not w3471;
w3489 <= not w3472 and w3488;
w3490 <= not A(972) and not w3473;
w3491 <= not w3489 and not w3490;
w3492 <= not w3487 and not w3491;
w3493 <= not w3483 and w3492;
w3494 <= not w3482 and w3493;
w3495 <= not w3482 and not w3483;
w3496 <= not w3492 and not w3495;
w3497 <= not w3494 and not w3496;
w3498 <= not w3487 and w3491;
w3499 <= w3487 and not w3491;
w3500 <= not w3498 and not w3499;
w3501 <= w3492 and not w3495;
w3502 <= not w3475 and not w3481;
w3503 <= not w3501 and not w3502;
w3504 <= not w3500 and not w3503;
w3505 <= not w3497 and not w3504;
w3506 <= not w3497 and not w3503;
w3507 <= A(976) and A(977);
w3508 <= A(976) and not A(977);
w3509 <= not A(976) and A(977);
w3510 <= not w3508 and not w3509;
w3511 <= A(978) and not w3510;
w3512 <= not w3507 and not w3511;
w3513 <= A(973) and A(974);
w3514 <= A(973) and not A(974);
w3515 <= not A(973) and A(974);
w3516 <= not w3514 and not w3515;
w3517 <= A(975) and not w3516;
w3518 <= not w3513 and not w3517;
w3519 <= not w3512 and w3518;
w3520 <= w3512 and not w3518;
w3521 <= not w3519 and not w3520;
w3522 <= A(975) and not w3514;
w3523 <= not w3515 and w3522;
w3524 <= not A(975) and not w3516;
w3525 <= not w3523 and not w3524;
w3526 <= A(978) and not w3508;
w3527 <= not w3509 and w3526;
w3528 <= not A(978) and not w3510;
w3529 <= not w3527 and not w3528;
w3530 <= not w3525 and not w3529;
w3531 <= not w3521 and w3530;
w3532 <= not w3512 and not w3518;
w3533 <= not w3531 and not w3532;
w3534 <= not w3519 and w3530;
w3535 <= not w3520 and w3534;
w3536 <= not w3521 and not w3530;
w3537 <= not w3535 and not w3536;
w3538 <= not w3533 and not w3537;
w3539 <= not w3525 and w3529;
w3540 <= w3525 and not w3529;
w3541 <= not w3539 and not w3540;
w3542 <= not w3500 and not w3541;
w3543 <= not w3538 and w3542;
w3544 <= not w3506 and w3543;
w3545 <= not w3533 and not w3541;
w3546 <= not w3537 and not w3545;
w3547 <= not w3544 and w3546;
w3548 <= w3544 and not w3546;
w3549 <= not w3547 and not w3548;
w3550 <= not w3505 and not w3549;
w3551 <= not w3544 and not w3546;
w3552 <= not w3537 and w3542;
w3553 <= not w3538 and w3552;
w3554 <= not w3506 and not w3545;
w3555 <= w3553 and w3554;
w3556 <= not w3551 and not w3555;
w3557 <= w3505 and not w3556;
w3558 <= not w3550 and not w3557;
w3559 <= A(982) and A(983);
w3560 <= A(982) and not A(983);
w3561 <= not A(982) and A(983);
w3562 <= not w3560 and not w3561;
w3563 <= A(984) and not w3562;
w3564 <= not w3559 and not w3563;
w3565 <= A(979) and A(980);
w3566 <= A(979) and not A(980);
w3567 <= not A(979) and A(980);
w3568 <= not w3566 and not w3567;
w3569 <= A(981) and not w3568;
w3570 <= not w3565 and not w3569;
w3571 <= w3564 and not w3570;
w3572 <= not w3564 and w3570;
w3573 <= A(981) and not w3566;
w3574 <= not w3567 and w3573;
w3575 <= not A(981) and not w3568;
w3576 <= not w3574 and not w3575;
w3577 <= A(984) and not w3560;
w3578 <= not w3561 and w3577;
w3579 <= not A(984) and not w3562;
w3580 <= not w3578 and not w3579;
w3581 <= not w3576 and not w3580;
w3582 <= not w3572 and w3581;
w3583 <= not w3571 and w3582;
w3584 <= not w3571 and not w3572;
w3585 <= not w3581 and not w3584;
w3586 <= not w3583 and not w3585;
w3587 <= not w3576 and w3580;
w3588 <= w3576 and not w3580;
w3589 <= not w3587 and not w3588;
w3590 <= w3581 and not w3584;
w3591 <= not w3564 and not w3570;
w3592 <= not w3590 and not w3591;
w3593 <= not w3589 and not w3592;
w3594 <= not w3586 and not w3593;
w3595 <= not w3586 and not w3592;
w3596 <= A(988) and A(989);
w3597 <= A(988) and not A(989);
w3598 <= not A(988) and A(989);
w3599 <= not w3597 and not w3598;
w3600 <= A(990) and not w3599;
w3601 <= not w3596 and not w3600;
w3602 <= A(985) and A(986);
w3603 <= A(985) and not A(986);
w3604 <= not A(985) and A(986);
w3605 <= not w3603 and not w3604;
w3606 <= A(987) and not w3605;
w3607 <= not w3602 and not w3606;
w3608 <= not w3601 and w3607;
w3609 <= w3601 and not w3607;
w3610 <= not w3608 and not w3609;
w3611 <= A(987) and not w3603;
w3612 <= not w3604 and w3611;
w3613 <= not A(987) and not w3605;
w3614 <= not w3612 and not w3613;
w3615 <= A(990) and not w3597;
w3616 <= not w3598 and w3615;
w3617 <= not A(990) and not w3599;
w3618 <= not w3616 and not w3617;
w3619 <= not w3614 and not w3618;
w3620 <= not w3610 and w3619;
w3621 <= not w3601 and not w3607;
w3622 <= not w3620 and not w3621;
w3623 <= not w3608 and w3619;
w3624 <= not w3609 and w3623;
w3625 <= not w3610 and not w3619;
w3626 <= not w3624 and not w3625;
w3627 <= not w3622 and not w3626;
w3628 <= not w3614 and w3618;
w3629 <= w3614 and not w3618;
w3630 <= not w3628 and not w3629;
w3631 <= not w3589 and not w3630;
w3632 <= not w3627 and w3631;
w3633 <= not w3595 and w3632;
w3634 <= not w3622 and not w3630;
w3635 <= not w3626 and not w3634;
w3636 <= not w3633 and not w3635;
w3637 <= not w3626 and w3631;
w3638 <= not w3627 and w3637;
w3639 <= not w3595 and not w3634;
w3640 <= w3638 and w3639;
w3641 <= not w3636 and not w3640;
w3642 <= w3594 and not w3641;
w3643 <= not w3633 and w3635;
w3644 <= w3633 and not w3635;
w3645 <= not w3643 and not w3644;
w3646 <= not w3594 and not w3645;
w3647 <= not w3627 and not w3630;
w3648 <= not w3589 and not w3595;
w3649 <= not w3647 and w3648;
w3650 <= w3647 and not w3648;
w3651 <= not w3649 and not w3650;
w3652 <= not w3538 and not w3541;
w3653 <= not w3500 and not w3506;
w3654 <= not w3652 and w3653;
w3655 <= w3652 and not w3653;
w3656 <= not w3654 and not w3655;
w3657 <= not w3651 and not w3656;
w3658 <= not w3646 and not w3657;
w3659 <= not w3642 and w3658;
w3660 <= not w3642 and not w3646;
w3661 <= w3657 and not w3660;
w3662 <= not w3659 and not w3661;
w3663 <= not w3558 and not w3662;
w3664 <= not w3646 and w3657;
w3665 <= not w3642 and w3664;
w3666 <= not w3657 and not w3660;
w3667 <= not w3665 and not w3666;
w3668 <= w3558 and not w3667;
w3669 <= not w3651 and w3656;
w3670 <= w3651 and not w3656;
w3671 <= not w3669 and not w3670;
w3672 <= not A(961) and A(962);
w3673 <= A(961) and not A(962);
w3674 <= A(963) and not w3673;
w3675 <= not w3672 and w3674;
w3676 <= not w3672 and not w3673;
w3677 <= not A(963) and not w3676;
w3678 <= not w3675 and not w3677;
w3679 <= not A(964) and A(965);
w3680 <= A(964) and not A(965);
w3681 <= A(966) and not w3680;
w3682 <= not w3679 and w3681;
w3683 <= not w3679 and not w3680;
w3684 <= not A(966) and not w3683;
w3685 <= not w3682 and not w3684;
w3686 <= not w3678 and w3685;
w3687 <= w3678 and not w3685;
w3688 <= not w3686 and not w3687;
w3689 <= A(964) and A(965);
w3690 <= A(966) and not w3683;
w3691 <= not w3689 and not w3690;
w3692 <= A(961) and A(962);
w3693 <= A(963) and not w3676;
w3694 <= not w3692 and not w3693;
w3695 <= not w3691 and w3694;
w3696 <= w3691 and not w3694;
w3697 <= not w3695 and not w3696;
w3698 <= not w3678 and not w3685;
w3699 <= not w3697 and w3698;
w3700 <= not w3691 and not w3694;
w3701 <= not w3699 and not w3700;
w3702 <= not w3695 and w3698;
w3703 <= not w3696 and w3702;
w3704 <= not w3697 and not w3698;
w3705 <= not w3703 and not w3704;
w3706 <= not w3701 and not w3705;
w3707 <= not w3688 and not w3706;
w3708 <= not A(955) and A(956);
w3709 <= A(955) and not A(956);
w3710 <= A(957) and not w3709;
w3711 <= not w3708 and w3710;
w3712 <= not w3708 and not w3709;
w3713 <= not A(957) and not w3712;
w3714 <= not w3711 and not w3713;
w3715 <= not A(958) and A(959);
w3716 <= A(958) and not A(959);
w3717 <= A(960) and not w3716;
w3718 <= not w3715 and w3717;
w3719 <= not w3715 and not w3716;
w3720 <= not A(960) and not w3719;
w3721 <= not w3718 and not w3720;
w3722 <= not w3714 and w3721;
w3723 <= w3714 and not w3721;
w3724 <= not w3722 and not w3723;
w3725 <= A(958) and A(959);
w3726 <= A(960) and not w3719;
w3727 <= not w3725 and not w3726;
w3728 <= A(955) and A(956);
w3729 <= A(957) and not w3712;
w3730 <= not w3728 and not w3729;
w3731 <= not w3727 and w3730;
w3732 <= w3727 and not w3730;
w3733 <= not w3731 and not w3732;
w3734 <= not w3714 and not w3721;
w3735 <= not w3733 and w3734;
w3736 <= not w3727 and not w3730;
w3737 <= not w3735 and not w3736;
w3738 <= not w3731 and w3734;
w3739 <= not w3732 and w3738;
w3740 <= not w3733 and not w3734;
w3741 <= not w3739 and not w3740;
w3742 <= not w3737 and not w3741;
w3743 <= not w3724 and not w3742;
w3744 <= not w3707 and w3743;
w3745 <= w3707 and not w3743;
w3746 <= not w3744 and not w3745;
w3747 <= not A(949) and A(950);
w3748 <= A(949) and not A(950);
w3749 <= A(951) and not w3748;
w3750 <= not w3747 and w3749;
w3751 <= not w3747 and not w3748;
w3752 <= not A(951) and not w3751;
w3753 <= not w3750 and not w3752;
w3754 <= not A(952) and A(953);
w3755 <= A(952) and not A(953);
w3756 <= A(954) and not w3755;
w3757 <= not w3754 and w3756;
w3758 <= not w3754 and not w3755;
w3759 <= not A(954) and not w3758;
w3760 <= not w3757 and not w3759;
w3761 <= not w3753 and w3760;
w3762 <= w3753 and not w3760;
w3763 <= not w3761 and not w3762;
w3764 <= A(952) and A(953);
w3765 <= A(954) and not w3758;
w3766 <= not w3764 and not w3765;
w3767 <= A(949) and A(950);
w3768 <= A(951) and not w3751;
w3769 <= not w3767 and not w3768;
w3770 <= not w3766 and w3769;
w3771 <= w3766 and not w3769;
w3772 <= not w3770 and not w3771;
w3773 <= not w3753 and not w3760;
w3774 <= not w3772 and w3773;
w3775 <= not w3766 and not w3769;
w3776 <= not w3774 and not w3775;
w3777 <= not w3770 and w3773;
w3778 <= not w3771 and w3777;
w3779 <= not w3772 and not w3773;
w3780 <= not w3778 and not w3779;
w3781 <= not w3776 and not w3780;
w3782 <= not w3763 and not w3781;
w3783 <= not A(943) and A(944);
w3784 <= A(943) and not A(944);
w3785 <= A(945) and not w3784;
w3786 <= not w3783 and w3785;
w3787 <= not w3783 and not w3784;
w3788 <= not A(945) and not w3787;
w3789 <= not w3786 and not w3788;
w3790 <= not A(946) and A(947);
w3791 <= A(946) and not A(947);
w3792 <= A(948) and not w3791;
w3793 <= not w3790 and w3792;
w3794 <= not w3790 and not w3791;
w3795 <= not A(948) and not w3794;
w3796 <= not w3793 and not w3795;
w3797 <= not w3789 and w3796;
w3798 <= w3789 and not w3796;
w3799 <= not w3797 and not w3798;
w3800 <= A(946) and A(947);
w3801 <= A(948) and not w3794;
w3802 <= not w3800 and not w3801;
w3803 <= A(943) and A(944);
w3804 <= A(945) and not w3787;
w3805 <= not w3803 and not w3804;
w3806 <= not w3802 and w3805;
w3807 <= w3802 and not w3805;
w3808 <= not w3806 and not w3807;
w3809 <= not w3789 and not w3796;
w3810 <= not w3808 and w3809;
w3811 <= not w3802 and not w3805;
w3812 <= not w3810 and not w3811;
w3813 <= not w3806 and w3809;
w3814 <= not w3807 and w3813;
w3815 <= not w3808 and not w3809;
w3816 <= not w3814 and not w3815;
w3817 <= not w3812 and not w3816;
w3818 <= not w3799 and not w3817;
w3819 <= not w3782 and w3818;
w3820 <= w3782 and not w3818;
w3821 <= not w3819 and not w3820;
w3822 <= not w3746 and w3821;
w3823 <= w3746 and not w3821;
w3824 <= not w3822 and not w3823;
w3825 <= not w3671 and not w3824;
w3826 <= not w3668 and w3825;
w3827 <= not w3663 and w3826;
w3828 <= not w3663 and not w3668;
w3829 <= not w3825 and not w3828;
w3830 <= not w3827 and not w3829;
w3831 <= not w3724 and not w3737;
w3832 <= not w3741 and not w3831;
w3833 <= not w3688 and not w3724;
w3834 <= not w3706 and w3833;
w3835 <= not w3742 and w3834;
w3836 <= not w3688 and not w3701;
w3837 <= not w3705 and not w3836;
w3838 <= not w3835 and not w3837;
w3839 <= not w3705 and w3833;
w3840 <= not w3706 and w3839;
w3841 <= not w3742 and not w3836;
w3842 <= w3840 and w3841;
w3843 <= not w3838 and not w3842;
w3844 <= w3832 and not w3843;
w3845 <= not w3835 and w3837;
w3846 <= w3835 and not w3837;
w3847 <= not w3845 and not w3846;
w3848 <= not w3832 and not w3847;
w3849 <= not w3746 and not w3821;
w3850 <= not w3848 and w3849;
w3851 <= not w3844 and w3850;
w3852 <= not w3844 and not w3848;
w3853 <= not w3849 and not w3852;
w3854 <= not w3851 and not w3853;
w3855 <= not w3799 and not w3812;
w3856 <= not w3816 and not w3855;
w3857 <= not w3763 and not w3799;
w3858 <= not w3781 and w3857;
w3859 <= not w3817 and w3858;
w3860 <= not w3763 and not w3776;
w3861 <= not w3780 and not w3860;
w3862 <= not w3859 and w3861;
w3863 <= w3859 and not w3861;
w3864 <= not w3862 and not w3863;
w3865 <= not w3856 and not w3864;
w3866 <= not w3859 and not w3861;
w3867 <= not w3780 and w3857;
w3868 <= not w3781 and w3867;
w3869 <= not w3817 and not w3860;
w3870 <= w3868 and w3869;
w3871 <= not w3866 and not w3870;
w3872 <= w3856 and not w3871;
w3873 <= not w3865 and not w3872;
w3874 <= not w3854 and w3873;
w3875 <= not w3848 and not w3849;
w3876 <= not w3844 and w3875;
w3877 <= w3849 and not w3852;
w3878 <= not w3876 and not w3877;
w3879 <= not w3873 and not w3878;
w3880 <= not w3874 and not w3879;
w3881 <= not w3830 and w3880;
w3882 <= not w3668 and not w3825;
w3883 <= not w3663 and w3882;
w3884 <= w3825 and not w3828;
w3885 <= not w3883 and not w3884;
w3886 <= not w3880 and not w3885;
w3887 <= not w3881 and not w3886;
w3888 <= A(10) and A(11);
w3889 <= A(10) and not A(11);
w3890 <= not A(10) and A(11);
w3891 <= not w3889 and not w3890;
w3892 <= A(12) and not w3891;
w3893 <= not w3888 and not w3892;
w3894 <= A(7) and A(8);
w3895 <= A(7) and not A(8);
w3896 <= not A(7) and A(8);
w3897 <= not w3895 and not w3896;
w3898 <= A(9) and not w3897;
w3899 <= not w3894 and not w3898;
w3900 <= w3893 and not w3899;
w3901 <= not w3893 and w3899;
w3902 <= A(9) and not w3895;
w3903 <= not w3896 and w3902;
w3904 <= not A(9) and not w3897;
w3905 <= not w3903 and not w3904;
w3906 <= A(12) and not w3889;
w3907 <= not w3890 and w3906;
w3908 <= not A(12) and not w3891;
w3909 <= not w3907 and not w3908;
w3910 <= not w3905 and not w3909;
w3911 <= not w3901 and w3910;
w3912 <= not w3900 and w3911;
w3913 <= not w3900 and not w3901;
w3914 <= not w3910 and not w3913;
w3915 <= not w3912 and not w3914;
w3916 <= not w3905 and w3909;
w3917 <= w3905 and not w3909;
w3918 <= not w3916 and not w3917;
w3919 <= w3910 and not w3913;
w3920 <= not w3893 and not w3899;
w3921 <= not w3919 and not w3920;
w3922 <= not w3918 and not w3921;
w3923 <= not w3915 and not w3922;
w3924 <= not w3915 and not w3921;
w3925 <= A(16) and A(17);
w3926 <= A(16) and not A(17);
w3927 <= not A(16) and A(17);
w3928 <= not w3926 and not w3927;
w3929 <= A(18) and not w3928;
w3930 <= not w3925 and not w3929;
w3931 <= A(13) and A(14);
w3932 <= A(13) and not A(14);
w3933 <= not A(13) and A(14);
w3934 <= not w3932 and not w3933;
w3935 <= A(15) and not w3934;
w3936 <= not w3931 and not w3935;
w3937 <= not w3930 and w3936;
w3938 <= w3930 and not w3936;
w3939 <= not w3937 and not w3938;
w3940 <= A(15) and not w3932;
w3941 <= not w3933 and w3940;
w3942 <= not A(15) and not w3934;
w3943 <= not w3941 and not w3942;
w3944 <= A(18) and not w3926;
w3945 <= not w3927 and w3944;
w3946 <= not A(18) and not w3928;
w3947 <= not w3945 and not w3946;
w3948 <= not w3943 and not w3947;
w3949 <= not w3939 and w3948;
w3950 <= not w3930 and not w3936;
w3951 <= not w3949 and not w3950;
w3952 <= not w3937 and w3948;
w3953 <= not w3938 and w3952;
w3954 <= not w3939 and not w3948;
w3955 <= not w3953 and not w3954;
w3956 <= not w3951 and not w3955;
w3957 <= not w3943 and w3947;
w3958 <= w3943 and not w3947;
w3959 <= not w3957 and not w3958;
w3960 <= not w3918 and not w3959;
w3961 <= not w3956 and w3960;
w3962 <= not w3924 and w3961;
w3963 <= not w3951 and not w3959;
w3964 <= not w3955 and not w3963;
w3965 <= not w3962 and w3964;
w3966 <= w3962 and not w3964;
w3967 <= not w3965 and not w3966;
w3968 <= not w3923 and not w3967;
w3969 <= not w3962 and not w3964;
w3970 <= not w3955 and w3960;
w3971 <= not w3956 and w3970;
w3972 <= not w3924 and not w3963;
w3973 <= w3971 and w3972;
w3974 <= not w3969 and not w3973;
w3975 <= w3923 and not w3974;
w3976 <= not w3968 and not w3975;
w3977 <= A(22) and A(23);
w3978 <= A(22) and not A(23);
w3979 <= not A(22) and A(23);
w3980 <= not w3978 and not w3979;
w3981 <= A(24) and not w3980;
w3982 <= not w3977 and not w3981;
w3983 <= A(19) and A(20);
w3984 <= A(19) and not A(20);
w3985 <= not A(19) and A(20);
w3986 <= not w3984 and not w3985;
w3987 <= A(21) and not w3986;
w3988 <= not w3983 and not w3987;
w3989 <= w3982 and not w3988;
w3990 <= not w3982 and w3988;
w3991 <= A(21) and not w3984;
w3992 <= not w3985 and w3991;
w3993 <= not A(21) and not w3986;
w3994 <= not w3992 and not w3993;
w3995 <= A(24) and not w3978;
w3996 <= not w3979 and w3995;
w3997 <= not A(24) and not w3980;
w3998 <= not w3996 and not w3997;
w3999 <= not w3994 and not w3998;
w4000 <= not w3990 and w3999;
w4001 <= not w3989 and w4000;
w4002 <= not w3989 and not w3990;
w4003 <= not w3999 and not w4002;
w4004 <= not w4001 and not w4003;
w4005 <= not w3994 and w3998;
w4006 <= w3994 and not w3998;
w4007 <= not w4005 and not w4006;
w4008 <= w3999 and not w4002;
w4009 <= not w3982 and not w3988;
w4010 <= not w4008 and not w4009;
w4011 <= not w4007 and not w4010;
w4012 <= not w4004 and not w4011;
w4013 <= not w4004 and not w4010;
w4014 <= A(28) and A(29);
w4015 <= A(28) and not A(29);
w4016 <= not A(28) and A(29);
w4017 <= not w4015 and not w4016;
w4018 <= A(30) and not w4017;
w4019 <= not w4014 and not w4018;
w4020 <= A(25) and A(26);
w4021 <= A(25) and not A(26);
w4022 <= not A(25) and A(26);
w4023 <= not w4021 and not w4022;
w4024 <= A(27) and not w4023;
w4025 <= not w4020 and not w4024;
w4026 <= not w4019 and w4025;
w4027 <= w4019 and not w4025;
w4028 <= not w4026 and not w4027;
w4029 <= A(27) and not w4021;
w4030 <= not w4022 and w4029;
w4031 <= not A(27) and not w4023;
w4032 <= not w4030 and not w4031;
w4033 <= A(30) and not w4015;
w4034 <= not w4016 and w4033;
w4035 <= not A(30) and not w4017;
w4036 <= not w4034 and not w4035;
w4037 <= not w4032 and not w4036;
w4038 <= not w4028 and w4037;
w4039 <= not w4019 and not w4025;
w4040 <= not w4038 and not w4039;
w4041 <= not w4026 and w4037;
w4042 <= not w4027 and w4041;
w4043 <= not w4028 and not w4037;
w4044 <= not w4042 and not w4043;
w4045 <= not w4040 and not w4044;
w4046 <= not w4032 and w4036;
w4047 <= w4032 and not w4036;
w4048 <= not w4046 and not w4047;
w4049 <= not w4007 and not w4048;
w4050 <= not w4045 and w4049;
w4051 <= not w4013 and w4050;
w4052 <= not w4040 and not w4048;
w4053 <= not w4044 and not w4052;
w4054 <= not w4051 and not w4053;
w4055 <= not w4044 and w4049;
w4056 <= not w4045 and w4055;
w4057 <= not w4013 and not w4052;
w4058 <= w4056 and w4057;
w4059 <= not w4054 and not w4058;
w4060 <= w4012 and not w4059;
w4061 <= not w4051 and w4053;
w4062 <= w4051 and not w4053;
w4063 <= not w4061 and not w4062;
w4064 <= not w4012 and not w4063;
w4065 <= not w4045 and not w4048;
w4066 <= not w4007 and not w4013;
w4067 <= not w4065 and w4066;
w4068 <= w4065 and not w4066;
w4069 <= not w4067 and not w4068;
w4070 <= not w3956 and not w3959;
w4071 <= not w3918 and not w3924;
w4072 <= not w4070 and w4071;
w4073 <= w4070 and not w4071;
w4074 <= not w4072 and not w4073;
w4075 <= not w4069 and not w4074;
w4076 <= not w4064 and not w4075;
w4077 <= not w4060 and w4076;
w4078 <= not w4060 and not w4064;
w4079 <= w4075 and not w4078;
w4080 <= not w4077 and not w4079;
w4081 <= not w3976 and not w4080;
w4082 <= not w4064 and w4075;
w4083 <= not w4060 and w4082;
w4084 <= not w4075 and not w4078;
w4085 <= not w4083 and not w4084;
w4086 <= w3976 and not w4085;
w4087 <= not w4069 and w4074;
w4088 <= w4069 and not w4074;
w4089 <= not w4087 and not w4088;
w4090 <= not A(991) and A(992);
w4091 <= A(991) and not A(992);
w4092 <= A(993) and not w4091;
w4093 <= not w4090 and w4092;
w4094 <= not w4090 and not w4091;
w4095 <= not A(993) and not w4094;
w4096 <= not w4093 and not w4095;
w4097 <= not A(994) and A(995);
w4098 <= A(994) and not A(995);
w4099 <= A(996) and not w4098;
w4100 <= not w4097 and w4099;
w4101 <= not w4097 and not w4098;
w4102 <= not A(996) and not w4101;
w4103 <= not w4100 and not w4102;
w4104 <= not w4096 and w4103;
w4105 <= w4096 and not w4103;
w4106 <= not w4104 and not w4105;
w4107 <= A(994) and A(995);
w4108 <= A(996) and not w4101;
w4109 <= not w4107 and not w4108;
w4110 <= A(991) and A(992);
w4111 <= A(993) and not w4094;
w4112 <= not w4110 and not w4111;
w4113 <= not w4109 and w4112;
w4114 <= w4109 and not w4112;
w4115 <= not w4113 and not w4114;
w4116 <= not w4096 and not w4103;
w4117 <= not w4115 and w4116;
w4118 <= not w4109 and not w4112;
w4119 <= not w4117 and not w4118;
w4120 <= not w4113 and w4116;
w4121 <= not w4114 and w4120;
w4122 <= not w4115 and not w4116;
w4123 <= not w4121 and not w4122;
w4124 <= not w4119 and not w4123;
w4125 <= not w4106 and not w4124;
w4126 <= A(3) and not A(4);
w4127 <= not A(3) and A(4);
w4128 <= A(5) and not w4127;
w4129 <= not w4126 and w4128;
w4130 <= not w4126 and not w4127;
w4131 <= not A(5) and not w4130;
w4132 <= not w4129 and not w4131;
w4133 <= not A(0) and A(1);
w4134 <= A(0) and not A(1);
w4135 <= not w4133 and not w4134;
w4136 <= not A(2) and not w4135;
w4137 <= A(2) and not w4133;
w4138 <= not w4134 and w4137;
w4139 <= A(6) and not w4138;
w4140 <= not w4136 and w4139;
w4141 <= not w4136 and not w4138;
w4142 <= not A(6) and not w4141;
w4143 <= not w4140 and not w4142;
w4144 <= w4132 and not w4143;
w4145 <= not w4132 and not w4140;
w4146 <= not w4142 and w4145;
w4147 <= not A(997) and A(998);
w4148 <= A(997) and not A(998);
w4149 <= A(999) and not w4148;
w4150 <= not w4147 and w4149;
w4151 <= not w4147 and not w4148;
w4152 <= not A(999) and not w4151;
w4153 <= not w4150 and not w4152;
w4154 <= not w4146 and not w4153;
w4155 <= not w4144 and w4154;
w4156 <= not w4144 and not w4146;
w4157 <= w4153 and not w4156;
w4158 <= not w4155 and not w4157;
w4159 <= w4125 and w4158;
w4160 <= not w4125 and not w4158;
w4161 <= not w4159 and not w4160;
w4162 <= not w4089 and not w4161;
w4163 <= not w4086 and w4162;
w4164 <= not w4081 and w4163;
w4165 <= not w4081 and not w4086;
w4166 <= not w4162 and not w4165;
w4167 <= not w4164 and not w4166;
w4168 <= not w4106 and not w4119;
w4169 <= not w4123 and not w4168;
w4170 <= not w4132 and not w4143;
w4171 <= A(6) and not w4141;
w4172 <= A(3) and A(4);
w4173 <= A(5) and not w4130;
w4174 <= not w4172 and not w4173;
w4175 <= A(0) and A(1);
w4176 <= A(2) and not w4135;
w4177 <= not w4175 and not w4176;
w4178 <= not w4174 and w4177;
w4179 <= w4174 and not w4177;
w4180 <= not w4178 and not w4179;
w4181 <= not w4171 and w4180;
w4182 <= not w4170 and w4181;
w4183 <= not w4170 and not w4171;
w4184 <= not w4180 and not w4183;
w4185 <= not w4182 and not w4184;
w4186 <= not w4153 and not w4156;
w4187 <= w4185 and w4186;
w4188 <= A(997) and A(998);
w4189 <= A(999) and not w4151;
w4190 <= not w4188 and not w4189;
w4191 <= not w4185 and not w4186;
w4192 <= w4190 and not w4191;
w4193 <= not w4187 and w4192;
w4194 <= not w4187 and not w4191;
w4195 <= not w4190 and not w4194;
w4196 <= w4125 and not w4158;
w4197 <= not w4195 and w4196;
w4198 <= not w4193 and w4197;
w4199 <= not w4193 and not w4195;
w4200 <= not w4196 and not w4199;
w4201 <= not w4198 and not w4200;
w4202 <= not w4169 and not w4201;
w4203 <= not w4195 and not w4196;
w4204 <= not w4193 and w4203;
w4205 <= w4196 and not w4199;
w4206 <= not w4204 and not w4205;
w4207 <= w4169 and not w4206;
w4208 <= not w4202 and not w4207;
w4209 <= not w4167 and w4208;
w4210 <= not w4086 and not w4162;
w4211 <= not w4081 and w4210;
w4212 <= w4162 and not w4165;
w4213 <= not w4211 and not w4212;
w4214 <= not w4208 and not w4213;
w4215 <= not w4209 and not w4214;
w4216 <= A(46) and A(47);
w4217 <= A(46) and not A(47);
w4218 <= not A(46) and A(47);
w4219 <= not w4217 and not w4218;
w4220 <= A(48) and not w4219;
w4221 <= not w4216 and not w4220;
w4222 <= A(43) and A(44);
w4223 <= A(43) and not A(44);
w4224 <= not A(43) and A(44);
w4225 <= not w4223 and not w4224;
w4226 <= A(45) and not w4225;
w4227 <= not w4222 and not w4226;
w4228 <= w4221 and not w4227;
w4229 <= not w4221 and w4227;
w4230 <= A(45) and not w4223;
w4231 <= not w4224 and w4230;
w4232 <= not A(45) and not w4225;
w4233 <= not w4231 and not w4232;
w4234 <= A(48) and not w4217;
w4235 <= not w4218 and w4234;
w4236 <= not A(48) and not w4219;
w4237 <= not w4235 and not w4236;
w4238 <= not w4233 and not w4237;
w4239 <= not w4229 and w4238;
w4240 <= not w4228 and w4239;
w4241 <= not w4228 and not w4229;
w4242 <= not w4238 and not w4241;
w4243 <= not w4240 and not w4242;
w4244 <= not w4233 and w4237;
w4245 <= w4233 and not w4237;
w4246 <= not w4244 and not w4245;
w4247 <= w4238 and not w4241;
w4248 <= not w4221 and not w4227;
w4249 <= not w4247 and not w4248;
w4250 <= not w4246 and not w4249;
w4251 <= not w4243 and not w4250;
w4252 <= not w4243 and not w4249;
w4253 <= A(52) and A(53);
w4254 <= A(52) and not A(53);
w4255 <= not A(52) and A(53);
w4256 <= not w4254 and not w4255;
w4257 <= A(54) and not w4256;
w4258 <= not w4253 and not w4257;
w4259 <= A(49) and A(50);
w4260 <= A(49) and not A(50);
w4261 <= not A(49) and A(50);
w4262 <= not w4260 and not w4261;
w4263 <= A(51) and not w4262;
w4264 <= not w4259 and not w4263;
w4265 <= not w4258 and w4264;
w4266 <= w4258 and not w4264;
w4267 <= not w4265 and not w4266;
w4268 <= A(51) and not w4260;
w4269 <= not w4261 and w4268;
w4270 <= not A(51) and not w4262;
w4271 <= not w4269 and not w4270;
w4272 <= A(54) and not w4254;
w4273 <= not w4255 and w4272;
w4274 <= not A(54) and not w4256;
w4275 <= not w4273 and not w4274;
w4276 <= not w4271 and not w4275;
w4277 <= not w4267 and w4276;
w4278 <= not w4258 and not w4264;
w4279 <= not w4277 and not w4278;
w4280 <= not w4265 and w4276;
w4281 <= not w4266 and w4280;
w4282 <= not w4267 and not w4276;
w4283 <= not w4281 and not w4282;
w4284 <= not w4279 and not w4283;
w4285 <= not w4271 and w4275;
w4286 <= w4271 and not w4275;
w4287 <= not w4285 and not w4286;
w4288 <= not w4246 and not w4287;
w4289 <= not w4284 and w4288;
w4290 <= not w4252 and w4289;
w4291 <= not w4279 and not w4287;
w4292 <= not w4283 and not w4291;
w4293 <= not w4290 and not w4292;
w4294 <= not w4283 and w4288;
w4295 <= not w4284 and w4294;
w4296 <= not w4252 and not w4291;
w4297 <= w4295 and w4296;
w4298 <= not w4293 and not w4297;
w4299 <= w4251 and not w4298;
w4300 <= not w4290 and w4292;
w4301 <= w4290 and not w4292;
w4302 <= not w4300 and not w4301;
w4303 <= not w4251 and not w4302;
w4304 <= not w4284 and not w4287;
w4305 <= not w4246 and not w4252;
w4306 <= not w4304 and w4305;
w4307 <= w4304 and not w4305;
w4308 <= not w4306 and not w4307;
w4309 <= not A(37) and A(38);
w4310 <= A(37) and not A(38);
w4311 <= A(39) and not w4310;
w4312 <= not w4309 and w4311;
w4313 <= not w4309 and not w4310;
w4314 <= not A(39) and not w4313;
w4315 <= not w4312 and not w4314;
w4316 <= not A(40) and A(41);
w4317 <= A(40) and not A(41);
w4318 <= A(42) and not w4317;
w4319 <= not w4316 and w4318;
w4320 <= not w4316 and not w4317;
w4321 <= not A(42) and not w4320;
w4322 <= not w4319 and not w4321;
w4323 <= not w4315 and w4322;
w4324 <= w4315 and not w4322;
w4325 <= not w4323 and not w4324;
w4326 <= A(40) and A(41);
w4327 <= A(42) and not w4320;
w4328 <= not w4326 and not w4327;
w4329 <= A(37) and A(38);
w4330 <= A(39) and not w4313;
w4331 <= not w4329 and not w4330;
w4332 <= not w4328 and w4331;
w4333 <= w4328 and not w4331;
w4334 <= not w4332 and not w4333;
w4335 <= not w4315 and not w4322;
w4336 <= not w4334 and w4335;
w4337 <= not w4328 and not w4331;
w4338 <= not w4336 and not w4337;
w4339 <= not w4332 and w4335;
w4340 <= not w4333 and w4339;
w4341 <= not w4334 and not w4335;
w4342 <= not w4340 and not w4341;
w4343 <= not w4338 and not w4342;
w4344 <= not w4325 and not w4343;
w4345 <= not A(31) and A(32);
w4346 <= A(31) and not A(32);
w4347 <= A(33) and not w4346;
w4348 <= not w4345 and w4347;
w4349 <= not w4345 and not w4346;
w4350 <= not A(33) and not w4349;
w4351 <= not w4348 and not w4350;
w4352 <= not A(34) and A(35);
w4353 <= A(34) and not A(35);
w4354 <= A(36) and not w4353;
w4355 <= not w4352 and w4354;
w4356 <= not w4352 and not w4353;
w4357 <= not A(36) and not w4356;
w4358 <= not w4355 and not w4357;
w4359 <= not w4351 and w4358;
w4360 <= w4351 and not w4358;
w4361 <= not w4359 and not w4360;
w4362 <= A(34) and A(35);
w4363 <= A(36) and not w4356;
w4364 <= not w4362 and not w4363;
w4365 <= A(31) and A(32);
w4366 <= A(33) and not w4349;
w4367 <= not w4365 and not w4366;
w4368 <= not w4364 and w4367;
w4369 <= w4364 and not w4367;
w4370 <= not w4368 and not w4369;
w4371 <= not w4351 and not w4358;
w4372 <= not w4370 and w4371;
w4373 <= not w4364 and not w4367;
w4374 <= not w4372 and not w4373;
w4375 <= not w4368 and w4371;
w4376 <= not w4369 and w4375;
w4377 <= not w4370 and not w4371;
w4378 <= not w4376 and not w4377;
w4379 <= not w4374 and not w4378;
w4380 <= not w4361 and not w4379;
w4381 <= not w4344 and w4380;
w4382 <= w4344 and not w4380;
w4383 <= not w4381 and not w4382;
w4384 <= not w4308 and not w4383;
w4385 <= not w4303 and w4384;
w4386 <= not w4299 and w4385;
w4387 <= not w4299 and not w4303;
w4388 <= not w4384 and not w4387;
w4389 <= not w4386 and not w4388;
w4390 <= not w4361 and not w4374;
w4391 <= not w4378 and not w4390;
w4392 <= not w4325 and not w4361;
w4393 <= not w4343 and w4392;
w4394 <= not w4379 and w4393;
w4395 <= not w4325 and not w4338;
w4396 <= not w4342 and not w4395;
w4397 <= not w4394 and w4396;
w4398 <= w4394 and not w4396;
w4399 <= not w4397 and not w4398;
w4400 <= not w4391 and not w4399;
w4401 <= not w4394 and not w4396;
w4402 <= not w4342 and w4392;
w4403 <= not w4343 and w4402;
w4404 <= not w4379 and not w4395;
w4405 <= w4403 and w4404;
w4406 <= not w4401 and not w4405;
w4407 <= w4391 and not w4406;
w4408 <= not w4400 and not w4407;
w4409 <= not w4389 and w4408;
w4410 <= not w4303 and not w4384;
w4411 <= not w4299 and w4410;
w4412 <= w4384 and not w4387;
w4413 <= not w4411 and not w4412;
w4414 <= not w4408 and not w4413;
w4415 <= not w4409 and not w4414;
w4416 <= A(58) and A(59);
w4417 <= A(58) and not A(59);
w4418 <= not A(58) and A(59);
w4419 <= not w4417 and not w4418;
w4420 <= A(60) and not w4419;
w4421 <= not w4416 and not w4420;
w4422 <= A(55) and A(56);
w4423 <= A(55) and not A(56);
w4424 <= not A(55) and A(56);
w4425 <= not w4423 and not w4424;
w4426 <= A(57) and not w4425;
w4427 <= not w4422 and not w4426;
w4428 <= w4421 and not w4427;
w4429 <= not w4421 and w4427;
w4430 <= A(57) and not w4423;
w4431 <= not w4424 and w4430;
w4432 <= not A(57) and not w4425;
w4433 <= not w4431 and not w4432;
w4434 <= A(60) and not w4417;
w4435 <= not w4418 and w4434;
w4436 <= not A(60) and not w4419;
w4437 <= not w4435 and not w4436;
w4438 <= not w4433 and not w4437;
w4439 <= not w4429 and w4438;
w4440 <= not w4428 and w4439;
w4441 <= not w4428 and not w4429;
w4442 <= not w4438 and not w4441;
w4443 <= not w4440 and not w4442;
w4444 <= not w4433 and w4437;
w4445 <= w4433 and not w4437;
w4446 <= not w4444 and not w4445;
w4447 <= w4438 and not w4441;
w4448 <= not w4421 and not w4427;
w4449 <= not w4447 and not w4448;
w4450 <= not w4446 and not w4449;
w4451 <= not w4443 and not w4450;
w4452 <= not w4443 and not w4449;
w4453 <= A(64) and A(65);
w4454 <= A(64) and not A(65);
w4455 <= not A(64) and A(65);
w4456 <= not w4454 and not w4455;
w4457 <= A(66) and not w4456;
w4458 <= not w4453 and not w4457;
w4459 <= A(61) and A(62);
w4460 <= A(61) and not A(62);
w4461 <= not A(61) and A(62);
w4462 <= not w4460 and not w4461;
w4463 <= A(63) and not w4462;
w4464 <= not w4459 and not w4463;
w4465 <= not w4458 and w4464;
w4466 <= w4458 and not w4464;
w4467 <= not w4465 and not w4466;
w4468 <= A(63) and not w4460;
w4469 <= not w4461 and w4468;
w4470 <= not A(63) and not w4462;
w4471 <= not w4469 and not w4470;
w4472 <= A(66) and not w4454;
w4473 <= not w4455 and w4472;
w4474 <= not A(66) and not w4456;
w4475 <= not w4473 and not w4474;
w4476 <= not w4471 and not w4475;
w4477 <= not w4467 and w4476;
w4478 <= not w4458 and not w4464;
w4479 <= not w4477 and not w4478;
w4480 <= not w4465 and w4476;
w4481 <= not w4466 and w4480;
w4482 <= not w4467 and not w4476;
w4483 <= not w4481 and not w4482;
w4484 <= not w4479 and not w4483;
w4485 <= not w4471 and w4475;
w4486 <= w4471 and not w4475;
w4487 <= not w4485 and not w4486;
w4488 <= not w4446 and not w4487;
w4489 <= not w4484 and w4488;
w4490 <= not w4452 and w4489;
w4491 <= not w4479 and not w4487;
w4492 <= not w4483 and not w4491;
w4493 <= not w4490 and w4492;
w4494 <= w4490 and not w4492;
w4495 <= not w4493 and not w4494;
w4496 <= not w4451 and not w4495;
w4497 <= not w4490 and not w4492;
w4498 <= not w4483 and w4488;
w4499 <= not w4484 and w4498;
w4500 <= not w4452 and not w4491;
w4501 <= w4499 and w4500;
w4502 <= not w4497 and not w4501;
w4503 <= w4451 and not w4502;
w4504 <= not w4496 and not w4503;
w4505 <= A(70) and A(71);
w4506 <= A(70) and not A(71);
w4507 <= not A(70) and A(71);
w4508 <= not w4506 and not w4507;
w4509 <= A(72) and not w4508;
w4510 <= not w4505 and not w4509;
w4511 <= A(67) and A(68);
w4512 <= A(67) and not A(68);
w4513 <= not A(67) and A(68);
w4514 <= not w4512 and not w4513;
w4515 <= A(69) and not w4514;
w4516 <= not w4511 and not w4515;
w4517 <= w4510 and not w4516;
w4518 <= not w4510 and w4516;
w4519 <= A(69) and not w4512;
w4520 <= not w4513 and w4519;
w4521 <= not A(69) and not w4514;
w4522 <= not w4520 and not w4521;
w4523 <= A(72) and not w4506;
w4524 <= not w4507 and w4523;
w4525 <= not A(72) and not w4508;
w4526 <= not w4524 and not w4525;
w4527 <= not w4522 and not w4526;
w4528 <= not w4518 and w4527;
w4529 <= not w4517 and w4528;
w4530 <= not w4517 and not w4518;
w4531 <= not w4527 and not w4530;
w4532 <= not w4529 and not w4531;
w4533 <= not w4522 and w4526;
w4534 <= w4522 and not w4526;
w4535 <= not w4533 and not w4534;
w4536 <= w4527 and not w4530;
w4537 <= not w4510 and not w4516;
w4538 <= not w4536 and not w4537;
w4539 <= not w4535 and not w4538;
w4540 <= not w4532 and not w4539;
w4541 <= not w4532 and not w4538;
w4542 <= A(76) and A(77);
w4543 <= A(76) and not A(77);
w4544 <= not A(76) and A(77);
w4545 <= not w4543 and not w4544;
w4546 <= A(78) and not w4545;
w4547 <= not w4542 and not w4546;
w4548 <= A(73) and A(74);
w4549 <= A(73) and not A(74);
w4550 <= not A(73) and A(74);
w4551 <= not w4549 and not w4550;
w4552 <= A(75) and not w4551;
w4553 <= not w4548 and not w4552;
w4554 <= not w4547 and w4553;
w4555 <= w4547 and not w4553;
w4556 <= not w4554 and not w4555;
w4557 <= A(75) and not w4549;
w4558 <= not w4550 and w4557;
w4559 <= not A(75) and not w4551;
w4560 <= not w4558 and not w4559;
w4561 <= A(78) and not w4543;
w4562 <= not w4544 and w4561;
w4563 <= not A(78) and not w4545;
w4564 <= not w4562 and not w4563;
w4565 <= not w4560 and not w4564;
w4566 <= not w4556 and w4565;
w4567 <= not w4547 and not w4553;
w4568 <= not w4566 and not w4567;
w4569 <= not w4554 and w4565;
w4570 <= not w4555 and w4569;
w4571 <= not w4556 and not w4565;
w4572 <= not w4570 and not w4571;
w4573 <= not w4568 and not w4572;
w4574 <= not w4560 and w4564;
w4575 <= w4560 and not w4564;
w4576 <= not w4574 and not w4575;
w4577 <= not w4535 and not w4576;
w4578 <= not w4573 and w4577;
w4579 <= not w4541 and w4578;
w4580 <= not w4568 and not w4576;
w4581 <= not w4572 and not w4580;
w4582 <= not w4579 and not w4581;
w4583 <= not w4572 and w4577;
w4584 <= not w4573 and w4583;
w4585 <= not w4541 and not w4580;
w4586 <= w4584 and w4585;
w4587 <= not w4582 and not w4586;
w4588 <= w4540 and not w4587;
w4589 <= not w4579 and w4581;
w4590 <= w4579 and not w4581;
w4591 <= not w4589 and not w4590;
w4592 <= not w4540 and not w4591;
w4593 <= not w4573 and not w4576;
w4594 <= not w4535 and not w4541;
w4595 <= not w4593 and w4594;
w4596 <= w4593 and not w4594;
w4597 <= not w4595 and not w4596;
w4598 <= not w4484 and not w4487;
w4599 <= not w4446 and not w4452;
w4600 <= not w4598 and w4599;
w4601 <= w4598 and not w4599;
w4602 <= not w4600 and not w4601;
w4603 <= not w4597 and not w4602;
w4604 <= not w4592 and not w4603;
w4605 <= not w4588 and w4604;
w4606 <= not w4588 and not w4592;
w4607 <= w4603 and not w4606;
w4608 <= not w4605 and not w4607;
w4609 <= not w4504 and not w4608;
w4610 <= not w4592 and w4603;
w4611 <= not w4588 and w4610;
w4612 <= not w4603 and not w4606;
w4613 <= not w4611 and not w4612;
w4614 <= w4504 and not w4613;
w4615 <= not w4597 and w4602;
w4616 <= w4597 and not w4602;
w4617 <= not w4615 and not w4616;
w4618 <= not w4308 and w4383;
w4619 <= w4308 and not w4383;
w4620 <= not w4618 and not w4619;
w4621 <= not w4617 and not w4620;
w4622 <= not w4614 and not w4621;
w4623 <= not w4609 and w4622;
w4624 <= not w4609 and not w4614;
w4625 <= w4621 and not w4624;
w4626 <= not w4623 and not w4625;
w4627 <= not w4415 and not w4626;
w4628 <= not w4614 and w4621;
w4629 <= not w4609 and w4628;
w4630 <= not w4621 and not w4624;
w4631 <= not w4629 and not w4630;
w4632 <= w4415 and not w4631;
w4633 <= not w4617 and w4620;
w4634 <= w4617 and not w4620;
w4635 <= not w4633 and not w4634;
w4636 <= not w4089 and w4161;
w4637 <= not w4087 and not w4161;
w4638 <= not w4088 and w4637;
w4639 <= not w4636 and not w4638;
w4640 <= not w4635 and not w4639;
w4641 <= not w4632 and not w4640;
w4642 <= not w4627 and w4641;
w4643 <= not w4627 and not w4632;
w4644 <= w4640 and not w4643;
w4645 <= not w4642 and not w4644;
w4646 <= not w4215 and not w4645;
w4647 <= not w4632 and w4640;
w4648 <= not w4627 and w4647;
w4649 <= not w4640 and not w4643;
w4650 <= not w4648 and not w4649;
w4651 <= w4215 and not w4650;
w4652 <= not w4635 and w4639;
w4653 <= w4635 and not w4639;
w4654 <= not w4652 and not w4653;
w4655 <= not w3671 and w3824;
w4656 <= w3671 and not w3824;
w4657 <= not w4655 and not w4656;
w4658 <= not w4654 and not w4657;
w4659 <= not w4651 and not w4658;
w4660 <= not w4646 and w4659;
w4661 <= not w4646 and not w4651;
w4662 <= w4658 and not w4661;
w4663 <= not w4660 and not w4662;
w4664 <= not w3887 and not w4663;
w4665 <= not w4651 and w4658;
w4666 <= not w4646 and w4665;
w4667 <= not w4658 and not w4661;
w4668 <= not w4666 and not w4667;
w4669 <= w3887 and not w4668;
w4670 <= not w4654 and w4657;
w4671 <= not w4652 and not w4657;
w4672 <= not w4653 and w4671;
w4673 <= not w4670 and not w4672;
w4674 <= not A(937) and A(938);
w4675 <= A(937) and not A(938);
w4676 <= A(939) and not w4675;
w4677 <= not w4674 and w4676;
w4678 <= not w4674 and not w4675;
w4679 <= not A(939) and not w4678;
w4680 <= not w4677 and not w4679;
w4681 <= not A(940) and A(941);
w4682 <= A(940) and not A(941);
w4683 <= A(942) and not w4682;
w4684 <= not w4681 and w4683;
w4685 <= not w4681 and not w4682;
w4686 <= not A(942) and not w4685;
w4687 <= not w4684 and not w4686;
w4688 <= not w4680 and w4687;
w4689 <= w4680 and not w4687;
w4690 <= not w4688 and not w4689;
w4691 <= A(940) and A(941);
w4692 <= A(942) and not w4685;
w4693 <= not w4691 and not w4692;
w4694 <= A(937) and A(938);
w4695 <= A(939) and not w4678;
w4696 <= not w4694 and not w4695;
w4697 <= not w4693 and w4696;
w4698 <= w4693 and not w4696;
w4699 <= not w4697 and not w4698;
w4700 <= not w4680 and not w4687;
w4701 <= not w4699 and w4700;
w4702 <= not w4693 and not w4696;
w4703 <= not w4701 and not w4702;
w4704 <= not w4697 and w4700;
w4705 <= not w4698 and w4704;
w4706 <= not w4699 and not w4700;
w4707 <= not w4705 and not w4706;
w4708 <= not w4703 and not w4707;
w4709 <= not w4690 and not w4708;
w4710 <= not A(931) and A(932);
w4711 <= A(931) and not A(932);
w4712 <= A(933) and not w4711;
w4713 <= not w4710 and w4712;
w4714 <= not w4710 and not w4711;
w4715 <= not A(933) and not w4714;
w4716 <= not w4713 and not w4715;
w4717 <= not A(934) and A(935);
w4718 <= A(934) and not A(935);
w4719 <= A(936) and not w4718;
w4720 <= not w4717 and w4719;
w4721 <= not w4717 and not w4718;
w4722 <= not A(936) and not w4721;
w4723 <= not w4720 and not w4722;
w4724 <= not w4716 and w4723;
w4725 <= w4716 and not w4723;
w4726 <= not w4724 and not w4725;
w4727 <= A(934) and A(935);
w4728 <= A(936) and not w4721;
w4729 <= not w4727 and not w4728;
w4730 <= A(931) and A(932);
w4731 <= A(933) and not w4714;
w4732 <= not w4730 and not w4731;
w4733 <= not w4729 and w4732;
w4734 <= w4729 and not w4732;
w4735 <= not w4733 and not w4734;
w4736 <= not w4716 and not w4723;
w4737 <= not w4735 and w4736;
w4738 <= not w4729 and not w4732;
w4739 <= not w4737 and not w4738;
w4740 <= not w4733 and w4736;
w4741 <= not w4734 and w4740;
w4742 <= not w4735 and not w4736;
w4743 <= not w4741 and not w4742;
w4744 <= not w4739 and not w4743;
w4745 <= not w4726 and not w4744;
w4746 <= not w4709 and w4745;
w4747 <= w4709 and not w4745;
w4748 <= not w4746 and not w4747;
w4749 <= not A(925) and A(926);
w4750 <= A(925) and not A(926);
w4751 <= A(927) and not w4750;
w4752 <= not w4749 and w4751;
w4753 <= not w4749 and not w4750;
w4754 <= not A(927) and not w4753;
w4755 <= not w4752 and not w4754;
w4756 <= not A(928) and A(929);
w4757 <= A(928) and not A(929);
w4758 <= A(930) and not w4757;
w4759 <= not w4756 and w4758;
w4760 <= not w4756 and not w4757;
w4761 <= not A(930) and not w4760;
w4762 <= not w4759 and not w4761;
w4763 <= not w4755 and w4762;
w4764 <= w4755 and not w4762;
w4765 <= not w4763 and not w4764;
w4766 <= A(928) and A(929);
w4767 <= A(930) and not w4760;
w4768 <= not w4766 and not w4767;
w4769 <= A(925) and A(926);
w4770 <= A(927) and not w4753;
w4771 <= not w4769 and not w4770;
w4772 <= not w4768 and w4771;
w4773 <= w4768 and not w4771;
w4774 <= not w4772 and not w4773;
w4775 <= not w4755 and not w4762;
w4776 <= not w4774 and w4775;
w4777 <= not w4768 and not w4771;
w4778 <= not w4776 and not w4777;
w4779 <= not w4772 and w4775;
w4780 <= not w4773 and w4779;
w4781 <= not w4774 and not w4775;
w4782 <= not w4780 and not w4781;
w4783 <= not w4778 and not w4782;
w4784 <= not w4765 and not w4783;
w4785 <= not A(919) and A(920);
w4786 <= A(919) and not A(920);
w4787 <= A(921) and not w4786;
w4788 <= not w4785 and w4787;
w4789 <= not w4785 and not w4786;
w4790 <= not A(921) and not w4789;
w4791 <= not w4788 and not w4790;
w4792 <= not A(922) and A(923);
w4793 <= A(922) and not A(923);
w4794 <= A(924) and not w4793;
w4795 <= not w4792 and w4794;
w4796 <= not w4792 and not w4793;
w4797 <= not A(924) and not w4796;
w4798 <= not w4795 and not w4797;
w4799 <= not w4791 and w4798;
w4800 <= w4791 and not w4798;
w4801 <= not w4799 and not w4800;
w4802 <= A(922) and A(923);
w4803 <= A(924) and not w4796;
w4804 <= not w4802 and not w4803;
w4805 <= A(919) and A(920);
w4806 <= A(921) and not w4789;
w4807 <= not w4805 and not w4806;
w4808 <= not w4804 and w4807;
w4809 <= w4804 and not w4807;
w4810 <= not w4808 and not w4809;
w4811 <= not w4791 and not w4798;
w4812 <= not w4810 and w4811;
w4813 <= not w4804 and not w4807;
w4814 <= not w4812 and not w4813;
w4815 <= not w4808 and w4811;
w4816 <= not w4809 and w4815;
w4817 <= not w4810 and not w4811;
w4818 <= not w4816 and not w4817;
w4819 <= not w4814 and not w4818;
w4820 <= not w4801 and not w4819;
w4821 <= not w4784 and w4820;
w4822 <= w4784 and not w4820;
w4823 <= not w4821 and not w4822;
w4824 <= not w4748 and w4823;
w4825 <= w4748 and not w4823;
w4826 <= not w4824 and not w4825;
w4827 <= not A(913) and A(914);
w4828 <= A(913) and not A(914);
w4829 <= A(915) and not w4828;
w4830 <= not w4827 and w4829;
w4831 <= not w4827 and not w4828;
w4832 <= not A(915) and not w4831;
w4833 <= not w4830 and not w4832;
w4834 <= not A(916) and A(917);
w4835 <= A(916) and not A(917);
w4836 <= A(918) and not w4835;
w4837 <= not w4834 and w4836;
w4838 <= not w4834 and not w4835;
w4839 <= not A(918) and not w4838;
w4840 <= not w4837 and not w4839;
w4841 <= not w4833 and w4840;
w4842 <= w4833 and not w4840;
w4843 <= not w4841 and not w4842;
w4844 <= A(916) and A(917);
w4845 <= A(918) and not w4838;
w4846 <= not w4844 and not w4845;
w4847 <= A(913) and A(914);
w4848 <= A(915) and not w4831;
w4849 <= not w4847 and not w4848;
w4850 <= not w4846 and w4849;
w4851 <= w4846 and not w4849;
w4852 <= not w4850 and not w4851;
w4853 <= not w4833 and not w4840;
w4854 <= not w4852 and w4853;
w4855 <= not w4846 and not w4849;
w4856 <= not w4854 and not w4855;
w4857 <= not w4850 and w4853;
w4858 <= not w4851 and w4857;
w4859 <= not w4852 and not w4853;
w4860 <= not w4858 and not w4859;
w4861 <= not w4856 and not w4860;
w4862 <= not w4843 and not w4861;
w4863 <= not A(907) and A(908);
w4864 <= A(907) and not A(908);
w4865 <= A(909) and not w4864;
w4866 <= not w4863 and w4865;
w4867 <= not w4863 and not w4864;
w4868 <= not A(909) and not w4867;
w4869 <= not w4866 and not w4868;
w4870 <= not A(910) and A(911);
w4871 <= A(910) and not A(911);
w4872 <= A(912) and not w4871;
w4873 <= not w4870 and w4872;
w4874 <= not w4870 and not w4871;
w4875 <= not A(912) and not w4874;
w4876 <= not w4873 and not w4875;
w4877 <= not w4869 and w4876;
w4878 <= w4869 and not w4876;
w4879 <= not w4877 and not w4878;
w4880 <= A(910) and A(911);
w4881 <= A(912) and not w4874;
w4882 <= not w4880 and not w4881;
w4883 <= A(907) and A(908);
w4884 <= A(909) and not w4867;
w4885 <= not w4883 and not w4884;
w4886 <= not w4882 and w4885;
w4887 <= w4882 and not w4885;
w4888 <= not w4886 and not w4887;
w4889 <= not w4869 and not w4876;
w4890 <= not w4888 and w4889;
w4891 <= not w4882 and not w4885;
w4892 <= not w4890 and not w4891;
w4893 <= not w4886 and w4889;
w4894 <= not w4887 and w4893;
w4895 <= not w4888 and not w4889;
w4896 <= not w4894 and not w4895;
w4897 <= not w4892 and not w4896;
w4898 <= not w4879 and not w4897;
w4899 <= not w4862 and w4898;
w4900 <= w4862 and not w4898;
w4901 <= not w4899 and not w4900;
w4902 <= not A(901) and A(902);
w4903 <= A(901) and not A(902);
w4904 <= A(903) and not w4903;
w4905 <= not w4902 and w4904;
w4906 <= not w4902 and not w4903;
w4907 <= not A(903) and not w4906;
w4908 <= not w4905 and not w4907;
w4909 <= not A(904) and A(905);
w4910 <= A(904) and not A(905);
w4911 <= A(906) and not w4910;
w4912 <= not w4909 and w4911;
w4913 <= not w4909 and not w4910;
w4914 <= not A(906) and not w4913;
w4915 <= not w4912 and not w4914;
w4916 <= not w4908 and w4915;
w4917 <= w4908 and not w4915;
w4918 <= not w4916 and not w4917;
w4919 <= A(904) and A(905);
w4920 <= A(906) and not w4913;
w4921 <= not w4919 and not w4920;
w4922 <= A(901) and A(902);
w4923 <= A(903) and not w4906;
w4924 <= not w4922 and not w4923;
w4925 <= not w4921 and w4924;
w4926 <= w4921 and not w4924;
w4927 <= not w4925 and not w4926;
w4928 <= not w4908 and not w4915;
w4929 <= not w4927 and w4928;
w4930 <= not w4921 and not w4924;
w4931 <= not w4929 and not w4930;
w4932 <= not w4925 and w4928;
w4933 <= not w4926 and w4932;
w4934 <= not w4927 and not w4928;
w4935 <= not w4933 and not w4934;
w4936 <= not w4931 and not w4935;
w4937 <= not w4918 and not w4936;
w4938 <= not A(895) and A(896);
w4939 <= A(895) and not A(896);
w4940 <= A(897) and not w4939;
w4941 <= not w4938 and w4940;
w4942 <= not w4938 and not w4939;
w4943 <= not A(897) and not w4942;
w4944 <= not w4941 and not w4943;
w4945 <= not A(898) and A(899);
w4946 <= A(898) and not A(899);
w4947 <= A(900) and not w4946;
w4948 <= not w4945 and w4947;
w4949 <= not w4945 and not w4946;
w4950 <= not A(900) and not w4949;
w4951 <= not w4948 and not w4950;
w4952 <= not w4944 and w4951;
w4953 <= w4944 and not w4951;
w4954 <= not w4952 and not w4953;
w4955 <= A(898) and A(899);
w4956 <= A(900) and not w4949;
w4957 <= not w4955 and not w4956;
w4958 <= A(895) and A(896);
w4959 <= A(897) and not w4942;
w4960 <= not w4958 and not w4959;
w4961 <= not w4957 and w4960;
w4962 <= w4957 and not w4960;
w4963 <= not w4961 and not w4962;
w4964 <= not w4944 and not w4951;
w4965 <= not w4963 and w4964;
w4966 <= not w4957 and not w4960;
w4967 <= not w4965 and not w4966;
w4968 <= not w4961 and w4964;
w4969 <= not w4962 and w4968;
w4970 <= not w4963 and not w4964;
w4971 <= not w4969 and not w4970;
w4972 <= not w4967 and not w4971;
w4973 <= not w4954 and not w4972;
w4974 <= not w4937 and w4973;
w4975 <= w4937 and not w4973;
w4976 <= not w4974 and not w4975;
w4977 <= not w4901 and w4976;
w4978 <= w4901 and not w4976;
w4979 <= not w4977 and not w4978;
w4980 <= not w4826 and w4979;
w4981 <= w4826 and not w4979;
w4982 <= not w4980 and not w4981;
w4983 <= not A(889) and A(890);
w4984 <= A(889) and not A(890);
w4985 <= A(891) and not w4984;
w4986 <= not w4983 and w4985;
w4987 <= not w4983 and not w4984;
w4988 <= not A(891) and not w4987;
w4989 <= not w4986 and not w4988;
w4990 <= not A(892) and A(893);
w4991 <= A(892) and not A(893);
w4992 <= A(894) and not w4991;
w4993 <= not w4990 and w4992;
w4994 <= not w4990 and not w4991;
w4995 <= not A(894) and not w4994;
w4996 <= not w4993 and not w4995;
w4997 <= not w4989 and w4996;
w4998 <= w4989 and not w4996;
w4999 <= not w4997 and not w4998;
w5000 <= A(892) and A(893);
w5001 <= A(894) and not w4994;
w5002 <= not w5000 and not w5001;
w5003 <= A(889) and A(890);
w5004 <= A(891) and not w4987;
w5005 <= not w5003 and not w5004;
w5006 <= not w5002 and w5005;
w5007 <= w5002 and not w5005;
w5008 <= not w5006 and not w5007;
w5009 <= not w4989 and not w4996;
w5010 <= not w5008 and w5009;
w5011 <= not w5002 and not w5005;
w5012 <= not w5010 and not w5011;
w5013 <= not w5006 and w5009;
w5014 <= not w5007 and w5013;
w5015 <= not w5008 and not w5009;
w5016 <= not w5014 and not w5015;
w5017 <= not w5012 and not w5016;
w5018 <= not w4999 and not w5017;
w5019 <= not A(883) and A(884);
w5020 <= A(883) and not A(884);
w5021 <= A(885) and not w5020;
w5022 <= not w5019 and w5021;
w5023 <= not w5019 and not w5020;
w5024 <= not A(885) and not w5023;
w5025 <= not w5022 and not w5024;
w5026 <= not A(886) and A(887);
w5027 <= A(886) and not A(887);
w5028 <= A(888) and not w5027;
w5029 <= not w5026 and w5028;
w5030 <= not w5026 and not w5027;
w5031 <= not A(888) and not w5030;
w5032 <= not w5029 and not w5031;
w5033 <= not w5025 and w5032;
w5034 <= w5025 and not w5032;
w5035 <= not w5033 and not w5034;
w5036 <= A(886) and A(887);
w5037 <= A(888) and not w5030;
w5038 <= not w5036 and not w5037;
w5039 <= A(883) and A(884);
w5040 <= A(885) and not w5023;
w5041 <= not w5039 and not w5040;
w5042 <= not w5038 and w5041;
w5043 <= w5038 and not w5041;
w5044 <= not w5042 and not w5043;
w5045 <= not w5025 and not w5032;
w5046 <= not w5044 and w5045;
w5047 <= not w5038 and not w5041;
w5048 <= not w5046 and not w5047;
w5049 <= not w5042 and w5045;
w5050 <= not w5043 and w5049;
w5051 <= not w5044 and not w5045;
w5052 <= not w5050 and not w5051;
w5053 <= not w5048 and not w5052;
w5054 <= not w5035 and not w5053;
w5055 <= not w5018 and w5054;
w5056 <= w5018 and not w5054;
w5057 <= not w5055 and not w5056;
w5058 <= not A(877) and A(878);
w5059 <= A(877) and not A(878);
w5060 <= A(879) and not w5059;
w5061 <= not w5058 and w5060;
w5062 <= not w5058 and not w5059;
w5063 <= not A(879) and not w5062;
w5064 <= not w5061 and not w5063;
w5065 <= not A(880) and A(881);
w5066 <= A(880) and not A(881);
w5067 <= A(882) and not w5066;
w5068 <= not w5065 and w5067;
w5069 <= not w5065 and not w5066;
w5070 <= not A(882) and not w5069;
w5071 <= not w5068 and not w5070;
w5072 <= not w5064 and w5071;
w5073 <= w5064 and not w5071;
w5074 <= not w5072 and not w5073;
w5075 <= A(880) and A(881);
w5076 <= A(882) and not w5069;
w5077 <= not w5075 and not w5076;
w5078 <= A(877) and A(878);
w5079 <= A(879) and not w5062;
w5080 <= not w5078 and not w5079;
w5081 <= not w5077 and w5080;
w5082 <= w5077 and not w5080;
w5083 <= not w5081 and not w5082;
w5084 <= not w5064 and not w5071;
w5085 <= not w5083 and w5084;
w5086 <= not w5077 and not w5080;
w5087 <= not w5085 and not w5086;
w5088 <= not w5081 and w5084;
w5089 <= not w5082 and w5088;
w5090 <= not w5083 and not w5084;
w5091 <= not w5089 and not w5090;
w5092 <= not w5087 and not w5091;
w5093 <= not w5074 and not w5092;
w5094 <= not A(871) and A(872);
w5095 <= A(871) and not A(872);
w5096 <= A(873) and not w5095;
w5097 <= not w5094 and w5096;
w5098 <= not w5094 and not w5095;
w5099 <= not A(873) and not w5098;
w5100 <= not w5097 and not w5099;
w5101 <= not A(874) and A(875);
w5102 <= A(874) and not A(875);
w5103 <= A(876) and not w5102;
w5104 <= not w5101 and w5103;
w5105 <= not w5101 and not w5102;
w5106 <= not A(876) and not w5105;
w5107 <= not w5104 and not w5106;
w5108 <= not w5100 and w5107;
w5109 <= w5100 and not w5107;
w5110 <= not w5108 and not w5109;
w5111 <= A(874) and A(875);
w5112 <= A(876) and not w5105;
w5113 <= not w5111 and not w5112;
w5114 <= A(871) and A(872);
w5115 <= A(873) and not w5098;
w5116 <= not w5114 and not w5115;
w5117 <= not w5113 and w5116;
w5118 <= w5113 and not w5116;
w5119 <= not w5117 and not w5118;
w5120 <= not w5100 and not w5107;
w5121 <= not w5119 and w5120;
w5122 <= not w5113 and not w5116;
w5123 <= not w5121 and not w5122;
w5124 <= not w5117 and w5120;
w5125 <= not w5118 and w5124;
w5126 <= not w5119 and not w5120;
w5127 <= not w5125 and not w5126;
w5128 <= not w5123 and not w5127;
w5129 <= not w5110 and not w5128;
w5130 <= not w5093 and w5129;
w5131 <= w5093 and not w5129;
w5132 <= not w5130 and not w5131;
w5133 <= not w5057 and w5132;
w5134 <= w5057 and not w5132;
w5135 <= not w5133 and not w5134;
w5136 <= not A(865) and A(866);
w5137 <= A(865) and not A(866);
w5138 <= A(867) and not w5137;
w5139 <= not w5136 and w5138;
w5140 <= not w5136 and not w5137;
w5141 <= not A(867) and not w5140;
w5142 <= not w5139 and not w5141;
w5143 <= not A(868) and A(869);
w5144 <= A(868) and not A(869);
w5145 <= A(870) and not w5144;
w5146 <= not w5143 and w5145;
w5147 <= not w5143 and not w5144;
w5148 <= not A(870) and not w5147;
w5149 <= not w5146 and not w5148;
w5150 <= not w5142 and w5149;
w5151 <= w5142 and not w5149;
w5152 <= not w5150 and not w5151;
w5153 <= A(868) and A(869);
w5154 <= A(870) and not w5147;
w5155 <= not w5153 and not w5154;
w5156 <= A(865) and A(866);
w5157 <= A(867) and not w5140;
w5158 <= not w5156 and not w5157;
w5159 <= not w5155 and w5158;
w5160 <= w5155 and not w5158;
w5161 <= not w5159 and not w5160;
w5162 <= not w5142 and not w5149;
w5163 <= not w5161 and w5162;
w5164 <= not w5155 and not w5158;
w5165 <= not w5163 and not w5164;
w5166 <= not w5159 and w5162;
w5167 <= not w5160 and w5166;
w5168 <= not w5161 and not w5162;
w5169 <= not w5167 and not w5168;
w5170 <= not w5165 and not w5169;
w5171 <= not w5152 and not w5170;
w5172 <= not A(859) and A(860);
w5173 <= A(859) and not A(860);
w5174 <= A(861) and not w5173;
w5175 <= not w5172 and w5174;
w5176 <= not w5172 and not w5173;
w5177 <= not A(861) and not w5176;
w5178 <= not w5175 and not w5177;
w5179 <= not A(862) and A(863);
w5180 <= A(862) and not A(863);
w5181 <= A(864) and not w5180;
w5182 <= not w5179 and w5181;
w5183 <= not w5179 and not w5180;
w5184 <= not A(864) and not w5183;
w5185 <= not w5182 and not w5184;
w5186 <= not w5178 and w5185;
w5187 <= w5178 and not w5185;
w5188 <= not w5186 and not w5187;
w5189 <= A(862) and A(863);
w5190 <= A(864) and not w5183;
w5191 <= not w5189 and not w5190;
w5192 <= A(859) and A(860);
w5193 <= A(861) and not w5176;
w5194 <= not w5192 and not w5193;
w5195 <= not w5191 and w5194;
w5196 <= w5191 and not w5194;
w5197 <= not w5195 and not w5196;
w5198 <= not w5178 and not w5185;
w5199 <= not w5197 and w5198;
w5200 <= not w5191 and not w5194;
w5201 <= not w5199 and not w5200;
w5202 <= not w5195 and w5198;
w5203 <= not w5196 and w5202;
w5204 <= not w5197 and not w5198;
w5205 <= not w5203 and not w5204;
w5206 <= not w5201 and not w5205;
w5207 <= not w5188 and not w5206;
w5208 <= not w5171 and w5207;
w5209 <= w5171 and not w5207;
w5210 <= not w5208 and not w5209;
w5211 <= not A(853) and A(854);
w5212 <= A(853) and not A(854);
w5213 <= A(855) and not w5212;
w5214 <= not w5211 and w5213;
w5215 <= not w5211 and not w5212;
w5216 <= not A(855) and not w5215;
w5217 <= not w5214 and not w5216;
w5218 <= not A(856) and A(857);
w5219 <= A(856) and not A(857);
w5220 <= A(858) and not w5219;
w5221 <= not w5218 and w5220;
w5222 <= not w5218 and not w5219;
w5223 <= not A(858) and not w5222;
w5224 <= not w5221 and not w5223;
w5225 <= not w5217 and w5224;
w5226 <= w5217 and not w5224;
w5227 <= not w5225 and not w5226;
w5228 <= A(856) and A(857);
w5229 <= A(858) and not w5222;
w5230 <= not w5228 and not w5229;
w5231 <= A(853) and A(854);
w5232 <= A(855) and not w5215;
w5233 <= not w5231 and not w5232;
w5234 <= not w5230 and w5233;
w5235 <= w5230 and not w5233;
w5236 <= not w5234 and not w5235;
w5237 <= not w5217 and not w5224;
w5238 <= not w5236 and w5237;
w5239 <= not w5230 and not w5233;
w5240 <= not w5238 and not w5239;
w5241 <= not w5234 and w5237;
w5242 <= not w5235 and w5241;
w5243 <= not w5236 and not w5237;
w5244 <= not w5242 and not w5243;
w5245 <= not w5240 and not w5244;
w5246 <= not w5227 and not w5245;
w5247 <= not A(847) and A(848);
w5248 <= A(847) and not A(848);
w5249 <= A(849) and not w5248;
w5250 <= not w5247 and w5249;
w5251 <= not w5247 and not w5248;
w5252 <= not A(849) and not w5251;
w5253 <= not w5250 and not w5252;
w5254 <= not A(850) and A(851);
w5255 <= A(850) and not A(851);
w5256 <= A(852) and not w5255;
w5257 <= not w5254 and w5256;
w5258 <= not w5254 and not w5255;
w5259 <= not A(852) and not w5258;
w5260 <= not w5257 and not w5259;
w5261 <= not w5253 and w5260;
w5262 <= w5253 and not w5260;
w5263 <= not w5261 and not w5262;
w5264 <= A(850) and A(851);
w5265 <= A(852) and not w5258;
w5266 <= not w5264 and not w5265;
w5267 <= A(847) and A(848);
w5268 <= A(849) and not w5251;
w5269 <= not w5267 and not w5268;
w5270 <= not w5266 and w5269;
w5271 <= w5266 and not w5269;
w5272 <= not w5270 and not w5271;
w5273 <= not w5253 and not w5260;
w5274 <= not w5272 and w5273;
w5275 <= not w5266 and not w5269;
w5276 <= not w5274 and not w5275;
w5277 <= not w5270 and w5273;
w5278 <= not w5271 and w5277;
w5279 <= not w5272 and not w5273;
w5280 <= not w5278 and not w5279;
w5281 <= not w5276 and not w5280;
w5282 <= not w5263 and not w5281;
w5283 <= not w5246 and w5282;
w5284 <= w5246 and not w5282;
w5285 <= not w5283 and not w5284;
w5286 <= not w5210 and w5285;
w5287 <= w5210 and not w5285;
w5288 <= not w5286 and not w5287;
w5289 <= not w5135 and w5288;
w5290 <= w5135 and not w5288;
w5291 <= not w5289 and not w5290;
w5292 <= not w4982 and w5291;
w5293 <= w4982 and not w5291;
w5294 <= not w5292 and not w5293;
w5295 <= not w4673 and not w5294;
w5296 <= not w4669 and w5295;
w5297 <= not w4664 and w5296;
w5298 <= not w4664 and not w4669;
w5299 <= not w5295 and not w5298;
w5300 <= not w5297 and not w5299;
w5301 <= not w4879 and not w4892;
w5302 <= not w4896 and not w5301;
w5303 <= not w4843 and not w4879;
w5304 <= not w4861 and w5303;
w5305 <= not w4897 and w5304;
w5306 <= not w4843 and not w4856;
w5307 <= not w4860 and not w5306;
w5308 <= not w5305 and not w5307;
w5309 <= not w4860 and w5303;
w5310 <= not w4861 and w5309;
w5311 <= not w4897 and not w5306;
w5312 <= w5310 and w5311;
w5313 <= not w5308 and not w5312;
w5314 <= w5302 and not w5313;
w5315 <= not w5305 and w5307;
w5316 <= w5305 and not w5307;
w5317 <= not w5315 and not w5316;
w5318 <= not w5302 and not w5317;
w5319 <= not w4901 and not w4976;
w5320 <= not w5318 and w5319;
w5321 <= not w5314 and w5320;
w5322 <= not w5314 and not w5318;
w5323 <= not w5319 and not w5322;
w5324 <= not w5321 and not w5323;
w5325 <= not w4954 and not w4967;
w5326 <= not w4971 and not w5325;
w5327 <= not w4918 and not w4954;
w5328 <= not w4936 and w5327;
w5329 <= not w4972 and w5328;
w5330 <= not w4918 and not w4931;
w5331 <= not w4935 and not w5330;
w5332 <= not w5329 and w5331;
w5333 <= w5329 and not w5331;
w5334 <= not w5332 and not w5333;
w5335 <= not w5326 and not w5334;
w5336 <= not w5329 and not w5331;
w5337 <= not w4935 and w5327;
w5338 <= not w4936 and w5337;
w5339 <= not w4972 and not w5330;
w5340 <= w5338 and w5339;
w5341 <= not w5336 and not w5340;
w5342 <= w5326 and not w5341;
w5343 <= not w5335 and not w5342;
w5344 <= not w5324 and w5343;
w5345 <= not w5318 and not w5319;
w5346 <= not w5314 and w5345;
w5347 <= w5319 and not w5322;
w5348 <= not w5346 and not w5347;
w5349 <= not w5343 and not w5348;
w5350 <= not w5344 and not w5349;
w5351 <= not w4801 and not w4814;
w5352 <= not w4818 and not w5351;
w5353 <= not w4765 and not w4801;
w5354 <= not w4783 and w5353;
w5355 <= not w4819 and w5354;
w5356 <= not w4765 and not w4778;
w5357 <= not w4782 and not w5356;
w5358 <= not w5355 and w5357;
w5359 <= w5355 and not w5357;
w5360 <= not w5358 and not w5359;
w5361 <= not w5352 and not w5360;
w5362 <= not w5355 and not w5357;
w5363 <= not w4782 and w5353;
w5364 <= not w4783 and w5363;
w5365 <= not w4819 and not w5356;
w5366 <= w5364 and w5365;
w5367 <= not w5362 and not w5366;
w5368 <= w5352 and not w5367;
w5369 <= not w5361 and not w5368;
w5370 <= not w4726 and not w4739;
w5371 <= not w4743 and not w5370;
w5372 <= not w4690 and not w4726;
w5373 <= not w4708 and w5372;
w5374 <= not w4744 and w5373;
w5375 <= not w4690 and not w4703;
w5376 <= not w4707 and not w5375;
w5377 <= not w5374 and not w5376;
w5378 <= not w4707 and w5372;
w5379 <= not w4708 and w5378;
w5380 <= not w4744 and not w5375;
w5381 <= w5379 and w5380;
w5382 <= not w5377 and not w5381;
w5383 <= w5371 and not w5382;
w5384 <= not w5374 and w5376;
w5385 <= w5374 and not w5376;
w5386 <= not w5384 and not w5385;
w5387 <= not w5371 and not w5386;
w5388 <= not w4748 and not w4823;
w5389 <= not w5387 and not w5388;
w5390 <= not w5383 and w5389;
w5391 <= not w5383 and not w5387;
w5392 <= w5388 and not w5391;
w5393 <= not w5390 and not w5392;
w5394 <= not w5369 and not w5393;
w5395 <= not w5387 and w5388;
w5396 <= not w5383 and w5395;
w5397 <= not w5388 and not w5391;
w5398 <= not w5396 and not w5397;
w5399 <= w5369 and not w5398;
w5400 <= not w4826 and not w4979;
w5401 <= not w5399 and not w5400;
w5402 <= not w5394 and w5401;
w5403 <= not w5394 and not w5399;
w5404 <= w5400 and not w5403;
w5405 <= not w5402 and not w5404;
w5406 <= not w5350 and not w5405;
w5407 <= not w5399 and w5400;
w5408 <= not w5394 and w5407;
w5409 <= not w5400 and not w5403;
w5410 <= not w5408 and not w5409;
w5411 <= w5350 and not w5410;
w5412 <= not w4982 and not w5291;
w5413 <= not w5411 and w5412;
w5414 <= not w5406 and w5413;
w5415 <= not w5406 and not w5411;
w5416 <= not w5412 and not w5415;
w5417 <= not w5414 and not w5416;
w5418 <= not w5110 and not w5123;
w5419 <= not w5127 and not w5418;
w5420 <= not w5074 and not w5110;
w5421 <= not w5092 and w5420;
w5422 <= not w5128 and w5421;
w5423 <= not w5074 and not w5087;
w5424 <= not w5091 and not w5423;
w5425 <= not w5422 and w5424;
w5426 <= w5422 and not w5424;
w5427 <= not w5425 and not w5426;
w5428 <= not w5419 and not w5427;
w5429 <= not w5422 and not w5424;
w5430 <= not w5091 and w5420;
w5431 <= not w5092 and w5430;
w5432 <= not w5128 and not w5423;
w5433 <= w5431 and w5432;
w5434 <= not w5429 and not w5433;
w5435 <= w5419 and not w5434;
w5436 <= not w5428 and not w5435;
w5437 <= not w5035 and not w5048;
w5438 <= not w5052 and not w5437;
w5439 <= not w4999 and not w5035;
w5440 <= not w5017 and w5439;
w5441 <= not w5053 and w5440;
w5442 <= not w4999 and not w5012;
w5443 <= not w5016 and not w5442;
w5444 <= not w5441 and not w5443;
w5445 <= not w5016 and w5439;
w5446 <= not w5017 and w5445;
w5447 <= not w5053 and not w5442;
w5448 <= w5446 and w5447;
w5449 <= not w5444 and not w5448;
w5450 <= w5438 and not w5449;
w5451 <= not w5441 and w5443;
w5452 <= w5441 and not w5443;
w5453 <= not w5451 and not w5452;
w5454 <= not w5438 and not w5453;
w5455 <= not w5057 and not w5132;
w5456 <= not w5454 and not w5455;
w5457 <= not w5450 and w5456;
w5458 <= not w5450 and not w5454;
w5459 <= w5455 and not w5458;
w5460 <= not w5457 and not w5459;
w5461 <= not w5436 and not w5460;
w5462 <= not w5454 and w5455;
w5463 <= not w5450 and w5462;
w5464 <= not w5455 and not w5458;
w5465 <= not w5463 and not w5464;
w5466 <= w5436 and not w5465;
w5467 <= not w5135 and not w5288;
w5468 <= not w5466 and w5467;
w5469 <= not w5461 and w5468;
w5470 <= not w5461 and not w5466;
w5471 <= not w5467 and not w5470;
w5472 <= not w5469 and not w5471;
w5473 <= not w5188 and not w5201;
w5474 <= not w5205 and not w5473;
w5475 <= not w5152 and not w5188;
w5476 <= not w5170 and w5475;
w5477 <= not w5206 and w5476;
w5478 <= not w5152 and not w5165;
w5479 <= not w5169 and not w5478;
w5480 <= not w5477 and not w5479;
w5481 <= not w5169 and w5475;
w5482 <= not w5170 and w5481;
w5483 <= not w5206 and not w5478;
w5484 <= w5482 and w5483;
w5485 <= not w5480 and not w5484;
w5486 <= w5474 and not w5485;
w5487 <= not w5477 and w5479;
w5488 <= w5477 and not w5479;
w5489 <= not w5487 and not w5488;
w5490 <= not w5474 and not w5489;
w5491 <= not w5210 and not w5285;
w5492 <= not w5490 and w5491;
w5493 <= not w5486 and w5492;
w5494 <= not w5486 and not w5490;
w5495 <= not w5491 and not w5494;
w5496 <= not w5493 and not w5495;
w5497 <= not w5263 and not w5276;
w5498 <= not w5280 and not w5497;
w5499 <= not w5227 and not w5263;
w5500 <= not w5245 and w5499;
w5501 <= not w5281 and w5500;
w5502 <= not w5227 and not w5240;
w5503 <= not w5244 and not w5502;
w5504 <= not w5501 and w5503;
w5505 <= w5501 and not w5503;
w5506 <= not w5504 and not w5505;
w5507 <= not w5498 and not w5506;
w5508 <= not w5501 and not w5503;
w5509 <= not w5244 and w5499;
w5510 <= not w5245 and w5509;
w5511 <= not w5281 and not w5502;
w5512 <= w5510 and w5511;
w5513 <= not w5508 and not w5512;
w5514 <= w5498 and not w5513;
w5515 <= not w5507 and not w5514;
w5516 <= not w5496 and w5515;
w5517 <= not w5490 and not w5491;
w5518 <= not w5486 and w5517;
w5519 <= w5491 and not w5494;
w5520 <= not w5518 and not w5519;
w5521 <= not w5515 and not w5520;
w5522 <= not w5516 and not w5521;
w5523 <= not w5472 and w5522;
w5524 <= not w5466 and not w5467;
w5525 <= not w5461 and w5524;
w5526 <= w5467 and not w5470;
w5527 <= not w5525 and not w5526;
w5528 <= not w5522 and not w5527;
w5529 <= not w5523 and not w5528;
w5530 <= not w5417 and w5529;
w5531 <= not w5411 and not w5412;
w5532 <= not w5406 and w5531;
w5533 <= w5412 and not w5415;
w5534 <= not w5532 and not w5533;
w5535 <= not w5529 and not w5534;
w5536 <= not w5530 and not w5535;
w5537 <= not w5300 and w5536;
w5538 <= not w4669 and not w5295;
w5539 <= not w4664 and w5538;
w5540 <= w5295 and not w5298;
w5541 <= not w5539 and not w5540;
w5542 <= not w5536 and not w5541;
w5543 <= not w5537 and not w5542;
w5544 <= A(202) and A(203);
w5545 <= A(202) and not A(203);
w5546 <= not A(202) and A(203);
w5547 <= not w5545 and not w5546;
w5548 <= A(204) and not w5547;
w5549 <= not w5544 and not w5548;
w5550 <= A(199) and A(200);
w5551 <= A(199) and not A(200);
w5552 <= not A(199) and A(200);
w5553 <= not w5551 and not w5552;
w5554 <= A(201) and not w5553;
w5555 <= not w5550 and not w5554;
w5556 <= w5549 and not w5555;
w5557 <= not w5549 and w5555;
w5558 <= A(201) and not w5551;
w5559 <= not w5552 and w5558;
w5560 <= not A(201) and not w5553;
w5561 <= not w5559 and not w5560;
w5562 <= A(204) and not w5545;
w5563 <= not w5546 and w5562;
w5564 <= not A(204) and not w5547;
w5565 <= not w5563 and not w5564;
w5566 <= not w5561 and not w5565;
w5567 <= not w5557 and w5566;
w5568 <= not w5556 and w5567;
w5569 <= not w5556 and not w5557;
w5570 <= not w5566 and not w5569;
w5571 <= not w5568 and not w5570;
w5572 <= not w5561 and w5565;
w5573 <= w5561 and not w5565;
w5574 <= not w5572 and not w5573;
w5575 <= w5566 and not w5569;
w5576 <= not w5549 and not w5555;
w5577 <= not w5575 and not w5576;
w5578 <= not w5574 and not w5577;
w5579 <= not w5571 and not w5578;
w5580 <= not w5571 and not w5577;
w5581 <= A(208) and A(209);
w5582 <= A(208) and not A(209);
w5583 <= not A(208) and A(209);
w5584 <= not w5582 and not w5583;
w5585 <= A(210) and not w5584;
w5586 <= not w5581 and not w5585;
w5587 <= A(205) and A(206);
w5588 <= A(205) and not A(206);
w5589 <= not A(205) and A(206);
w5590 <= not w5588 and not w5589;
w5591 <= A(207) and not w5590;
w5592 <= not w5587 and not w5591;
w5593 <= not w5586 and w5592;
w5594 <= w5586 and not w5592;
w5595 <= not w5593 and not w5594;
w5596 <= A(207) and not w5588;
w5597 <= not w5589 and w5596;
w5598 <= not A(207) and not w5590;
w5599 <= not w5597 and not w5598;
w5600 <= A(210) and not w5582;
w5601 <= not w5583 and w5600;
w5602 <= not A(210) and not w5584;
w5603 <= not w5601 and not w5602;
w5604 <= not w5599 and not w5603;
w5605 <= not w5595 and w5604;
w5606 <= not w5586 and not w5592;
w5607 <= not w5605 and not w5606;
w5608 <= not w5593 and w5604;
w5609 <= not w5594 and w5608;
w5610 <= not w5595 and not w5604;
w5611 <= not w5609 and not w5610;
w5612 <= not w5607 and not w5611;
w5613 <= not w5599 and w5603;
w5614 <= w5599 and not w5603;
w5615 <= not w5613 and not w5614;
w5616 <= not w5574 and not w5615;
w5617 <= not w5612 and w5616;
w5618 <= not w5580 and w5617;
w5619 <= not w5607 and not w5615;
w5620 <= not w5611 and not w5619;
w5621 <= not w5618 and w5620;
w5622 <= w5618 and not w5620;
w5623 <= not w5621 and not w5622;
w5624 <= not w5579 and not w5623;
w5625 <= not w5618 and not w5620;
w5626 <= not w5611 and w5616;
w5627 <= not w5612 and w5626;
w5628 <= not w5580 and not w5619;
w5629 <= w5627 and w5628;
w5630 <= not w5625 and not w5629;
w5631 <= w5579 and not w5630;
w5632 <= not w5624 and not w5631;
w5633 <= A(214) and A(215);
w5634 <= A(214) and not A(215);
w5635 <= not A(214) and A(215);
w5636 <= not w5634 and not w5635;
w5637 <= A(216) and not w5636;
w5638 <= not w5633 and not w5637;
w5639 <= A(211) and A(212);
w5640 <= A(211) and not A(212);
w5641 <= not A(211) and A(212);
w5642 <= not w5640 and not w5641;
w5643 <= A(213) and not w5642;
w5644 <= not w5639 and not w5643;
w5645 <= w5638 and not w5644;
w5646 <= not w5638 and w5644;
w5647 <= A(213) and not w5640;
w5648 <= not w5641 and w5647;
w5649 <= not A(213) and not w5642;
w5650 <= not w5648 and not w5649;
w5651 <= A(216) and not w5634;
w5652 <= not w5635 and w5651;
w5653 <= not A(216) and not w5636;
w5654 <= not w5652 and not w5653;
w5655 <= not w5650 and not w5654;
w5656 <= not w5646 and w5655;
w5657 <= not w5645 and w5656;
w5658 <= not w5645 and not w5646;
w5659 <= not w5655 and not w5658;
w5660 <= not w5657 and not w5659;
w5661 <= not w5650 and w5654;
w5662 <= w5650 and not w5654;
w5663 <= not w5661 and not w5662;
w5664 <= w5655 and not w5658;
w5665 <= not w5638 and not w5644;
w5666 <= not w5664 and not w5665;
w5667 <= not w5663 and not w5666;
w5668 <= not w5660 and not w5667;
w5669 <= not w5660 and not w5666;
w5670 <= A(220) and A(221);
w5671 <= A(220) and not A(221);
w5672 <= not A(220) and A(221);
w5673 <= not w5671 and not w5672;
w5674 <= A(222) and not w5673;
w5675 <= not w5670 and not w5674;
w5676 <= A(217) and A(218);
w5677 <= A(217) and not A(218);
w5678 <= not A(217) and A(218);
w5679 <= not w5677 and not w5678;
w5680 <= A(219) and not w5679;
w5681 <= not w5676 and not w5680;
w5682 <= not w5675 and w5681;
w5683 <= w5675 and not w5681;
w5684 <= not w5682 and not w5683;
w5685 <= A(219) and not w5677;
w5686 <= not w5678 and w5685;
w5687 <= not A(219) and not w5679;
w5688 <= not w5686 and not w5687;
w5689 <= A(222) and not w5671;
w5690 <= not w5672 and w5689;
w5691 <= not A(222) and not w5673;
w5692 <= not w5690 and not w5691;
w5693 <= not w5688 and not w5692;
w5694 <= not w5684 and w5693;
w5695 <= not w5675 and not w5681;
w5696 <= not w5694 and not w5695;
w5697 <= not w5682 and w5693;
w5698 <= not w5683 and w5697;
w5699 <= not w5684 and not w5693;
w5700 <= not w5698 and not w5699;
w5701 <= not w5696 and not w5700;
w5702 <= not w5688 and w5692;
w5703 <= w5688 and not w5692;
w5704 <= not w5702 and not w5703;
w5705 <= not w5663 and not w5704;
w5706 <= not w5701 and w5705;
w5707 <= not w5669 and w5706;
w5708 <= not w5696 and not w5704;
w5709 <= not w5700 and not w5708;
w5710 <= not w5707 and not w5709;
w5711 <= not w5700 and w5705;
w5712 <= not w5701 and w5711;
w5713 <= not w5669 and not w5708;
w5714 <= w5712 and w5713;
w5715 <= not w5710 and not w5714;
w5716 <= w5668 and not w5715;
w5717 <= not w5707 and w5709;
w5718 <= w5707 and not w5709;
w5719 <= not w5717 and not w5718;
w5720 <= not w5668 and not w5719;
w5721 <= not w5701 and not w5704;
w5722 <= not w5663 and not w5669;
w5723 <= not w5721 and w5722;
w5724 <= w5721 and not w5722;
w5725 <= not w5723 and not w5724;
w5726 <= not w5612 and not w5615;
w5727 <= not w5574 and not w5580;
w5728 <= not w5726 and w5727;
w5729 <= w5726 and not w5727;
w5730 <= not w5728 and not w5729;
w5731 <= not w5725 and not w5730;
w5732 <= not w5720 and not w5731;
w5733 <= not w5716 and w5732;
w5734 <= not w5716 and not w5720;
w5735 <= w5731 and not w5734;
w5736 <= not w5733 and not w5735;
w5737 <= not w5632 and not w5736;
w5738 <= not w5720 and w5731;
w5739 <= not w5716 and w5738;
w5740 <= not w5731 and not w5734;
w5741 <= not w5739 and not w5740;
w5742 <= w5632 and not w5741;
w5743 <= not w5725 and w5730;
w5744 <= w5725 and not w5730;
w5745 <= not w5743 and not w5744;
w5746 <= not A(193) and A(194);
w5747 <= A(193) and not A(194);
w5748 <= A(195) and not w5747;
w5749 <= not w5746 and w5748;
w5750 <= not w5746 and not w5747;
w5751 <= not A(195) and not w5750;
w5752 <= not w5749 and not w5751;
w5753 <= not A(196) and A(197);
w5754 <= A(196) and not A(197);
w5755 <= A(198) and not w5754;
w5756 <= not w5753 and w5755;
w5757 <= not w5753 and not w5754;
w5758 <= not A(198) and not w5757;
w5759 <= not w5756 and not w5758;
w5760 <= not w5752 and w5759;
w5761 <= w5752 and not w5759;
w5762 <= not w5760 and not w5761;
w5763 <= A(196) and A(197);
w5764 <= A(198) and not w5757;
w5765 <= not w5763 and not w5764;
w5766 <= A(193) and A(194);
w5767 <= A(195) and not w5750;
w5768 <= not w5766 and not w5767;
w5769 <= not w5765 and w5768;
w5770 <= w5765 and not w5768;
w5771 <= not w5769 and not w5770;
w5772 <= not w5752 and not w5759;
w5773 <= not w5771 and w5772;
w5774 <= not w5765 and not w5768;
w5775 <= not w5773 and not w5774;
w5776 <= not w5769 and w5772;
w5777 <= not w5770 and w5776;
w5778 <= not w5771 and not w5772;
w5779 <= not w5777 and not w5778;
w5780 <= not w5775 and not w5779;
w5781 <= not w5762 and not w5780;
w5782 <= not A(187) and A(188);
w5783 <= A(187) and not A(188);
w5784 <= A(189) and not w5783;
w5785 <= not w5782 and w5784;
w5786 <= not w5782 and not w5783;
w5787 <= not A(189) and not w5786;
w5788 <= not w5785 and not w5787;
w5789 <= not A(190) and A(191);
w5790 <= A(190) and not A(191);
w5791 <= A(192) and not w5790;
w5792 <= not w5789 and w5791;
w5793 <= not w5789 and not w5790;
w5794 <= not A(192) and not w5793;
w5795 <= not w5792 and not w5794;
w5796 <= not w5788 and w5795;
w5797 <= w5788 and not w5795;
w5798 <= not w5796 and not w5797;
w5799 <= A(190) and A(191);
w5800 <= A(192) and not w5793;
w5801 <= not w5799 and not w5800;
w5802 <= A(187) and A(188);
w5803 <= A(189) and not w5786;
w5804 <= not w5802 and not w5803;
w5805 <= not w5801 and w5804;
w5806 <= w5801 and not w5804;
w5807 <= not w5805 and not w5806;
w5808 <= not w5788 and not w5795;
w5809 <= not w5807 and w5808;
w5810 <= not w5801 and not w5804;
w5811 <= not w5809 and not w5810;
w5812 <= not w5805 and w5808;
w5813 <= not w5806 and w5812;
w5814 <= not w5807 and not w5808;
w5815 <= not w5813 and not w5814;
w5816 <= not w5811 and not w5815;
w5817 <= not w5798 and not w5816;
w5818 <= not w5781 and w5817;
w5819 <= w5781 and not w5817;
w5820 <= not w5818 and not w5819;
w5821 <= not A(181) and A(182);
w5822 <= A(181) and not A(182);
w5823 <= A(183) and not w5822;
w5824 <= not w5821 and w5823;
w5825 <= not w5821 and not w5822;
w5826 <= not A(183) and not w5825;
w5827 <= not w5824 and not w5826;
w5828 <= not A(184) and A(185);
w5829 <= A(184) and not A(185);
w5830 <= A(186) and not w5829;
w5831 <= not w5828 and w5830;
w5832 <= not w5828 and not w5829;
w5833 <= not A(186) and not w5832;
w5834 <= not w5831 and not w5833;
w5835 <= not w5827 and w5834;
w5836 <= w5827 and not w5834;
w5837 <= not w5835 and not w5836;
w5838 <= A(184) and A(185);
w5839 <= A(186) and not w5832;
w5840 <= not w5838 and not w5839;
w5841 <= A(181) and A(182);
w5842 <= A(183) and not w5825;
w5843 <= not w5841 and not w5842;
w5844 <= not w5840 and w5843;
w5845 <= w5840 and not w5843;
w5846 <= not w5844 and not w5845;
w5847 <= not w5827 and not w5834;
w5848 <= not w5846 and w5847;
w5849 <= not w5840 and not w5843;
w5850 <= not w5848 and not w5849;
w5851 <= not w5844 and w5847;
w5852 <= not w5845 and w5851;
w5853 <= not w5846 and not w5847;
w5854 <= not w5852 and not w5853;
w5855 <= not w5850 and not w5854;
w5856 <= not w5837 and not w5855;
w5857 <= not A(175) and A(176);
w5858 <= A(175) and not A(176);
w5859 <= A(177) and not w5858;
w5860 <= not w5857 and w5859;
w5861 <= not w5857 and not w5858;
w5862 <= not A(177) and not w5861;
w5863 <= not w5860 and not w5862;
w5864 <= not A(178) and A(179);
w5865 <= A(178) and not A(179);
w5866 <= A(180) and not w5865;
w5867 <= not w5864 and w5866;
w5868 <= not w5864 and not w5865;
w5869 <= not A(180) and not w5868;
w5870 <= not w5867 and not w5869;
w5871 <= not w5863 and w5870;
w5872 <= w5863 and not w5870;
w5873 <= not w5871 and not w5872;
w5874 <= A(178) and A(179);
w5875 <= A(180) and not w5868;
w5876 <= not w5874 and not w5875;
w5877 <= A(175) and A(176);
w5878 <= A(177) and not w5861;
w5879 <= not w5877 and not w5878;
w5880 <= not w5876 and w5879;
w5881 <= w5876 and not w5879;
w5882 <= not w5880 and not w5881;
w5883 <= not w5863 and not w5870;
w5884 <= not w5882 and w5883;
w5885 <= not w5876 and not w5879;
w5886 <= not w5884 and not w5885;
w5887 <= not w5880 and w5883;
w5888 <= not w5881 and w5887;
w5889 <= not w5882 and not w5883;
w5890 <= not w5888 and not w5889;
w5891 <= not w5886 and not w5890;
w5892 <= not w5873 and not w5891;
w5893 <= not w5856 and w5892;
w5894 <= w5856 and not w5892;
w5895 <= not w5893 and not w5894;
w5896 <= not w5820 and w5895;
w5897 <= w5820 and not w5895;
w5898 <= not w5896 and not w5897;
w5899 <= not w5745 and not w5898;
w5900 <= not w5742 and w5899;
w5901 <= not w5737 and w5900;
w5902 <= not w5737 and not w5742;
w5903 <= not w5899 and not w5902;
w5904 <= not w5901 and not w5903;
w5905 <= not w5798 and not w5811;
w5906 <= not w5815 and not w5905;
w5907 <= not w5762 and not w5798;
w5908 <= not w5780 and w5907;
w5909 <= not w5816 and w5908;
w5910 <= not w5762 and not w5775;
w5911 <= not w5779 and not w5910;
w5912 <= not w5909 and not w5911;
w5913 <= not w5779 and w5907;
w5914 <= not w5780 and w5913;
w5915 <= not w5816 and not w5910;
w5916 <= w5914 and w5915;
w5917 <= not w5912 and not w5916;
w5918 <= w5906 and not w5917;
w5919 <= not w5909 and w5911;
w5920 <= w5909 and not w5911;
w5921 <= not w5919 and not w5920;
w5922 <= not w5906 and not w5921;
w5923 <= not w5820 and not w5895;
w5924 <= not w5922 and w5923;
w5925 <= not w5918 and w5924;
w5926 <= not w5918 and not w5922;
w5927 <= not w5923 and not w5926;
w5928 <= not w5925 and not w5927;
w5929 <= not w5873 and not w5886;
w5930 <= not w5890 and not w5929;
w5931 <= not w5837 and not w5873;
w5932 <= not w5855 and w5931;
w5933 <= not w5891 and w5932;
w5934 <= not w5837 and not w5850;
w5935 <= not w5854 and not w5934;
w5936 <= not w5933 and w5935;
w5937 <= w5933 and not w5935;
w5938 <= not w5936 and not w5937;
w5939 <= not w5930 and not w5938;
w5940 <= not w5933 and not w5935;
w5941 <= not w5854 and w5931;
w5942 <= not w5855 and w5941;
w5943 <= not w5891 and not w5934;
w5944 <= w5942 and w5943;
w5945 <= not w5940 and not w5944;
w5946 <= w5930 and not w5945;
w5947 <= not w5939 and not w5946;
w5948 <= not w5928 and w5947;
w5949 <= not w5922 and not w5923;
w5950 <= not w5918 and w5949;
w5951 <= w5923 and not w5926;
w5952 <= not w5950 and not w5951;
w5953 <= not w5947 and not w5952;
w5954 <= not w5948 and not w5953;
w5955 <= not w5904 and w5954;
w5956 <= not w5742 and not w5899;
w5957 <= not w5737 and w5956;
w5958 <= w5899 and not w5902;
w5959 <= not w5957 and not w5958;
w5960 <= not w5954 and not w5959;
w5961 <= not w5955 and not w5960;
w5962 <= A(238) and A(239);
w5963 <= A(238) and not A(239);
w5964 <= not A(238) and A(239);
w5965 <= not w5963 and not w5964;
w5966 <= A(240) and not w5965;
w5967 <= not w5962 and not w5966;
w5968 <= A(235) and A(236);
w5969 <= A(235) and not A(236);
w5970 <= not A(235) and A(236);
w5971 <= not w5969 and not w5970;
w5972 <= A(237) and not w5971;
w5973 <= not w5968 and not w5972;
w5974 <= w5967 and not w5973;
w5975 <= not w5967 and w5973;
w5976 <= A(237) and not w5969;
w5977 <= not w5970 and w5976;
w5978 <= not A(237) and not w5971;
w5979 <= not w5977 and not w5978;
w5980 <= A(240) and not w5963;
w5981 <= not w5964 and w5980;
w5982 <= not A(240) and not w5965;
w5983 <= not w5981 and not w5982;
w5984 <= not w5979 and not w5983;
w5985 <= not w5975 and w5984;
w5986 <= not w5974 and w5985;
w5987 <= not w5974 and not w5975;
w5988 <= not w5984 and not w5987;
w5989 <= not w5986 and not w5988;
w5990 <= not w5979 and w5983;
w5991 <= w5979 and not w5983;
w5992 <= not w5990 and not w5991;
w5993 <= w5984 and not w5987;
w5994 <= not w5967 and not w5973;
w5995 <= not w5993 and not w5994;
w5996 <= not w5992 and not w5995;
w5997 <= not w5989 and not w5996;
w5998 <= not w5989 and not w5995;
w5999 <= A(244) and A(245);
w6000 <= A(244) and not A(245);
w6001 <= not A(244) and A(245);
w6002 <= not w6000 and not w6001;
w6003 <= A(246) and not w6002;
w6004 <= not w5999 and not w6003;
w6005 <= A(241) and A(242);
w6006 <= A(241) and not A(242);
w6007 <= not A(241) and A(242);
w6008 <= not w6006 and not w6007;
w6009 <= A(243) and not w6008;
w6010 <= not w6005 and not w6009;
w6011 <= not w6004 and w6010;
w6012 <= w6004 and not w6010;
w6013 <= not w6011 and not w6012;
w6014 <= A(243) and not w6006;
w6015 <= not w6007 and w6014;
w6016 <= not A(243) and not w6008;
w6017 <= not w6015 and not w6016;
w6018 <= A(246) and not w6000;
w6019 <= not w6001 and w6018;
w6020 <= not A(246) and not w6002;
w6021 <= not w6019 and not w6020;
w6022 <= not w6017 and not w6021;
w6023 <= not w6013 and w6022;
w6024 <= not w6004 and not w6010;
w6025 <= not w6023 and not w6024;
w6026 <= not w6011 and w6022;
w6027 <= not w6012 and w6026;
w6028 <= not w6013 and not w6022;
w6029 <= not w6027 and not w6028;
w6030 <= not w6025 and not w6029;
w6031 <= not w6017 and w6021;
w6032 <= w6017 and not w6021;
w6033 <= not w6031 and not w6032;
w6034 <= not w5992 and not w6033;
w6035 <= not w6030 and w6034;
w6036 <= not w5998 and w6035;
w6037 <= not w6025 and not w6033;
w6038 <= not w6029 and not w6037;
w6039 <= not w6036 and not w6038;
w6040 <= not w6029 and w6034;
w6041 <= not w6030 and w6040;
w6042 <= not w5998 and not w6037;
w6043 <= w6041 and w6042;
w6044 <= not w6039 and not w6043;
w6045 <= w5997 and not w6044;
w6046 <= not w6036 and w6038;
w6047 <= w6036 and not w6038;
w6048 <= not w6046 and not w6047;
w6049 <= not w5997 and not w6048;
w6050 <= not w6030 and not w6033;
w6051 <= not w5992 and not w5998;
w6052 <= not w6050 and w6051;
w6053 <= w6050 and not w6051;
w6054 <= not w6052 and not w6053;
w6055 <= not A(229) and A(230);
w6056 <= A(229) and not A(230);
w6057 <= A(231) and not w6056;
w6058 <= not w6055 and w6057;
w6059 <= not w6055 and not w6056;
w6060 <= not A(231) and not w6059;
w6061 <= not w6058 and not w6060;
w6062 <= not A(232) and A(233);
w6063 <= A(232) and not A(233);
w6064 <= A(234) and not w6063;
w6065 <= not w6062 and w6064;
w6066 <= not w6062 and not w6063;
w6067 <= not A(234) and not w6066;
w6068 <= not w6065 and not w6067;
w6069 <= not w6061 and w6068;
w6070 <= w6061 and not w6068;
w6071 <= not w6069 and not w6070;
w6072 <= A(232) and A(233);
w6073 <= A(234) and not w6066;
w6074 <= not w6072 and not w6073;
w6075 <= A(229) and A(230);
w6076 <= A(231) and not w6059;
w6077 <= not w6075 and not w6076;
w6078 <= not w6074 and w6077;
w6079 <= w6074 and not w6077;
w6080 <= not w6078 and not w6079;
w6081 <= not w6061 and not w6068;
w6082 <= not w6080 and w6081;
w6083 <= not w6074 and not w6077;
w6084 <= not w6082 and not w6083;
w6085 <= not w6078 and w6081;
w6086 <= not w6079 and w6085;
w6087 <= not w6080 and not w6081;
w6088 <= not w6086 and not w6087;
w6089 <= not w6084 and not w6088;
w6090 <= not w6071 and not w6089;
w6091 <= not A(223) and A(224);
w6092 <= A(223) and not A(224);
w6093 <= A(225) and not w6092;
w6094 <= not w6091 and w6093;
w6095 <= not w6091 and not w6092;
w6096 <= not A(225) and not w6095;
w6097 <= not w6094 and not w6096;
w6098 <= not A(226) and A(227);
w6099 <= A(226) and not A(227);
w6100 <= A(228) and not w6099;
w6101 <= not w6098 and w6100;
w6102 <= not w6098 and not w6099;
w6103 <= not A(228) and not w6102;
w6104 <= not w6101 and not w6103;
w6105 <= not w6097 and w6104;
w6106 <= w6097 and not w6104;
w6107 <= not w6105 and not w6106;
w6108 <= A(226) and A(227);
w6109 <= A(228) and not w6102;
w6110 <= not w6108 and not w6109;
w6111 <= A(223) and A(224);
w6112 <= A(225) and not w6095;
w6113 <= not w6111 and not w6112;
w6114 <= not w6110 and w6113;
w6115 <= w6110 and not w6113;
w6116 <= not w6114 and not w6115;
w6117 <= not w6097 and not w6104;
w6118 <= not w6116 and w6117;
w6119 <= not w6110 and not w6113;
w6120 <= not w6118 and not w6119;
w6121 <= not w6114 and w6117;
w6122 <= not w6115 and w6121;
w6123 <= not w6116 and not w6117;
w6124 <= not w6122 and not w6123;
w6125 <= not w6120 and not w6124;
w6126 <= not w6107 and not w6125;
w6127 <= not w6090 and w6126;
w6128 <= w6090 and not w6126;
w6129 <= not w6127 and not w6128;
w6130 <= not w6054 and not w6129;
w6131 <= not w6049 and w6130;
w6132 <= not w6045 and w6131;
w6133 <= not w6045 and not w6049;
w6134 <= not w6130 and not w6133;
w6135 <= not w6132 and not w6134;
w6136 <= not w6107 and not w6120;
w6137 <= not w6124 and not w6136;
w6138 <= not w6071 and not w6107;
w6139 <= not w6089 and w6138;
w6140 <= not w6125 and w6139;
w6141 <= not w6071 and not w6084;
w6142 <= not w6088 and not w6141;
w6143 <= not w6140 and w6142;
w6144 <= w6140 and not w6142;
w6145 <= not w6143 and not w6144;
w6146 <= not w6137 and not w6145;
w6147 <= not w6140 and not w6142;
w6148 <= not w6088 and w6138;
w6149 <= not w6089 and w6148;
w6150 <= not w6125 and not w6141;
w6151 <= w6149 and w6150;
w6152 <= not w6147 and not w6151;
w6153 <= w6137 and not w6152;
w6154 <= not w6146 and not w6153;
w6155 <= not w6135 and w6154;
w6156 <= not w6049 and not w6130;
w6157 <= not w6045 and w6156;
w6158 <= w6130 and not w6133;
w6159 <= not w6157 and not w6158;
w6160 <= not w6154 and not w6159;
w6161 <= not w6155 and not w6160;
w6162 <= A(250) and A(251);
w6163 <= A(250) and not A(251);
w6164 <= not A(250) and A(251);
w6165 <= not w6163 and not w6164;
w6166 <= A(252) and not w6165;
w6167 <= not w6162 and not w6166;
w6168 <= A(247) and A(248);
w6169 <= A(247) and not A(248);
w6170 <= not A(247) and A(248);
w6171 <= not w6169 and not w6170;
w6172 <= A(249) and not w6171;
w6173 <= not w6168 and not w6172;
w6174 <= w6167 and not w6173;
w6175 <= not w6167 and w6173;
w6176 <= A(249) and not w6169;
w6177 <= not w6170 and w6176;
w6178 <= not A(249) and not w6171;
w6179 <= not w6177 and not w6178;
w6180 <= A(252) and not w6163;
w6181 <= not w6164 and w6180;
w6182 <= not A(252) and not w6165;
w6183 <= not w6181 and not w6182;
w6184 <= not w6179 and not w6183;
w6185 <= not w6175 and w6184;
w6186 <= not w6174 and w6185;
w6187 <= not w6174 and not w6175;
w6188 <= not w6184 and not w6187;
w6189 <= not w6186 and not w6188;
w6190 <= not w6179 and w6183;
w6191 <= w6179 and not w6183;
w6192 <= not w6190 and not w6191;
w6193 <= w6184 and not w6187;
w6194 <= not w6167 and not w6173;
w6195 <= not w6193 and not w6194;
w6196 <= not w6192 and not w6195;
w6197 <= not w6189 and not w6196;
w6198 <= not w6189 and not w6195;
w6199 <= A(256) and A(257);
w6200 <= A(256) and not A(257);
w6201 <= not A(256) and A(257);
w6202 <= not w6200 and not w6201;
w6203 <= A(258) and not w6202;
w6204 <= not w6199 and not w6203;
w6205 <= A(253) and A(254);
w6206 <= A(253) and not A(254);
w6207 <= not A(253) and A(254);
w6208 <= not w6206 and not w6207;
w6209 <= A(255) and not w6208;
w6210 <= not w6205 and not w6209;
w6211 <= not w6204 and w6210;
w6212 <= w6204 and not w6210;
w6213 <= not w6211 and not w6212;
w6214 <= A(255) and not w6206;
w6215 <= not w6207 and w6214;
w6216 <= not A(255) and not w6208;
w6217 <= not w6215 and not w6216;
w6218 <= A(258) and not w6200;
w6219 <= not w6201 and w6218;
w6220 <= not A(258) and not w6202;
w6221 <= not w6219 and not w6220;
w6222 <= not w6217 and not w6221;
w6223 <= not w6213 and w6222;
w6224 <= not w6204 and not w6210;
w6225 <= not w6223 and not w6224;
w6226 <= not w6211 and w6222;
w6227 <= not w6212 and w6226;
w6228 <= not w6213 and not w6222;
w6229 <= not w6227 and not w6228;
w6230 <= not w6225 and not w6229;
w6231 <= not w6217 and w6221;
w6232 <= w6217 and not w6221;
w6233 <= not w6231 and not w6232;
w6234 <= not w6192 and not w6233;
w6235 <= not w6230 and w6234;
w6236 <= not w6198 and w6235;
w6237 <= not w6225 and not w6233;
w6238 <= not w6229 and not w6237;
w6239 <= not w6236 and w6238;
w6240 <= w6236 and not w6238;
w6241 <= not w6239 and not w6240;
w6242 <= not w6197 and not w6241;
w6243 <= not w6236 and not w6238;
w6244 <= not w6229 and w6234;
w6245 <= not w6230 and w6244;
w6246 <= not w6198 and not w6237;
w6247 <= w6245 and w6246;
w6248 <= not w6243 and not w6247;
w6249 <= w6197 and not w6248;
w6250 <= not w6242 and not w6249;
w6251 <= A(262) and A(263);
w6252 <= A(262) and not A(263);
w6253 <= not A(262) and A(263);
w6254 <= not w6252 and not w6253;
w6255 <= A(264) and not w6254;
w6256 <= not w6251 and not w6255;
w6257 <= A(259) and A(260);
w6258 <= A(259) and not A(260);
w6259 <= not A(259) and A(260);
w6260 <= not w6258 and not w6259;
w6261 <= A(261) and not w6260;
w6262 <= not w6257 and not w6261;
w6263 <= w6256 and not w6262;
w6264 <= not w6256 and w6262;
w6265 <= A(261) and not w6258;
w6266 <= not w6259 and w6265;
w6267 <= not A(261) and not w6260;
w6268 <= not w6266 and not w6267;
w6269 <= A(264) and not w6252;
w6270 <= not w6253 and w6269;
w6271 <= not A(264) and not w6254;
w6272 <= not w6270 and not w6271;
w6273 <= not w6268 and not w6272;
w6274 <= not w6264 and w6273;
w6275 <= not w6263 and w6274;
w6276 <= not w6263 and not w6264;
w6277 <= not w6273 and not w6276;
w6278 <= not w6275 and not w6277;
w6279 <= not w6268 and w6272;
w6280 <= w6268 and not w6272;
w6281 <= not w6279 and not w6280;
w6282 <= w6273 and not w6276;
w6283 <= not w6256 and not w6262;
w6284 <= not w6282 and not w6283;
w6285 <= not w6281 and not w6284;
w6286 <= not w6278 and not w6285;
w6287 <= not w6278 and not w6284;
w6288 <= A(268) and A(269);
w6289 <= A(268) and not A(269);
w6290 <= not A(268) and A(269);
w6291 <= not w6289 and not w6290;
w6292 <= A(270) and not w6291;
w6293 <= not w6288 and not w6292;
w6294 <= A(265) and A(266);
w6295 <= A(265) and not A(266);
w6296 <= not A(265) and A(266);
w6297 <= not w6295 and not w6296;
w6298 <= A(267) and not w6297;
w6299 <= not w6294 and not w6298;
w6300 <= not w6293 and w6299;
w6301 <= w6293 and not w6299;
w6302 <= not w6300 and not w6301;
w6303 <= A(267) and not w6295;
w6304 <= not w6296 and w6303;
w6305 <= not A(267) and not w6297;
w6306 <= not w6304 and not w6305;
w6307 <= A(270) and not w6289;
w6308 <= not w6290 and w6307;
w6309 <= not A(270) and not w6291;
w6310 <= not w6308 and not w6309;
w6311 <= not w6306 and not w6310;
w6312 <= not w6302 and w6311;
w6313 <= not w6293 and not w6299;
w6314 <= not w6312 and not w6313;
w6315 <= not w6300 and w6311;
w6316 <= not w6301 and w6315;
w6317 <= not w6302 and not w6311;
w6318 <= not w6316 and not w6317;
w6319 <= not w6314 and not w6318;
w6320 <= not w6306 and w6310;
w6321 <= w6306 and not w6310;
w6322 <= not w6320 and not w6321;
w6323 <= not w6281 and not w6322;
w6324 <= not w6319 and w6323;
w6325 <= not w6287 and w6324;
w6326 <= not w6314 and not w6322;
w6327 <= not w6318 and not w6326;
w6328 <= not w6325 and not w6327;
w6329 <= not w6318 and w6323;
w6330 <= not w6319 and w6329;
w6331 <= not w6287 and not w6326;
w6332 <= w6330 and w6331;
w6333 <= not w6328 and not w6332;
w6334 <= w6286 and not w6333;
w6335 <= not w6325 and w6327;
w6336 <= w6325 and not w6327;
w6337 <= not w6335 and not w6336;
w6338 <= not w6286 and not w6337;
w6339 <= not w6319 and not w6322;
w6340 <= not w6281 and not w6287;
w6341 <= not w6339 and w6340;
w6342 <= w6339 and not w6340;
w6343 <= not w6341 and not w6342;
w6344 <= not w6230 and not w6233;
w6345 <= not w6192 and not w6198;
w6346 <= not w6344 and w6345;
w6347 <= w6344 and not w6345;
w6348 <= not w6346 and not w6347;
w6349 <= not w6343 and not w6348;
w6350 <= not w6338 and not w6349;
w6351 <= not w6334 and w6350;
w6352 <= not w6334 and not w6338;
w6353 <= w6349 and not w6352;
w6354 <= not w6351 and not w6353;
w6355 <= not w6250 and not w6354;
w6356 <= not w6338 and w6349;
w6357 <= not w6334 and w6356;
w6358 <= not w6349 and not w6352;
w6359 <= not w6357 and not w6358;
w6360 <= w6250 and not w6359;
w6361 <= not w6343 and w6348;
w6362 <= w6343 and not w6348;
w6363 <= not w6361 and not w6362;
w6364 <= not w6054 and w6129;
w6365 <= w6054 and not w6129;
w6366 <= not w6364 and not w6365;
w6367 <= not w6363 and not w6366;
w6368 <= not w6360 and not w6367;
w6369 <= not w6355 and w6368;
w6370 <= not w6355 and not w6360;
w6371 <= w6367 and not w6370;
w6372 <= not w6369 and not w6371;
w6373 <= not w6161 and not w6372;
w6374 <= not w6360 and w6367;
w6375 <= not w6355 and w6374;
w6376 <= not w6367 and not w6370;
w6377 <= not w6375 and not w6376;
w6378 <= w6161 and not w6377;
w6379 <= not w6363 and w6366;
w6380 <= w6363 and not w6366;
w6381 <= not w6379 and not w6380;
w6382 <= not w5745 and w5898;
w6383 <= w5745 and not w5898;
w6384 <= not w6382 and not w6383;
w6385 <= not w6381 and not w6384;
w6386 <= not w6378 and not w6385;
w6387 <= not w6373 and w6386;
w6388 <= not w6373 and not w6378;
w6389 <= w6385 and not w6388;
w6390 <= not w6387 and not w6389;
w6391 <= not w5961 and not w6390;
w6392 <= not w6378 and w6385;
w6393 <= not w6373 and w6392;
w6394 <= not w6385 and not w6388;
w6395 <= not w6393 and not w6394;
w6396 <= w5961 and not w6395;
w6397 <= not w6381 and w6384;
w6398 <= w6381 and not w6384;
w6399 <= not w6397 and not w6398;
w6400 <= not A(169) and A(170);
w6401 <= A(169) and not A(170);
w6402 <= A(171) and not w6401;
w6403 <= not w6400 and w6402;
w6404 <= not w6400 and not w6401;
w6405 <= not A(171) and not w6404;
w6406 <= not w6403 and not w6405;
w6407 <= not A(172) and A(173);
w6408 <= A(172) and not A(173);
w6409 <= A(174) and not w6408;
w6410 <= not w6407 and w6409;
w6411 <= not w6407 and not w6408;
w6412 <= not A(174) and not w6411;
w6413 <= not w6410 and not w6412;
w6414 <= not w6406 and w6413;
w6415 <= w6406 and not w6413;
w6416 <= not w6414 and not w6415;
w6417 <= A(172) and A(173);
w6418 <= A(174) and not w6411;
w6419 <= not w6417 and not w6418;
w6420 <= A(169) and A(170);
w6421 <= A(171) and not w6404;
w6422 <= not w6420 and not w6421;
w6423 <= not w6419 and w6422;
w6424 <= w6419 and not w6422;
w6425 <= not w6423 and not w6424;
w6426 <= not w6406 and not w6413;
w6427 <= not w6425 and w6426;
w6428 <= not w6419 and not w6422;
w6429 <= not w6427 and not w6428;
w6430 <= not w6423 and w6426;
w6431 <= not w6424 and w6430;
w6432 <= not w6425 and not w6426;
w6433 <= not w6431 and not w6432;
w6434 <= not w6429 and not w6433;
w6435 <= not w6416 and not w6434;
w6436 <= not A(163) and A(164);
w6437 <= A(163) and not A(164);
w6438 <= A(165) and not w6437;
w6439 <= not w6436 and w6438;
w6440 <= not w6436 and not w6437;
w6441 <= not A(165) and not w6440;
w6442 <= not w6439 and not w6441;
w6443 <= not A(166) and A(167);
w6444 <= A(166) and not A(167);
w6445 <= A(168) and not w6444;
w6446 <= not w6443 and w6445;
w6447 <= not w6443 and not w6444;
w6448 <= not A(168) and not w6447;
w6449 <= not w6446 and not w6448;
w6450 <= not w6442 and w6449;
w6451 <= w6442 and not w6449;
w6452 <= not w6450 and not w6451;
w6453 <= A(166) and A(167);
w6454 <= A(168) and not w6447;
w6455 <= not w6453 and not w6454;
w6456 <= A(163) and A(164);
w6457 <= A(165) and not w6440;
w6458 <= not w6456 and not w6457;
w6459 <= not w6455 and w6458;
w6460 <= w6455 and not w6458;
w6461 <= not w6459 and not w6460;
w6462 <= not w6442 and not w6449;
w6463 <= not w6461 and w6462;
w6464 <= not w6455 and not w6458;
w6465 <= not w6463 and not w6464;
w6466 <= not w6459 and w6462;
w6467 <= not w6460 and w6466;
w6468 <= not w6461 and not w6462;
w6469 <= not w6467 and not w6468;
w6470 <= not w6465 and not w6469;
w6471 <= not w6452 and not w6470;
w6472 <= not w6435 and w6471;
w6473 <= w6435 and not w6471;
w6474 <= not w6472 and not w6473;
w6475 <= not A(157) and A(158);
w6476 <= A(157) and not A(158);
w6477 <= A(159) and not w6476;
w6478 <= not w6475 and w6477;
w6479 <= not w6475 and not w6476;
w6480 <= not A(159) and not w6479;
w6481 <= not w6478 and not w6480;
w6482 <= not A(160) and A(161);
w6483 <= A(160) and not A(161);
w6484 <= A(162) and not w6483;
w6485 <= not w6482 and w6484;
w6486 <= not w6482 and not w6483;
w6487 <= not A(162) and not w6486;
w6488 <= not w6485 and not w6487;
w6489 <= not w6481 and w6488;
w6490 <= w6481 and not w6488;
w6491 <= not w6489 and not w6490;
w6492 <= A(160) and A(161);
w6493 <= A(162) and not w6486;
w6494 <= not w6492 and not w6493;
w6495 <= A(157) and A(158);
w6496 <= A(159) and not w6479;
w6497 <= not w6495 and not w6496;
w6498 <= not w6494 and w6497;
w6499 <= w6494 and not w6497;
w6500 <= not w6498 and not w6499;
w6501 <= not w6481 and not w6488;
w6502 <= not w6500 and w6501;
w6503 <= not w6494 and not w6497;
w6504 <= not w6502 and not w6503;
w6505 <= not w6498 and w6501;
w6506 <= not w6499 and w6505;
w6507 <= not w6500 and not w6501;
w6508 <= not w6506 and not w6507;
w6509 <= not w6504 and not w6508;
w6510 <= not w6491 and not w6509;
w6511 <= not A(151) and A(152);
w6512 <= A(151) and not A(152);
w6513 <= A(153) and not w6512;
w6514 <= not w6511 and w6513;
w6515 <= not w6511 and not w6512;
w6516 <= not A(153) and not w6515;
w6517 <= not w6514 and not w6516;
w6518 <= not A(154) and A(155);
w6519 <= A(154) and not A(155);
w6520 <= A(156) and not w6519;
w6521 <= not w6518 and w6520;
w6522 <= not w6518 and not w6519;
w6523 <= not A(156) and not w6522;
w6524 <= not w6521 and not w6523;
w6525 <= not w6517 and w6524;
w6526 <= w6517 and not w6524;
w6527 <= not w6525 and not w6526;
w6528 <= A(154) and A(155);
w6529 <= A(156) and not w6522;
w6530 <= not w6528 and not w6529;
w6531 <= A(151) and A(152);
w6532 <= A(153) and not w6515;
w6533 <= not w6531 and not w6532;
w6534 <= not w6530 and w6533;
w6535 <= w6530 and not w6533;
w6536 <= not w6534 and not w6535;
w6537 <= not w6517 and not w6524;
w6538 <= not w6536 and w6537;
w6539 <= not w6530 and not w6533;
w6540 <= not w6538 and not w6539;
w6541 <= not w6534 and w6537;
w6542 <= not w6535 and w6541;
w6543 <= not w6536 and not w6537;
w6544 <= not w6542 and not w6543;
w6545 <= not w6540 and not w6544;
w6546 <= not w6527 and not w6545;
w6547 <= not w6510 and w6546;
w6548 <= w6510 and not w6546;
w6549 <= not w6547 and not w6548;
w6550 <= not w6474 and w6549;
w6551 <= w6474 and not w6549;
w6552 <= not w6550 and not w6551;
w6553 <= not A(145) and A(146);
w6554 <= A(145) and not A(146);
w6555 <= A(147) and not w6554;
w6556 <= not w6553 and w6555;
w6557 <= not w6553 and not w6554;
w6558 <= not A(147) and not w6557;
w6559 <= not w6556 and not w6558;
w6560 <= not A(148) and A(149);
w6561 <= A(148) and not A(149);
w6562 <= A(150) and not w6561;
w6563 <= not w6560 and w6562;
w6564 <= not w6560 and not w6561;
w6565 <= not A(150) and not w6564;
w6566 <= not w6563 and not w6565;
w6567 <= not w6559 and w6566;
w6568 <= w6559 and not w6566;
w6569 <= not w6567 and not w6568;
w6570 <= A(148) and A(149);
w6571 <= A(150) and not w6564;
w6572 <= not w6570 and not w6571;
w6573 <= A(145) and A(146);
w6574 <= A(147) and not w6557;
w6575 <= not w6573 and not w6574;
w6576 <= not w6572 and w6575;
w6577 <= w6572 and not w6575;
w6578 <= not w6576 and not w6577;
w6579 <= not w6559 and not w6566;
w6580 <= not w6578 and w6579;
w6581 <= not w6572 and not w6575;
w6582 <= not w6580 and not w6581;
w6583 <= not w6576 and w6579;
w6584 <= not w6577 and w6583;
w6585 <= not w6578 and not w6579;
w6586 <= not w6584 and not w6585;
w6587 <= not w6582 and not w6586;
w6588 <= not w6569 and not w6587;
w6589 <= not A(139) and A(140);
w6590 <= A(139) and not A(140);
w6591 <= A(141) and not w6590;
w6592 <= not w6589 and w6591;
w6593 <= not w6589 and not w6590;
w6594 <= not A(141) and not w6593;
w6595 <= not w6592 and not w6594;
w6596 <= not A(142) and A(143);
w6597 <= A(142) and not A(143);
w6598 <= A(144) and not w6597;
w6599 <= not w6596 and w6598;
w6600 <= not w6596 and not w6597;
w6601 <= not A(144) and not w6600;
w6602 <= not w6599 and not w6601;
w6603 <= not w6595 and w6602;
w6604 <= w6595 and not w6602;
w6605 <= not w6603 and not w6604;
w6606 <= A(142) and A(143);
w6607 <= A(144) and not w6600;
w6608 <= not w6606 and not w6607;
w6609 <= A(139) and A(140);
w6610 <= A(141) and not w6593;
w6611 <= not w6609 and not w6610;
w6612 <= not w6608 and w6611;
w6613 <= w6608 and not w6611;
w6614 <= not w6612 and not w6613;
w6615 <= not w6595 and not w6602;
w6616 <= not w6614 and w6615;
w6617 <= not w6608 and not w6611;
w6618 <= not w6616 and not w6617;
w6619 <= not w6612 and w6615;
w6620 <= not w6613 and w6619;
w6621 <= not w6614 and not w6615;
w6622 <= not w6620 and not w6621;
w6623 <= not w6618 and not w6622;
w6624 <= not w6605 and not w6623;
w6625 <= not w6588 and w6624;
w6626 <= w6588 and not w6624;
w6627 <= not w6625 and not w6626;
w6628 <= not A(133) and A(134);
w6629 <= A(133) and not A(134);
w6630 <= A(135) and not w6629;
w6631 <= not w6628 and w6630;
w6632 <= not w6628 and not w6629;
w6633 <= not A(135) and not w6632;
w6634 <= not w6631 and not w6633;
w6635 <= not A(136) and A(137);
w6636 <= A(136) and not A(137);
w6637 <= A(138) and not w6636;
w6638 <= not w6635 and w6637;
w6639 <= not w6635 and not w6636;
w6640 <= not A(138) and not w6639;
w6641 <= not w6638 and not w6640;
w6642 <= not w6634 and w6641;
w6643 <= w6634 and not w6641;
w6644 <= not w6642 and not w6643;
w6645 <= A(136) and A(137);
w6646 <= A(138) and not w6639;
w6647 <= not w6645 and not w6646;
w6648 <= A(133) and A(134);
w6649 <= A(135) and not w6632;
w6650 <= not w6648 and not w6649;
w6651 <= not w6647 and w6650;
w6652 <= w6647 and not w6650;
w6653 <= not w6651 and not w6652;
w6654 <= not w6634 and not w6641;
w6655 <= not w6653 and w6654;
w6656 <= not w6647 and not w6650;
w6657 <= not w6655 and not w6656;
w6658 <= not w6651 and w6654;
w6659 <= not w6652 and w6658;
w6660 <= not w6653 and not w6654;
w6661 <= not w6659 and not w6660;
w6662 <= not w6657 and not w6661;
w6663 <= not w6644 and not w6662;
w6664 <= not A(127) and A(128);
w6665 <= A(127) and not A(128);
w6666 <= A(129) and not w6665;
w6667 <= not w6664 and w6666;
w6668 <= not w6664 and not w6665;
w6669 <= not A(129) and not w6668;
w6670 <= not w6667 and not w6669;
w6671 <= not A(130) and A(131);
w6672 <= A(130) and not A(131);
w6673 <= A(132) and not w6672;
w6674 <= not w6671 and w6673;
w6675 <= not w6671 and not w6672;
w6676 <= not A(132) and not w6675;
w6677 <= not w6674 and not w6676;
w6678 <= not w6670 and w6677;
w6679 <= w6670 and not w6677;
w6680 <= not w6678 and not w6679;
w6681 <= A(130) and A(131);
w6682 <= A(132) and not w6675;
w6683 <= not w6681 and not w6682;
w6684 <= A(127) and A(128);
w6685 <= A(129) and not w6668;
w6686 <= not w6684 and not w6685;
w6687 <= not w6683 and w6686;
w6688 <= w6683 and not w6686;
w6689 <= not w6687 and not w6688;
w6690 <= not w6670 and not w6677;
w6691 <= not w6689 and w6690;
w6692 <= not w6683 and not w6686;
w6693 <= not w6691 and not w6692;
w6694 <= not w6687 and w6690;
w6695 <= not w6688 and w6694;
w6696 <= not w6689 and not w6690;
w6697 <= not w6695 and not w6696;
w6698 <= not w6693 and not w6697;
w6699 <= not w6680 and not w6698;
w6700 <= not w6663 and w6699;
w6701 <= w6663 and not w6699;
w6702 <= not w6700 and not w6701;
w6703 <= not w6627 and w6702;
w6704 <= w6627 and not w6702;
w6705 <= not w6703 and not w6704;
w6706 <= not w6552 and w6705;
w6707 <= w6552 and not w6705;
w6708 <= not w6706 and not w6707;
w6709 <= not A(121) and A(122);
w6710 <= A(121) and not A(122);
w6711 <= A(123) and not w6710;
w6712 <= not w6709 and w6711;
w6713 <= not w6709 and not w6710;
w6714 <= not A(123) and not w6713;
w6715 <= not w6712 and not w6714;
w6716 <= not A(124) and A(125);
w6717 <= A(124) and not A(125);
w6718 <= A(126) and not w6717;
w6719 <= not w6716 and w6718;
w6720 <= not w6716 and not w6717;
w6721 <= not A(126) and not w6720;
w6722 <= not w6719 and not w6721;
w6723 <= not w6715 and w6722;
w6724 <= w6715 and not w6722;
w6725 <= not w6723 and not w6724;
w6726 <= A(124) and A(125);
w6727 <= A(126) and not w6720;
w6728 <= not w6726 and not w6727;
w6729 <= A(121) and A(122);
w6730 <= A(123) and not w6713;
w6731 <= not w6729 and not w6730;
w6732 <= not w6728 and w6731;
w6733 <= w6728 and not w6731;
w6734 <= not w6732 and not w6733;
w6735 <= not w6715 and not w6722;
w6736 <= not w6734 and w6735;
w6737 <= not w6728 and not w6731;
w6738 <= not w6736 and not w6737;
w6739 <= not w6732 and w6735;
w6740 <= not w6733 and w6739;
w6741 <= not w6734 and not w6735;
w6742 <= not w6740 and not w6741;
w6743 <= not w6738 and not w6742;
w6744 <= not w6725 and not w6743;
w6745 <= not A(115) and A(116);
w6746 <= A(115) and not A(116);
w6747 <= A(117) and not w6746;
w6748 <= not w6745 and w6747;
w6749 <= not w6745 and not w6746;
w6750 <= not A(117) and not w6749;
w6751 <= not w6748 and not w6750;
w6752 <= not A(118) and A(119);
w6753 <= A(118) and not A(119);
w6754 <= A(120) and not w6753;
w6755 <= not w6752 and w6754;
w6756 <= not w6752 and not w6753;
w6757 <= not A(120) and not w6756;
w6758 <= not w6755 and not w6757;
w6759 <= not w6751 and w6758;
w6760 <= w6751 and not w6758;
w6761 <= not w6759 and not w6760;
w6762 <= A(118) and A(119);
w6763 <= A(120) and not w6756;
w6764 <= not w6762 and not w6763;
w6765 <= A(115) and A(116);
w6766 <= A(117) and not w6749;
w6767 <= not w6765 and not w6766;
w6768 <= not w6764 and w6767;
w6769 <= w6764 and not w6767;
w6770 <= not w6768 and not w6769;
w6771 <= not w6751 and not w6758;
w6772 <= not w6770 and w6771;
w6773 <= not w6764 and not w6767;
w6774 <= not w6772 and not w6773;
w6775 <= not w6768 and w6771;
w6776 <= not w6769 and w6775;
w6777 <= not w6770 and not w6771;
w6778 <= not w6776 and not w6777;
w6779 <= not w6774 and not w6778;
w6780 <= not w6761 and not w6779;
w6781 <= not w6744 and w6780;
w6782 <= w6744 and not w6780;
w6783 <= not w6781 and not w6782;
w6784 <= not A(109) and A(110);
w6785 <= A(109) and not A(110);
w6786 <= A(111) and not w6785;
w6787 <= not w6784 and w6786;
w6788 <= not w6784 and not w6785;
w6789 <= not A(111) and not w6788;
w6790 <= not w6787 and not w6789;
w6791 <= not A(112) and A(113);
w6792 <= A(112) and not A(113);
w6793 <= A(114) and not w6792;
w6794 <= not w6791 and w6793;
w6795 <= not w6791 and not w6792;
w6796 <= not A(114) and not w6795;
w6797 <= not w6794 and not w6796;
w6798 <= not w6790 and w6797;
w6799 <= w6790 and not w6797;
w6800 <= not w6798 and not w6799;
w6801 <= A(112) and A(113);
w6802 <= A(114) and not w6795;
w6803 <= not w6801 and not w6802;
w6804 <= A(109) and A(110);
w6805 <= A(111) and not w6788;
w6806 <= not w6804 and not w6805;
w6807 <= not w6803 and w6806;
w6808 <= w6803 and not w6806;
w6809 <= not w6807 and not w6808;
w6810 <= not w6790 and not w6797;
w6811 <= not w6809 and w6810;
w6812 <= not w6803 and not w6806;
w6813 <= not w6811 and not w6812;
w6814 <= not w6807 and w6810;
w6815 <= not w6808 and w6814;
w6816 <= not w6809 and not w6810;
w6817 <= not w6815 and not w6816;
w6818 <= not w6813 and not w6817;
w6819 <= not w6800 and not w6818;
w6820 <= not A(103) and A(104);
w6821 <= A(103) and not A(104);
w6822 <= A(105) and not w6821;
w6823 <= not w6820 and w6822;
w6824 <= not w6820 and not w6821;
w6825 <= not A(105) and not w6824;
w6826 <= not w6823 and not w6825;
w6827 <= not A(106) and A(107);
w6828 <= A(106) and not A(107);
w6829 <= A(108) and not w6828;
w6830 <= not w6827 and w6829;
w6831 <= not w6827 and not w6828;
w6832 <= not A(108) and not w6831;
w6833 <= not w6830 and not w6832;
w6834 <= not w6826 and w6833;
w6835 <= w6826 and not w6833;
w6836 <= not w6834 and not w6835;
w6837 <= A(106) and A(107);
w6838 <= A(108) and not w6831;
w6839 <= not w6837 and not w6838;
w6840 <= A(103) and A(104);
w6841 <= A(105) and not w6824;
w6842 <= not w6840 and not w6841;
w6843 <= not w6839 and w6842;
w6844 <= w6839 and not w6842;
w6845 <= not w6843 and not w6844;
w6846 <= not w6826 and not w6833;
w6847 <= not w6845 and w6846;
w6848 <= not w6839 and not w6842;
w6849 <= not w6847 and not w6848;
w6850 <= not w6843 and w6846;
w6851 <= not w6844 and w6850;
w6852 <= not w6845 and not w6846;
w6853 <= not w6851 and not w6852;
w6854 <= not w6849 and not w6853;
w6855 <= not w6836 and not w6854;
w6856 <= not w6819 and w6855;
w6857 <= w6819 and not w6855;
w6858 <= not w6856 and not w6857;
w6859 <= not w6783 and w6858;
w6860 <= w6783 and not w6858;
w6861 <= not w6859 and not w6860;
w6862 <= not A(97) and A(98);
w6863 <= A(97) and not A(98);
w6864 <= A(99) and not w6863;
w6865 <= not w6862 and w6864;
w6866 <= not w6862 and not w6863;
w6867 <= not A(99) and not w6866;
w6868 <= not w6865 and not w6867;
w6869 <= not A(100) and A(101);
w6870 <= A(100) and not A(101);
w6871 <= A(102) and not w6870;
w6872 <= not w6869 and w6871;
w6873 <= not w6869 and not w6870;
w6874 <= not A(102) and not w6873;
w6875 <= not w6872 and not w6874;
w6876 <= not w6868 and w6875;
w6877 <= w6868 and not w6875;
w6878 <= not w6876 and not w6877;
w6879 <= A(100) and A(101);
w6880 <= A(102) and not w6873;
w6881 <= not w6879 and not w6880;
w6882 <= A(97) and A(98);
w6883 <= A(99) and not w6866;
w6884 <= not w6882 and not w6883;
w6885 <= not w6881 and w6884;
w6886 <= w6881 and not w6884;
w6887 <= not w6885 and not w6886;
w6888 <= not w6868 and not w6875;
w6889 <= not w6887 and w6888;
w6890 <= not w6881 and not w6884;
w6891 <= not w6889 and not w6890;
w6892 <= not w6885 and w6888;
w6893 <= not w6886 and w6892;
w6894 <= not w6887 and not w6888;
w6895 <= not w6893 and not w6894;
w6896 <= not w6891 and not w6895;
w6897 <= not w6878 and not w6896;
w6898 <= not A(91) and A(92);
w6899 <= A(91) and not A(92);
w6900 <= A(93) and not w6899;
w6901 <= not w6898 and w6900;
w6902 <= not w6898 and not w6899;
w6903 <= not A(93) and not w6902;
w6904 <= not w6901 and not w6903;
w6905 <= not A(94) and A(95);
w6906 <= A(94) and not A(95);
w6907 <= A(96) and not w6906;
w6908 <= not w6905 and w6907;
w6909 <= not w6905 and not w6906;
w6910 <= not A(96) and not w6909;
w6911 <= not w6908 and not w6910;
w6912 <= not w6904 and w6911;
w6913 <= w6904 and not w6911;
w6914 <= not w6912 and not w6913;
w6915 <= A(94) and A(95);
w6916 <= A(96) and not w6909;
w6917 <= not w6915 and not w6916;
w6918 <= A(91) and A(92);
w6919 <= A(93) and not w6902;
w6920 <= not w6918 and not w6919;
w6921 <= not w6917 and w6920;
w6922 <= w6917 and not w6920;
w6923 <= not w6921 and not w6922;
w6924 <= not w6904 and not w6911;
w6925 <= not w6923 and w6924;
w6926 <= not w6917 and not w6920;
w6927 <= not w6925 and not w6926;
w6928 <= not w6921 and w6924;
w6929 <= not w6922 and w6928;
w6930 <= not w6923 and not w6924;
w6931 <= not w6929 and not w6930;
w6932 <= not w6927 and not w6931;
w6933 <= not w6914 and not w6932;
w6934 <= not w6897 and w6933;
w6935 <= w6897 and not w6933;
w6936 <= not w6934 and not w6935;
w6937 <= not A(85) and A(86);
w6938 <= A(85) and not A(86);
w6939 <= A(87) and not w6938;
w6940 <= not w6937 and w6939;
w6941 <= not w6937 and not w6938;
w6942 <= not A(87) and not w6941;
w6943 <= not w6940 and not w6942;
w6944 <= not A(88) and A(89);
w6945 <= A(88) and not A(89);
w6946 <= A(90) and not w6945;
w6947 <= not w6944 and w6946;
w6948 <= not w6944 and not w6945;
w6949 <= not A(90) and not w6948;
w6950 <= not w6947 and not w6949;
w6951 <= not w6943 and w6950;
w6952 <= w6943 and not w6950;
w6953 <= not w6951 and not w6952;
w6954 <= A(88) and A(89);
w6955 <= A(90) and not w6948;
w6956 <= not w6954 and not w6955;
w6957 <= A(85) and A(86);
w6958 <= A(87) and not w6941;
w6959 <= not w6957 and not w6958;
w6960 <= not w6956 and w6959;
w6961 <= w6956 and not w6959;
w6962 <= not w6960 and not w6961;
w6963 <= not w6943 and not w6950;
w6964 <= not w6962 and w6963;
w6965 <= not w6956 and not w6959;
w6966 <= not w6964 and not w6965;
w6967 <= not w6960 and w6963;
w6968 <= not w6961 and w6967;
w6969 <= not w6962 and not w6963;
w6970 <= not w6968 and not w6969;
w6971 <= not w6966 and not w6970;
w6972 <= not w6953 and not w6971;
w6973 <= not A(79) and A(80);
w6974 <= A(79) and not A(80);
w6975 <= A(81) and not w6974;
w6976 <= not w6973 and w6975;
w6977 <= not w6973 and not w6974;
w6978 <= not A(81) and not w6977;
w6979 <= not w6976 and not w6978;
w6980 <= not A(82) and A(83);
w6981 <= A(82) and not A(83);
w6982 <= A(84) and not w6981;
w6983 <= not w6980 and w6982;
w6984 <= not w6980 and not w6981;
w6985 <= not A(84) and not w6984;
w6986 <= not w6983 and not w6985;
w6987 <= not w6979 and w6986;
w6988 <= w6979 and not w6986;
w6989 <= not w6987 and not w6988;
w6990 <= A(82) and A(83);
w6991 <= A(84) and not w6984;
w6992 <= not w6990 and not w6991;
w6993 <= A(79) and A(80);
w6994 <= A(81) and not w6977;
w6995 <= not w6993 and not w6994;
w6996 <= not w6992 and w6995;
w6997 <= w6992 and not w6995;
w6998 <= not w6996 and not w6997;
w6999 <= not w6979 and not w6986;
w7000 <= not w6998 and w6999;
w7001 <= not w6992 and not w6995;
w7002 <= not w7000 and not w7001;
w7003 <= not w6996 and w6999;
w7004 <= not w6997 and w7003;
w7005 <= not w6998 and not w6999;
w7006 <= not w7004 and not w7005;
w7007 <= not w7002 and not w7006;
w7008 <= not w6989 and not w7007;
w7009 <= not w6972 and w7008;
w7010 <= w6972 and not w7008;
w7011 <= not w7009 and not w7010;
w7012 <= not w6936 and w7011;
w7013 <= w6936 and not w7011;
w7014 <= not w7012 and not w7013;
w7015 <= not w6861 and w7014;
w7016 <= w6861 and not w7014;
w7017 <= not w7015 and not w7016;
w7018 <= not w6708 and w7017;
w7019 <= w6708 and not w7017;
w7020 <= not w7018 and not w7019;
w7021 <= not w6399 and not w7020;
w7022 <= not w6396 and w7021;
w7023 <= not w6391 and w7022;
w7024 <= not w6391 and not w6396;
w7025 <= not w7021 and not w7024;
w7026 <= not w7023 and not w7025;
w7027 <= not w6605 and not w6618;
w7028 <= not w6622 and not w7027;
w7029 <= not w6569 and not w6605;
w7030 <= not w6587 and w7029;
w7031 <= not w6623 and w7030;
w7032 <= not w6569 and not w6582;
w7033 <= not w6586 and not w7032;
w7034 <= not w7031 and not w7033;
w7035 <= not w6586 and w7029;
w7036 <= not w6587 and w7035;
w7037 <= not w6623 and not w7032;
w7038 <= w7036 and w7037;
w7039 <= not w7034 and not w7038;
w7040 <= w7028 and not w7039;
w7041 <= not w7031 and w7033;
w7042 <= w7031 and not w7033;
w7043 <= not w7041 and not w7042;
w7044 <= not w7028 and not w7043;
w7045 <= not w6627 and not w6702;
w7046 <= not w7044 and w7045;
w7047 <= not w7040 and w7046;
w7048 <= not w7040 and not w7044;
w7049 <= not w7045 and not w7048;
w7050 <= not w7047 and not w7049;
w7051 <= not w6680 and not w6693;
w7052 <= not w6697 and not w7051;
w7053 <= not w6644 and not w6680;
w7054 <= not w6662 and w7053;
w7055 <= not w6698 and w7054;
w7056 <= not w6644 and not w6657;
w7057 <= not w6661 and not w7056;
w7058 <= not w7055 and w7057;
w7059 <= w7055 and not w7057;
w7060 <= not w7058 and not w7059;
w7061 <= not w7052 and not w7060;
w7062 <= not w7055 and not w7057;
w7063 <= not w6661 and w7053;
w7064 <= not w6662 and w7063;
w7065 <= not w6698 and not w7056;
w7066 <= w7064 and w7065;
w7067 <= not w7062 and not w7066;
w7068 <= w7052 and not w7067;
w7069 <= not w7061 and not w7068;
w7070 <= not w7050 and w7069;
w7071 <= not w7044 and not w7045;
w7072 <= not w7040 and w7071;
w7073 <= w7045 and not w7048;
w7074 <= not w7072 and not w7073;
w7075 <= not w7069 and not w7074;
w7076 <= not w7070 and not w7075;
w7077 <= not w6527 and not w6540;
w7078 <= not w6544 and not w7077;
w7079 <= not w6491 and not w6527;
w7080 <= not w6509 and w7079;
w7081 <= not w6545 and w7080;
w7082 <= not w6491 and not w6504;
w7083 <= not w6508 and not w7082;
w7084 <= not w7081 and w7083;
w7085 <= w7081 and not w7083;
w7086 <= not w7084 and not w7085;
w7087 <= not w7078 and not w7086;
w7088 <= not w7081 and not w7083;
w7089 <= not w6508 and w7079;
w7090 <= not w6509 and w7089;
w7091 <= not w6545 and not w7082;
w7092 <= w7090 and w7091;
w7093 <= not w7088 and not w7092;
w7094 <= w7078 and not w7093;
w7095 <= not w7087 and not w7094;
w7096 <= not w6452 and not w6465;
w7097 <= not w6469 and not w7096;
w7098 <= not w6416 and not w6452;
w7099 <= not w6434 and w7098;
w7100 <= not w6470 and w7099;
w7101 <= not w6416 and not w6429;
w7102 <= not w6433 and not w7101;
w7103 <= not w7100 and not w7102;
w7104 <= not w6433 and w7098;
w7105 <= not w6434 and w7104;
w7106 <= not w6470 and not w7101;
w7107 <= w7105 and w7106;
w7108 <= not w7103 and not w7107;
w7109 <= w7097 and not w7108;
w7110 <= not w7100 and w7102;
w7111 <= w7100 and not w7102;
w7112 <= not w7110 and not w7111;
w7113 <= not w7097 and not w7112;
w7114 <= not w6474 and not w6549;
w7115 <= not w7113 and not w7114;
w7116 <= not w7109 and w7115;
w7117 <= not w7109 and not w7113;
w7118 <= w7114 and not w7117;
w7119 <= not w7116 and not w7118;
w7120 <= not w7095 and not w7119;
w7121 <= not w7113 and w7114;
w7122 <= not w7109 and w7121;
w7123 <= not w7114 and not w7117;
w7124 <= not w7122 and not w7123;
w7125 <= w7095 and not w7124;
w7126 <= not w6552 and not w6705;
w7127 <= not w7125 and not w7126;
w7128 <= not w7120 and w7127;
w7129 <= not w7120 and not w7125;
w7130 <= w7126 and not w7129;
w7131 <= not w7128 and not w7130;
w7132 <= not w7076 and not w7131;
w7133 <= not w7125 and w7126;
w7134 <= not w7120 and w7133;
w7135 <= not w7126 and not w7129;
w7136 <= not w7134 and not w7135;
w7137 <= w7076 and not w7136;
w7138 <= not w6708 and not w7017;
w7139 <= not w7137 and w7138;
w7140 <= not w7132 and w7139;
w7141 <= not w7132 and not w7137;
w7142 <= not w7138 and not w7141;
w7143 <= not w7140 and not w7142;
w7144 <= not w6836 and not w6849;
w7145 <= not w6853 and not w7144;
w7146 <= not w6800 and not w6836;
w7147 <= not w6818 and w7146;
w7148 <= not w6854 and w7147;
w7149 <= not w6800 and not w6813;
w7150 <= not w6817 and not w7149;
w7151 <= not w7148 and w7150;
w7152 <= w7148 and not w7150;
w7153 <= not w7151 and not w7152;
w7154 <= not w7145 and not w7153;
w7155 <= not w7148 and not w7150;
w7156 <= not w6817 and w7146;
w7157 <= not w6818 and w7156;
w7158 <= not w6854 and not w7149;
w7159 <= w7157 and w7158;
w7160 <= not w7155 and not w7159;
w7161 <= w7145 and not w7160;
w7162 <= not w7154 and not w7161;
w7163 <= not w6761 and not w6774;
w7164 <= not w6778 and not w7163;
w7165 <= not w6725 and not w6761;
w7166 <= not w6743 and w7165;
w7167 <= not w6779 and w7166;
w7168 <= not w6725 and not w6738;
w7169 <= not w6742 and not w7168;
w7170 <= not w7167 and not w7169;
w7171 <= not w6742 and w7165;
w7172 <= not w6743 and w7171;
w7173 <= not w6779 and not w7168;
w7174 <= w7172 and w7173;
w7175 <= not w7170 and not w7174;
w7176 <= w7164 and not w7175;
w7177 <= not w7167 and w7169;
w7178 <= w7167 and not w7169;
w7179 <= not w7177 and not w7178;
w7180 <= not w7164 and not w7179;
w7181 <= not w6783 and not w6858;
w7182 <= not w7180 and not w7181;
w7183 <= not w7176 and w7182;
w7184 <= not w7176 and not w7180;
w7185 <= w7181 and not w7184;
w7186 <= not w7183 and not w7185;
w7187 <= not w7162 and not w7186;
w7188 <= not w7180 and w7181;
w7189 <= not w7176 and w7188;
w7190 <= not w7181 and not w7184;
w7191 <= not w7189 and not w7190;
w7192 <= w7162 and not w7191;
w7193 <= not w6861 and not w7014;
w7194 <= not w7192 and w7193;
w7195 <= not w7187 and w7194;
w7196 <= not w7187 and not w7192;
w7197 <= not w7193 and not w7196;
w7198 <= not w7195 and not w7197;
w7199 <= not w6914 and not w6927;
w7200 <= not w6931 and not w7199;
w7201 <= not w6878 and not w6914;
w7202 <= not w6896 and w7201;
w7203 <= not w6932 and w7202;
w7204 <= not w6878 and not w6891;
w7205 <= not w6895 and not w7204;
w7206 <= not w7203 and not w7205;
w7207 <= not w6895 and w7201;
w7208 <= not w6896 and w7207;
w7209 <= not w6932 and not w7204;
w7210 <= w7208 and w7209;
w7211 <= not w7206 and not w7210;
w7212 <= w7200 and not w7211;
w7213 <= not w7203 and w7205;
w7214 <= w7203 and not w7205;
w7215 <= not w7213 and not w7214;
w7216 <= not w7200 and not w7215;
w7217 <= not w6936 and not w7011;
w7218 <= not w7216 and w7217;
w7219 <= not w7212 and w7218;
w7220 <= not w7212 and not w7216;
w7221 <= not w7217 and not w7220;
w7222 <= not w7219 and not w7221;
w7223 <= not w6989 and not w7002;
w7224 <= not w7006 and not w7223;
w7225 <= not w6953 and not w6989;
w7226 <= not w6971 and w7225;
w7227 <= not w7007 and w7226;
w7228 <= not w6953 and not w6966;
w7229 <= not w6970 and not w7228;
w7230 <= not w7227 and w7229;
w7231 <= w7227 and not w7229;
w7232 <= not w7230 and not w7231;
w7233 <= not w7224 and not w7232;
w7234 <= not w7227 and not w7229;
w7235 <= not w6970 and w7225;
w7236 <= not w6971 and w7235;
w7237 <= not w7007 and not w7228;
w7238 <= w7236 and w7237;
w7239 <= not w7234 and not w7238;
w7240 <= w7224 and not w7239;
w7241 <= not w7233 and not w7240;
w7242 <= not w7222 and w7241;
w7243 <= not w7216 and not w7217;
w7244 <= not w7212 and w7243;
w7245 <= w7217 and not w7220;
w7246 <= not w7244 and not w7245;
w7247 <= not w7241 and not w7246;
w7248 <= not w7242 and not w7247;
w7249 <= not w7198 and w7248;
w7250 <= not w7192 and not w7193;
w7251 <= not w7187 and w7250;
w7252 <= w7193 and not w7196;
w7253 <= not w7251 and not w7252;
w7254 <= not w7248 and not w7253;
w7255 <= not w7249 and not w7254;
w7256 <= not w7143 and w7255;
w7257 <= not w7137 and not w7138;
w7258 <= not w7132 and w7257;
w7259 <= w7138 and not w7141;
w7260 <= not w7258 and not w7259;
w7261 <= not w7255 and not w7260;
w7262 <= not w7256 and not w7261;
w7263 <= not w7026 and w7262;
w7264 <= not w6396 and not w7021;
w7265 <= not w6391 and w7264;
w7266 <= w7021 and not w7024;
w7267 <= not w7265 and not w7266;
w7268 <= not w7262 and not w7267;
w7269 <= not w7263 and not w7268;
w7270 <= A(334) and A(335);
w7271 <= A(334) and not A(335);
w7272 <= not A(334) and A(335);
w7273 <= not w7271 and not w7272;
w7274 <= A(336) and not w7273;
w7275 <= not w7270 and not w7274;
w7276 <= A(331) and A(332);
w7277 <= A(331) and not A(332);
w7278 <= not A(331) and A(332);
w7279 <= not w7277 and not w7278;
w7280 <= A(333) and not w7279;
w7281 <= not w7276 and not w7280;
w7282 <= w7275 and not w7281;
w7283 <= not w7275 and w7281;
w7284 <= A(333) and not w7277;
w7285 <= not w7278 and w7284;
w7286 <= not A(333) and not w7279;
w7287 <= not w7285 and not w7286;
w7288 <= A(336) and not w7271;
w7289 <= not w7272 and w7288;
w7290 <= not A(336) and not w7273;
w7291 <= not w7289 and not w7290;
w7292 <= not w7287 and not w7291;
w7293 <= not w7283 and w7292;
w7294 <= not w7282 and w7293;
w7295 <= not w7282 and not w7283;
w7296 <= not w7292 and not w7295;
w7297 <= not w7294 and not w7296;
w7298 <= not w7287 and w7291;
w7299 <= w7287 and not w7291;
w7300 <= not w7298 and not w7299;
w7301 <= w7292 and not w7295;
w7302 <= not w7275 and not w7281;
w7303 <= not w7301 and not w7302;
w7304 <= not w7300 and not w7303;
w7305 <= not w7297 and not w7304;
w7306 <= not w7297 and not w7303;
w7307 <= A(340) and A(341);
w7308 <= A(340) and not A(341);
w7309 <= not A(340) and A(341);
w7310 <= not w7308 and not w7309;
w7311 <= A(342) and not w7310;
w7312 <= not w7307 and not w7311;
w7313 <= A(337) and A(338);
w7314 <= A(337) and not A(338);
w7315 <= not A(337) and A(338);
w7316 <= not w7314 and not w7315;
w7317 <= A(339) and not w7316;
w7318 <= not w7313 and not w7317;
w7319 <= not w7312 and w7318;
w7320 <= w7312 and not w7318;
w7321 <= not w7319 and not w7320;
w7322 <= A(339) and not w7314;
w7323 <= not w7315 and w7322;
w7324 <= not A(339) and not w7316;
w7325 <= not w7323 and not w7324;
w7326 <= A(342) and not w7308;
w7327 <= not w7309 and w7326;
w7328 <= not A(342) and not w7310;
w7329 <= not w7327 and not w7328;
w7330 <= not w7325 and not w7329;
w7331 <= not w7321 and w7330;
w7332 <= not w7312 and not w7318;
w7333 <= not w7331 and not w7332;
w7334 <= not w7319 and w7330;
w7335 <= not w7320 and w7334;
w7336 <= not w7321 and not w7330;
w7337 <= not w7335 and not w7336;
w7338 <= not w7333 and not w7337;
w7339 <= not w7325 and w7329;
w7340 <= w7325 and not w7329;
w7341 <= not w7339 and not w7340;
w7342 <= not w7300 and not w7341;
w7343 <= not w7338 and w7342;
w7344 <= not w7306 and w7343;
w7345 <= not w7333 and not w7341;
w7346 <= not w7337 and not w7345;
w7347 <= not w7344 and not w7346;
w7348 <= not w7337 and w7342;
w7349 <= not w7338 and w7348;
w7350 <= not w7306 and not w7345;
w7351 <= w7349 and w7350;
w7352 <= not w7347 and not w7351;
w7353 <= w7305 and not w7352;
w7354 <= not w7344 and w7346;
w7355 <= w7344 and not w7346;
w7356 <= not w7354 and not w7355;
w7357 <= not w7305 and not w7356;
w7358 <= not w7338 and not w7341;
w7359 <= not w7300 and not w7306;
w7360 <= not w7358 and w7359;
w7361 <= w7358 and not w7359;
w7362 <= not w7360 and not w7361;
w7363 <= not A(325) and A(326);
w7364 <= A(325) and not A(326);
w7365 <= A(327) and not w7364;
w7366 <= not w7363 and w7365;
w7367 <= not w7363 and not w7364;
w7368 <= not A(327) and not w7367;
w7369 <= not w7366 and not w7368;
w7370 <= not A(328) and A(329);
w7371 <= A(328) and not A(329);
w7372 <= A(330) and not w7371;
w7373 <= not w7370 and w7372;
w7374 <= not w7370 and not w7371;
w7375 <= not A(330) and not w7374;
w7376 <= not w7373 and not w7375;
w7377 <= not w7369 and w7376;
w7378 <= w7369 and not w7376;
w7379 <= not w7377 and not w7378;
w7380 <= A(328) and A(329);
w7381 <= A(330) and not w7374;
w7382 <= not w7380 and not w7381;
w7383 <= A(325) and A(326);
w7384 <= A(327) and not w7367;
w7385 <= not w7383 and not w7384;
w7386 <= not w7382 and w7385;
w7387 <= w7382 and not w7385;
w7388 <= not w7386 and not w7387;
w7389 <= not w7369 and not w7376;
w7390 <= not w7388 and w7389;
w7391 <= not w7382 and not w7385;
w7392 <= not w7390 and not w7391;
w7393 <= not w7386 and w7389;
w7394 <= not w7387 and w7393;
w7395 <= not w7388 and not w7389;
w7396 <= not w7394 and not w7395;
w7397 <= not w7392 and not w7396;
w7398 <= not w7379 and not w7397;
w7399 <= not A(319) and A(320);
w7400 <= A(319) and not A(320);
w7401 <= A(321) and not w7400;
w7402 <= not w7399 and w7401;
w7403 <= not w7399 and not w7400;
w7404 <= not A(321) and not w7403;
w7405 <= not w7402 and not w7404;
w7406 <= not A(322) and A(323);
w7407 <= A(322) and not A(323);
w7408 <= A(324) and not w7407;
w7409 <= not w7406 and w7408;
w7410 <= not w7406 and not w7407;
w7411 <= not A(324) and not w7410;
w7412 <= not w7409 and not w7411;
w7413 <= not w7405 and w7412;
w7414 <= w7405 and not w7412;
w7415 <= not w7413 and not w7414;
w7416 <= A(322) and A(323);
w7417 <= A(324) and not w7410;
w7418 <= not w7416 and not w7417;
w7419 <= A(319) and A(320);
w7420 <= A(321) and not w7403;
w7421 <= not w7419 and not w7420;
w7422 <= not w7418 and w7421;
w7423 <= w7418 and not w7421;
w7424 <= not w7422 and not w7423;
w7425 <= not w7405 and not w7412;
w7426 <= not w7424 and w7425;
w7427 <= not w7418 and not w7421;
w7428 <= not w7426 and not w7427;
w7429 <= not w7422 and w7425;
w7430 <= not w7423 and w7429;
w7431 <= not w7424 and not w7425;
w7432 <= not w7430 and not w7431;
w7433 <= not w7428 and not w7432;
w7434 <= not w7415 and not w7433;
w7435 <= not w7398 and w7434;
w7436 <= w7398 and not w7434;
w7437 <= not w7435 and not w7436;
w7438 <= not w7362 and not w7437;
w7439 <= not w7357 and w7438;
w7440 <= not w7353 and w7439;
w7441 <= not w7353 and not w7357;
w7442 <= not w7438 and not w7441;
w7443 <= not w7440 and not w7442;
w7444 <= not w7415 and not w7428;
w7445 <= not w7432 and not w7444;
w7446 <= not w7379 and not w7415;
w7447 <= not w7397 and w7446;
w7448 <= not w7433 and w7447;
w7449 <= not w7379 and not w7392;
w7450 <= not w7396 and not w7449;
w7451 <= not w7448 and w7450;
w7452 <= w7448 and not w7450;
w7453 <= not w7451 and not w7452;
w7454 <= not w7445 and not w7453;
w7455 <= not w7448 and not w7450;
w7456 <= not w7396 and w7446;
w7457 <= not w7397 and w7456;
w7458 <= not w7433 and not w7449;
w7459 <= w7457 and w7458;
w7460 <= not w7455 and not w7459;
w7461 <= w7445 and not w7460;
w7462 <= not w7454 and not w7461;
w7463 <= not w7443 and w7462;
w7464 <= not w7357 and not w7438;
w7465 <= not w7353 and w7464;
w7466 <= w7438 and not w7441;
w7467 <= not w7465 and not w7466;
w7468 <= not w7462 and not w7467;
w7469 <= not w7463 and not w7468;
w7470 <= A(346) and A(347);
w7471 <= A(346) and not A(347);
w7472 <= not A(346) and A(347);
w7473 <= not w7471 and not w7472;
w7474 <= A(348) and not w7473;
w7475 <= not w7470 and not w7474;
w7476 <= A(343) and A(344);
w7477 <= A(343) and not A(344);
w7478 <= not A(343) and A(344);
w7479 <= not w7477 and not w7478;
w7480 <= A(345) and not w7479;
w7481 <= not w7476 and not w7480;
w7482 <= w7475 and not w7481;
w7483 <= not w7475 and w7481;
w7484 <= A(345) and not w7477;
w7485 <= not w7478 and w7484;
w7486 <= not A(345) and not w7479;
w7487 <= not w7485 and not w7486;
w7488 <= A(348) and not w7471;
w7489 <= not w7472 and w7488;
w7490 <= not A(348) and not w7473;
w7491 <= not w7489 and not w7490;
w7492 <= not w7487 and not w7491;
w7493 <= not w7483 and w7492;
w7494 <= not w7482 and w7493;
w7495 <= not w7482 and not w7483;
w7496 <= not w7492 and not w7495;
w7497 <= not w7494 and not w7496;
w7498 <= not w7487 and w7491;
w7499 <= w7487 and not w7491;
w7500 <= not w7498 and not w7499;
w7501 <= w7492 and not w7495;
w7502 <= not w7475 and not w7481;
w7503 <= not w7501 and not w7502;
w7504 <= not w7500 and not w7503;
w7505 <= not w7497 and not w7504;
w7506 <= not w7497 and not w7503;
w7507 <= A(352) and A(353);
w7508 <= A(352) and not A(353);
w7509 <= not A(352) and A(353);
w7510 <= not w7508 and not w7509;
w7511 <= A(354) and not w7510;
w7512 <= not w7507 and not w7511;
w7513 <= A(349) and A(350);
w7514 <= A(349) and not A(350);
w7515 <= not A(349) and A(350);
w7516 <= not w7514 and not w7515;
w7517 <= A(351) and not w7516;
w7518 <= not w7513 and not w7517;
w7519 <= not w7512 and w7518;
w7520 <= w7512 and not w7518;
w7521 <= not w7519 and not w7520;
w7522 <= A(351) and not w7514;
w7523 <= not w7515 and w7522;
w7524 <= not A(351) and not w7516;
w7525 <= not w7523 and not w7524;
w7526 <= A(354) and not w7508;
w7527 <= not w7509 and w7526;
w7528 <= not A(354) and not w7510;
w7529 <= not w7527 and not w7528;
w7530 <= not w7525 and not w7529;
w7531 <= not w7521 and w7530;
w7532 <= not w7512 and not w7518;
w7533 <= not w7531 and not w7532;
w7534 <= not w7519 and w7530;
w7535 <= not w7520 and w7534;
w7536 <= not w7521 and not w7530;
w7537 <= not w7535 and not w7536;
w7538 <= not w7533 and not w7537;
w7539 <= not w7525 and w7529;
w7540 <= w7525 and not w7529;
w7541 <= not w7539 and not w7540;
w7542 <= not w7500 and not w7541;
w7543 <= not w7538 and w7542;
w7544 <= not w7506 and w7543;
w7545 <= not w7533 and not w7541;
w7546 <= not w7537 and not w7545;
w7547 <= not w7544 and w7546;
w7548 <= w7544 and not w7546;
w7549 <= not w7547 and not w7548;
w7550 <= not w7505 and not w7549;
w7551 <= not w7544 and not w7546;
w7552 <= not w7537 and w7542;
w7553 <= not w7538 and w7552;
w7554 <= not w7506 and not w7545;
w7555 <= w7553 and w7554;
w7556 <= not w7551 and not w7555;
w7557 <= w7505 and not w7556;
w7558 <= not w7550 and not w7557;
w7559 <= A(358) and A(359);
w7560 <= A(358) and not A(359);
w7561 <= not A(358) and A(359);
w7562 <= not w7560 and not w7561;
w7563 <= A(360) and not w7562;
w7564 <= not w7559 and not w7563;
w7565 <= A(355) and A(356);
w7566 <= A(355) and not A(356);
w7567 <= not A(355) and A(356);
w7568 <= not w7566 and not w7567;
w7569 <= A(357) and not w7568;
w7570 <= not w7565 and not w7569;
w7571 <= w7564 and not w7570;
w7572 <= not w7564 and w7570;
w7573 <= A(357) and not w7566;
w7574 <= not w7567 and w7573;
w7575 <= not A(357) and not w7568;
w7576 <= not w7574 and not w7575;
w7577 <= A(360) and not w7560;
w7578 <= not w7561 and w7577;
w7579 <= not A(360) and not w7562;
w7580 <= not w7578 and not w7579;
w7581 <= not w7576 and not w7580;
w7582 <= not w7572 and w7581;
w7583 <= not w7571 and w7582;
w7584 <= not w7571 and not w7572;
w7585 <= not w7581 and not w7584;
w7586 <= not w7583 and not w7585;
w7587 <= not w7576 and w7580;
w7588 <= w7576 and not w7580;
w7589 <= not w7587 and not w7588;
w7590 <= w7581 and not w7584;
w7591 <= not w7564 and not w7570;
w7592 <= not w7590 and not w7591;
w7593 <= not w7589 and not w7592;
w7594 <= not w7586 and not w7593;
w7595 <= not w7586 and not w7592;
w7596 <= A(364) and A(365);
w7597 <= A(364) and not A(365);
w7598 <= not A(364) and A(365);
w7599 <= not w7597 and not w7598;
w7600 <= A(366) and not w7599;
w7601 <= not w7596 and not w7600;
w7602 <= A(361) and A(362);
w7603 <= A(361) and not A(362);
w7604 <= not A(361) and A(362);
w7605 <= not w7603 and not w7604;
w7606 <= A(363) and not w7605;
w7607 <= not w7602 and not w7606;
w7608 <= not w7601 and w7607;
w7609 <= w7601 and not w7607;
w7610 <= not w7608 and not w7609;
w7611 <= A(363) and not w7603;
w7612 <= not w7604 and w7611;
w7613 <= not A(363) and not w7605;
w7614 <= not w7612 and not w7613;
w7615 <= A(366) and not w7597;
w7616 <= not w7598 and w7615;
w7617 <= not A(366) and not w7599;
w7618 <= not w7616 and not w7617;
w7619 <= not w7614 and not w7618;
w7620 <= not w7610 and w7619;
w7621 <= not w7601 and not w7607;
w7622 <= not w7620 and not w7621;
w7623 <= not w7608 and w7619;
w7624 <= not w7609 and w7623;
w7625 <= not w7610 and not w7619;
w7626 <= not w7624 and not w7625;
w7627 <= not w7622 and not w7626;
w7628 <= not w7614 and w7618;
w7629 <= w7614 and not w7618;
w7630 <= not w7628 and not w7629;
w7631 <= not w7589 and not w7630;
w7632 <= not w7627 and w7631;
w7633 <= not w7595 and w7632;
w7634 <= not w7622 and not w7630;
w7635 <= not w7626 and not w7634;
w7636 <= not w7633 and not w7635;
w7637 <= not w7626 and w7631;
w7638 <= not w7627 and w7637;
w7639 <= not w7595 and not w7634;
w7640 <= w7638 and w7639;
w7641 <= not w7636 and not w7640;
w7642 <= w7594 and not w7641;
w7643 <= not w7633 and w7635;
w7644 <= w7633 and not w7635;
w7645 <= not w7643 and not w7644;
w7646 <= not w7594 and not w7645;
w7647 <= not w7627 and not w7630;
w7648 <= not w7589 and not w7595;
w7649 <= not w7647 and w7648;
w7650 <= w7647 and not w7648;
w7651 <= not w7649 and not w7650;
w7652 <= not w7538 and not w7541;
w7653 <= not w7500 and not w7506;
w7654 <= not w7652 and w7653;
w7655 <= w7652 and not w7653;
w7656 <= not w7654 and not w7655;
w7657 <= not w7651 and not w7656;
w7658 <= not w7646 and not w7657;
w7659 <= not w7642 and w7658;
w7660 <= not w7642 and not w7646;
w7661 <= w7657 and not w7660;
w7662 <= not w7659 and not w7661;
w7663 <= not w7558 and not w7662;
w7664 <= not w7646 and w7657;
w7665 <= not w7642 and w7664;
w7666 <= not w7657 and not w7660;
w7667 <= not w7665 and not w7666;
w7668 <= w7558 and not w7667;
w7669 <= not w7651 and w7656;
w7670 <= w7651 and not w7656;
w7671 <= not w7669 and not w7670;
w7672 <= not w7362 and w7437;
w7673 <= w7362 and not w7437;
w7674 <= not w7672 and not w7673;
w7675 <= not w7671 and not w7674;
w7676 <= not w7668 and not w7675;
w7677 <= not w7663 and w7676;
w7678 <= not w7663 and not w7668;
w7679 <= w7675 and not w7678;
w7680 <= not w7677 and not w7679;
w7681 <= not w7469 and not w7680;
w7682 <= not w7668 and w7675;
w7683 <= not w7663 and w7682;
w7684 <= not w7675 and not w7678;
w7685 <= not w7683 and not w7684;
w7686 <= w7469 and not w7685;
w7687 <= not w7671 and w7674;
w7688 <= w7671 and not w7674;
w7689 <= not w7687 and not w7688;
w7690 <= not A(313) and A(314);
w7691 <= A(313) and not A(314);
w7692 <= A(315) and not w7691;
w7693 <= not w7690 and w7692;
w7694 <= not w7690 and not w7691;
w7695 <= not A(315) and not w7694;
w7696 <= not w7693 and not w7695;
w7697 <= not A(316) and A(317);
w7698 <= A(316) and not A(317);
w7699 <= A(318) and not w7698;
w7700 <= not w7697 and w7699;
w7701 <= not w7697 and not w7698;
w7702 <= not A(318) and not w7701;
w7703 <= not w7700 and not w7702;
w7704 <= not w7696 and w7703;
w7705 <= w7696 and not w7703;
w7706 <= not w7704 and not w7705;
w7707 <= A(316) and A(317);
w7708 <= A(318) and not w7701;
w7709 <= not w7707 and not w7708;
w7710 <= A(313) and A(314);
w7711 <= A(315) and not w7694;
w7712 <= not w7710 and not w7711;
w7713 <= not w7709 and w7712;
w7714 <= w7709 and not w7712;
w7715 <= not w7713 and not w7714;
w7716 <= not w7696 and not w7703;
w7717 <= not w7715 and w7716;
w7718 <= not w7709 and not w7712;
w7719 <= not w7717 and not w7718;
w7720 <= not w7713 and w7716;
w7721 <= not w7714 and w7720;
w7722 <= not w7715 and not w7716;
w7723 <= not w7721 and not w7722;
w7724 <= not w7719 and not w7723;
w7725 <= not w7706 and not w7724;
w7726 <= not A(307) and A(308);
w7727 <= A(307) and not A(308);
w7728 <= A(309) and not w7727;
w7729 <= not w7726 and w7728;
w7730 <= not w7726 and not w7727;
w7731 <= not A(309) and not w7730;
w7732 <= not w7729 and not w7731;
w7733 <= not A(310) and A(311);
w7734 <= A(310) and not A(311);
w7735 <= A(312) and not w7734;
w7736 <= not w7733 and w7735;
w7737 <= not w7733 and not w7734;
w7738 <= not A(312) and not w7737;
w7739 <= not w7736 and not w7738;
w7740 <= not w7732 and w7739;
w7741 <= w7732 and not w7739;
w7742 <= not w7740 and not w7741;
w7743 <= A(310) and A(311);
w7744 <= A(312) and not w7737;
w7745 <= not w7743 and not w7744;
w7746 <= A(307) and A(308);
w7747 <= A(309) and not w7730;
w7748 <= not w7746 and not w7747;
w7749 <= not w7745 and w7748;
w7750 <= w7745 and not w7748;
w7751 <= not w7749 and not w7750;
w7752 <= not w7732 and not w7739;
w7753 <= not w7751 and w7752;
w7754 <= not w7745 and not w7748;
w7755 <= not w7753 and not w7754;
w7756 <= not w7749 and w7752;
w7757 <= not w7750 and w7756;
w7758 <= not w7751 and not w7752;
w7759 <= not w7757 and not w7758;
w7760 <= not w7755 and not w7759;
w7761 <= not w7742 and not w7760;
w7762 <= not w7725 and w7761;
w7763 <= w7725 and not w7761;
w7764 <= not w7762 and not w7763;
w7765 <= not A(301) and A(302);
w7766 <= A(301) and not A(302);
w7767 <= A(303) and not w7766;
w7768 <= not w7765 and w7767;
w7769 <= not w7765 and not w7766;
w7770 <= not A(303) and not w7769;
w7771 <= not w7768 and not w7770;
w7772 <= not A(304) and A(305);
w7773 <= A(304) and not A(305);
w7774 <= A(306) and not w7773;
w7775 <= not w7772 and w7774;
w7776 <= not w7772 and not w7773;
w7777 <= not A(306) and not w7776;
w7778 <= not w7775 and not w7777;
w7779 <= not w7771 and w7778;
w7780 <= w7771 and not w7778;
w7781 <= not w7779 and not w7780;
w7782 <= A(304) and A(305);
w7783 <= A(306) and not w7776;
w7784 <= not w7782 and not w7783;
w7785 <= A(301) and A(302);
w7786 <= A(303) and not w7769;
w7787 <= not w7785 and not w7786;
w7788 <= not w7784 and w7787;
w7789 <= w7784 and not w7787;
w7790 <= not w7788 and not w7789;
w7791 <= not w7771 and not w7778;
w7792 <= not w7790 and w7791;
w7793 <= not w7784 and not w7787;
w7794 <= not w7792 and not w7793;
w7795 <= not w7788 and w7791;
w7796 <= not w7789 and w7795;
w7797 <= not w7790 and not w7791;
w7798 <= not w7796 and not w7797;
w7799 <= not w7794 and not w7798;
w7800 <= not w7781 and not w7799;
w7801 <= not A(295) and A(296);
w7802 <= A(295) and not A(296);
w7803 <= A(297) and not w7802;
w7804 <= not w7801 and w7803;
w7805 <= not w7801 and not w7802;
w7806 <= not A(297) and not w7805;
w7807 <= not w7804 and not w7806;
w7808 <= not A(298) and A(299);
w7809 <= A(298) and not A(299);
w7810 <= A(300) and not w7809;
w7811 <= not w7808 and w7810;
w7812 <= not w7808 and not w7809;
w7813 <= not A(300) and not w7812;
w7814 <= not w7811 and not w7813;
w7815 <= not w7807 and w7814;
w7816 <= w7807 and not w7814;
w7817 <= not w7815 and not w7816;
w7818 <= A(298) and A(299);
w7819 <= A(300) and not w7812;
w7820 <= not w7818 and not w7819;
w7821 <= A(295) and A(296);
w7822 <= A(297) and not w7805;
w7823 <= not w7821 and not w7822;
w7824 <= not w7820 and w7823;
w7825 <= w7820 and not w7823;
w7826 <= not w7824 and not w7825;
w7827 <= not w7807 and not w7814;
w7828 <= not w7826 and w7827;
w7829 <= not w7820 and not w7823;
w7830 <= not w7828 and not w7829;
w7831 <= not w7824 and w7827;
w7832 <= not w7825 and w7831;
w7833 <= not w7826 and not w7827;
w7834 <= not w7832 and not w7833;
w7835 <= not w7830 and not w7834;
w7836 <= not w7817 and not w7835;
w7837 <= not w7800 and w7836;
w7838 <= w7800 and not w7836;
w7839 <= not w7837 and not w7838;
w7840 <= not w7764 and w7839;
w7841 <= w7764 and not w7839;
w7842 <= not w7840 and not w7841;
w7843 <= not A(289) and A(290);
w7844 <= A(289) and not A(290);
w7845 <= A(291) and not w7844;
w7846 <= not w7843 and w7845;
w7847 <= not w7843 and not w7844;
w7848 <= not A(291) and not w7847;
w7849 <= not w7846 and not w7848;
w7850 <= not A(292) and A(293);
w7851 <= A(292) and not A(293);
w7852 <= A(294) and not w7851;
w7853 <= not w7850 and w7852;
w7854 <= not w7850 and not w7851;
w7855 <= not A(294) and not w7854;
w7856 <= not w7853 and not w7855;
w7857 <= not w7849 and w7856;
w7858 <= w7849 and not w7856;
w7859 <= not w7857 and not w7858;
w7860 <= A(292) and A(293);
w7861 <= A(294) and not w7854;
w7862 <= not w7860 and not w7861;
w7863 <= A(289) and A(290);
w7864 <= A(291) and not w7847;
w7865 <= not w7863 and not w7864;
w7866 <= not w7862 and w7865;
w7867 <= w7862 and not w7865;
w7868 <= not w7866 and not w7867;
w7869 <= not w7849 and not w7856;
w7870 <= not w7868 and w7869;
w7871 <= not w7862 and not w7865;
w7872 <= not w7870 and not w7871;
w7873 <= not w7866 and w7869;
w7874 <= not w7867 and w7873;
w7875 <= not w7868 and not w7869;
w7876 <= not w7874 and not w7875;
w7877 <= not w7872 and not w7876;
w7878 <= not w7859 and not w7877;
w7879 <= not A(283) and A(284);
w7880 <= A(283) and not A(284);
w7881 <= A(285) and not w7880;
w7882 <= not w7879 and w7881;
w7883 <= not w7879 and not w7880;
w7884 <= not A(285) and not w7883;
w7885 <= not w7882 and not w7884;
w7886 <= not A(286) and A(287);
w7887 <= A(286) and not A(287);
w7888 <= A(288) and not w7887;
w7889 <= not w7886 and w7888;
w7890 <= not w7886 and not w7887;
w7891 <= not A(288) and not w7890;
w7892 <= not w7889 and not w7891;
w7893 <= not w7885 and w7892;
w7894 <= w7885 and not w7892;
w7895 <= not w7893 and not w7894;
w7896 <= A(286) and A(287);
w7897 <= A(288) and not w7890;
w7898 <= not w7896 and not w7897;
w7899 <= A(283) and A(284);
w7900 <= A(285) and not w7883;
w7901 <= not w7899 and not w7900;
w7902 <= not w7898 and w7901;
w7903 <= w7898 and not w7901;
w7904 <= not w7902 and not w7903;
w7905 <= not w7885 and not w7892;
w7906 <= not w7904 and w7905;
w7907 <= not w7898 and not w7901;
w7908 <= not w7906 and not w7907;
w7909 <= not w7902 and w7905;
w7910 <= not w7903 and w7909;
w7911 <= not w7904 and not w7905;
w7912 <= not w7910 and not w7911;
w7913 <= not w7908 and not w7912;
w7914 <= not w7895 and not w7913;
w7915 <= not w7878 and w7914;
w7916 <= w7878 and not w7914;
w7917 <= not w7915 and not w7916;
w7918 <= not A(277) and A(278);
w7919 <= A(277) and not A(278);
w7920 <= A(279) and not w7919;
w7921 <= not w7918 and w7920;
w7922 <= not w7918 and not w7919;
w7923 <= not A(279) and not w7922;
w7924 <= not w7921 and not w7923;
w7925 <= not A(280) and A(281);
w7926 <= A(280) and not A(281);
w7927 <= A(282) and not w7926;
w7928 <= not w7925 and w7927;
w7929 <= not w7925 and not w7926;
w7930 <= not A(282) and not w7929;
w7931 <= not w7928 and not w7930;
w7932 <= not w7924 and w7931;
w7933 <= w7924 and not w7931;
w7934 <= not w7932 and not w7933;
w7935 <= A(280) and A(281);
w7936 <= A(282) and not w7929;
w7937 <= not w7935 and not w7936;
w7938 <= A(277) and A(278);
w7939 <= A(279) and not w7922;
w7940 <= not w7938 and not w7939;
w7941 <= not w7937 and w7940;
w7942 <= w7937 and not w7940;
w7943 <= not w7941 and not w7942;
w7944 <= not w7924 and not w7931;
w7945 <= not w7943 and w7944;
w7946 <= not w7937 and not w7940;
w7947 <= not w7945 and not w7946;
w7948 <= not w7941 and w7944;
w7949 <= not w7942 and w7948;
w7950 <= not w7943 and not w7944;
w7951 <= not w7949 and not w7950;
w7952 <= not w7947 and not w7951;
w7953 <= not w7934 and not w7952;
w7954 <= not A(271) and A(272);
w7955 <= A(271) and not A(272);
w7956 <= A(273) and not w7955;
w7957 <= not w7954 and w7956;
w7958 <= not w7954 and not w7955;
w7959 <= not A(273) and not w7958;
w7960 <= not w7957 and not w7959;
w7961 <= not A(274) and A(275);
w7962 <= A(274) and not A(275);
w7963 <= A(276) and not w7962;
w7964 <= not w7961 and w7963;
w7965 <= not w7961 and not w7962;
w7966 <= not A(276) and not w7965;
w7967 <= not w7964 and not w7966;
w7968 <= not w7960 and w7967;
w7969 <= w7960 and not w7967;
w7970 <= not w7968 and not w7969;
w7971 <= A(274) and A(275);
w7972 <= A(276) and not w7965;
w7973 <= not w7971 and not w7972;
w7974 <= A(271) and A(272);
w7975 <= A(273) and not w7958;
w7976 <= not w7974 and not w7975;
w7977 <= not w7973 and w7976;
w7978 <= w7973 and not w7976;
w7979 <= not w7977 and not w7978;
w7980 <= not w7960 and not w7967;
w7981 <= not w7979 and w7980;
w7982 <= not w7973 and not w7976;
w7983 <= not w7981 and not w7982;
w7984 <= not w7977 and w7980;
w7985 <= not w7978 and w7984;
w7986 <= not w7979 and not w7980;
w7987 <= not w7985 and not w7986;
w7988 <= not w7983 and not w7987;
w7989 <= not w7970 and not w7988;
w7990 <= not w7953 and w7989;
w7991 <= w7953 and not w7989;
w7992 <= not w7990 and not w7991;
w7993 <= not w7917 and w7992;
w7994 <= w7917 and not w7992;
w7995 <= not w7993 and not w7994;
w7996 <= not w7842 and w7995;
w7997 <= w7842 and not w7995;
w7998 <= not w7996 and not w7997;
w7999 <= not w7689 and not w7998;
w8000 <= not w7686 and w7999;
w8001 <= not w7681 and w8000;
w8002 <= not w7681 and not w7686;
w8003 <= not w7999 and not w8002;
w8004 <= not w8001 and not w8003;
w8005 <= not w7817 and not w7830;
w8006 <= not w7834 and not w8005;
w8007 <= not w7781 and not w7817;
w8008 <= not w7799 and w8007;
w8009 <= not w7835 and w8008;
w8010 <= not w7781 and not w7794;
w8011 <= not w7798 and not w8010;
w8012 <= not w8009 and w8011;
w8013 <= w8009 and not w8011;
w8014 <= not w8012 and not w8013;
w8015 <= not w8006 and not w8014;
w8016 <= not w8009 and not w8011;
w8017 <= not w7798 and w8007;
w8018 <= not w7799 and w8017;
w8019 <= not w7835 and not w8010;
w8020 <= w8018 and w8019;
w8021 <= not w8016 and not w8020;
w8022 <= w8006 and not w8021;
w8023 <= not w8015 and not w8022;
w8024 <= not w7742 and not w7755;
w8025 <= not w7759 and not w8024;
w8026 <= not w7706 and not w7742;
w8027 <= not w7724 and w8026;
w8028 <= not w7760 and w8027;
w8029 <= not w7706 and not w7719;
w8030 <= not w7723 and not w8029;
w8031 <= not w8028 and not w8030;
w8032 <= not w7723 and w8026;
w8033 <= not w7724 and w8032;
w8034 <= not w7760 and not w8029;
w8035 <= w8033 and w8034;
w8036 <= not w8031 and not w8035;
w8037 <= w8025 and not w8036;
w8038 <= not w8028 and w8030;
w8039 <= w8028 and not w8030;
w8040 <= not w8038 and not w8039;
w8041 <= not w8025 and not w8040;
w8042 <= not w7764 and not w7839;
w8043 <= not w8041 and not w8042;
w8044 <= not w8037 and w8043;
w8045 <= not w8037 and not w8041;
w8046 <= w8042 and not w8045;
w8047 <= not w8044 and not w8046;
w8048 <= not w8023 and not w8047;
w8049 <= not w8041 and w8042;
w8050 <= not w8037 and w8049;
w8051 <= not w8042 and not w8045;
w8052 <= not w8050 and not w8051;
w8053 <= w8023 and not w8052;
w8054 <= not w7842 and not w7995;
w8055 <= not w8053 and w8054;
w8056 <= not w8048 and w8055;
w8057 <= not w8048 and not w8053;
w8058 <= not w8054 and not w8057;
w8059 <= not w8056 and not w8058;
w8060 <= not w7895 and not w7908;
w8061 <= not w7912 and not w8060;
w8062 <= not w7859 and not w7895;
w8063 <= not w7877 and w8062;
w8064 <= not w7913 and w8063;
w8065 <= not w7859 and not w7872;
w8066 <= not w7876 and not w8065;
w8067 <= not w8064 and not w8066;
w8068 <= not w7876 and w8062;
w8069 <= not w7877 and w8068;
w8070 <= not w7913 and not w8065;
w8071 <= w8069 and w8070;
w8072 <= not w8067 and not w8071;
w8073 <= w8061 and not w8072;
w8074 <= not w8064 and w8066;
w8075 <= w8064 and not w8066;
w8076 <= not w8074 and not w8075;
w8077 <= not w8061 and not w8076;
w8078 <= not w7917 and not w7992;
w8079 <= not w8077 and w8078;
w8080 <= not w8073 and w8079;
w8081 <= not w8073 and not w8077;
w8082 <= not w8078 and not w8081;
w8083 <= not w8080 and not w8082;
w8084 <= not w7970 and not w7983;
w8085 <= not w7987 and not w8084;
w8086 <= not w7934 and not w7970;
w8087 <= not w7952 and w8086;
w8088 <= not w7988 and w8087;
w8089 <= not w7934 and not w7947;
w8090 <= not w7951 and not w8089;
w8091 <= not w8088 and w8090;
w8092 <= w8088 and not w8090;
w8093 <= not w8091 and not w8092;
w8094 <= not w8085 and not w8093;
w8095 <= not w8088 and not w8090;
w8096 <= not w7951 and w8086;
w8097 <= not w7952 and w8096;
w8098 <= not w7988 and not w8089;
w8099 <= w8097 and w8098;
w8100 <= not w8095 and not w8099;
w8101 <= w8085 and not w8100;
w8102 <= not w8094 and not w8101;
w8103 <= not w8083 and w8102;
w8104 <= not w8077 and not w8078;
w8105 <= not w8073 and w8104;
w8106 <= w8078 and not w8081;
w8107 <= not w8105 and not w8106;
w8108 <= not w8102 and not w8107;
w8109 <= not w8103 and not w8108;
w8110 <= not w8059 and w8109;
w8111 <= not w8053 and not w8054;
w8112 <= not w8048 and w8111;
w8113 <= w8054 and not w8057;
w8114 <= not w8112 and not w8113;
w8115 <= not w8109 and not w8114;
w8116 <= not w8110 and not w8115;
w8117 <= not w8004 and w8116;
w8118 <= not w7686 and not w7999;
w8119 <= not w7681 and w8118;
w8120 <= w7999 and not w8002;
w8121 <= not w8119 and not w8120;
w8122 <= not w8116 and not w8121;
w8123 <= not w8117 and not w8122;
w8124 <= A(394) and A(395);
w8125 <= A(394) and not A(395);
w8126 <= not A(394) and A(395);
w8127 <= not w8125 and not w8126;
w8128 <= A(396) and not w8127;
w8129 <= not w8124 and not w8128;
w8130 <= A(391) and A(392);
w8131 <= A(391) and not A(392);
w8132 <= not A(391) and A(392);
w8133 <= not w8131 and not w8132;
w8134 <= A(393) and not w8133;
w8135 <= not w8130 and not w8134;
w8136 <= w8129 and not w8135;
w8137 <= not w8129 and w8135;
w8138 <= A(393) and not w8131;
w8139 <= not w8132 and w8138;
w8140 <= not A(393) and not w8133;
w8141 <= not w8139 and not w8140;
w8142 <= A(396) and not w8125;
w8143 <= not w8126 and w8142;
w8144 <= not A(396) and not w8127;
w8145 <= not w8143 and not w8144;
w8146 <= not w8141 and not w8145;
w8147 <= not w8137 and w8146;
w8148 <= not w8136 and w8147;
w8149 <= not w8136 and not w8137;
w8150 <= not w8146 and not w8149;
w8151 <= not w8148 and not w8150;
w8152 <= not w8141 and w8145;
w8153 <= w8141 and not w8145;
w8154 <= not w8152 and not w8153;
w8155 <= w8146 and not w8149;
w8156 <= not w8129 and not w8135;
w8157 <= not w8155 and not w8156;
w8158 <= not w8154 and not w8157;
w8159 <= not w8151 and not w8158;
w8160 <= not w8151 and not w8157;
w8161 <= A(400) and A(401);
w8162 <= A(400) and not A(401);
w8163 <= not A(400) and A(401);
w8164 <= not w8162 and not w8163;
w8165 <= A(402) and not w8164;
w8166 <= not w8161 and not w8165;
w8167 <= A(397) and A(398);
w8168 <= A(397) and not A(398);
w8169 <= not A(397) and A(398);
w8170 <= not w8168 and not w8169;
w8171 <= A(399) and not w8170;
w8172 <= not w8167 and not w8171;
w8173 <= not w8166 and w8172;
w8174 <= w8166 and not w8172;
w8175 <= not w8173 and not w8174;
w8176 <= A(399) and not w8168;
w8177 <= not w8169 and w8176;
w8178 <= not A(399) and not w8170;
w8179 <= not w8177 and not w8178;
w8180 <= A(402) and not w8162;
w8181 <= not w8163 and w8180;
w8182 <= not A(402) and not w8164;
w8183 <= not w8181 and not w8182;
w8184 <= not w8179 and not w8183;
w8185 <= not w8175 and w8184;
w8186 <= not w8166 and not w8172;
w8187 <= not w8185 and not w8186;
w8188 <= not w8173 and w8184;
w8189 <= not w8174 and w8188;
w8190 <= not w8175 and not w8184;
w8191 <= not w8189 and not w8190;
w8192 <= not w8187 and not w8191;
w8193 <= not w8179 and w8183;
w8194 <= w8179 and not w8183;
w8195 <= not w8193 and not w8194;
w8196 <= not w8154 and not w8195;
w8197 <= not w8192 and w8196;
w8198 <= not w8160 and w8197;
w8199 <= not w8187 and not w8195;
w8200 <= not w8191 and not w8199;
w8201 <= not w8198 and w8200;
w8202 <= w8198 and not w8200;
w8203 <= not w8201 and not w8202;
w8204 <= not w8159 and not w8203;
w8205 <= not w8198 and not w8200;
w8206 <= not w8191 and w8196;
w8207 <= not w8192 and w8206;
w8208 <= not w8160 and not w8199;
w8209 <= w8207 and w8208;
w8210 <= not w8205 and not w8209;
w8211 <= w8159 and not w8210;
w8212 <= not w8204 and not w8211;
w8213 <= A(406) and A(407);
w8214 <= A(406) and not A(407);
w8215 <= not A(406) and A(407);
w8216 <= not w8214 and not w8215;
w8217 <= A(408) and not w8216;
w8218 <= not w8213 and not w8217;
w8219 <= A(403) and A(404);
w8220 <= A(403) and not A(404);
w8221 <= not A(403) and A(404);
w8222 <= not w8220 and not w8221;
w8223 <= A(405) and not w8222;
w8224 <= not w8219 and not w8223;
w8225 <= w8218 and not w8224;
w8226 <= not w8218 and w8224;
w8227 <= A(405) and not w8220;
w8228 <= not w8221 and w8227;
w8229 <= not A(405) and not w8222;
w8230 <= not w8228 and not w8229;
w8231 <= A(408) and not w8214;
w8232 <= not w8215 and w8231;
w8233 <= not A(408) and not w8216;
w8234 <= not w8232 and not w8233;
w8235 <= not w8230 and not w8234;
w8236 <= not w8226 and w8235;
w8237 <= not w8225 and w8236;
w8238 <= not w8225 and not w8226;
w8239 <= not w8235 and not w8238;
w8240 <= not w8237 and not w8239;
w8241 <= not w8230 and w8234;
w8242 <= w8230 and not w8234;
w8243 <= not w8241 and not w8242;
w8244 <= w8235 and not w8238;
w8245 <= not w8218 and not w8224;
w8246 <= not w8244 and not w8245;
w8247 <= not w8243 and not w8246;
w8248 <= not w8240 and not w8247;
w8249 <= not w8240 and not w8246;
w8250 <= A(412) and A(413);
w8251 <= A(412) and not A(413);
w8252 <= not A(412) and A(413);
w8253 <= not w8251 and not w8252;
w8254 <= A(414) and not w8253;
w8255 <= not w8250 and not w8254;
w8256 <= A(409) and A(410);
w8257 <= A(409) and not A(410);
w8258 <= not A(409) and A(410);
w8259 <= not w8257 and not w8258;
w8260 <= A(411) and not w8259;
w8261 <= not w8256 and not w8260;
w8262 <= not w8255 and w8261;
w8263 <= w8255 and not w8261;
w8264 <= not w8262 and not w8263;
w8265 <= A(411) and not w8257;
w8266 <= not w8258 and w8265;
w8267 <= not A(411) and not w8259;
w8268 <= not w8266 and not w8267;
w8269 <= A(414) and not w8251;
w8270 <= not w8252 and w8269;
w8271 <= not A(414) and not w8253;
w8272 <= not w8270 and not w8271;
w8273 <= not w8268 and not w8272;
w8274 <= not w8264 and w8273;
w8275 <= not w8255 and not w8261;
w8276 <= not w8274 and not w8275;
w8277 <= not w8262 and w8273;
w8278 <= not w8263 and w8277;
w8279 <= not w8264 and not w8273;
w8280 <= not w8278 and not w8279;
w8281 <= not w8276 and not w8280;
w8282 <= not w8268 and w8272;
w8283 <= w8268 and not w8272;
w8284 <= not w8282 and not w8283;
w8285 <= not w8243 and not w8284;
w8286 <= not w8281 and w8285;
w8287 <= not w8249 and w8286;
w8288 <= not w8276 and not w8284;
w8289 <= not w8280 and not w8288;
w8290 <= not w8287 and not w8289;
w8291 <= not w8280 and w8285;
w8292 <= not w8281 and w8291;
w8293 <= not w8249 and not w8288;
w8294 <= w8292 and w8293;
w8295 <= not w8290 and not w8294;
w8296 <= w8248 and not w8295;
w8297 <= not w8287 and w8289;
w8298 <= w8287 and not w8289;
w8299 <= not w8297 and not w8298;
w8300 <= not w8248 and not w8299;
w8301 <= not w8281 and not w8284;
w8302 <= not w8243 and not w8249;
w8303 <= not w8301 and w8302;
w8304 <= w8301 and not w8302;
w8305 <= not w8303 and not w8304;
w8306 <= not w8192 and not w8195;
w8307 <= not w8154 and not w8160;
w8308 <= not w8306 and w8307;
w8309 <= w8306 and not w8307;
w8310 <= not w8308 and not w8309;
w8311 <= not w8305 and not w8310;
w8312 <= not w8300 and not w8311;
w8313 <= not w8296 and w8312;
w8314 <= not w8296 and not w8300;
w8315 <= w8311 and not w8314;
w8316 <= not w8313 and not w8315;
w8317 <= not w8212 and not w8316;
w8318 <= not w8300 and w8311;
w8319 <= not w8296 and w8318;
w8320 <= not w8311 and not w8314;
w8321 <= not w8319 and not w8320;
w8322 <= w8212 and not w8321;
w8323 <= not w8305 and w8310;
w8324 <= w8305 and not w8310;
w8325 <= not w8323 and not w8324;
w8326 <= not A(385) and A(386);
w8327 <= A(385) and not A(386);
w8328 <= A(387) and not w8327;
w8329 <= not w8326 and w8328;
w8330 <= not w8326 and not w8327;
w8331 <= not A(387) and not w8330;
w8332 <= not w8329 and not w8331;
w8333 <= not A(388) and A(389);
w8334 <= A(388) and not A(389);
w8335 <= A(390) and not w8334;
w8336 <= not w8333 and w8335;
w8337 <= not w8333 and not w8334;
w8338 <= not A(390) and not w8337;
w8339 <= not w8336 and not w8338;
w8340 <= not w8332 and w8339;
w8341 <= w8332 and not w8339;
w8342 <= not w8340 and not w8341;
w8343 <= A(388) and A(389);
w8344 <= A(390) and not w8337;
w8345 <= not w8343 and not w8344;
w8346 <= A(385) and A(386);
w8347 <= A(387) and not w8330;
w8348 <= not w8346 and not w8347;
w8349 <= not w8345 and w8348;
w8350 <= w8345 and not w8348;
w8351 <= not w8349 and not w8350;
w8352 <= not w8332 and not w8339;
w8353 <= not w8351 and w8352;
w8354 <= not w8345 and not w8348;
w8355 <= not w8353 and not w8354;
w8356 <= not w8349 and w8352;
w8357 <= not w8350 and w8356;
w8358 <= not w8351 and not w8352;
w8359 <= not w8357 and not w8358;
w8360 <= not w8355 and not w8359;
w8361 <= not w8342 and not w8360;
w8362 <= not A(379) and A(380);
w8363 <= A(379) and not A(380);
w8364 <= A(381) and not w8363;
w8365 <= not w8362 and w8364;
w8366 <= not w8362 and not w8363;
w8367 <= not A(381) and not w8366;
w8368 <= not w8365 and not w8367;
w8369 <= not A(382) and A(383);
w8370 <= A(382) and not A(383);
w8371 <= A(384) and not w8370;
w8372 <= not w8369 and w8371;
w8373 <= not w8369 and not w8370;
w8374 <= not A(384) and not w8373;
w8375 <= not w8372 and not w8374;
w8376 <= not w8368 and w8375;
w8377 <= w8368 and not w8375;
w8378 <= not w8376 and not w8377;
w8379 <= A(382) and A(383);
w8380 <= A(384) and not w8373;
w8381 <= not w8379 and not w8380;
w8382 <= A(379) and A(380);
w8383 <= A(381) and not w8366;
w8384 <= not w8382 and not w8383;
w8385 <= not w8381 and w8384;
w8386 <= w8381 and not w8384;
w8387 <= not w8385 and not w8386;
w8388 <= not w8368 and not w8375;
w8389 <= not w8387 and w8388;
w8390 <= not w8381 and not w8384;
w8391 <= not w8389 and not w8390;
w8392 <= not w8385 and w8388;
w8393 <= not w8386 and w8392;
w8394 <= not w8387 and not w8388;
w8395 <= not w8393 and not w8394;
w8396 <= not w8391 and not w8395;
w8397 <= not w8378 and not w8396;
w8398 <= not w8361 and w8397;
w8399 <= w8361 and not w8397;
w8400 <= not w8398 and not w8399;
w8401 <= not A(373) and A(374);
w8402 <= A(373) and not A(374);
w8403 <= A(375) and not w8402;
w8404 <= not w8401 and w8403;
w8405 <= not w8401 and not w8402;
w8406 <= not A(375) and not w8405;
w8407 <= not w8404 and not w8406;
w8408 <= not A(376) and A(377);
w8409 <= A(376) and not A(377);
w8410 <= A(378) and not w8409;
w8411 <= not w8408 and w8410;
w8412 <= not w8408 and not w8409;
w8413 <= not A(378) and not w8412;
w8414 <= not w8411 and not w8413;
w8415 <= not w8407 and w8414;
w8416 <= w8407 and not w8414;
w8417 <= not w8415 and not w8416;
w8418 <= A(376) and A(377);
w8419 <= A(378) and not w8412;
w8420 <= not w8418 and not w8419;
w8421 <= A(373) and A(374);
w8422 <= A(375) and not w8405;
w8423 <= not w8421 and not w8422;
w8424 <= not w8420 and w8423;
w8425 <= w8420 and not w8423;
w8426 <= not w8424 and not w8425;
w8427 <= not w8407 and not w8414;
w8428 <= not w8426 and w8427;
w8429 <= not w8420 and not w8423;
w8430 <= not w8428 and not w8429;
w8431 <= not w8424 and w8427;
w8432 <= not w8425 and w8431;
w8433 <= not w8426 and not w8427;
w8434 <= not w8432 and not w8433;
w8435 <= not w8430 and not w8434;
w8436 <= not w8417 and not w8435;
w8437 <= not A(367) and A(368);
w8438 <= A(367) and not A(368);
w8439 <= A(369) and not w8438;
w8440 <= not w8437 and w8439;
w8441 <= not w8437 and not w8438;
w8442 <= not A(369) and not w8441;
w8443 <= not w8440 and not w8442;
w8444 <= not A(370) and A(371);
w8445 <= A(370) and not A(371);
w8446 <= A(372) and not w8445;
w8447 <= not w8444 and w8446;
w8448 <= not w8444 and not w8445;
w8449 <= not A(372) and not w8448;
w8450 <= not w8447 and not w8449;
w8451 <= not w8443 and w8450;
w8452 <= w8443 and not w8450;
w8453 <= not w8451 and not w8452;
w8454 <= A(370) and A(371);
w8455 <= A(372) and not w8448;
w8456 <= not w8454 and not w8455;
w8457 <= A(367) and A(368);
w8458 <= A(369) and not w8441;
w8459 <= not w8457 and not w8458;
w8460 <= not w8456 and w8459;
w8461 <= w8456 and not w8459;
w8462 <= not w8460 and not w8461;
w8463 <= not w8443 and not w8450;
w8464 <= not w8462 and w8463;
w8465 <= not w8456 and not w8459;
w8466 <= not w8464 and not w8465;
w8467 <= not w8460 and w8463;
w8468 <= not w8461 and w8467;
w8469 <= not w8462 and not w8463;
w8470 <= not w8468 and not w8469;
w8471 <= not w8466 and not w8470;
w8472 <= not w8453 and not w8471;
w8473 <= not w8436 and w8472;
w8474 <= w8436 and not w8472;
w8475 <= not w8473 and not w8474;
w8476 <= not w8400 and w8475;
w8477 <= w8400 and not w8475;
w8478 <= not w8476 and not w8477;
w8479 <= not w8325 and not w8478;
w8480 <= not w8322 and w8479;
w8481 <= not w8317 and w8480;
w8482 <= not w8317 and not w8322;
w8483 <= not w8479 and not w8482;
w8484 <= not w8481 and not w8483;
w8485 <= not w8378 and not w8391;
w8486 <= not w8395 and not w8485;
w8487 <= not w8342 and not w8378;
w8488 <= not w8360 and w8487;
w8489 <= not w8396 and w8488;
w8490 <= not w8342 and not w8355;
w8491 <= not w8359 and not w8490;
w8492 <= not w8489 and not w8491;
w8493 <= not w8359 and w8487;
w8494 <= not w8360 and w8493;
w8495 <= not w8396 and not w8490;
w8496 <= w8494 and w8495;
w8497 <= not w8492 and not w8496;
w8498 <= w8486 and not w8497;
w8499 <= not w8489 and w8491;
w8500 <= w8489 and not w8491;
w8501 <= not w8499 and not w8500;
w8502 <= not w8486 and not w8501;
w8503 <= not w8400 and not w8475;
w8504 <= not w8502 and w8503;
w8505 <= not w8498 and w8504;
w8506 <= not w8498 and not w8502;
w8507 <= not w8503 and not w8506;
w8508 <= not w8505 and not w8507;
w8509 <= not w8453 and not w8466;
w8510 <= not w8470 and not w8509;
w8511 <= not w8417 and not w8453;
w8512 <= not w8435 and w8511;
w8513 <= not w8471 and w8512;
w8514 <= not w8417 and not w8430;
w8515 <= not w8434 and not w8514;
w8516 <= not w8513 and w8515;
w8517 <= w8513 and not w8515;
w8518 <= not w8516 and not w8517;
w8519 <= not w8510 and not w8518;
w8520 <= not w8513 and not w8515;
w8521 <= not w8434 and w8511;
w8522 <= not w8435 and w8521;
w8523 <= not w8471 and not w8514;
w8524 <= w8522 and w8523;
w8525 <= not w8520 and not w8524;
w8526 <= w8510 and not w8525;
w8527 <= not w8519 and not w8526;
w8528 <= not w8508 and w8527;
w8529 <= not w8502 and not w8503;
w8530 <= not w8498 and w8529;
w8531 <= w8503 and not w8506;
w8532 <= not w8530 and not w8531;
w8533 <= not w8527 and not w8532;
w8534 <= not w8528 and not w8533;
w8535 <= not w8484 and w8534;
w8536 <= not w8322 and not w8479;
w8537 <= not w8317 and w8536;
w8538 <= w8479 and not w8482;
w8539 <= not w8537 and not w8538;
w8540 <= not w8534 and not w8539;
w8541 <= not w8535 and not w8540;
w8542 <= A(430) and A(431);
w8543 <= A(430) and not A(431);
w8544 <= not A(430) and A(431);
w8545 <= not w8543 and not w8544;
w8546 <= A(432) and not w8545;
w8547 <= not w8542 and not w8546;
w8548 <= A(427) and A(428);
w8549 <= A(427) and not A(428);
w8550 <= not A(427) and A(428);
w8551 <= not w8549 and not w8550;
w8552 <= A(429) and not w8551;
w8553 <= not w8548 and not w8552;
w8554 <= w8547 and not w8553;
w8555 <= not w8547 and w8553;
w8556 <= A(429) and not w8549;
w8557 <= not w8550 and w8556;
w8558 <= not A(429) and not w8551;
w8559 <= not w8557 and not w8558;
w8560 <= A(432) and not w8543;
w8561 <= not w8544 and w8560;
w8562 <= not A(432) and not w8545;
w8563 <= not w8561 and not w8562;
w8564 <= not w8559 and not w8563;
w8565 <= not w8555 and w8564;
w8566 <= not w8554 and w8565;
w8567 <= not w8554 and not w8555;
w8568 <= not w8564 and not w8567;
w8569 <= not w8566 and not w8568;
w8570 <= not w8559 and w8563;
w8571 <= w8559 and not w8563;
w8572 <= not w8570 and not w8571;
w8573 <= w8564 and not w8567;
w8574 <= not w8547 and not w8553;
w8575 <= not w8573 and not w8574;
w8576 <= not w8572 and not w8575;
w8577 <= not w8569 and not w8576;
w8578 <= not w8569 and not w8575;
w8579 <= A(436) and A(437);
w8580 <= A(436) and not A(437);
w8581 <= not A(436) and A(437);
w8582 <= not w8580 and not w8581;
w8583 <= A(438) and not w8582;
w8584 <= not w8579 and not w8583;
w8585 <= A(433) and A(434);
w8586 <= A(433) and not A(434);
w8587 <= not A(433) and A(434);
w8588 <= not w8586 and not w8587;
w8589 <= A(435) and not w8588;
w8590 <= not w8585 and not w8589;
w8591 <= not w8584 and w8590;
w8592 <= w8584 and not w8590;
w8593 <= not w8591 and not w8592;
w8594 <= A(435) and not w8586;
w8595 <= not w8587 and w8594;
w8596 <= not A(435) and not w8588;
w8597 <= not w8595 and not w8596;
w8598 <= A(438) and not w8580;
w8599 <= not w8581 and w8598;
w8600 <= not A(438) and not w8582;
w8601 <= not w8599 and not w8600;
w8602 <= not w8597 and not w8601;
w8603 <= not w8593 and w8602;
w8604 <= not w8584 and not w8590;
w8605 <= not w8603 and not w8604;
w8606 <= not w8591 and w8602;
w8607 <= not w8592 and w8606;
w8608 <= not w8593 and not w8602;
w8609 <= not w8607 and not w8608;
w8610 <= not w8605 and not w8609;
w8611 <= not w8597 and w8601;
w8612 <= w8597 and not w8601;
w8613 <= not w8611 and not w8612;
w8614 <= not w8572 and not w8613;
w8615 <= not w8610 and w8614;
w8616 <= not w8578 and w8615;
w8617 <= not w8605 and not w8613;
w8618 <= not w8609 and not w8617;
w8619 <= not w8616 and not w8618;
w8620 <= not w8609 and w8614;
w8621 <= not w8610 and w8620;
w8622 <= not w8578 and not w8617;
w8623 <= w8621 and w8622;
w8624 <= not w8619 and not w8623;
w8625 <= w8577 and not w8624;
w8626 <= not w8616 and w8618;
w8627 <= w8616 and not w8618;
w8628 <= not w8626 and not w8627;
w8629 <= not w8577 and not w8628;
w8630 <= not w8610 and not w8613;
w8631 <= not w8572 and not w8578;
w8632 <= not w8630 and w8631;
w8633 <= w8630 and not w8631;
w8634 <= not w8632 and not w8633;
w8635 <= not A(421) and A(422);
w8636 <= A(421) and not A(422);
w8637 <= A(423) and not w8636;
w8638 <= not w8635 and w8637;
w8639 <= not w8635 and not w8636;
w8640 <= not A(423) and not w8639;
w8641 <= not w8638 and not w8640;
w8642 <= not A(424) and A(425);
w8643 <= A(424) and not A(425);
w8644 <= A(426) and not w8643;
w8645 <= not w8642 and w8644;
w8646 <= not w8642 and not w8643;
w8647 <= not A(426) and not w8646;
w8648 <= not w8645 and not w8647;
w8649 <= not w8641 and w8648;
w8650 <= w8641 and not w8648;
w8651 <= not w8649 and not w8650;
w8652 <= A(424) and A(425);
w8653 <= A(426) and not w8646;
w8654 <= not w8652 and not w8653;
w8655 <= A(421) and A(422);
w8656 <= A(423) and not w8639;
w8657 <= not w8655 and not w8656;
w8658 <= not w8654 and w8657;
w8659 <= w8654 and not w8657;
w8660 <= not w8658 and not w8659;
w8661 <= not w8641 and not w8648;
w8662 <= not w8660 and w8661;
w8663 <= not w8654 and not w8657;
w8664 <= not w8662 and not w8663;
w8665 <= not w8658 and w8661;
w8666 <= not w8659 and w8665;
w8667 <= not w8660 and not w8661;
w8668 <= not w8666 and not w8667;
w8669 <= not w8664 and not w8668;
w8670 <= not w8651 and not w8669;
w8671 <= not A(415) and A(416);
w8672 <= A(415) and not A(416);
w8673 <= A(417) and not w8672;
w8674 <= not w8671 and w8673;
w8675 <= not w8671 and not w8672;
w8676 <= not A(417) and not w8675;
w8677 <= not w8674 and not w8676;
w8678 <= not A(418) and A(419);
w8679 <= A(418) and not A(419);
w8680 <= A(420) and not w8679;
w8681 <= not w8678 and w8680;
w8682 <= not w8678 and not w8679;
w8683 <= not A(420) and not w8682;
w8684 <= not w8681 and not w8683;
w8685 <= not w8677 and w8684;
w8686 <= w8677 and not w8684;
w8687 <= not w8685 and not w8686;
w8688 <= A(418) and A(419);
w8689 <= A(420) and not w8682;
w8690 <= not w8688 and not w8689;
w8691 <= A(415) and A(416);
w8692 <= A(417) and not w8675;
w8693 <= not w8691 and not w8692;
w8694 <= not w8690 and w8693;
w8695 <= w8690 and not w8693;
w8696 <= not w8694 and not w8695;
w8697 <= not w8677 and not w8684;
w8698 <= not w8696 and w8697;
w8699 <= not w8690 and not w8693;
w8700 <= not w8698 and not w8699;
w8701 <= not w8694 and w8697;
w8702 <= not w8695 and w8701;
w8703 <= not w8696 and not w8697;
w8704 <= not w8702 and not w8703;
w8705 <= not w8700 and not w8704;
w8706 <= not w8687 and not w8705;
w8707 <= not w8670 and w8706;
w8708 <= w8670 and not w8706;
w8709 <= not w8707 and not w8708;
w8710 <= not w8634 and not w8709;
w8711 <= not w8629 and w8710;
w8712 <= not w8625 and w8711;
w8713 <= not w8625 and not w8629;
w8714 <= not w8710 and not w8713;
w8715 <= not w8712 and not w8714;
w8716 <= not w8687 and not w8700;
w8717 <= not w8704 and not w8716;
w8718 <= not w8651 and not w8687;
w8719 <= not w8669 and w8718;
w8720 <= not w8705 and w8719;
w8721 <= not w8651 and not w8664;
w8722 <= not w8668 and not w8721;
w8723 <= not w8720 and w8722;
w8724 <= w8720 and not w8722;
w8725 <= not w8723 and not w8724;
w8726 <= not w8717 and not w8725;
w8727 <= not w8720 and not w8722;
w8728 <= not w8668 and w8718;
w8729 <= not w8669 and w8728;
w8730 <= not w8705 and not w8721;
w8731 <= w8729 and w8730;
w8732 <= not w8727 and not w8731;
w8733 <= w8717 and not w8732;
w8734 <= not w8726 and not w8733;
w8735 <= not w8715 and w8734;
w8736 <= not w8629 and not w8710;
w8737 <= not w8625 and w8736;
w8738 <= w8710 and not w8713;
w8739 <= not w8737 and not w8738;
w8740 <= not w8734 and not w8739;
w8741 <= not w8735 and not w8740;
w8742 <= A(442) and A(443);
w8743 <= A(442) and not A(443);
w8744 <= not A(442) and A(443);
w8745 <= not w8743 and not w8744;
w8746 <= A(444) and not w8745;
w8747 <= not w8742 and not w8746;
w8748 <= A(439) and A(440);
w8749 <= A(439) and not A(440);
w8750 <= not A(439) and A(440);
w8751 <= not w8749 and not w8750;
w8752 <= A(441) and not w8751;
w8753 <= not w8748 and not w8752;
w8754 <= w8747 and not w8753;
w8755 <= not w8747 and w8753;
w8756 <= A(441) and not w8749;
w8757 <= not w8750 and w8756;
w8758 <= not A(441) and not w8751;
w8759 <= not w8757 and not w8758;
w8760 <= A(444) and not w8743;
w8761 <= not w8744 and w8760;
w8762 <= not A(444) and not w8745;
w8763 <= not w8761 and not w8762;
w8764 <= not w8759 and not w8763;
w8765 <= not w8755 and w8764;
w8766 <= not w8754 and w8765;
w8767 <= not w8754 and not w8755;
w8768 <= not w8764 and not w8767;
w8769 <= not w8766 and not w8768;
w8770 <= not w8759 and w8763;
w8771 <= w8759 and not w8763;
w8772 <= not w8770 and not w8771;
w8773 <= w8764 and not w8767;
w8774 <= not w8747 and not w8753;
w8775 <= not w8773 and not w8774;
w8776 <= not w8772 and not w8775;
w8777 <= not w8769 and not w8776;
w8778 <= not w8769 and not w8775;
w8779 <= A(448) and A(449);
w8780 <= A(448) and not A(449);
w8781 <= not A(448) and A(449);
w8782 <= not w8780 and not w8781;
w8783 <= A(450) and not w8782;
w8784 <= not w8779 and not w8783;
w8785 <= A(445) and A(446);
w8786 <= A(445) and not A(446);
w8787 <= not A(445) and A(446);
w8788 <= not w8786 and not w8787;
w8789 <= A(447) and not w8788;
w8790 <= not w8785 and not w8789;
w8791 <= not w8784 and w8790;
w8792 <= w8784 and not w8790;
w8793 <= not w8791 and not w8792;
w8794 <= A(447) and not w8786;
w8795 <= not w8787 and w8794;
w8796 <= not A(447) and not w8788;
w8797 <= not w8795 and not w8796;
w8798 <= A(450) and not w8780;
w8799 <= not w8781 and w8798;
w8800 <= not A(450) and not w8782;
w8801 <= not w8799 and not w8800;
w8802 <= not w8797 and not w8801;
w8803 <= not w8793 and w8802;
w8804 <= not w8784 and not w8790;
w8805 <= not w8803 and not w8804;
w8806 <= not w8791 and w8802;
w8807 <= not w8792 and w8806;
w8808 <= not w8793 and not w8802;
w8809 <= not w8807 and not w8808;
w8810 <= not w8805 and not w8809;
w8811 <= not w8797 and w8801;
w8812 <= w8797 and not w8801;
w8813 <= not w8811 and not w8812;
w8814 <= not w8772 and not w8813;
w8815 <= not w8810 and w8814;
w8816 <= not w8778 and w8815;
w8817 <= not w8805 and not w8813;
w8818 <= not w8809 and not w8817;
w8819 <= not w8816 and w8818;
w8820 <= w8816 and not w8818;
w8821 <= not w8819 and not w8820;
w8822 <= not w8777 and not w8821;
w8823 <= not w8816 and not w8818;
w8824 <= not w8809 and w8814;
w8825 <= not w8810 and w8824;
w8826 <= not w8778 and not w8817;
w8827 <= w8825 and w8826;
w8828 <= not w8823 and not w8827;
w8829 <= w8777 and not w8828;
w8830 <= not w8822 and not w8829;
w8831 <= A(454) and A(455);
w8832 <= A(454) and not A(455);
w8833 <= not A(454) and A(455);
w8834 <= not w8832 and not w8833;
w8835 <= A(456) and not w8834;
w8836 <= not w8831 and not w8835;
w8837 <= A(451) and A(452);
w8838 <= A(451) and not A(452);
w8839 <= not A(451) and A(452);
w8840 <= not w8838 and not w8839;
w8841 <= A(453) and not w8840;
w8842 <= not w8837 and not w8841;
w8843 <= w8836 and not w8842;
w8844 <= not w8836 and w8842;
w8845 <= A(453) and not w8838;
w8846 <= not w8839 and w8845;
w8847 <= not A(453) and not w8840;
w8848 <= not w8846 and not w8847;
w8849 <= A(456) and not w8832;
w8850 <= not w8833 and w8849;
w8851 <= not A(456) and not w8834;
w8852 <= not w8850 and not w8851;
w8853 <= not w8848 and not w8852;
w8854 <= not w8844 and w8853;
w8855 <= not w8843 and w8854;
w8856 <= not w8843 and not w8844;
w8857 <= not w8853 and not w8856;
w8858 <= not w8855 and not w8857;
w8859 <= not w8848 and w8852;
w8860 <= w8848 and not w8852;
w8861 <= not w8859 and not w8860;
w8862 <= w8853 and not w8856;
w8863 <= not w8836 and not w8842;
w8864 <= not w8862 and not w8863;
w8865 <= not w8861 and not w8864;
w8866 <= not w8858 and not w8865;
w8867 <= not w8858 and not w8864;
w8868 <= A(460) and A(461);
w8869 <= A(460) and not A(461);
w8870 <= not A(460) and A(461);
w8871 <= not w8869 and not w8870;
w8872 <= A(462) and not w8871;
w8873 <= not w8868 and not w8872;
w8874 <= A(457) and A(458);
w8875 <= A(457) and not A(458);
w8876 <= not A(457) and A(458);
w8877 <= not w8875 and not w8876;
w8878 <= A(459) and not w8877;
w8879 <= not w8874 and not w8878;
w8880 <= not w8873 and w8879;
w8881 <= w8873 and not w8879;
w8882 <= not w8880 and not w8881;
w8883 <= A(459) and not w8875;
w8884 <= not w8876 and w8883;
w8885 <= not A(459) and not w8877;
w8886 <= not w8884 and not w8885;
w8887 <= A(462) and not w8869;
w8888 <= not w8870 and w8887;
w8889 <= not A(462) and not w8871;
w8890 <= not w8888 and not w8889;
w8891 <= not w8886 and not w8890;
w8892 <= not w8882 and w8891;
w8893 <= not w8873 and not w8879;
w8894 <= not w8892 and not w8893;
w8895 <= not w8880 and w8891;
w8896 <= not w8881 and w8895;
w8897 <= not w8882 and not w8891;
w8898 <= not w8896 and not w8897;
w8899 <= not w8894 and not w8898;
w8900 <= not w8886 and w8890;
w8901 <= w8886 and not w8890;
w8902 <= not w8900 and not w8901;
w8903 <= not w8861 and not w8902;
w8904 <= not w8899 and w8903;
w8905 <= not w8867 and w8904;
w8906 <= not w8894 and not w8902;
w8907 <= not w8898 and not w8906;
w8908 <= not w8905 and not w8907;
w8909 <= not w8898 and w8903;
w8910 <= not w8899 and w8909;
w8911 <= not w8867 and not w8906;
w8912 <= w8910 and w8911;
w8913 <= not w8908 and not w8912;
w8914 <= w8866 and not w8913;
w8915 <= not w8905 and w8907;
w8916 <= w8905 and not w8907;
w8917 <= not w8915 and not w8916;
w8918 <= not w8866 and not w8917;
w8919 <= not w8899 and not w8902;
w8920 <= not w8861 and not w8867;
w8921 <= not w8919 and w8920;
w8922 <= w8919 and not w8920;
w8923 <= not w8921 and not w8922;
w8924 <= not w8810 and not w8813;
w8925 <= not w8772 and not w8778;
w8926 <= not w8924 and w8925;
w8927 <= w8924 and not w8925;
w8928 <= not w8926 and not w8927;
w8929 <= not w8923 and not w8928;
w8930 <= not w8918 and not w8929;
w8931 <= not w8914 and w8930;
w8932 <= not w8914 and not w8918;
w8933 <= w8929 and not w8932;
w8934 <= not w8931 and not w8933;
w8935 <= not w8830 and not w8934;
w8936 <= not w8918 and w8929;
w8937 <= not w8914 and w8936;
w8938 <= not w8929 and not w8932;
w8939 <= not w8937 and not w8938;
w8940 <= w8830 and not w8939;
w8941 <= not w8923 and w8928;
w8942 <= w8923 and not w8928;
w8943 <= not w8941 and not w8942;
w8944 <= not w8634 and w8709;
w8945 <= w8634 and not w8709;
w8946 <= not w8944 and not w8945;
w8947 <= not w8943 and not w8946;
w8948 <= not w8940 and not w8947;
w8949 <= not w8935 and w8948;
w8950 <= not w8935 and not w8940;
w8951 <= w8947 and not w8950;
w8952 <= not w8949 and not w8951;
w8953 <= not w8741 and not w8952;
w8954 <= not w8940 and w8947;
w8955 <= not w8935 and w8954;
w8956 <= not w8947 and not w8950;
w8957 <= not w8955 and not w8956;
w8958 <= w8741 and not w8957;
w8959 <= not w8943 and w8946;
w8960 <= w8943 and not w8946;
w8961 <= not w8959 and not w8960;
w8962 <= not w8325 and w8478;
w8963 <= w8325 and not w8478;
w8964 <= not w8962 and not w8963;
w8965 <= not w8961 and not w8964;
w8966 <= not w8958 and not w8965;
w8967 <= not w8953 and w8966;
w8968 <= not w8953 and not w8958;
w8969 <= w8965 and not w8968;
w8970 <= not w8967 and not w8969;
w8971 <= not w8541 and not w8970;
w8972 <= not w8958 and w8965;
w8973 <= not w8953 and w8972;
w8974 <= not w8965 and not w8968;
w8975 <= not w8973 and not w8974;
w8976 <= w8541 and not w8975;
w8977 <= not w8961 and w8964;
w8978 <= w8961 and not w8964;
w8979 <= not w8977 and not w8978;
w8980 <= not w7689 and w7998;
w8981 <= w7689 and not w7998;
w8982 <= not w8980 and not w8981;
w8983 <= not w8979 and not w8982;
w8984 <= not w8976 and not w8983;
w8985 <= not w8971 and w8984;
w8986 <= not w8971 and not w8976;
w8987 <= w8983 and not w8986;
w8988 <= not w8985 and not w8987;
w8989 <= not w8123 and not w8988;
w8990 <= not w8976 and w8983;
w8991 <= not w8971 and w8990;
w8992 <= not w8983 and not w8986;
w8993 <= not w8991 and not w8992;
w8994 <= w8123 and not w8993;
w8995 <= not w8979 and w8982;
w8996 <= w8979 and not w8982;
w8997 <= not w8995 and not w8996;
w8998 <= not w6399 and w7020;
w8999 <= w6399 and not w7020;
w9000 <= not w8998 and not w8999;
w9001 <= not w8997 and not w9000;
w9002 <= not w8994 and not w9001;
w9003 <= not w8989 and w9002;
w9004 <= not w8989 and not w8994;
w9005 <= w9001 and not w9004;
w9006 <= not w9003 and not w9005;
w9007 <= not w7269 and not w9006;
w9008 <= not w8994 and w9001;
w9009 <= not w8989 and w9008;
w9010 <= not w9001 and not w9004;
w9011 <= not w9009 and not w9010;
w9012 <= w7269 and not w9011;
w9013 <= not w8997 and w9000;
w9014 <= w8997 and not w9000;
w9015 <= not w9013 and not w9014;
w9016 <= not w4673 and w5294;
w9017 <= not w4670 and not w5294;
w9018 <= not w4672 and w9017;
w9019 <= not w9016 and not w9018;
w9020 <= not w9015 and not w9019;
w9021 <= not w9012 and not w9020;
w9022 <= not w9007 and w9021;
w9023 <= not w9007 and not w9012;
w9024 <= w9020 and not w9023;
w9025 <= not w9022 and not w9024;
w9026 <= not w5543 and not w9025;
w9027 <= not w2969 and w2972;
w9028 <= w2969 and not w2972;
w9029 <= not w9027 and not w9028;
w9030 <= not w9015 and w9019;
w9031 <= w9015 and not w9019;
w9032 <= not w9030 and not w9031;
w9033 <= not w9029 and not w9032;
w9034 <= not w9012 and w9020;
w9035 <= not w9007 and w9034;
w9036 <= not w9020 and not w9023;
w9037 <= not w9035 and not w9036;
w9038 <= w5543 and not w9037;
w9039 <= not w9033 and not w9038;
w9040 <= not w9026 and w9039;
w9041 <= not w3469 and not w9040;
w9042 <= not w9026 and not w9038;
w9043 <= w9033 and not w9042;
w9044 <= not w9041 and not w9043;
w9045 <= not w5543 and not w9022;
w9046 <= not w9024 and not w9045;
w9047 <= not w5536 and not w5539;
w9048 <= not w5540 and not w9047;
w9049 <= not w3887 and not w4660;
w9050 <= not w4662 and not w9049;
w9051 <= not w4215 and not w4642;
w9052 <= not w4644 and not w9051;
w9053 <= not w4208 and not w4211;
w9054 <= not w4212 and not w9053;
w9055 <= w4169 and not w4204;
w9056 <= not w4205 and not w9055;
w9057 <= not w4190 and not w4191;
w9058 <= not w4187 and not w9057;
w9059 <= not w4174 and not w4177;
w9060 <= not w4184 and not w9059;
w9061 <= not w9058 and w9060;
w9062 <= not w4187 and not w9060;
w9063 <= not w9057 and w9062;
w9064 <= not w4106 and not w4123;
w9065 <= not w4119 and not w9064;
w9066 <= not w9063 and w9065;
w9067 <= not w9061 and w9066;
w9068 <= not w9061 and not w9063;
w9069 <= not w9065 and not w9068;
w9070 <= not w9067 and not w9069;
w9071 <= not w9056 and not w9070;
w9072 <= not w4205 and not w9067;
w9073 <= not w9055 and w9072;
w9074 <= not w9069 and w9073;
w9075 <= not w9071 and not w9074;
w9076 <= not w3976 and not w4077;
w9077 <= not w4079 and not w9076;
w9078 <= w3923 and not w3969;
w9079 <= not w3973 and not w9078;
w9080 <= not w3955 and not w3959;
w9081 <= not w3951 and not w9080;
w9082 <= not w3915 and not w3918;
w9083 <= not w3921 and not w9082;
w9084 <= not w9081 and w9083;
w9085 <= w9081 and not w9083;
w9086 <= not w9084 and not w9085;
w9087 <= not w9079 and not w9086;
w9088 <= not w3973 and not w9084;
w9089 <= not w9085 and w9088;
w9090 <= not w9078 and w9089;
w9091 <= not w9087 and not w9090;
w9092 <= w4012 and not w4054;
w9093 <= not w4058 and not w9092;
w9094 <= not w4044 and not w4048;
w9095 <= not w4040 and not w9094;
w9096 <= not w4004 and not w4007;
w9097 <= not w4010 and not w9096;
w9098 <= not w9095 and w9097;
w9099 <= w9095 and not w9097;
w9100 <= not w9098 and not w9099;
w9101 <= not w9093 and not w9100;
w9102 <= not w4058 and not w9098;
w9103 <= not w9099 and w9102;
w9104 <= not w9092 and w9103;
w9105 <= not w9101 and not w9104;
w9106 <= not w9091 and w9105;
w9107 <= w9091 and not w9105;
w9108 <= not w9106 and not w9107;
w9109 <= not w9077 and not w9108;
w9110 <= w9077 and w9108;
w9111 <= not w9109 and not w9110;
w9112 <= not w9075 and w9111;
w9113 <= w9075 and not w9111;
w9114 <= not w9112 and not w9113;
w9115 <= not w9054 and not w9114;
w9116 <= w9054 and w9114;
w9117 <= not w9115 and not w9116;
w9118 <= not w4415 and not w4623;
w9119 <= not w4625 and not w9118;
w9120 <= not w4408 and not w4411;
w9121 <= not w4412 and not w9120;
w9122 <= w4391 and not w4401;
w9123 <= not w4405 and not w9122;
w9124 <= not w4325 and not w4342;
w9125 <= not w4338 and not w9124;
w9126 <= not w4361 and not w4378;
w9127 <= not w4374 and not w9126;
w9128 <= not w9125 and w9127;
w9129 <= w9125 and not w9127;
w9130 <= not w9128 and not w9129;
w9131 <= not w9123 and not w9130;
w9132 <= not w4405 and not w9128;
w9133 <= not w9129 and w9132;
w9134 <= not w9122 and w9133;
w9135 <= not w9131 and not w9134;
w9136 <= w4251 and not w4293;
w9137 <= not w4297 and not w9136;
w9138 <= not w4283 and not w4287;
w9139 <= not w4279 and not w9138;
w9140 <= not w4243 and not w4246;
w9141 <= not w4249 and not w9140;
w9142 <= not w9139 and w9141;
w9143 <= w9139 and not w9141;
w9144 <= not w9142 and not w9143;
w9145 <= not w9137 and not w9144;
w9146 <= not w4297 and not w9142;
w9147 <= not w9143 and w9146;
w9148 <= not w9136 and w9147;
w9149 <= not w9145 and not w9148;
w9150 <= not w9135 and w9149;
w9151 <= w9135 and not w9149;
w9152 <= not w9150 and not w9151;
w9153 <= not w9121 and not w9152;
w9154 <= w9121 and w9152;
w9155 <= not w9153 and not w9154;
w9156 <= not w4504 and not w4605;
w9157 <= not w4607 and not w9156;
w9158 <= w4451 and not w4497;
w9159 <= not w4501 and not w9158;
w9160 <= not w4483 and not w4487;
w9161 <= not w4479 and not w9160;
w9162 <= not w4443 and not w4446;
w9163 <= not w4449 and not w9162;
w9164 <= not w9161 and w9163;
w9165 <= w9161 and not w9163;
w9166 <= not w9164 and not w9165;
w9167 <= not w9159 and not w9166;
w9168 <= not w4501 and not w9164;
w9169 <= not w9165 and w9168;
w9170 <= not w9158 and w9169;
w9171 <= not w9167 and not w9170;
w9172 <= w4540 and not w4582;
w9173 <= not w4586 and not w9172;
w9174 <= not w4572 and not w4576;
w9175 <= not w4568 and not w9174;
w9176 <= not w4532 and not w4535;
w9177 <= not w4538 and not w9176;
w9178 <= not w9175 and w9177;
w9179 <= w9175 and not w9177;
w9180 <= not w9178 and not w9179;
w9181 <= not w9173 and not w9180;
w9182 <= not w4586 and not w9178;
w9183 <= not w9179 and w9182;
w9184 <= not w9172 and w9183;
w9185 <= not w9181 and not w9184;
w9186 <= not w9171 and w9185;
w9187 <= w9171 and not w9185;
w9188 <= not w9186 and not w9187;
w9189 <= not w9157 and not w9188;
w9190 <= w9157 and w9188;
w9191 <= not w9189 and not w9190;
w9192 <= not w9155 and w9191;
w9193 <= w9155 and not w9191;
w9194 <= not w9192 and not w9193;
w9195 <= not w9119 and not w9194;
w9196 <= w9119 and w9194;
w9197 <= not w9195 and not w9196;
w9198 <= not w9117 and w9197;
w9199 <= w9117 and not w9197;
w9200 <= not w9198 and not w9199;
w9201 <= w9052 and w9200;
w9202 <= not w9052 and not w9200;
w9203 <= not w3880 and not w3883;
w9204 <= not w3884 and not w9203;
w9205 <= not w3873 and not w3876;
w9206 <= not w3877 and not w9205;
w9207 <= w3856 and not w3866;
w9208 <= not w3870 and not w9207;
w9209 <= not w3763 and not w3780;
w9210 <= not w3776 and not w9209;
w9211 <= not w3799 and not w3816;
w9212 <= not w3812 and not w9211;
w9213 <= not w9210 and w9212;
w9214 <= w9210 and not w9212;
w9215 <= not w9213 and not w9214;
w9216 <= not w9208 and not w9215;
w9217 <= not w3870 and not w9213;
w9218 <= not w9214 and w9217;
w9219 <= not w9207 and w9218;
w9220 <= not w9216 and not w9219;
w9221 <= w3832 and not w3838;
w9222 <= not w3842 and not w9221;
w9223 <= not w3688 and not w3705;
w9224 <= not w3701 and not w9223;
w9225 <= not w3724 and not w3741;
w9226 <= not w3737 and not w9225;
w9227 <= not w9224 and w9226;
w9228 <= w9224 and not w9226;
w9229 <= not w9227 and not w9228;
w9230 <= not w9222 and not w9229;
w9231 <= not w3842 and not w9227;
w9232 <= not w9228 and w9231;
w9233 <= not w9221 and w9232;
w9234 <= not w9230 and not w9233;
w9235 <= not w9220 and w9234;
w9236 <= w9220 and not w9234;
w9237 <= not w9235 and not w9236;
w9238 <= not w9206 and not w9237;
w9239 <= w9206 and w9237;
w9240 <= not w9238 and not w9239;
w9241 <= not w3558 and not w3659;
w9242 <= not w3661 and not w9241;
w9243 <= w3505 and not w3551;
w9244 <= not w3555 and not w9243;
w9245 <= not w3537 and not w3541;
w9246 <= not w3533 and not w9245;
w9247 <= not w3497 and not w3500;
w9248 <= not w3503 and not w9247;
w9249 <= not w9246 and w9248;
w9250 <= w9246 and not w9248;
w9251 <= not w9249 and not w9250;
w9252 <= not w9244 and not w9251;
w9253 <= not w3555 and not w9249;
w9254 <= not w9250 and w9253;
w9255 <= not w9243 and w9254;
w9256 <= not w9252 and not w9255;
w9257 <= w3594 and not w3636;
w9258 <= not w3640 and not w9257;
w9259 <= not w3626 and not w3630;
w9260 <= not w3622 and not w9259;
w9261 <= not w3586 and not w3589;
w9262 <= not w3592 and not w9261;
w9263 <= not w9260 and w9262;
w9264 <= w9260 and not w9262;
w9265 <= not w9263 and not w9264;
w9266 <= not w9258 and not w9265;
w9267 <= not w3640 and not w9263;
w9268 <= not w9264 and w9267;
w9269 <= not w9257 and w9268;
w9270 <= not w9266 and not w9269;
w9271 <= not w9256 and w9270;
w9272 <= w9256 and not w9270;
w9273 <= not w9271 and not w9272;
w9274 <= not w9242 and not w9273;
w9275 <= w9242 and w9273;
w9276 <= not w9274 and not w9275;
w9277 <= not w9240 and w9276;
w9278 <= w9240 and not w9276;
w9279 <= not w9277 and not w9278;
w9280 <= not w9204 and not w9279;
w9281 <= w9204 and w9279;
w9282 <= not w9280 and not w9281;
w9283 <= not w9202 and not w9282;
w9284 <= not w9201 and w9283;
w9285 <= not w9201 and not w9202;
w9286 <= w9282 and not w9285;
w9287 <= not w9284 and not w9286;
w9288 <= w9050 and w9287;
w9289 <= not w9050 and not w9287;
w9290 <= not w5529 and not w5532;
w9291 <= not w5533 and not w9290;
w9292 <= not w5522 and not w5525;
w9293 <= not w5526 and not w9292;
w9294 <= not w5515 and not w5518;
w9295 <= not w5519 and not w9294;
w9296 <= w5498 and not w5508;
w9297 <= not w5512 and not w9296;
w9298 <= not w5227 and not w5244;
w9299 <= not w5240 and not w9298;
w9300 <= not w5263 and not w5280;
w9301 <= not w5276 and not w9300;
w9302 <= not w9299 and w9301;
w9303 <= w9299 and not w9301;
w9304 <= not w9302 and not w9303;
w9305 <= not w9297 and not w9304;
w9306 <= not w5512 and not w9302;
w9307 <= not w9303 and w9306;
w9308 <= not w9296 and w9307;
w9309 <= not w9305 and not w9308;
w9310 <= w5474 and not w5480;
w9311 <= not w5484 and not w9310;
w9312 <= not w5152 and not w5169;
w9313 <= not w5165 and not w9312;
w9314 <= not w5188 and not w5205;
w9315 <= not w5201 and not w9314;
w9316 <= not w9313 and w9315;
w9317 <= w9313 and not w9315;
w9318 <= not w9316 and not w9317;
w9319 <= not w9311 and not w9318;
w9320 <= not w5484 and not w9316;
w9321 <= not w9317 and w9320;
w9322 <= not w9310 and w9321;
w9323 <= not w9319 and not w9322;
w9324 <= not w9309 and w9323;
w9325 <= w9309 and not w9323;
w9326 <= not w9324 and not w9325;
w9327 <= not w9295 and not w9326;
w9328 <= w9295 and w9326;
w9329 <= not w9327 and not w9328;
w9330 <= not w5436 and not w5457;
w9331 <= not w5459 and not w9330;
w9332 <= w5419 and not w5429;
w9333 <= not w5433 and not w9332;
w9334 <= not w5074 and not w5091;
w9335 <= not w5087 and not w9334;
w9336 <= not w5110 and not w5127;
w9337 <= not w5123 and not w9336;
w9338 <= not w9335 and w9337;
w9339 <= w9335 and not w9337;
w9340 <= not w9338 and not w9339;
w9341 <= not w9333 and not w9340;
w9342 <= not w5433 and not w9338;
w9343 <= not w9339 and w9342;
w9344 <= not w9332 and w9343;
w9345 <= not w9341 and not w9344;
w9346 <= w5438 and not w5444;
w9347 <= not w5448 and not w9346;
w9348 <= not w4999 and not w5016;
w9349 <= not w5012 and not w9348;
w9350 <= not w5035 and not w5052;
w9351 <= not w5048 and not w9350;
w9352 <= not w9349 and w9351;
w9353 <= w9349 and not w9351;
w9354 <= not w9352 and not w9353;
w9355 <= not w9347 and not w9354;
w9356 <= not w5448 and not w9352;
w9357 <= not w9353 and w9356;
w9358 <= not w9346 and w9357;
w9359 <= not w9355 and not w9358;
w9360 <= not w9345 and w9359;
w9361 <= w9345 and not w9359;
w9362 <= not w9360 and not w9361;
w9363 <= not w9331 and not w9362;
w9364 <= w9331 and w9362;
w9365 <= not w9363 and not w9364;
w9366 <= not w9329 and w9365;
w9367 <= w9329 and not w9365;
w9368 <= not w9366 and not w9367;
w9369 <= not w9293 and not w9368;
w9370 <= w9293 and w9368;
w9371 <= not w9369 and not w9370;
w9372 <= not w5350 and not w5402;
w9373 <= not w5404 and not w9372;
w9374 <= not w5343 and not w5346;
w9375 <= not w5347 and not w9374;
w9376 <= w5326 and not w5336;
w9377 <= not w5340 and not w9376;
w9378 <= not w4918 and not w4935;
w9379 <= not w4931 and not w9378;
w9380 <= not w4954 and not w4971;
w9381 <= not w4967 and not w9380;
w9382 <= not w9379 and w9381;
w9383 <= w9379 and not w9381;
w9384 <= not w9382 and not w9383;
w9385 <= not w9377 and not w9384;
w9386 <= not w5340 and not w9382;
w9387 <= not w9383 and w9386;
w9388 <= not w9376 and w9387;
w9389 <= not w9385 and not w9388;
w9390 <= w5302 and not w5308;
w9391 <= not w5312 and not w9390;
w9392 <= not w4843 and not w4860;
w9393 <= not w4856 and not w9392;
w9394 <= not w4879 and not w4896;
w9395 <= not w4892 and not w9394;
w9396 <= not w9393 and w9395;
w9397 <= w9393 and not w9395;
w9398 <= not w9396 and not w9397;
w9399 <= not w9391 and not w9398;
w9400 <= not w5312 and not w9396;
w9401 <= not w9397 and w9400;
w9402 <= not w9390 and w9401;
w9403 <= not w9399 and not w9402;
w9404 <= not w9389 and w9403;
w9405 <= w9389 and not w9403;
w9406 <= not w9404 and not w9405;
w9407 <= not w9375 and not w9406;
w9408 <= w9375 and w9406;
w9409 <= not w9407 and not w9408;
w9410 <= not w5369 and not w5390;
w9411 <= not w5392 and not w9410;
w9412 <= w5352 and not w5362;
w9413 <= not w5366 and not w9412;
w9414 <= not w4765 and not w4782;
w9415 <= not w4778 and not w9414;
w9416 <= not w4801 and not w4818;
w9417 <= not w4814 and not w9416;
w9418 <= not w9415 and w9417;
w9419 <= w9415 and not w9417;
w9420 <= not w9418 and not w9419;
w9421 <= not w9413 and not w9420;
w9422 <= not w5366 and not w9418;
w9423 <= not w9419 and w9422;
w9424 <= not w9412 and w9423;
w9425 <= not w9421 and not w9424;
w9426 <= w5371 and not w5377;
w9427 <= not w5381 and not w9426;
w9428 <= not w4690 and not w4707;
w9429 <= not w4703 and not w9428;
w9430 <= not w4726 and not w4743;
w9431 <= not w4739 and not w9430;
w9432 <= not w9429 and w9431;
w9433 <= w9429 and not w9431;
w9434 <= not w9432 and not w9433;
w9435 <= not w9427 and not w9434;
w9436 <= not w5381 and not w9432;
w9437 <= not w9433 and w9436;
w9438 <= not w9426 and w9437;
w9439 <= not w9435 and not w9438;
w9440 <= not w9425 and w9439;
w9441 <= w9425 and not w9439;
w9442 <= not w9440 and not w9441;
w9443 <= not w9411 and not w9442;
w9444 <= w9411 and w9442;
w9445 <= not w9443 and not w9444;
w9446 <= not w9409 and w9445;
w9447 <= w9409 and not w9445;
w9448 <= not w9446 and not w9447;
w9449 <= not w9373 and not w9448;
w9450 <= w9373 and w9448;
w9451 <= not w9449 and not w9450;
w9452 <= not w9371 and w9451;
w9453 <= w9371 and not w9451;
w9454 <= not w9452 and not w9453;
w9455 <= not w9291 and not w9454;
w9456 <= w9291 and w9454;
w9457 <= not w9455 and not w9456;
w9458 <= not w9289 and not w9457;
w9459 <= not w9288 and w9458;
w9460 <= not w9288 and not w9289;
w9461 <= w9457 and not w9460;
w9462 <= not w9459 and not w9461;
w9463 <= not w9048 and not w9462;
w9464 <= w9048 and w9462;
w9465 <= not w9463 and not w9464;
w9466 <= not w7269 and not w9003;
w9467 <= not w9005 and not w9466;
w9468 <= not w7262 and not w7265;
w9469 <= not w7266 and not w9468;
w9470 <= not w7255 and not w7258;
w9471 <= not w7259 and not w9470;
w9472 <= not w7248 and not w7251;
w9473 <= not w7252 and not w9472;
w9474 <= not w7241 and not w7244;
w9475 <= not w7245 and not w9474;
w9476 <= w7224 and not w7234;
w9477 <= not w7238 and not w9476;
w9478 <= not w6953 and not w6970;
w9479 <= not w6966 and not w9478;
w9480 <= not w6989 and not w7006;
w9481 <= not w7002 and not w9480;
w9482 <= not w9479 and w9481;
w9483 <= w9479 and not w9481;
w9484 <= not w9482 and not w9483;
w9485 <= not w9477 and not w9484;
w9486 <= not w7238 and not w9482;
w9487 <= not w9483 and w9486;
w9488 <= not w9476 and w9487;
w9489 <= not w9485 and not w9488;
w9490 <= w7200 and not w7206;
w9491 <= not w7210 and not w9490;
w9492 <= not w6878 and not w6895;
w9493 <= not w6891 and not w9492;
w9494 <= not w6914 and not w6931;
w9495 <= not w6927 and not w9494;
w9496 <= not w9493 and w9495;
w9497 <= w9493 and not w9495;
w9498 <= not w9496 and not w9497;
w9499 <= not w9491 and not w9498;
w9500 <= not w7210 and not w9496;
w9501 <= not w9497 and w9500;
w9502 <= not w9490 and w9501;
w9503 <= not w9499 and not w9502;
w9504 <= not w9489 and w9503;
w9505 <= w9489 and not w9503;
w9506 <= not w9504 and not w9505;
w9507 <= not w9475 and not w9506;
w9508 <= w9475 and w9506;
w9509 <= not w9507 and not w9508;
w9510 <= not w7162 and not w7183;
w9511 <= not w7185 and not w9510;
w9512 <= w7145 and not w7155;
w9513 <= not w7159 and not w9512;
w9514 <= not w6800 and not w6817;
w9515 <= not w6813 and not w9514;
w9516 <= not w6836 and not w6853;
w9517 <= not w6849 and not w9516;
w9518 <= not w9515 and w9517;
w9519 <= w9515 and not w9517;
w9520 <= not w9518 and not w9519;
w9521 <= not w9513 and not w9520;
w9522 <= not w7159 and not w9518;
w9523 <= not w9519 and w9522;
w9524 <= not w9512 and w9523;
w9525 <= not w9521 and not w9524;
w9526 <= w7164 and not w7170;
w9527 <= not w7174 and not w9526;
w9528 <= not w6725 and not w6742;
w9529 <= not w6738 and not w9528;
w9530 <= not w6761 and not w6778;
w9531 <= not w6774 and not w9530;
w9532 <= not w9529 and w9531;
w9533 <= w9529 and not w9531;
w9534 <= not w9532 and not w9533;
w9535 <= not w9527 and not w9534;
w9536 <= not w7174 and not w9532;
w9537 <= not w9533 and w9536;
w9538 <= not w9526 and w9537;
w9539 <= not w9535 and not w9538;
w9540 <= not w9525 and w9539;
w9541 <= w9525 and not w9539;
w9542 <= not w9540 and not w9541;
w9543 <= not w9511 and not w9542;
w9544 <= w9511 and w9542;
w9545 <= not w9543 and not w9544;
w9546 <= not w9509 and w9545;
w9547 <= w9509 and not w9545;
w9548 <= not w9546 and not w9547;
w9549 <= not w9473 and not w9548;
w9550 <= w9473 and w9548;
w9551 <= not w9549 and not w9550;
w9552 <= not w7076 and not w7128;
w9553 <= not w7130 and not w9552;
w9554 <= not w7069 and not w7072;
w9555 <= not w7073 and not w9554;
w9556 <= w7052 and not w7062;
w9557 <= not w7066 and not w9556;
w9558 <= not w6644 and not w6661;
w9559 <= not w6657 and not w9558;
w9560 <= not w6680 and not w6697;
w9561 <= not w6693 and not w9560;
w9562 <= not w9559 and w9561;
w9563 <= w9559 and not w9561;
w9564 <= not w9562 and not w9563;
w9565 <= not w9557 and not w9564;
w9566 <= not w7066 and not w9562;
w9567 <= not w9563 and w9566;
w9568 <= not w9556 and w9567;
w9569 <= not w9565 and not w9568;
w9570 <= w7028 and not w7034;
w9571 <= not w7038 and not w9570;
w9572 <= not w6569 and not w6586;
w9573 <= not w6582 and not w9572;
w9574 <= not w6605 and not w6622;
w9575 <= not w6618 and not w9574;
w9576 <= not w9573 and w9575;
w9577 <= w9573 and not w9575;
w9578 <= not w9576 and not w9577;
w9579 <= not w9571 and not w9578;
w9580 <= not w7038 and not w9576;
w9581 <= not w9577 and w9580;
w9582 <= not w9570 and w9581;
w9583 <= not w9579 and not w9582;
w9584 <= not w9569 and w9583;
w9585 <= w9569 and not w9583;
w9586 <= not w9584 and not w9585;
w9587 <= not w9555 and not w9586;
w9588 <= w9555 and w9586;
w9589 <= not w9587 and not w9588;
w9590 <= not w7095 and not w7116;
w9591 <= not w7118 and not w9590;
w9592 <= w7078 and not w7088;
w9593 <= not w7092 and not w9592;
w9594 <= not w6491 and not w6508;
w9595 <= not w6504 and not w9594;
w9596 <= not w6527 and not w6544;
w9597 <= not w6540 and not w9596;
w9598 <= not w9595 and w9597;
w9599 <= w9595 and not w9597;
w9600 <= not w9598 and not w9599;
w9601 <= not w9593 and not w9600;
w9602 <= not w7092 and not w9598;
w9603 <= not w9599 and w9602;
w9604 <= not w9592 and w9603;
w9605 <= not w9601 and not w9604;
w9606 <= w7097 and not w7103;
w9607 <= not w7107 and not w9606;
w9608 <= not w6416 and not w6433;
w9609 <= not w6429 and not w9608;
w9610 <= not w6452 and not w6469;
w9611 <= not w6465 and not w9610;
w9612 <= not w9609 and w9611;
w9613 <= w9609 and not w9611;
w9614 <= not w9612 and not w9613;
w9615 <= not w9607 and not w9614;
w9616 <= not w7107 and not w9612;
w9617 <= not w9613 and w9616;
w9618 <= not w9606 and w9617;
w9619 <= not w9615 and not w9618;
w9620 <= not w9605 and w9619;
w9621 <= w9605 and not w9619;
w9622 <= not w9620 and not w9621;
w9623 <= not w9591 and not w9622;
w9624 <= w9591 and w9622;
w9625 <= not w9623 and not w9624;
w9626 <= not w9589 and w9625;
w9627 <= w9589 and not w9625;
w9628 <= not w9626 and not w9627;
w9629 <= not w9553 and not w9628;
w9630 <= w9553 and w9628;
w9631 <= not w9629 and not w9630;
w9632 <= not w9551 and w9631;
w9633 <= w9551 and not w9631;
w9634 <= not w9632 and not w9633;
w9635 <= not w9471 and not w9634;
w9636 <= w9471 and w9634;
w9637 <= not w9635 and not w9636;
w9638 <= not w5961 and not w6387;
w9639 <= not w6389 and not w9638;
w9640 <= not w5954 and not w5957;
w9641 <= not w5958 and not w9640;
w9642 <= not w5947 and not w5950;
w9643 <= not w5951 and not w9642;
w9644 <= w5930 and not w5940;
w9645 <= not w5944 and not w9644;
w9646 <= not w5837 and not w5854;
w9647 <= not w5850 and not w9646;
w9648 <= not w5873 and not w5890;
w9649 <= not w5886 and not w9648;
w9650 <= not w9647 and w9649;
w9651 <= w9647 and not w9649;
w9652 <= not w9650 and not w9651;
w9653 <= not w9645 and not w9652;
w9654 <= not w5944 and not w9650;
w9655 <= not w9651 and w9654;
w9656 <= not w9644 and w9655;
w9657 <= not w9653 and not w9656;
w9658 <= w5906 and not w5912;
w9659 <= not w5916 and not w9658;
w9660 <= not w5762 and not w5779;
w9661 <= not w5775 and not w9660;
w9662 <= not w5798 and not w5815;
w9663 <= not w5811 and not w9662;
w9664 <= not w9661 and w9663;
w9665 <= w9661 and not w9663;
w9666 <= not w9664 and not w9665;
w9667 <= not w9659 and not w9666;
w9668 <= not w5916 and not w9664;
w9669 <= not w9665 and w9668;
w9670 <= not w9658 and w9669;
w9671 <= not w9667 and not w9670;
w9672 <= not w9657 and w9671;
w9673 <= w9657 and not w9671;
w9674 <= not w9672 and not w9673;
w9675 <= not w9643 and not w9674;
w9676 <= w9643 and w9674;
w9677 <= not w9675 and not w9676;
w9678 <= not w5632 and not w5733;
w9679 <= not w5735 and not w9678;
w9680 <= w5579 and not w5625;
w9681 <= not w5629 and not w9680;
w9682 <= not w5611 and not w5615;
w9683 <= not w5607 and not w9682;
w9684 <= not w5571 and not w5574;
w9685 <= not w5577 and not w9684;
w9686 <= not w9683 and w9685;
w9687 <= w9683 and not w9685;
w9688 <= not w9686 and not w9687;
w9689 <= not w9681 and not w9688;
w9690 <= not w5629 and not w9686;
w9691 <= not w9687 and w9690;
w9692 <= not w9680 and w9691;
w9693 <= not w9689 and not w9692;
w9694 <= w5668 and not w5710;
w9695 <= not w5714 and not w9694;
w9696 <= not w5700 and not w5704;
w9697 <= not w5696 and not w9696;
w9698 <= not w5660 and not w5663;
w9699 <= not w5666 and not w9698;
w9700 <= not w9697 and w9699;
w9701 <= w9697 and not w9699;
w9702 <= not w9700 and not w9701;
w9703 <= not w9695 and not w9702;
w9704 <= not w5714 and not w9700;
w9705 <= not w9701 and w9704;
w9706 <= not w9694 and w9705;
w9707 <= not w9703 and not w9706;
w9708 <= not w9693 and w9707;
w9709 <= w9693 and not w9707;
w9710 <= not w9708 and not w9709;
w9711 <= not w9679 and not w9710;
w9712 <= w9679 and w9710;
w9713 <= not w9711 and not w9712;
w9714 <= not w9677 and w9713;
w9715 <= w9677 and not w9713;
w9716 <= not w9714 and not w9715;
w9717 <= not w9641 and not w9716;
w9718 <= w9641 and w9716;
w9719 <= not w9717 and not w9718;
w9720 <= not w6161 and not w6369;
w9721 <= not w6371 and not w9720;
w9722 <= not w6154 and not w6157;
w9723 <= not w6158 and not w9722;
w9724 <= w6137 and not w6147;
w9725 <= not w6151 and not w9724;
w9726 <= not w6071 and not w6088;
w9727 <= not w6084 and not w9726;
w9728 <= not w6107 and not w6124;
w9729 <= not w6120 and not w9728;
w9730 <= not w9727 and w9729;
w9731 <= w9727 and not w9729;
w9732 <= not w9730 and not w9731;
w9733 <= not w9725 and not w9732;
w9734 <= not w6151 and not w9730;
w9735 <= not w9731 and w9734;
w9736 <= not w9724 and w9735;
w9737 <= not w9733 and not w9736;
w9738 <= w5997 and not w6039;
w9739 <= not w6043 and not w9738;
w9740 <= not w6029 and not w6033;
w9741 <= not w6025 and not w9740;
w9742 <= not w5989 and not w5992;
w9743 <= not w5995 and not w9742;
w9744 <= not w9741 and w9743;
w9745 <= w9741 and not w9743;
w9746 <= not w9744 and not w9745;
w9747 <= not w9739 and not w9746;
w9748 <= not w6043 and not w9744;
w9749 <= not w9745 and w9748;
w9750 <= not w9738 and w9749;
w9751 <= not w9747 and not w9750;
w9752 <= not w9737 and w9751;
w9753 <= w9737 and not w9751;
w9754 <= not w9752 and not w9753;
w9755 <= not w9723 and not w9754;
w9756 <= w9723 and w9754;
w9757 <= not w9755 and not w9756;
w9758 <= not w6250 and not w6351;
w9759 <= not w6353 and not w9758;
w9760 <= w6197 and not w6243;
w9761 <= not w6247 and not w9760;
w9762 <= not w6229 and not w6233;
w9763 <= not w6225 and not w9762;
w9764 <= not w6189 and not w6192;
w9765 <= not w6195 and not w9764;
w9766 <= not w9763 and w9765;
w9767 <= w9763 and not w9765;
w9768 <= not w9766 and not w9767;
w9769 <= not w9761 and not w9768;
w9770 <= not w6247 and not w9766;
w9771 <= not w9767 and w9770;
w9772 <= not w9760 and w9771;
w9773 <= not w9769 and not w9772;
w9774 <= w6286 and not w6328;
w9775 <= not w6332 and not w9774;
w9776 <= not w6318 and not w6322;
w9777 <= not w6314 and not w9776;
w9778 <= not w6278 and not w6281;
w9779 <= not w6284 and not w9778;
w9780 <= not w9777 and w9779;
w9781 <= w9777 and not w9779;
w9782 <= not w9780 and not w9781;
w9783 <= not w9775 and not w9782;
w9784 <= not w6332 and not w9780;
w9785 <= not w9781 and w9784;
w9786 <= not w9774 and w9785;
w9787 <= not w9783 and not w9786;
w9788 <= not w9773 and w9787;
w9789 <= w9773 and not w9787;
w9790 <= not w9788 and not w9789;
w9791 <= not w9759 and not w9790;
w9792 <= w9759 and w9790;
w9793 <= not w9791 and not w9792;
w9794 <= not w9757 and w9793;
w9795 <= w9757 and not w9793;
w9796 <= not w9794 and not w9795;
w9797 <= not w9721 and not w9796;
w9798 <= w9721 and w9796;
w9799 <= not w9797 and not w9798;
w9800 <= not w9719 and w9799;
w9801 <= w9719 and not w9799;
w9802 <= not w9800 and not w9801;
w9803 <= not w9639 and not w9802;
w9804 <= w9639 and w9802;
w9805 <= not w9803 and not w9804;
w9806 <= not w9637 and w9805;
w9807 <= w9637 and not w9805;
w9808 <= not w9806 and not w9807;
w9809 <= not w9469 and not w9808;
w9810 <= w9469 and w9808;
w9811 <= not w9809 and not w9810;
w9812 <= not w8123 and not w8985;
w9813 <= not w8987 and not w9812;
w9814 <= not w8116 and not w8119;
w9815 <= not w8120 and not w9814;
w9816 <= not w8109 and not w8112;
w9817 <= not w8113 and not w9816;
w9818 <= not w8102 and not w8105;
w9819 <= not w8106 and not w9818;
w9820 <= w8085 and not w8095;
w9821 <= not w8099 and not w9820;
w9822 <= not w7934 and not w7951;
w9823 <= not w7947 and not w9822;
w9824 <= not w7970 and not w7987;
w9825 <= not w7983 and not w9824;
w9826 <= not w9823 and w9825;
w9827 <= w9823 and not w9825;
w9828 <= not w9826 and not w9827;
w9829 <= not w9821 and not w9828;
w9830 <= not w8099 and not w9826;
w9831 <= not w9827 and w9830;
w9832 <= not w9820 and w9831;
w9833 <= not w9829 and not w9832;
w9834 <= w8061 and not w8067;
w9835 <= not w8071 and not w9834;
w9836 <= not w7859 and not w7876;
w9837 <= not w7872 and not w9836;
w9838 <= not w7895 and not w7912;
w9839 <= not w7908 and not w9838;
w9840 <= not w9837 and w9839;
w9841 <= w9837 and not w9839;
w9842 <= not w9840 and not w9841;
w9843 <= not w9835 and not w9842;
w9844 <= not w8071 and not w9840;
w9845 <= not w9841 and w9844;
w9846 <= not w9834 and w9845;
w9847 <= not w9843 and not w9846;
w9848 <= not w9833 and w9847;
w9849 <= w9833 and not w9847;
w9850 <= not w9848 and not w9849;
w9851 <= not w9819 and not w9850;
w9852 <= w9819 and w9850;
w9853 <= not w9851 and not w9852;
w9854 <= not w8023 and not w8044;
w9855 <= not w8046 and not w9854;
w9856 <= w8006 and not w8016;
w9857 <= not w8020 and not w9856;
w9858 <= not w7781 and not w7798;
w9859 <= not w7794 and not w9858;
w9860 <= not w7817 and not w7834;
w9861 <= not w7830 and not w9860;
w9862 <= not w9859 and w9861;
w9863 <= w9859 and not w9861;
w9864 <= not w9862 and not w9863;
w9865 <= not w9857 and not w9864;
w9866 <= not w8020 and not w9862;
w9867 <= not w9863 and w9866;
w9868 <= not w9856 and w9867;
w9869 <= not w9865 and not w9868;
w9870 <= w8025 and not w8031;
w9871 <= not w8035 and not w9870;
w9872 <= not w7706 and not w7723;
w9873 <= not w7719 and not w9872;
w9874 <= not w7742 and not w7759;
w9875 <= not w7755 and not w9874;
w9876 <= not w9873 and w9875;
w9877 <= w9873 and not w9875;
w9878 <= not w9876 and not w9877;
w9879 <= not w9871 and not w9878;
w9880 <= not w8035 and not w9876;
w9881 <= not w9877 and w9880;
w9882 <= not w9870 and w9881;
w9883 <= not w9879 and not w9882;
w9884 <= not w9869 and w9883;
w9885 <= w9869 and not w9883;
w9886 <= not w9884 and not w9885;
w9887 <= not w9855 and not w9886;
w9888 <= w9855 and w9886;
w9889 <= not w9887 and not w9888;
w9890 <= not w9853 and w9889;
w9891 <= w9853 and not w9889;
w9892 <= not w9890 and not w9891;
w9893 <= not w9817 and not w9892;
w9894 <= w9817 and w9892;
w9895 <= not w9893 and not w9894;
w9896 <= not w7469 and not w7677;
w9897 <= not w7679 and not w9896;
w9898 <= not w7462 and not w7465;
w9899 <= not w7466 and not w9898;
w9900 <= w7445 and not w7455;
w9901 <= not w7459 and not w9900;
w9902 <= not w7379 and not w7396;
w9903 <= not w7392 and not w9902;
w9904 <= not w7415 and not w7432;
w9905 <= not w7428 and not w9904;
w9906 <= not w9903 and w9905;
w9907 <= w9903 and not w9905;
w9908 <= not w9906 and not w9907;
w9909 <= not w9901 and not w9908;
w9910 <= not w7459 and not w9906;
w9911 <= not w9907 and w9910;
w9912 <= not w9900 and w9911;
w9913 <= not w9909 and not w9912;
w9914 <= w7305 and not w7347;
w9915 <= not w7351 and not w9914;
w9916 <= not w7337 and not w7341;
w9917 <= not w7333 and not w9916;
w9918 <= not w7297 and not w7300;
w9919 <= not w7303 and not w9918;
w9920 <= not w9917 and w9919;
w9921 <= w9917 and not w9919;
w9922 <= not w9920 and not w9921;
w9923 <= not w9915 and not w9922;
w9924 <= not w7351 and not w9920;
w9925 <= not w9921 and w9924;
w9926 <= not w9914 and w9925;
w9927 <= not w9923 and not w9926;
w9928 <= not w9913 and w9927;
w9929 <= w9913 and not w9927;
w9930 <= not w9928 and not w9929;
w9931 <= not w9899 and not w9930;
w9932 <= w9899 and w9930;
w9933 <= not w9931 and not w9932;
w9934 <= not w7558 and not w7659;
w9935 <= not w7661 and not w9934;
w9936 <= w7505 and not w7551;
w9937 <= not w7555 and not w9936;
w9938 <= not w7537 and not w7541;
w9939 <= not w7533 and not w9938;
w9940 <= not w7497 and not w7500;
w9941 <= not w7503 and not w9940;
w9942 <= not w9939 and w9941;
w9943 <= w9939 and not w9941;
w9944 <= not w9942 and not w9943;
w9945 <= not w9937 and not w9944;
w9946 <= not w7555 and not w9942;
w9947 <= not w9943 and w9946;
w9948 <= not w9936 and w9947;
w9949 <= not w9945 and not w9948;
w9950 <= w7594 and not w7636;
w9951 <= not w7640 and not w9950;
w9952 <= not w7626 and not w7630;
w9953 <= not w7622 and not w9952;
w9954 <= not w7586 and not w7589;
w9955 <= not w7592 and not w9954;
w9956 <= not w9953 and w9955;
w9957 <= w9953 and not w9955;
w9958 <= not w9956 and not w9957;
w9959 <= not w9951 and not w9958;
w9960 <= not w7640 and not w9956;
w9961 <= not w9957 and w9960;
w9962 <= not w9950 and w9961;
w9963 <= not w9959 and not w9962;
w9964 <= not w9949 and w9963;
w9965 <= w9949 and not w9963;
w9966 <= not w9964 and not w9965;
w9967 <= not w9935 and not w9966;
w9968 <= w9935 and w9966;
w9969 <= not w9967 and not w9968;
w9970 <= not w9933 and w9969;
w9971 <= w9933 and not w9969;
w9972 <= not w9970 and not w9971;
w9973 <= not w9897 and not w9972;
w9974 <= w9897 and w9972;
w9975 <= not w9973 and not w9974;
w9976 <= not w9895 and w9975;
w9977 <= w9895 and not w9975;
w9978 <= not w9976 and not w9977;
w9979 <= not w9815 and not w9978;
w9980 <= w9815 and w9978;
w9981 <= not w9979 and not w9980;
w9982 <= not w8541 and not w8967;
w9983 <= not w8969 and not w9982;
w9984 <= not w8534 and not w8537;
w9985 <= not w8538 and not w9984;
w9986 <= not w8527 and not w8530;
w9987 <= not w8531 and not w9986;
w9988 <= w8510 and not w8520;
w9989 <= not w8524 and not w9988;
w9990 <= not w8417 and not w8434;
w9991 <= not w8430 and not w9990;
w9992 <= not w8453 and not w8470;
w9993 <= not w8466 and not w9992;
w9994 <= not w9991 and w9993;
w9995 <= w9991 and not w9993;
w9996 <= not w9994 and not w9995;
w9997 <= not w9989 and not w9996;
w9998 <= not w8524 and not w9994;
w9999 <= not w9995 and w9998;
w10000 <= not w9988 and w9999;
w10001 <= not w9997 and not w10000;
w10002 <= w8486 and not w8492;
w10003 <= not w8496 and not w10002;
w10004 <= not w8342 and not w8359;
w10005 <= not w8355 and not w10004;
w10006 <= not w8378 and not w8395;
w10007 <= not w8391 and not w10006;
w10008 <= not w10005 and w10007;
w10009 <= w10005 and not w10007;
w10010 <= not w10008 and not w10009;
w10011 <= not w10003 and not w10010;
w10012 <= not w8496 and not w10008;
w10013 <= not w10009 and w10012;
w10014 <= not w10002 and w10013;
w10015 <= not w10011 and not w10014;
w10016 <= not w10001 and w10015;
w10017 <= w10001 and not w10015;
w10018 <= not w10016 and not w10017;
w10019 <= not w9987 and not w10018;
w10020 <= w9987 and w10018;
w10021 <= not w10019 and not w10020;
w10022 <= not w8212 and not w8313;
w10023 <= not w8315 and not w10022;
w10024 <= w8159 and not w8205;
w10025 <= not w8209 and not w10024;
w10026 <= not w8191 and not w8195;
w10027 <= not w8187 and not w10026;
w10028 <= not w8151 and not w8154;
w10029 <= not w8157 and not w10028;
w10030 <= not w10027 and w10029;
w10031 <= w10027 and not w10029;
w10032 <= not w10030 and not w10031;
w10033 <= not w10025 and not w10032;
w10034 <= not w8209 and not w10030;
w10035 <= not w10031 and w10034;
w10036 <= not w10024 and w10035;
w10037 <= not w10033 and not w10036;
w10038 <= w8248 and not w8290;
w10039 <= not w8294 and not w10038;
w10040 <= not w8280 and not w8284;
w10041 <= not w8276 and not w10040;
w10042 <= not w8240 and not w8243;
w10043 <= not w8246 and not w10042;
w10044 <= not w10041 and w10043;
w10045 <= w10041 and not w10043;
w10046 <= not w10044 and not w10045;
w10047 <= not w10039 and not w10046;
w10048 <= not w8294 and not w10044;
w10049 <= not w10045 and w10048;
w10050 <= not w10038 and w10049;
w10051 <= not w10047 and not w10050;
w10052 <= not w10037 and w10051;
w10053 <= w10037 and not w10051;
w10054 <= not w10052 and not w10053;
w10055 <= not w10023 and not w10054;
w10056 <= w10023 and w10054;
w10057 <= not w10055 and not w10056;
w10058 <= not w10021 and w10057;
w10059 <= w10021 and not w10057;
w10060 <= not w10058 and not w10059;
w10061 <= not w9985 and not w10060;
w10062 <= w9985 and w10060;
w10063 <= not w10061 and not w10062;
w10064 <= not w8741 and not w8949;
w10065 <= not w8951 and not w10064;
w10066 <= not w8734 and not w8737;
w10067 <= not w8738 and not w10066;
w10068 <= w8717 and not w8727;
w10069 <= not w8731 and not w10068;
w10070 <= not w8651 and not w8668;
w10071 <= not w8664 and not w10070;
w10072 <= not w8687 and not w8704;
w10073 <= not w8700 and not w10072;
w10074 <= not w10071 and w10073;
w10075 <= w10071 and not w10073;
w10076 <= not w10074 and not w10075;
w10077 <= not w10069 and not w10076;
w10078 <= not w8731 and not w10074;
w10079 <= not w10075 and w10078;
w10080 <= not w10068 and w10079;
w10081 <= not w10077 and not w10080;
w10082 <= w8577 and not w8619;
w10083 <= not w8623 and not w10082;
w10084 <= not w8609 and not w8613;
w10085 <= not w8605 and not w10084;
w10086 <= not w8569 and not w8572;
w10087 <= not w8575 and not w10086;
w10088 <= not w10085 and w10087;
w10089 <= w10085 and not w10087;
w10090 <= not w10088 and not w10089;
w10091 <= not w10083 and not w10090;
w10092 <= not w8623 and not w10088;
w10093 <= not w10089 and w10092;
w10094 <= not w10082 and w10093;
w10095 <= not w10091 and not w10094;
w10096 <= not w10081 and w10095;
w10097 <= w10081 and not w10095;
w10098 <= not w10096 and not w10097;
w10099 <= not w10067 and not w10098;
w10100 <= w10067 and w10098;
w10101 <= not w10099 and not w10100;
w10102 <= not w8830 and not w8931;
w10103 <= not w8933 and not w10102;
w10104 <= w8777 and not w8823;
w10105 <= not w8827 and not w10104;
w10106 <= not w8809 and not w8813;
w10107 <= not w8805 and not w10106;
w10108 <= not w8769 and not w8772;
w10109 <= not w8775 and not w10108;
w10110 <= not w10107 and w10109;
w10111 <= w10107 and not w10109;
w10112 <= not w10110 and not w10111;
w10113 <= not w10105 and not w10112;
w10114 <= not w8827 and not w10110;
w10115 <= not w10111 and w10114;
w10116 <= not w10104 and w10115;
w10117 <= not w10113 and not w10116;
w10118 <= w8866 and not w8908;
w10119 <= not w8912 and not w10118;
w10120 <= not w8898 and not w8902;
w10121 <= not w8894 and not w10120;
w10122 <= not w8858 and not w8861;
w10123 <= not w8864 and not w10122;
w10124 <= not w10121 and w10123;
w10125 <= w10121 and not w10123;
w10126 <= not w10124 and not w10125;
w10127 <= not w10119 and not w10126;
w10128 <= not w8912 and not w10124;
w10129 <= not w10125 and w10128;
w10130 <= not w10118 and w10129;
w10131 <= not w10127 and not w10130;
w10132 <= not w10117 and w10131;
w10133 <= w10117 and not w10131;
w10134 <= not w10132 and not w10133;
w10135 <= not w10103 and not w10134;
w10136 <= w10103 and w10134;
w10137 <= not w10135 and not w10136;
w10138 <= not w10101 and w10137;
w10139 <= w10101 and not w10137;
w10140 <= not w10138 and not w10139;
w10141 <= not w10065 and not w10140;
w10142 <= w10065 and w10140;
w10143 <= not w10141 and not w10142;
w10144 <= not w10063 and w10143;
w10145 <= w10063 and not w10143;
w10146 <= not w10144 and not w10145;
w10147 <= not w9983 and not w10146;
w10148 <= w9983 and w10146;
w10149 <= not w10147 and not w10148;
w10150 <= not w9981 and w10149;
w10151 <= w9981 and not w10149;
w10152 <= not w10150 and not w10151;
w10153 <= not w9813 and not w10152;
w10154 <= w9813 and w10152;
w10155 <= not w10153 and not w10154;
w10156 <= not w9811 and w10155;
w10157 <= w9811 and not w10155;
w10158 <= not w10156 and not w10157;
w10159 <= not w9467 and not w10158;
w10160 <= w9467 and w10158;
w10161 <= not w10159 and not w10160;
w10162 <= not w9465 and w10161;
w10163 <= w9465 and not w10161;
w10164 <= not w10162 and not w10163;
w10165 <= not w9046 and not w10164;
w10166 <= w9046 and w10164;
w10167 <= not w10165 and not w10166;
w10168 <= not w3462 and not w3465;
w10169 <= not w3466 and not w10168;
w10170 <= not w3455 and not w3458;
w10171 <= not w3459 and not w10170;
w10172 <= not w3448 and not w3451;
w10173 <= not w3452 and not w10172;
w10174 <= not w3441 and not w3444;
w10175 <= not w3445 and not w10174;
w10176 <= not w3434 and not w3437;
w10177 <= not w3438 and not w10176;
w10178 <= w3417 and not w3427;
w10179 <= not w3431 and not w10178;
w10180 <= not w1741 and not w1758;
w10181 <= not w1754 and not w10180;
w10182 <= not w1777 and not w1791;
w10183 <= not w1794 and not w10182;
w10184 <= not w10181 and w10183;
w10185 <= w10181 and not w10183;
w10186 <= not w10184 and not w10185;
w10187 <= not w10179 and not w10186;
w10188 <= not w3431 and not w10184;
w10189 <= not w10185 and w10188;
w10190 <= not w10178 and w10189;
w10191 <= not w10187 and not w10190;
w10192 <= w3393 and not w3399;
w10193 <= not w3403 and not w10192;
w10194 <= not w1816 and not w1833;
w10195 <= not w1829 and not w10194;
w10196 <= not w1852 and not w1869;
w10197 <= not w1865 and not w10196;
w10198 <= not w10195 and w10197;
w10199 <= w10195 and not w10197;
w10200 <= not w10198 and not w10199;
w10201 <= not w10193 and not w10200;
w10202 <= not w3403 and not w10198;
w10203 <= not w10199 and w10202;
w10204 <= not w10192 and w10203;
w10205 <= not w10201 and not w10204;
w10206 <= not w10191 and w10205;
w10207 <= w10191 and not w10205;
w10208 <= not w10206 and not w10207;
w10209 <= not w10177 and not w10208;
w10210 <= w10177 and w10208;
w10211 <= not w10209 and not w10210;
w10212 <= not w3355 and not w3376;
w10213 <= not w3378 and not w10212;
w10214 <= w3338 and not w3348;
w10215 <= not w3352 and not w10214;
w10216 <= not w1969 and not w1986;
w10217 <= not w1982 and not w10216;
w10218 <= not w2005 and not w2022;
w10219 <= not w2018 and not w10218;
w10220 <= not w10217 and w10219;
w10221 <= w10217 and not w10219;
w10222 <= not w10220 and not w10221;
w10223 <= not w10215 and not w10222;
w10224 <= not w3352 and not w10220;
w10225 <= not w10221 and w10224;
w10226 <= not w10214 and w10225;
w10227 <= not w10223 and not w10226;
w10228 <= w3357 and not w3363;
w10229 <= not w3367 and not w10228;
w10230 <= not w1894 and not w1911;
w10231 <= not w1907 and not w10230;
w10232 <= not w1930 and not w1947;
w10233 <= not w1943 and not w10232;
w10234 <= not w10231 and w10233;
w10235 <= w10231 and not w10233;
w10236 <= not w10234 and not w10235;
w10237 <= not w10229 and not w10236;
w10238 <= not w3367 and not w10234;
w10239 <= not w10235 and w10238;
w10240 <= not w10228 and w10239;
w10241 <= not w10237 and not w10240;
w10242 <= not w10227 and w10241;
w10243 <= w10227 and not w10241;
w10244 <= not w10242 and not w10243;
w10245 <= not w10213 and not w10244;
w10246 <= w10213 and w10244;
w10247 <= not w10245 and not w10246;
w10248 <= not w10211 and w10247;
w10249 <= w10211 and not w10247;
w10250 <= not w10248 and not w10249;
w10251 <= not w10175 and not w10250;
w10252 <= w10175 and w10250;
w10253 <= not w10251 and not w10252;
w10254 <= not w3269 and not w3321;
w10255 <= not w3323 and not w10254;
w10256 <= not w3262 and not w3265;
w10257 <= not w3266 and not w10256;
w10258 <= w3245 and not w3255;
w10259 <= not w3259 and not w10258;
w10260 <= not w2278 and not w2295;
w10261 <= not w2291 and not w10260;
w10262 <= not w2314 and not w2331;
w10263 <= not w2327 and not w10262;
w10264 <= not w10261 and w10263;
w10265 <= w10261 and not w10263;
w10266 <= not w10264 and not w10265;
w10267 <= not w10259 and not w10266;
w10268 <= not w3259 and not w10264;
w10269 <= not w10265 and w10268;
w10270 <= not w10258 and w10269;
w10271 <= not w10267 and not w10270;
w10272 <= w3221 and not w3227;
w10273 <= not w3231 and not w10272;
w10274 <= not w2203 and not w2220;
w10275 <= not w2216 and not w10274;
w10276 <= not w2239 and not w2256;
w10277 <= not w2252 and not w10276;
w10278 <= not w10275 and w10277;
w10279 <= w10275 and not w10277;
w10280 <= not w10278 and not w10279;
w10281 <= not w10273 and not w10280;
w10282 <= not w3231 and not w10278;
w10283 <= not w10279 and w10282;
w10284 <= not w10272 and w10283;
w10285 <= not w10281 and not w10284;
w10286 <= not w10271 and w10285;
w10287 <= w10271 and not w10285;
w10288 <= not w10286 and not w10287;
w10289 <= not w10257 and not w10288;
w10290 <= w10257 and w10288;
w10291 <= not w10289 and not w10290;
w10292 <= not w3288 and not w3309;
w10293 <= not w3311 and not w10292;
w10294 <= w3271 and not w3281;
w10295 <= not w3285 and not w10294;
w10296 <= not w2125 and not w2142;
w10297 <= not w2138 and not w10296;
w10298 <= not w2161 and not w2178;
w10299 <= not w2174 and not w10298;
w10300 <= not w10297 and w10299;
w10301 <= w10297 and not w10299;
w10302 <= not w10300 and not w10301;
w10303 <= not w10295 and not w10302;
w10304 <= not w3285 and not w10300;
w10305 <= not w10301 and w10304;
w10306 <= not w10294 and w10305;
w10307 <= not w10303 and not w10306;
w10308 <= w3290 and not w3296;
w10309 <= not w3300 and not w10308;
w10310 <= not w2050 and not w2067;
w10311 <= not w2063 and not w10310;
w10312 <= not w2086 and not w2103;
w10313 <= not w2099 and not w10312;
w10314 <= not w10311 and w10313;
w10315 <= w10311 and not w10313;
w10316 <= not w10314 and not w10315;
w10317 <= not w10309 and not w10316;
w10318 <= not w3300 and not w10314;
w10319 <= not w10315 and w10318;
w10320 <= not w10308 and w10319;
w10321 <= not w10317 and not w10320;
w10322 <= not w10307 and w10321;
w10323 <= w10307 and not w10321;
w10324 <= not w10322 and not w10323;
w10325 <= not w10293 and not w10324;
w10326 <= w10293 and w10324;
w10327 <= not w10325 and not w10326;
w10328 <= not w10291 and w10327;
w10329 <= w10291 and not w10327;
w10330 <= not w10328 and not w10329;
w10331 <= not w10255 and not w10330;
w10332 <= w10255 and w10330;
w10333 <= not w10331 and not w10332;
w10334 <= not w10253 and w10333;
w10335 <= w10253 and not w10333;
w10336 <= not w10334 and not w10335;
w10337 <= not w10173 and not w10336;
w10338 <= w10173 and w10336;
w10339 <= not w10337 and not w10338;
w10340 <= not w3090 and not w3204;
w10341 <= not w3206 and not w10340;
w10342 <= not w3083 and not w3086;
w10343 <= not w3087 and not w10342;
w10344 <= not w3076 and not w3079;
w10345 <= not w3080 and not w10344;
w10346 <= w3059 and not w3069;
w10347 <= not w3073 and not w10346;
w10348 <= not w2899 and not w2916;
w10349 <= not w2912 and not w10348;
w10350 <= not w2935 and not w2952;
w10351 <= not w2948 and not w10350;
w10352 <= not w10349 and w10351;
w10353 <= w10349 and not w10351;
w10354 <= not w10352 and not w10353;
w10355 <= not w10347 and not w10354;
w10356 <= not w3073 and not w10352;
w10357 <= not w10353 and w10356;
w10358 <= not w10346 and w10357;
w10359 <= not w10355 and not w10358;
w10360 <= w3035 and not w3041;
w10361 <= not w3045 and not w10360;
w10362 <= not w2824 and not w2841;
w10363 <= not w2837 and not w10362;
w10364 <= not w2860 and not w2877;
w10365 <= not w2873 and not w10364;
w10366 <= not w10363 and w10365;
w10367 <= w10363 and not w10365;
w10368 <= not w10366 and not w10367;
w10369 <= not w10361 and not w10368;
w10370 <= not w3045 and not w10366;
w10371 <= not w10367 and w10370;
w10372 <= not w10360 and w10371;
w10373 <= not w10369 and not w10372;
w10374 <= not w10359 and w10373;
w10375 <= w10359 and not w10373;
w10376 <= not w10374 and not w10375;
w10377 <= not w10345 and not w10376;
w10378 <= w10345 and w10376;
w10379 <= not w10377 and not w10378;
w10380 <= not w2997 and not w3018;
w10381 <= not w3020 and not w10380;
w10382 <= w2980 and not w2990;
w10383 <= not w2994 and not w10382;
w10384 <= not w2746 and not w2763;
w10385 <= not w2759 and not w10384;
w10386 <= not w2782 and not w2799;
w10387 <= not w2795 and not w10386;
w10388 <= not w10385 and w10387;
w10389 <= w10385 and not w10387;
w10390 <= not w10388 and not w10389;
w10391 <= not w10383 and not w10390;
w10392 <= not w2994 and not w10388;
w10393 <= not w10389 and w10392;
w10394 <= not w10382 and w10393;
w10395 <= not w10391 and not w10394;
w10396 <= w2999 and not w3005;
w10397 <= not w3009 and not w10396;
w10398 <= not w2671 and not w2688;
w10399 <= not w2684 and not w10398;
w10400 <= not w2707 and not w2724;
w10401 <= not w2720 and not w10400;
w10402 <= not w10399 and w10401;
w10403 <= w10399 and not w10401;
w10404 <= not w10402 and not w10403;
w10405 <= not w10397 and not w10404;
w10406 <= not w3009 and not w10402;
w10407 <= not w10403 and w10406;
w10408 <= not w10396 and w10407;
w10409 <= not w10405 and not w10408;
w10410 <= not w10395 and w10409;
w10411 <= w10395 and not w10409;
w10412 <= not w10410 and not w10411;
w10413 <= not w10381 and not w10412;
w10414 <= w10381 and w10412;
w10415 <= not w10413 and not w10414;
w10416 <= not w10379 and w10415;
w10417 <= w10379 and not w10415;
w10418 <= not w10416 and not w10417;
w10419 <= not w10343 and not w10418;
w10420 <= w10343 and w10418;
w10421 <= not w10419 and not w10420;
w10422 <= not w3140 and not w3192;
w10423 <= not w3194 and not w10422;
w10424 <= not w3133 and not w3136;
w10425 <= not w3137 and not w10424;
w10426 <= w3116 and not w3126;
w10427 <= not w3130 and not w10426;
w10428 <= not w2590 and not w2607;
w10429 <= not w2603 and not w10428;
w10430 <= not w2626 and not w2643;
w10431 <= not w2639 and not w10430;
w10432 <= not w10429 and w10431;
w10433 <= w10429 and not w10431;
w10434 <= not w10432 and not w10433;
w10435 <= not w10427 and not w10434;
w10436 <= not w3130 and not w10432;
w10437 <= not w10433 and w10436;
w10438 <= not w10426 and w10437;
w10439 <= not w10435 and not w10438;
w10440 <= w3092 and not w3098;
w10441 <= not w3102 and not w10440;
w10442 <= not w2515 and not w2532;
w10443 <= not w2528 and not w10442;
w10444 <= not w2551 and not w2568;
w10445 <= not w2564 and not w10444;
w10446 <= not w10443 and w10445;
w10447 <= w10443 and not w10445;
w10448 <= not w10446 and not w10447;
w10449 <= not w10441 and not w10448;
w10450 <= not w3102 and not w10446;
w10451 <= not w10447 and w10450;
w10452 <= not w10440 and w10451;
w10453 <= not w10449 and not w10452;
w10454 <= not w10439 and w10453;
w10455 <= w10439 and not w10453;
w10456 <= not w10454 and not w10455;
w10457 <= not w10425 and not w10456;
w10458 <= w10425 and w10456;
w10459 <= not w10457 and not w10458;
w10460 <= not w3159 and not w3180;
w10461 <= not w3182 and not w10460;
w10462 <= w3142 and not w3152;
w10463 <= not w3156 and not w10462;
w10464 <= not w2437 and not w2454;
w10465 <= not w2450 and not w10464;
w10466 <= not w2473 and not w2490;
w10467 <= not w2486 and not w10466;
w10468 <= not w10465 and w10467;
w10469 <= w10465 and not w10467;
w10470 <= not w10468 and not w10469;
w10471 <= not w10463 and not w10470;
w10472 <= not w3156 and not w10468;
w10473 <= not w10469 and w10472;
w10474 <= not w10462 and w10473;
w10475 <= not w10471 and not w10474;
w10476 <= w3161 and not w3167;
w10477 <= not w3171 and not w10476;
w10478 <= not w2362 and not w2379;
w10479 <= not w2375 and not w10478;
w10480 <= not w2398 and not w2415;
w10481 <= not w2411 and not w10480;
w10482 <= not w10479 and w10481;
w10483 <= w10479 and not w10481;
w10484 <= not w10482 and not w10483;
w10485 <= not w10477 and not w10484;
w10486 <= not w3171 and not w10482;
w10487 <= not w10483 and w10486;
w10488 <= not w10476 and w10487;
w10489 <= not w10485 and not w10488;
w10490 <= not w10475 and w10489;
w10491 <= w10475 and not w10489;
w10492 <= not w10490 and not w10491;
w10493 <= not w10461 and not w10492;
w10494 <= w10461 and w10492;
w10495 <= not w10493 and not w10494;
w10496 <= not w10459 and w10495;
w10497 <= w10459 and not w10495;
w10498 <= not w10496 and not w10497;
w10499 <= not w10423 and not w10498;
w10500 <= w10423 and w10498;
w10501 <= not w10499 and not w10500;
w10502 <= not w10421 and w10501;
w10503 <= w10421 and not w10501;
w10504 <= not w10502 and not w10503;
w10505 <= not w10341 and not w10504;
w10506 <= w10341 and w10504;
w10507 <= not w10505 and not w10506;
w10508 <= not w10339 and w10507;
w10509 <= w10339 and not w10507;
w10510 <= not w10508 and not w10509;
w10511 <= not w10171 and not w10510;
w10512 <= w10171 and w10510;
w10513 <= not w10511 and not w10512;
w10514 <= not w853 and not w1715;
w10515 <= not w1717 and not w10514;
w10516 <= not w846 and not w849;
w10517 <= not w850 and not w10516;
w10518 <= not w839 and not w842;
w10519 <= not w843 and not w10518;
w10520 <= not w832 and not w835;
w10521 <= not w836 and not w10520;
w10522 <= w815 and not w825;
w10523 <= not w829 and not w10522;
w10524 <= not w664 and not w681;
w10525 <= not w677 and not w10524;
w10526 <= not w700 and not w717;
w10527 <= not w713 and not w10526;
w10528 <= not w10525 and w10527;
w10529 <= w10525 and not w10527;
w10530 <= not w10528 and not w10529;
w10531 <= not w10523 and not w10530;
w10532 <= not w829 and not w10528;
w10533 <= not w10529 and w10532;
w10534 <= not w10522 and w10533;
w10535 <= not w10531 and not w10534;
w10536 <= w791 and not w797;
w10537 <= not w801 and not w10536;
w10538 <= not w589 and not w606;
w10539 <= not w602 and not w10538;
w10540 <= not w625 and not w642;
w10541 <= not w638 and not w10540;
w10542 <= not w10539 and w10541;
w10543 <= w10539 and not w10541;
w10544 <= not w10542 and not w10543;
w10545 <= not w10537 and not w10544;
w10546 <= not w801 and not w10542;
w10547 <= not w10543 and w10546;
w10548 <= not w10536 and w10547;
w10549 <= not w10545 and not w10548;
w10550 <= not w10535 and w10549;
w10551 <= w10535 and not w10549;
w10552 <= not w10550 and not w10551;
w10553 <= not w10521 and not w10552;
w10554 <= w10521 and w10552;
w10555 <= not w10553 and not w10554;
w10556 <= not w753 and not w774;
w10557 <= not w776 and not w10556;
w10558 <= w736 and not w746;
w10559 <= not w750 and not w10558;
w10560 <= not w511 and not w528;
w10561 <= not w524 and not w10560;
w10562 <= not w547 and not w564;
w10563 <= not w560 and not w10562;
w10564 <= not w10561 and w10563;
w10565 <= w10561 and not w10563;
w10566 <= not w10564 and not w10565;
w10567 <= not w10559 and not w10566;
w10568 <= not w750 and not w10564;
w10569 <= not w10565 and w10568;
w10570 <= not w10558 and w10569;
w10571 <= not w10567 and not w10570;
w10572 <= w755 and not w761;
w10573 <= not w765 and not w10572;
w10574 <= not w436 and not w453;
w10575 <= not w449 and not w10574;
w10576 <= not w472 and not w489;
w10577 <= not w485 and not w10576;
w10578 <= not w10575 and w10577;
w10579 <= w10575 and not w10577;
w10580 <= not w10578 and not w10579;
w10581 <= not w10573 and not w10580;
w10582 <= not w765 and not w10578;
w10583 <= not w10579 and w10582;
w10584 <= not w10572 and w10583;
w10585 <= not w10581 and not w10584;
w10586 <= not w10571 and w10585;
w10587 <= w10571 and not w10585;
w10588 <= not w10586 and not w10587;
w10589 <= not w10557 and not w10588;
w10590 <= w10557 and w10588;
w10591 <= not w10589 and not w10590;
w10592 <= not w10555 and w10591;
w10593 <= w10555 and not w10591;
w10594 <= not w10592 and not w10593;
w10595 <= not w10519 and not w10594;
w10596 <= w10519 and w10594;
w10597 <= not w10595 and not w10596;
w10598 <= not w199 and not w407;
w10599 <= not w409 and not w10598;
w10600 <= not w192 and not w195;
w10601 <= not w196 and not w10600;
w10602 <= w175 and not w185;
w10603 <= not w189 and not w10602;
w10604 <= not w109 and not w126;
w10605 <= not w122 and not w10604;
w10606 <= not w145 and not w162;
w10607 <= not w158 and not w10606;
w10608 <= not w10605 and w10607;
w10609 <= w10605 and not w10607;
w10610 <= not w10608 and not w10609;
w10611 <= not w10603 and not w10610;
w10612 <= not w189 and not w10608;
w10613 <= not w10609 and w10612;
w10614 <= not w10602 and w10613;
w10615 <= not w10611 and not w10614;
w10616 <= w35 and not w77;
w10617 <= not w81 and not w10616;
w10618 <= not w67 and not w71;
w10619 <= not w63 and not w10618;
w10620 <= not w27 and not w30;
w10621 <= not w33 and not w10620;
w10622 <= not w10619 and w10621;
w10623 <= w10619 and not w10621;
w10624 <= not w10622 and not w10623;
w10625 <= not w10617 and not w10624;
w10626 <= not w81 and not w10622;
w10627 <= not w10623 and w10626;
w10628 <= not w10616 and w10627;
w10629 <= not w10625 and not w10628;
w10630 <= not w10615 and w10629;
w10631 <= w10615 and not w10629;
w10632 <= not w10630 and not w10631;
w10633 <= not w10601 and not w10632;
w10634 <= w10601 and w10632;
w10635 <= not w10633 and not w10634;
w10636 <= not w288 and not w389;
w10637 <= not w391 and not w10636;
w10638 <= w235 and not w281;
w10639 <= not w285 and not w10638;
w10640 <= not w267 and not w271;
w10641 <= not w263 and not w10640;
w10642 <= not w227 and not w230;
w10643 <= not w233 and not w10642;
w10644 <= not w10641 and w10643;
w10645 <= w10641 and not w10643;
w10646 <= not w10644 and not w10645;
w10647 <= not w10639 and not w10646;
w10648 <= not w285 and not w10644;
w10649 <= not w10645 and w10648;
w10650 <= not w10638 and w10649;
w10651 <= not w10647 and not w10650;
w10652 <= w324 and not w366;
w10653 <= not w370 and not w10652;
w10654 <= not w356 and not w360;
w10655 <= not w352 and not w10654;
w10656 <= not w316 and not w319;
w10657 <= not w322 and not w10656;
w10658 <= not w10655 and w10657;
w10659 <= w10655 and not w10657;
w10660 <= not w10658 and not w10659;
w10661 <= not w10653 and not w10660;
w10662 <= not w370 and not w10658;
w10663 <= not w10659 and w10662;
w10664 <= not w10652 and w10663;
w10665 <= not w10661 and not w10664;
w10666 <= not w10651 and w10665;
w10667 <= w10651 and not w10665;
w10668 <= not w10666 and not w10667;
w10669 <= not w10637 and not w10668;
w10670 <= w10637 and w10668;
w10671 <= not w10669 and not w10670;
w10672 <= not w10635 and w10671;
w10673 <= w10635 and not w10671;
w10674 <= not w10672 and not w10673;
w10675 <= not w10599 and not w10674;
w10676 <= w10599 and w10674;
w10677 <= not w10675 and not w10676;
w10678 <= not w10597 and w10677;
w10679 <= w10597 and not w10677;
w10680 <= not w10678 and not w10679;
w10681 <= not w10517 and not w10680;
w10682 <= w10517 and w10680;
w10683 <= not w10681 and not w10682;
w10684 <= not w1271 and not w1697;
w10685 <= not w1699 and not w10684;
w10686 <= not w1264 and not w1267;
w10687 <= not w1268 and not w10686;
w10688 <= not w1257 and not w1260;
w10689 <= not w1261 and not w10688;
w10690 <= w1240 and not w1250;
w10691 <= not w1254 and not w10690;
w10692 <= not w1147 and not w1164;
w10693 <= not w1160 and not w10692;
w10694 <= not w1183 and not w1200;
w10695 <= not w1196 and not w10694;
w10696 <= not w10693 and w10695;
w10697 <= w10693 and not w10695;
w10698 <= not w10696 and not w10697;
w10699 <= not w10691 and not w10698;
w10700 <= not w1254 and not w10696;
w10701 <= not w10697 and w10700;
w10702 <= not w10690 and w10701;
w10703 <= not w10699 and not w10702;
w10704 <= w1216 and not w1222;
w10705 <= not w1226 and not w10704;
w10706 <= not w1072 and not w1089;
w10707 <= not w1085 and not w10706;
w10708 <= not w1108 and not w1125;
w10709 <= not w1121 and not w10708;
w10710 <= not w10707 and w10709;
w10711 <= w10707 and not w10709;
w10712 <= not w10710 and not w10711;
w10713 <= not w10705 and not w10712;
w10714 <= not w1226 and not w10710;
w10715 <= not w10711 and w10714;
w10716 <= not w10704 and w10715;
w10717 <= not w10713 and not w10716;
w10718 <= not w10703 and w10717;
w10719 <= w10703 and not w10717;
w10720 <= not w10718 and not w10719;
w10721 <= not w10689 and not w10720;
w10722 <= w10689 and w10720;
w10723 <= not w10721 and not w10722;
w10724 <= not w942 and not w1043;
w10725 <= not w1045 and not w10724;
w10726 <= w889 and not w935;
w10727 <= not w939 and not w10726;
w10728 <= not w921 and not w925;
w10729 <= not w917 and not w10728;
w10730 <= not w881 and not w884;
w10731 <= not w887 and not w10730;
w10732 <= not w10729 and w10731;
w10733 <= w10729 and not w10731;
w10734 <= not w10732 and not w10733;
w10735 <= not w10727 and not w10734;
w10736 <= not w939 and not w10732;
w10737 <= not w10733 and w10736;
w10738 <= not w10726 and w10737;
w10739 <= not w10735 and not w10738;
w10740 <= w978 and not w1020;
w10741 <= not w1024 and not w10740;
w10742 <= not w1010 and not w1014;
w10743 <= not w1006 and not w10742;
w10744 <= not w970 and not w973;
w10745 <= not w976 and not w10744;
w10746 <= not w10743 and w10745;
w10747 <= w10743 and not w10745;
w10748 <= not w10746 and not w10747;
w10749 <= not w10741 and not w10748;
w10750 <= not w1024 and not w10746;
w10751 <= not w10747 and w10750;
w10752 <= not w10740 and w10751;
w10753 <= not w10749 and not w10752;
w10754 <= not w10739 and w10753;
w10755 <= w10739 and not w10753;
w10756 <= not w10754 and not w10755;
w10757 <= not w10725 and not w10756;
w10758 <= w10725 and w10756;
w10759 <= not w10757 and not w10758;
w10760 <= not w10723 and w10759;
w10761 <= w10723 and not w10759;
w10762 <= not w10760 and not w10761;
w10763 <= not w10687 and not w10762;
w10764 <= w10687 and w10762;
w10765 <= not w10763 and not w10764;
w10766 <= not w1471 and not w1679;
w10767 <= not w1681 and not w10766;
w10768 <= not w1464 and not w1467;
w10769 <= not w1468 and not w10768;
w10770 <= w1447 and not w1457;
w10771 <= not w1461 and not w10770;
w10772 <= not w1381 and not w1398;
w10773 <= not w1394 and not w10772;
w10774 <= not w1417 and not w1434;
w10775 <= not w1430 and not w10774;
w10776 <= not w10773 and w10775;
w10777 <= w10773 and not w10775;
w10778 <= not w10776 and not w10777;
w10779 <= not w10771 and not w10778;
w10780 <= not w1461 and not w10776;
w10781 <= not w10777 and w10780;
w10782 <= not w10770 and w10781;
w10783 <= not w10779 and not w10782;
w10784 <= w1307 and not w1349;
w10785 <= not w1353 and not w10784;
w10786 <= not w1339 and not w1343;
w10787 <= not w1335 and not w10786;
w10788 <= not w1299 and not w1302;
w10789 <= not w1305 and not w10788;
w10790 <= not w10787 and w10789;
w10791 <= w10787 and not w10789;
w10792 <= not w10790 and not w10791;
w10793 <= not w10785 and not w10792;
w10794 <= not w1353 and not w10790;
w10795 <= not w10791 and w10794;
w10796 <= not w10784 and w10795;
w10797 <= not w10793 and not w10796;
w10798 <= not w10783 and w10797;
w10799 <= w10783 and not w10797;
w10800 <= not w10798 and not w10799;
w10801 <= not w10769 and not w10800;
w10802 <= w10769 and w10800;
w10803 <= not w10801 and not w10802;
w10804 <= not w1560 and not w1661;
w10805 <= not w1663 and not w10804;
w10806 <= w1507 and not w1553;
w10807 <= not w1557 and not w10806;
w10808 <= not w1539 and not w1543;
w10809 <= not w1535 and not w10808;
w10810 <= not w1499 and not w1502;
w10811 <= not w1505 and not w10810;
w10812 <= not w10809 and w10811;
w10813 <= w10809 and not w10811;
w10814 <= not w10812 and not w10813;
w10815 <= not w10807 and not w10814;
w10816 <= not w1557 and not w10812;
w10817 <= not w10813 and w10816;
w10818 <= not w10806 and w10817;
w10819 <= not w10815 and not w10818;
w10820 <= w1596 and not w1638;
w10821 <= not w1642 and not w10820;
w10822 <= not w1628 and not w1632;
w10823 <= not w1624 and not w10822;
w10824 <= not w1588 and not w1591;
w10825 <= not w1594 and not w10824;
w10826 <= not w10823 and w10825;
w10827 <= w10823 and not w10825;
w10828 <= not w10826 and not w10827;
w10829 <= not w10821 and not w10828;
w10830 <= not w1642 and not w10826;
w10831 <= not w10827 and w10830;
w10832 <= not w10820 and w10831;
w10833 <= not w10829 and not w10832;
w10834 <= not w10819 and w10833;
w10835 <= w10819 and not w10833;
w10836 <= not w10834 and not w10835;
w10837 <= not w10805 and not w10836;
w10838 <= w10805 and w10836;
w10839 <= not w10837 and not w10838;
w10840 <= not w10803 and w10839;
w10841 <= w10803 and not w10839;
w10842 <= not w10840 and not w10841;
w10843 <= not w10767 and not w10842;
w10844 <= w10767 and w10842;
w10845 <= not w10843 and not w10844;
w10846 <= not w10765 and w10845;
w10847 <= w10765 and not w10845;
w10848 <= not w10846 and not w10847;
w10849 <= not w10685 and not w10848;
w10850 <= w10685 and w10848;
w10851 <= not w10849 and not w10850;
w10852 <= not w10683 and w10851;
w10853 <= w10683 and not w10851;
w10854 <= not w10852 and not w10853;
w10855 <= not w10515 and not w10854;
w10856 <= w10515 and w10854;
w10857 <= not w10855 and not w10856;
w10858 <= not w10513 and w10857;
w10859 <= w10513 and not w10857;
w10860 <= not w10858 and not w10859;
w10861 <= not w10169 and not w10860;
w10862 <= w10169 and w10860;
w10863 <= not w10861 and not w10862;
w10864 <= not w10167 and not w10863;
w10865 <= not w9044 and not w10864;
w10866 <= not w10165 and w10863;
w10867 <= not w10166 and w10866;
w10868 <= not w10865 and not w10867;
w10869 <= not w9465 and not w10161;
w10870 <= not w9046 and not w10869;
w10871 <= w9465 and w10161;
w10872 <= not w10870 and not w10871;
w10873 <= not w9811 and not w10155;
w10874 <= not w9467 and not w10873;
w10875 <= w9811 and w10155;
w10876 <= not w10874 and not w10875;
w10877 <= not w9981 and not w10149;
w10878 <= not w9813 and not w10877;
w10879 <= w9981 and w10149;
w10880 <= not w10878 and not w10879;
w10881 <= not w10063 and not w10143;
w10882 <= not w9983 and not w10881;
w10883 <= w10063 and w10143;
w10884 <= not w10882 and not w10883;
w10885 <= not w10101 and not w10137;
w10886 <= not w10065 and not w10885;
w10887 <= w10101 and w10137;
w10888 <= not w10886 and not w10887;
w10889 <= not w10117 and not w10131;
w10890 <= not w10103 and not w10889;
w10891 <= not w10116 and not w10130;
w10892 <= not w10127 and w10891;
w10893 <= not w10113 and w10892;
w10894 <= not w10890 and not w10893;
w10895 <= not w8912 and not w10121;
w10896 <= not w10118 and w10895;
w10897 <= w10123 and not w10896;
w10898 <= not w10119 and w10121;
w10899 <= not w10897 and not w10898;
w10900 <= not w8827 and not w10107;
w10901 <= not w10104 and w10900;
w10902 <= w10109 and not w10901;
w10903 <= not w10105 and w10107;
w10904 <= not w10902 and not w10903;
w10905 <= not w10899 and w10904;
w10906 <= w10899 and not w10904;
w10907 <= not w10905 and not w10906;
w10908 <= not w10894 and not w10907;
w10909 <= not w10893 and not w10905;
w10910 <= not w10906 and w10909;
w10911 <= not w10890 and w10910;
w10912 <= not w10908 and not w10911;
w10913 <= not w10081 and not w10095;
w10914 <= not w10067 and not w10913;
w10915 <= not w10080 and not w10094;
w10916 <= not w10091 and w10915;
w10917 <= not w10077 and w10916;
w10918 <= not w10914 and not w10917;
w10919 <= not w8623 and not w10085;
w10920 <= not w10082 and w10919;
w10921 <= w10087 and not w10920;
w10922 <= not w10083 and w10085;
w10923 <= not w10921 and not w10922;
w10924 <= not w8731 and not w10071;
w10925 <= not w10068 and w10924;
w10926 <= w10073 and not w10925;
w10927 <= not w10069 and w10071;
w10928 <= not w10926 and not w10927;
w10929 <= not w10923 and w10928;
w10930 <= w10923 and not w10928;
w10931 <= not w10929 and not w10930;
w10932 <= not w10918 and not w10931;
w10933 <= not w10917 and not w10929;
w10934 <= not w10930 and w10933;
w10935 <= not w10914 and w10934;
w10936 <= not w10932 and not w10935;
w10937 <= not w10912 and w10936;
w10938 <= w10912 and not w10936;
w10939 <= not w10937 and not w10938;
w10940 <= not w10888 and not w10939;
w10941 <= w10888 and w10939;
w10942 <= not w10940 and not w10941;
w10943 <= not w10021 and not w10057;
w10944 <= not w9985 and not w10943;
w10945 <= w10021 and w10057;
w10946 <= not w10944 and not w10945;
w10947 <= not w10037 and not w10051;
w10948 <= not w10023 and not w10947;
w10949 <= not w10036 and not w10050;
w10950 <= not w10047 and w10949;
w10951 <= not w10033 and w10950;
w10952 <= not w10948 and not w10951;
w10953 <= not w8294 and not w10041;
w10954 <= not w10038 and w10953;
w10955 <= w10043 and not w10954;
w10956 <= not w10039 and w10041;
w10957 <= not w10955 and not w10956;
w10958 <= not w8209 and not w10027;
w10959 <= not w10024 and w10958;
w10960 <= w10029 and not w10959;
w10961 <= not w10025 and w10027;
w10962 <= not w10960 and not w10961;
w10963 <= not w10957 and w10962;
w10964 <= w10957 and not w10962;
w10965 <= not w10963 and not w10964;
w10966 <= not w10952 and not w10965;
w10967 <= not w10951 and not w10963;
w10968 <= not w10964 and w10967;
w10969 <= not w10948 and w10968;
w10970 <= not w10966 and not w10969;
w10971 <= not w10001 and not w10015;
w10972 <= not w9987 and not w10971;
w10973 <= not w10000 and not w10014;
w10974 <= not w10011 and w10973;
w10975 <= not w9997 and w10974;
w10976 <= not w10972 and not w10975;
w10977 <= not w8496 and not w10005;
w10978 <= not w10002 and w10977;
w10979 <= w10007 and not w10978;
w10980 <= not w10003 and w10005;
w10981 <= not w10979 and not w10980;
w10982 <= not w8524 and not w9991;
w10983 <= not w9988 and w10982;
w10984 <= w9993 and not w10983;
w10985 <= not w9989 and w9991;
w10986 <= not w10984 and not w10985;
w10987 <= not w10981 and w10986;
w10988 <= w10981 and not w10986;
w10989 <= not w10987 and not w10988;
w10990 <= not w10976 and not w10989;
w10991 <= not w10975 and not w10987;
w10992 <= not w10988 and w10991;
w10993 <= not w10972 and w10992;
w10994 <= not w10990 and not w10993;
w10995 <= not w10970 and w10994;
w10996 <= w10970 and not w10994;
w10997 <= not w10995 and not w10996;
w10998 <= not w10946 and not w10997;
w10999 <= w10946 and w10997;
w11000 <= not w10998 and not w10999;
w11001 <= not w10942 and w11000;
w11002 <= w10942 and not w11000;
w11003 <= not w11001 and not w11002;
w11004 <= not w10884 and not w11003;
w11005 <= w10884 and w11003;
w11006 <= not w11004 and not w11005;
w11007 <= not w9895 and not w9975;
w11008 <= not w9815 and not w11007;
w11009 <= w9895 and w9975;
w11010 <= not w11008 and not w11009;
w11011 <= not w9933 and not w9969;
w11012 <= not w9897 and not w11011;
w11013 <= w9933 and w9969;
w11014 <= not w11012 and not w11013;
w11015 <= not w9949 and not w9963;
w11016 <= not w9935 and not w11015;
w11017 <= not w9948 and not w9962;
w11018 <= not w9959 and w11017;
w11019 <= not w9945 and w11018;
w11020 <= not w11016 and not w11019;
w11021 <= not w7640 and not w9953;
w11022 <= not w9950 and w11021;
w11023 <= w9955 and not w11022;
w11024 <= not w9951 and w9953;
w11025 <= not w11023 and not w11024;
w11026 <= not w7555 and not w9939;
w11027 <= not w9936 and w11026;
w11028 <= w9941 and not w11027;
w11029 <= not w9937 and w9939;
w11030 <= not w11028 and not w11029;
w11031 <= not w11025 and w11030;
w11032 <= w11025 and not w11030;
w11033 <= not w11031 and not w11032;
w11034 <= not w11020 and not w11033;
w11035 <= not w11019 and not w11031;
w11036 <= not w11032 and w11035;
w11037 <= not w11016 and w11036;
w11038 <= not w11034 and not w11037;
w11039 <= not w9913 and not w9927;
w11040 <= not w9899 and not w11039;
w11041 <= not w9912 and not w9926;
w11042 <= not w9923 and w11041;
w11043 <= not w9909 and w11042;
w11044 <= not w11040 and not w11043;
w11045 <= not w7351 and not w9917;
w11046 <= not w9914 and w11045;
w11047 <= w9919 and not w11046;
w11048 <= not w9915 and w9917;
w11049 <= not w11047 and not w11048;
w11050 <= not w7459 and not w9903;
w11051 <= not w9900 and w11050;
w11052 <= w9905 and not w11051;
w11053 <= not w9901 and w9903;
w11054 <= not w11052 and not w11053;
w11055 <= not w11049 and w11054;
w11056 <= w11049 and not w11054;
w11057 <= not w11055 and not w11056;
w11058 <= not w11044 and not w11057;
w11059 <= not w11043 and not w11055;
w11060 <= not w11056 and w11059;
w11061 <= not w11040 and w11060;
w11062 <= not w11058 and not w11061;
w11063 <= not w11038 and w11062;
w11064 <= w11038 and not w11062;
w11065 <= not w11063 and not w11064;
w11066 <= not w11014 and not w11065;
w11067 <= w11014 and w11065;
w11068 <= not w11066 and not w11067;
w11069 <= not w9853 and not w9889;
w11070 <= not w9817 and not w11069;
w11071 <= w9853 and w9889;
w11072 <= not w11070 and not w11071;
w11073 <= not w9869 and not w9883;
w11074 <= not w9855 and not w11073;
w11075 <= not w9868 and not w9882;
w11076 <= not w9879 and w11075;
w11077 <= not w9865 and w11076;
w11078 <= not w11074 and not w11077;
w11079 <= not w8035 and not w9873;
w11080 <= not w9870 and w11079;
w11081 <= w9875 and not w11080;
w11082 <= not w9871 and w9873;
w11083 <= not w11081 and not w11082;
w11084 <= not w8020 and not w9859;
w11085 <= not w9856 and w11084;
w11086 <= w9861 and not w11085;
w11087 <= not w9857 and w9859;
w11088 <= not w11086 and not w11087;
w11089 <= not w11083 and w11088;
w11090 <= w11083 and not w11088;
w11091 <= not w11089 and not w11090;
w11092 <= not w11078 and not w11091;
w11093 <= not w11077 and not w11089;
w11094 <= not w11090 and w11093;
w11095 <= not w11074 and w11094;
w11096 <= not w11092 and not w11095;
w11097 <= not w9833 and not w9847;
w11098 <= not w9819 and not w11097;
w11099 <= not w9832 and not w9846;
w11100 <= not w9843 and w11099;
w11101 <= not w9829 and w11100;
w11102 <= not w11098 and not w11101;
w11103 <= not w8071 and not w9837;
w11104 <= not w9834 and w11103;
w11105 <= w9839 and not w11104;
w11106 <= not w9835 and w9837;
w11107 <= not w11105 and not w11106;
w11108 <= not w8099 and not w9823;
w11109 <= not w9820 and w11108;
w11110 <= w9825 and not w11109;
w11111 <= not w9821 and w9823;
w11112 <= not w11110 and not w11111;
w11113 <= not w11107 and w11112;
w11114 <= w11107 and not w11112;
w11115 <= not w11113 and not w11114;
w11116 <= not w11102 and not w11115;
w11117 <= not w11101 and not w11113;
w11118 <= not w11114 and w11117;
w11119 <= not w11098 and w11118;
w11120 <= not w11116 and not w11119;
w11121 <= not w11096 and w11120;
w11122 <= w11096 and not w11120;
w11123 <= not w11121 and not w11122;
w11124 <= not w11072 and not w11123;
w11125 <= w11072 and w11123;
w11126 <= not w11124 and not w11125;
w11127 <= not w11068 and w11126;
w11128 <= w11068 and not w11126;
w11129 <= not w11127 and not w11128;
w11130 <= not w11010 and not w11129;
w11131 <= w11010 and w11129;
w11132 <= not w11130 and not w11131;
w11133 <= not w11006 and w11132;
w11134 <= w11006 and not w11132;
w11135 <= not w11133 and not w11134;
w11136 <= not w10880 and not w11135;
w11137 <= w10880 and w11135;
w11138 <= not w11136 and not w11137;
w11139 <= not w9637 and not w9805;
w11140 <= not w9469 and not w11139;
w11141 <= w9637 and w9805;
w11142 <= not w11140 and not w11141;
w11143 <= not w9719 and not w9799;
w11144 <= not w9639 and not w11143;
w11145 <= w9719 and w9799;
w11146 <= not w11144 and not w11145;
w11147 <= not w9757 and not w9793;
w11148 <= not w9721 and not w11147;
w11149 <= w9757 and w9793;
w11150 <= not w11148 and not w11149;
w11151 <= not w9773 and not w9787;
w11152 <= not w9759 and not w11151;
w11153 <= not w9772 and not w9786;
w11154 <= not w9783 and w11153;
w11155 <= not w9769 and w11154;
w11156 <= not w11152 and not w11155;
w11157 <= not w6332 and not w9777;
w11158 <= not w9774 and w11157;
w11159 <= w9779 and not w11158;
w11160 <= not w9775 and w9777;
w11161 <= not w11159 and not w11160;
w11162 <= not w6247 and not w9763;
w11163 <= not w9760 and w11162;
w11164 <= w9765 and not w11163;
w11165 <= not w9761 and w9763;
w11166 <= not w11164 and not w11165;
w11167 <= not w11161 and w11166;
w11168 <= w11161 and not w11166;
w11169 <= not w11167 and not w11168;
w11170 <= not w11156 and not w11169;
w11171 <= not w11155 and not w11167;
w11172 <= not w11168 and w11171;
w11173 <= not w11152 and w11172;
w11174 <= not w11170 and not w11173;
w11175 <= not w9737 and not w9751;
w11176 <= not w9723 and not w11175;
w11177 <= not w9736 and not w9750;
w11178 <= not w9747 and w11177;
w11179 <= not w9733 and w11178;
w11180 <= not w11176 and not w11179;
w11181 <= not w6043 and not w9741;
w11182 <= not w9738 and w11181;
w11183 <= w9743 and not w11182;
w11184 <= not w9739 and w9741;
w11185 <= not w11183 and not w11184;
w11186 <= not w6151 and not w9727;
w11187 <= not w9724 and w11186;
w11188 <= w9729 and not w11187;
w11189 <= not w9725 and w9727;
w11190 <= not w11188 and not w11189;
w11191 <= not w11185 and w11190;
w11192 <= w11185 and not w11190;
w11193 <= not w11191 and not w11192;
w11194 <= not w11180 and not w11193;
w11195 <= not w11179 and not w11191;
w11196 <= not w11192 and w11195;
w11197 <= not w11176 and w11196;
w11198 <= not w11194 and not w11197;
w11199 <= not w11174 and w11198;
w11200 <= w11174 and not w11198;
w11201 <= not w11199 and not w11200;
w11202 <= not w11150 and not w11201;
w11203 <= w11150 and w11201;
w11204 <= not w11202 and not w11203;
w11205 <= not w9677 and not w9713;
w11206 <= not w9641 and not w11205;
w11207 <= w9677 and w9713;
w11208 <= not w11206 and not w11207;
w11209 <= not w9693 and not w9707;
w11210 <= not w9679 and not w11209;
w11211 <= not w9692 and not w9706;
w11212 <= not w9703 and w11211;
w11213 <= not w9689 and w11212;
w11214 <= not w11210 and not w11213;
w11215 <= not w5714 and not w9697;
w11216 <= not w9694 and w11215;
w11217 <= w9699 and not w11216;
w11218 <= not w9695 and w9697;
w11219 <= not w11217 and not w11218;
w11220 <= not w5629 and not w9683;
w11221 <= not w9680 and w11220;
w11222 <= w9685 and not w11221;
w11223 <= not w9681 and w9683;
w11224 <= not w11222 and not w11223;
w11225 <= not w11219 and w11224;
w11226 <= w11219 and not w11224;
w11227 <= not w11225 and not w11226;
w11228 <= not w11214 and not w11227;
w11229 <= not w11213 and not w11225;
w11230 <= not w11226 and w11229;
w11231 <= not w11210 and w11230;
w11232 <= not w11228 and not w11231;
w11233 <= not w9657 and not w9671;
w11234 <= not w9643 and not w11233;
w11235 <= not w9656 and not w9670;
w11236 <= not w9667 and w11235;
w11237 <= not w9653 and w11236;
w11238 <= not w11234 and not w11237;
w11239 <= not w5916 and not w9661;
w11240 <= not w9658 and w11239;
w11241 <= w9663 and not w11240;
w11242 <= not w9659 and w9661;
w11243 <= not w11241 and not w11242;
w11244 <= not w5944 and not w9647;
w11245 <= not w9644 and w11244;
w11246 <= w9649 and not w11245;
w11247 <= not w9645 and w9647;
w11248 <= not w11246 and not w11247;
w11249 <= not w11243 and w11248;
w11250 <= w11243 and not w11248;
w11251 <= not w11249 and not w11250;
w11252 <= not w11238 and not w11251;
w11253 <= not w11237 and not w11249;
w11254 <= not w11250 and w11253;
w11255 <= not w11234 and w11254;
w11256 <= not w11252 and not w11255;
w11257 <= not w11232 and w11256;
w11258 <= w11232 and not w11256;
w11259 <= not w11257 and not w11258;
w11260 <= not w11208 and not w11259;
w11261 <= w11208 and w11259;
w11262 <= not w11260 and not w11261;
w11263 <= not w11204 and w11262;
w11264 <= w11204 and not w11262;
w11265 <= not w11263 and not w11264;
w11266 <= not w11146 and not w11265;
w11267 <= w11146 and w11265;
w11268 <= not w11266 and not w11267;
w11269 <= not w9551 and not w9631;
w11270 <= not w9471 and not w11269;
w11271 <= w9551 and w9631;
w11272 <= not w11270 and not w11271;
w11273 <= not w9589 and not w9625;
w11274 <= not w9553 and not w11273;
w11275 <= w9589 and w9625;
w11276 <= not w11274 and not w11275;
w11277 <= not w9605 and not w9619;
w11278 <= not w9591 and not w11277;
w11279 <= not w9604 and not w9618;
w11280 <= not w9615 and w11279;
w11281 <= not w9601 and w11280;
w11282 <= not w11278 and not w11281;
w11283 <= not w7107 and not w9609;
w11284 <= not w9606 and w11283;
w11285 <= w9611 and not w11284;
w11286 <= not w9607 and w9609;
w11287 <= not w11285 and not w11286;
w11288 <= not w7092 and not w9595;
w11289 <= not w9592 and w11288;
w11290 <= w9597 and not w11289;
w11291 <= not w9593 and w9595;
w11292 <= not w11290 and not w11291;
w11293 <= not w11287 and w11292;
w11294 <= w11287 and not w11292;
w11295 <= not w11293 and not w11294;
w11296 <= not w11282 and not w11295;
w11297 <= not w11281 and not w11293;
w11298 <= not w11294 and w11297;
w11299 <= not w11278 and w11298;
w11300 <= not w11296 and not w11299;
w11301 <= not w9569 and not w9583;
w11302 <= not w9555 and not w11301;
w11303 <= not w9568 and not w9582;
w11304 <= not w9579 and w11303;
w11305 <= not w9565 and w11304;
w11306 <= not w11302 and not w11305;
w11307 <= not w7038 and not w9573;
w11308 <= not w9570 and w11307;
w11309 <= w9575 and not w11308;
w11310 <= not w9571 and w9573;
w11311 <= not w11309 and not w11310;
w11312 <= not w7066 and not w9559;
w11313 <= not w9556 and w11312;
w11314 <= w9561 and not w11313;
w11315 <= not w9557 and w9559;
w11316 <= not w11314 and not w11315;
w11317 <= not w11311 and w11316;
w11318 <= w11311 and not w11316;
w11319 <= not w11317 and not w11318;
w11320 <= not w11306 and not w11319;
w11321 <= not w11305 and not w11317;
w11322 <= not w11318 and w11321;
w11323 <= not w11302 and w11322;
w11324 <= not w11320 and not w11323;
w11325 <= not w11300 and w11324;
w11326 <= w11300 and not w11324;
w11327 <= not w11325 and not w11326;
w11328 <= not w11276 and not w11327;
w11329 <= w11276 and w11327;
w11330 <= not w11328 and not w11329;
w11331 <= not w9509 and not w9545;
w11332 <= not w9473 and not w11331;
w11333 <= w9509 and w9545;
w11334 <= not w11332 and not w11333;
w11335 <= not w9525 and not w9539;
w11336 <= not w9511 and not w11335;
w11337 <= not w9524 and not w9538;
w11338 <= not w9535 and w11337;
w11339 <= not w9521 and w11338;
w11340 <= not w11336 and not w11339;
w11341 <= not w7174 and not w9529;
w11342 <= not w9526 and w11341;
w11343 <= w9531 and not w11342;
w11344 <= not w9527 and w9529;
w11345 <= not w11343 and not w11344;
w11346 <= not w7159 and not w9515;
w11347 <= not w9512 and w11346;
w11348 <= w9517 and not w11347;
w11349 <= not w9513 and w9515;
w11350 <= not w11348 and not w11349;
w11351 <= not w11345 and w11350;
w11352 <= w11345 and not w11350;
w11353 <= not w11351 and not w11352;
w11354 <= not w11340 and not w11353;
w11355 <= not w11339 and not w11351;
w11356 <= not w11352 and w11355;
w11357 <= not w11336 and w11356;
w11358 <= not w11354 and not w11357;
w11359 <= not w9489 and not w9503;
w11360 <= not w9475 and not w11359;
w11361 <= not w9488 and not w9502;
w11362 <= not w9499 and w11361;
w11363 <= not w9485 and w11362;
w11364 <= not w11360 and not w11363;
w11365 <= not w7210 and not w9493;
w11366 <= not w9490 and w11365;
w11367 <= w9495 and not w11366;
w11368 <= not w9491 and w9493;
w11369 <= not w11367 and not w11368;
w11370 <= not w7238 and not w9479;
w11371 <= not w9476 and w11370;
w11372 <= w9481 and not w11371;
w11373 <= not w9477 and w9479;
w11374 <= not w11372 and not w11373;
w11375 <= not w11369 and w11374;
w11376 <= w11369 and not w11374;
w11377 <= not w11375 and not w11376;
w11378 <= not w11364 and not w11377;
w11379 <= not w11363 and not w11375;
w11380 <= not w11376 and w11379;
w11381 <= not w11360 and w11380;
w11382 <= not w11378 and not w11381;
w11383 <= not w11358 and w11382;
w11384 <= w11358 and not w11382;
w11385 <= not w11383 and not w11384;
w11386 <= not w11334 and not w11385;
w11387 <= w11334 and w11385;
w11388 <= not w11386 and not w11387;
w11389 <= not w11330 and w11388;
w11390 <= w11330 and not w11388;
w11391 <= not w11389 and not w11390;
w11392 <= not w11272 and not w11391;
w11393 <= w11272 and w11391;
w11394 <= not w11392 and not w11393;
w11395 <= not w11268 and w11394;
w11396 <= w11268 and not w11394;
w11397 <= not w11395 and not w11396;
w11398 <= not w11142 and not w11397;
w11399 <= w11142 and w11397;
w11400 <= not w11398 and not w11399;
w11401 <= not w11138 and w11400;
w11402 <= w11138 and not w11400;
w11403 <= not w11401 and not w11402;
w11404 <= not w10876 and not w11403;
w11405 <= w10876 and w11403;
w11406 <= not w11404 and not w11405;
w11407 <= not w9457 and not w9460;
w11408 <= not w9048 and not w11407;
w11409 <= not w9289 and w9457;
w11410 <= not w9288 and w11409;
w11411 <= not w11408 and not w11410;
w11412 <= not w9282 and not w9285;
w11413 <= not w9050 and not w11412;
w11414 <= not w9202 and w9282;
w11415 <= not w9201 and w11414;
w11416 <= not w11413 and not w11415;
w11417 <= not w9117 and not w9197;
w11418 <= not w9052 and not w11417;
w11419 <= w9117 and w9197;
w11420 <= not w11418 and not w11419;
w11421 <= not w9155 and not w9191;
w11422 <= not w9119 and not w11421;
w11423 <= w9155 and w9191;
w11424 <= not w11422 and not w11423;
w11425 <= not w9171 and not w9185;
w11426 <= not w9157 and not w11425;
w11427 <= not w9170 and not w9184;
w11428 <= not w9181 and w11427;
w11429 <= not w9167 and w11428;
w11430 <= not w11426 and not w11429;
w11431 <= not w4586 and not w9175;
w11432 <= not w9172 and w11431;
w11433 <= w9177 and not w11432;
w11434 <= not w9173 and w9175;
w11435 <= not w11433 and not w11434;
w11436 <= not w4501 and not w9161;
w11437 <= not w9158 and w11436;
w11438 <= w9163 and not w11437;
w11439 <= not w9159 and w9161;
w11440 <= not w11438 and not w11439;
w11441 <= not w11435 and w11440;
w11442 <= w11435 and not w11440;
w11443 <= not w11441 and not w11442;
w11444 <= not w11430 and not w11443;
w11445 <= not w11429 and not w11441;
w11446 <= not w11442 and w11445;
w11447 <= not w11426 and w11446;
w11448 <= not w11444 and not w11447;
w11449 <= not w9135 and not w9149;
w11450 <= not w9121 and not w11449;
w11451 <= not w9134 and not w9148;
w11452 <= not w9145 and w11451;
w11453 <= not w9131 and w11452;
w11454 <= not w11450 and not w11453;
w11455 <= not w4297 and not w9139;
w11456 <= not w9136 and w11455;
w11457 <= w9141 and not w11456;
w11458 <= not w9137 and w9139;
w11459 <= not w11457 and not w11458;
w11460 <= not w4405 and not w9125;
w11461 <= not w9122 and w11460;
w11462 <= w9127 and not w11461;
w11463 <= not w9123 and w9125;
w11464 <= not w11462 and not w11463;
w11465 <= not w11459 and w11464;
w11466 <= w11459 and not w11464;
w11467 <= not w11465 and not w11466;
w11468 <= not w11454 and not w11467;
w11469 <= not w11453 and not w11465;
w11470 <= not w11466 and w11469;
w11471 <= not w11450 and w11470;
w11472 <= not w11468 and not w11471;
w11473 <= not w11448 and w11472;
w11474 <= w11448 and not w11472;
w11475 <= not w11473 and not w11474;
w11476 <= not w11424 and not w11475;
w11477 <= w11424 and w11475;
w11478 <= not w11476 and not w11477;
w11479 <= not w9075 and not w9111;
w11480 <= not w9054 and not w11479;
w11481 <= w9075 and not w9109;
w11482 <= not w9110 and w11481;
w11483 <= not w11480 and not w11482;
w11484 <= not w4205 and w9068;
w11485 <= not w9055 and w11484;
w11486 <= w9065 and not w11485;
w11487 <= not w9056 and not w9068;
w11488 <= not w11486 and not w11487;
w11489 <= not w9058 and not w9060;
w11490 <= not w11488 and w11489;
w11491 <= not w11486 and not w11489;
w11492 <= not w11487 and w11491;
w11493 <= not w11490 and not w11492;
w11494 <= not w9091 and not w9105;
w11495 <= not w9077 and not w11494;
w11496 <= not w9090 and not w9104;
w11497 <= not w9101 and w11496;
w11498 <= not w9087 and w11497;
w11499 <= not w11495 and not w11498;
w11500 <= not w4058 and not w9095;
w11501 <= not w9092 and w11500;
w11502 <= w9097 and not w11501;
w11503 <= not w9093 and w9095;
w11504 <= not w11502 and not w11503;
w11505 <= not w3973 and not w9081;
w11506 <= not w9078 and w11505;
w11507 <= w9083 and not w11506;
w11508 <= not w9079 and w9081;
w11509 <= not w11507 and not w11508;
w11510 <= not w11504 and w11509;
w11511 <= w11504 and not w11509;
w11512 <= not w11510 and not w11511;
w11513 <= not w11499 and not w11512;
w11514 <= not w11498 and not w11510;
w11515 <= not w11511 and w11514;
w11516 <= not w11495 and w11515;
w11517 <= not w11513 and not w11516;
w11518 <= not w11493 and not w11517;
w11519 <= w11493 and w11517;
w11520 <= not w11518 and not w11519;
w11521 <= not w11483 and w11520;
w11522 <= w11483 and not w11520;
w11523 <= not w11521 and not w11522;
w11524 <= not w11478 and w11523;
w11525 <= w11478 and not w11523;
w11526 <= not w11524 and not w11525;
w11527 <= not w11420 and not w11526;
w11528 <= w11420 and w11526;
w11529 <= not w11527 and not w11528;
w11530 <= not w9240 and not w9276;
w11531 <= not w9204 and not w11530;
w11532 <= w9240 and w9276;
w11533 <= not w11531 and not w11532;
w11534 <= not w9256 and not w9270;
w11535 <= not w9242 and not w11534;
w11536 <= not w9255 and not w9269;
w11537 <= not w9266 and w11536;
w11538 <= not w9252 and w11537;
w11539 <= not w11535 and not w11538;
w11540 <= not w3640 and not w9260;
w11541 <= not w9257 and w11540;
w11542 <= w9262 and not w11541;
w11543 <= not w9258 and w9260;
w11544 <= not w11542 and not w11543;
w11545 <= not w3555 and not w9246;
w11546 <= not w9243 and w11545;
w11547 <= w9248 and not w11546;
w11548 <= not w9244 and w9246;
w11549 <= not w11547 and not w11548;
w11550 <= not w11544 and w11549;
w11551 <= w11544 and not w11549;
w11552 <= not w11550 and not w11551;
w11553 <= not w11539 and not w11552;
w11554 <= not w11538 and not w11550;
w11555 <= not w11551 and w11554;
w11556 <= not w11535 and w11555;
w11557 <= not w11553 and not w11556;
w11558 <= not w9220 and not w9234;
w11559 <= not w9206 and not w11558;
w11560 <= not w9219 and not w9233;
w11561 <= not w9230 and w11560;
w11562 <= not w9216 and w11561;
w11563 <= not w11559 and not w11562;
w11564 <= not w3842 and not w9224;
w11565 <= not w9221 and w11564;
w11566 <= w9226 and not w11565;
w11567 <= not w9222 and w9224;
w11568 <= not w11566 and not w11567;
w11569 <= not w3870 and not w9210;
w11570 <= not w9207 and w11569;
w11571 <= w9212 and not w11570;
w11572 <= not w9208 and w9210;
w11573 <= not w11571 and not w11572;
w11574 <= not w11568 and w11573;
w11575 <= w11568 and not w11573;
w11576 <= not w11574 and not w11575;
w11577 <= not w11563 and not w11576;
w11578 <= not w11562 and not w11574;
w11579 <= not w11575 and w11578;
w11580 <= not w11559 and w11579;
w11581 <= not w11577 and not w11580;
w11582 <= not w11557 and w11581;
w11583 <= w11557 and not w11581;
w11584 <= not w11582 and not w11583;
w11585 <= not w11533 and not w11584;
w11586 <= w11533 and w11584;
w11587 <= not w11585 and not w11586;
w11588 <= not w11529 and w11587;
w11589 <= not w11527 and not w11587;
w11590 <= not w11528 and w11589;
w11591 <= not w11588 and not w11590;
w11592 <= not w11416 and not w11591;
w11593 <= w11416 and w11591;
w11594 <= not w11592 and not w11593;
w11595 <= not w9371 and not w9451;
w11596 <= not w9291 and not w11595;
w11597 <= w9371 and w9451;
w11598 <= not w11596 and not w11597;
w11599 <= not w9409 and not w9445;
w11600 <= not w9373 and not w11599;
w11601 <= w9409 and w9445;
w11602 <= not w11600 and not w11601;
w11603 <= not w9425 and not w9439;
w11604 <= not w9411 and not w11603;
w11605 <= not w9424 and not w9438;
w11606 <= not w9435 and w11605;
w11607 <= not w9421 and w11606;
w11608 <= not w11604 and not w11607;
w11609 <= not w5381 and not w9429;
w11610 <= not w9426 and w11609;
w11611 <= w9431 and not w11610;
w11612 <= not w9427 and w9429;
w11613 <= not w11611 and not w11612;
w11614 <= not w5366 and not w9415;
w11615 <= not w9412 and w11614;
w11616 <= w9417 and not w11615;
w11617 <= not w9413 and w9415;
w11618 <= not w11616 and not w11617;
w11619 <= not w11613 and w11618;
w11620 <= w11613 and not w11618;
w11621 <= not w11619 and not w11620;
w11622 <= not w11608 and not w11621;
w11623 <= not w11607 and not w11619;
w11624 <= not w11620 and w11623;
w11625 <= not w11604 and w11624;
w11626 <= not w11622 and not w11625;
w11627 <= not w9389 and not w9403;
w11628 <= not w9375 and not w11627;
w11629 <= not w9388 and not w9402;
w11630 <= not w9399 and w11629;
w11631 <= not w9385 and w11630;
w11632 <= not w11628 and not w11631;
w11633 <= not w5312 and not w9393;
w11634 <= not w9390 and w11633;
w11635 <= w9395 and not w11634;
w11636 <= not w9391 and w9393;
w11637 <= not w11635 and not w11636;
w11638 <= not w5340 and not w9379;
w11639 <= not w9376 and w11638;
w11640 <= w9381 and not w11639;
w11641 <= not w9377 and w9379;
w11642 <= not w11640 and not w11641;
w11643 <= not w11637 and w11642;
w11644 <= w11637 and not w11642;
w11645 <= not w11643 and not w11644;
w11646 <= not w11632 and not w11645;
w11647 <= not w11631 and not w11643;
w11648 <= not w11644 and w11647;
w11649 <= not w11628 and w11648;
w11650 <= not w11646 and not w11649;
w11651 <= not w11626 and w11650;
w11652 <= w11626 and not w11650;
w11653 <= not w11651 and not w11652;
w11654 <= not w11602 and not w11653;
w11655 <= w11602 and w11653;
w11656 <= not w11654 and not w11655;
w11657 <= not w9329 and not w9365;
w11658 <= not w9293 and not w11657;
w11659 <= w9329 and w9365;
w11660 <= not w11658 and not w11659;
w11661 <= not w9345 and not w9359;
w11662 <= not w9331 and not w11661;
w11663 <= not w9344 and not w9358;
w11664 <= not w9355 and w11663;
w11665 <= not w9341 and w11664;
w11666 <= not w11662 and not w11665;
w11667 <= not w5448 and not w9349;
w11668 <= not w9346 and w11667;
w11669 <= w9351 and not w11668;
w11670 <= not w9347 and w9349;
w11671 <= not w11669 and not w11670;
w11672 <= not w5433 and not w9335;
w11673 <= not w9332 and w11672;
w11674 <= w9337 and not w11673;
w11675 <= not w9333 and w9335;
w11676 <= not w11674 and not w11675;
w11677 <= not w11671 and w11676;
w11678 <= w11671 and not w11676;
w11679 <= not w11677 and not w11678;
w11680 <= not w11666 and not w11679;
w11681 <= not w11665 and not w11677;
w11682 <= not w11678 and w11681;
w11683 <= not w11662 and w11682;
w11684 <= not w11680 and not w11683;
w11685 <= not w9309 and not w9323;
w11686 <= not w9295 and not w11685;
w11687 <= not w9308 and not w9322;
w11688 <= not w9319 and w11687;
w11689 <= not w9305 and w11688;
w11690 <= not w11686 and not w11689;
w11691 <= not w5484 and not w9313;
w11692 <= not w9310 and w11691;
w11693 <= w9315 and not w11692;
w11694 <= not w9311 and w9313;
w11695 <= not w11693 and not w11694;
w11696 <= not w5512 and not w9299;
w11697 <= not w9296 and w11696;
w11698 <= w9301 and not w11697;
w11699 <= not w9297 and w9299;
w11700 <= not w11698 and not w11699;
w11701 <= not w11695 and w11700;
w11702 <= w11695 and not w11700;
w11703 <= not w11701 and not w11702;
w11704 <= not w11690 and not w11703;
w11705 <= not w11689 and not w11701;
w11706 <= not w11702 and w11705;
w11707 <= not w11686 and w11706;
w11708 <= not w11704 and not w11707;
w11709 <= not w11684 and w11708;
w11710 <= w11684 and not w11708;
w11711 <= not w11709 and not w11710;
w11712 <= not w11660 and not w11711;
w11713 <= w11660 and w11711;
w11714 <= not w11712 and not w11713;
w11715 <= not w11656 and w11714;
w11716 <= w11656 and not w11714;
w11717 <= not w11715 and not w11716;
w11718 <= not w11598 and not w11717;
w11719 <= w11598 and w11717;
w11720 <= not w11718 and not w11719;
w11721 <= not w11594 and w11720;
w11722 <= not w11592 and not w11720;
w11723 <= not w11593 and w11722;
w11724 <= not w11721 and not w11723;
w11725 <= not w11411 and not w11724;
w11726 <= w11411 and w11724;
w11727 <= not w11725 and not w11726;
w11728 <= not w11406 and w11727;
w11729 <= w11406 and not w11727;
w11730 <= not w11728 and not w11729;
w11731 <= not w10872 and not w11730;
w11732 <= w10872 and w11730;
w11733 <= not w11731 and not w11732;
w11734 <= not w10513 and not w10857;
w11735 <= not w10169 and not w11734;
w11736 <= w10513 and w10857;
w11737 <= not w11735 and not w11736;
w11738 <= not w10683 and not w10851;
w11739 <= not w10515 and not w11738;
w11740 <= w10683 and w10851;
w11741 <= not w11739 and not w11740;
w11742 <= not w10765 and not w10845;
w11743 <= not w10685 and not w11742;
w11744 <= w10765 and w10845;
w11745 <= not w11743 and not w11744;
w11746 <= not w10803 and not w10839;
w11747 <= not w10767 and not w11746;
w11748 <= w10803 and w10839;
w11749 <= not w11747 and not w11748;
w11750 <= not w10819 and not w10833;
w11751 <= not w10805 and not w11750;
w11752 <= not w10818 and not w10832;
w11753 <= not w10829 and w11752;
w11754 <= not w10815 and w11753;
w11755 <= not w11751 and not w11754;
w11756 <= not w1642 and not w10823;
w11757 <= not w10820 and w11756;
w11758 <= w10825 and not w11757;
w11759 <= not w10821 and w10823;
w11760 <= not w11758 and not w11759;
w11761 <= not w1557 and not w10809;
w11762 <= not w10806 and w11761;
w11763 <= w10811 and not w11762;
w11764 <= not w10807 and w10809;
w11765 <= not w11763 and not w11764;
w11766 <= not w11760 and w11765;
w11767 <= w11760 and not w11765;
w11768 <= not w11766 and not w11767;
w11769 <= not w11755 and not w11768;
w11770 <= not w11754 and not w11766;
w11771 <= not w11767 and w11770;
w11772 <= not w11751 and w11771;
w11773 <= not w11769 and not w11772;
w11774 <= not w10783 and not w10797;
w11775 <= not w10769 and not w11774;
w11776 <= not w10782 and not w10796;
w11777 <= not w10793 and w11776;
w11778 <= not w10779 and w11777;
w11779 <= not w11775 and not w11778;
w11780 <= not w1353 and not w10787;
w11781 <= not w10784 and w11780;
w11782 <= w10789 and not w11781;
w11783 <= not w10785 and w10787;
w11784 <= not w11782 and not w11783;
w11785 <= not w1461 and not w10773;
w11786 <= not w10770 and w11785;
w11787 <= w10775 and not w11786;
w11788 <= not w10771 and w10773;
w11789 <= not w11787 and not w11788;
w11790 <= not w11784 and w11789;
w11791 <= w11784 and not w11789;
w11792 <= not w11790 and not w11791;
w11793 <= not w11779 and not w11792;
w11794 <= not w11778 and not w11790;
w11795 <= not w11791 and w11794;
w11796 <= not w11775 and w11795;
w11797 <= not w11793 and not w11796;
w11798 <= not w11773 and w11797;
w11799 <= w11773 and not w11797;
w11800 <= not w11798 and not w11799;
w11801 <= not w11749 and not w11800;
w11802 <= w11749 and w11800;
w11803 <= not w11801 and not w11802;
w11804 <= not w10723 and not w10759;
w11805 <= not w10687 and not w11804;
w11806 <= w10723 and w10759;
w11807 <= not w11805 and not w11806;
w11808 <= not w10739 and not w10753;
w11809 <= not w10725 and not w11808;
w11810 <= not w10738 and not w10752;
w11811 <= not w10749 and w11810;
w11812 <= not w10735 and w11811;
w11813 <= not w11809 and not w11812;
w11814 <= not w1024 and not w10743;
w11815 <= not w10740 and w11814;
w11816 <= w10745 and not w11815;
w11817 <= not w10741 and w10743;
w11818 <= not w11816 and not w11817;
w11819 <= not w939 and not w10729;
w11820 <= not w10726 and w11819;
w11821 <= w10731 and not w11820;
w11822 <= not w10727 and w10729;
w11823 <= not w11821 and not w11822;
w11824 <= not w11818 and w11823;
w11825 <= w11818 and not w11823;
w11826 <= not w11824 and not w11825;
w11827 <= not w11813 and not w11826;
w11828 <= not w11812 and not w11824;
w11829 <= not w11825 and w11828;
w11830 <= not w11809 and w11829;
w11831 <= not w11827 and not w11830;
w11832 <= not w10703 and not w10717;
w11833 <= not w10689 and not w11832;
w11834 <= not w10702 and not w10716;
w11835 <= not w10713 and w11834;
w11836 <= not w10699 and w11835;
w11837 <= not w11833 and not w11836;
w11838 <= not w1226 and not w10707;
w11839 <= not w10704 and w11838;
w11840 <= w10709 and not w11839;
w11841 <= not w10705 and w10707;
w11842 <= not w11840 and not w11841;
w11843 <= not w1254 and not w10693;
w11844 <= not w10690 and w11843;
w11845 <= w10695 and not w11844;
w11846 <= not w10691 and w10693;
w11847 <= not w11845 and not w11846;
w11848 <= not w11842 and w11847;
w11849 <= w11842 and not w11847;
w11850 <= not w11848 and not w11849;
w11851 <= not w11837 and not w11850;
w11852 <= not w11836 and not w11848;
w11853 <= not w11849 and w11852;
w11854 <= not w11833 and w11853;
w11855 <= not w11851 and not w11854;
w11856 <= not w11831 and w11855;
w11857 <= w11831 and not w11855;
w11858 <= not w11856 and not w11857;
w11859 <= not w11807 and not w11858;
w11860 <= w11807 and w11858;
w11861 <= not w11859 and not w11860;
w11862 <= not w11803 and w11861;
w11863 <= w11803 and not w11861;
w11864 <= not w11862 and not w11863;
w11865 <= not w11745 and not w11864;
w11866 <= w11745 and w11864;
w11867 <= not w11865 and not w11866;
w11868 <= not w10597 and not w10677;
w11869 <= not w10517 and not w11868;
w11870 <= w10597 and w10677;
w11871 <= not w11869 and not w11870;
w11872 <= not w10635 and not w10671;
w11873 <= not w10599 and not w11872;
w11874 <= w10635 and w10671;
w11875 <= not w11873 and not w11874;
w11876 <= not w10651 and not w10665;
w11877 <= not w10637 and not w11876;
w11878 <= not w10650 and not w10664;
w11879 <= not w10661 and w11878;
w11880 <= not w10647 and w11879;
w11881 <= not w11877 and not w11880;
w11882 <= not w370 and not w10655;
w11883 <= not w10652 and w11882;
w11884 <= w10657 and not w11883;
w11885 <= not w10653 and w10655;
w11886 <= not w11884 and not w11885;
w11887 <= not w285 and not w10641;
w11888 <= not w10638 and w11887;
w11889 <= w10643 and not w11888;
w11890 <= not w10639 and w10641;
w11891 <= not w11889 and not w11890;
w11892 <= not w11886 and w11891;
w11893 <= w11886 and not w11891;
w11894 <= not w11892 and not w11893;
w11895 <= not w11881 and not w11894;
w11896 <= not w11880 and not w11892;
w11897 <= not w11893 and w11896;
w11898 <= not w11877 and w11897;
w11899 <= not w11895 and not w11898;
w11900 <= not w10615 and not w10629;
w11901 <= not w10601 and not w11900;
w11902 <= not w10614 and not w10628;
w11903 <= not w10625 and w11902;
w11904 <= not w10611 and w11903;
w11905 <= not w11901 and not w11904;
w11906 <= not w81 and not w10619;
w11907 <= not w10616 and w11906;
w11908 <= w10621 and not w11907;
w11909 <= not w10617 and w10619;
w11910 <= not w11908 and not w11909;
w11911 <= not w189 and not w10605;
w11912 <= not w10602 and w11911;
w11913 <= w10607 and not w11912;
w11914 <= not w10603 and w10605;
w11915 <= not w11913 and not w11914;
w11916 <= not w11910 and w11915;
w11917 <= w11910 and not w11915;
w11918 <= not w11916 and not w11917;
w11919 <= not w11905 and not w11918;
w11920 <= not w11904 and not w11916;
w11921 <= not w11917 and w11920;
w11922 <= not w11901 and w11921;
w11923 <= not w11919 and not w11922;
w11924 <= not w11899 and w11923;
w11925 <= w11899 and not w11923;
w11926 <= not w11924 and not w11925;
w11927 <= not w11875 and not w11926;
w11928 <= w11875 and w11926;
w11929 <= not w11927 and not w11928;
w11930 <= not w10555 and not w10591;
w11931 <= not w10519 and not w11930;
w11932 <= w10555 and w10591;
w11933 <= not w11931 and not w11932;
w11934 <= not w10571 and not w10585;
w11935 <= not w10557 and not w11934;
w11936 <= not w10570 and not w10584;
w11937 <= not w10581 and w11936;
w11938 <= not w10567 and w11937;
w11939 <= not w11935 and not w11938;
w11940 <= not w765 and not w10575;
w11941 <= not w10572 and w11940;
w11942 <= w10577 and not w11941;
w11943 <= not w10573 and w10575;
w11944 <= not w11942 and not w11943;
w11945 <= not w750 and not w10561;
w11946 <= not w10558 and w11945;
w11947 <= w10563 and not w11946;
w11948 <= not w10559 and w10561;
w11949 <= not w11947 and not w11948;
w11950 <= not w11944 and w11949;
w11951 <= w11944 and not w11949;
w11952 <= not w11950 and not w11951;
w11953 <= not w11939 and not w11952;
w11954 <= not w11938 and not w11950;
w11955 <= not w11951 and w11954;
w11956 <= not w11935 and w11955;
w11957 <= not w11953 and not w11956;
w11958 <= not w10535 and not w10549;
w11959 <= not w10521 and not w11958;
w11960 <= not w10534 and not w10548;
w11961 <= not w10545 and w11960;
w11962 <= not w10531 and w11961;
w11963 <= not w11959 and not w11962;
w11964 <= not w801 and not w10539;
w11965 <= not w10536 and w11964;
w11966 <= w10541 and not w11965;
w11967 <= not w10537 and w10539;
w11968 <= not w11966 and not w11967;
w11969 <= not w829 and not w10525;
w11970 <= not w10522 and w11969;
w11971 <= w10527 and not w11970;
w11972 <= not w10523 and w10525;
w11973 <= not w11971 and not w11972;
w11974 <= not w11968 and w11973;
w11975 <= w11968 and not w11973;
w11976 <= not w11974 and not w11975;
w11977 <= not w11963 and not w11976;
w11978 <= not w11962 and not w11974;
w11979 <= not w11975 and w11978;
w11980 <= not w11959 and w11979;
w11981 <= not w11977 and not w11980;
w11982 <= not w11957 and w11981;
w11983 <= w11957 and not w11981;
w11984 <= not w11982 and not w11983;
w11985 <= not w11933 and not w11984;
w11986 <= w11933 and w11984;
w11987 <= not w11985 and not w11986;
w11988 <= not w11929 and w11987;
w11989 <= w11929 and not w11987;
w11990 <= not w11988 and not w11989;
w11991 <= not w11871 and not w11990;
w11992 <= w11871 and w11990;
w11993 <= not w11991 and not w11992;
w11994 <= not w11867 and w11993;
w11995 <= w11867 and not w11993;
w11996 <= not w11994 and not w11995;
w11997 <= not w11741 and not w11996;
w11998 <= w11741 and w11996;
w11999 <= not w11997 and not w11998;
w12000 <= not w10339 and not w10507;
w12001 <= not w10171 and not w12000;
w12002 <= w10339 and w10507;
w12003 <= not w12001 and not w12002;
w12004 <= not w10421 and not w10501;
w12005 <= not w10341 and not w12004;
w12006 <= w10421 and w10501;
w12007 <= not w12005 and not w12006;
w12008 <= not w10459 and not w10495;
w12009 <= not w10423 and not w12008;
w12010 <= w10459 and w10495;
w12011 <= not w12009 and not w12010;
w12012 <= not w10475 and not w10489;
w12013 <= not w10461 and not w12012;
w12014 <= not w10474 and not w10488;
w12015 <= not w10485 and w12014;
w12016 <= not w10471 and w12015;
w12017 <= not w12013 and not w12016;
w12018 <= not w3171 and not w10479;
w12019 <= not w10476 and w12018;
w12020 <= w10481 and not w12019;
w12021 <= not w10477 and w10479;
w12022 <= not w12020 and not w12021;
w12023 <= not w3156 and not w10465;
w12024 <= not w10462 and w12023;
w12025 <= w10467 and not w12024;
w12026 <= not w10463 and w10465;
w12027 <= not w12025 and not w12026;
w12028 <= not w12022 and w12027;
w12029 <= w12022 and not w12027;
w12030 <= not w12028 and not w12029;
w12031 <= not w12017 and not w12030;
w12032 <= not w12016 and not w12028;
w12033 <= not w12029 and w12032;
w12034 <= not w12013 and w12033;
w12035 <= not w12031 and not w12034;
w12036 <= not w10439 and not w10453;
w12037 <= not w10425 and not w12036;
w12038 <= not w10438 and not w10452;
w12039 <= not w10449 and w12038;
w12040 <= not w10435 and w12039;
w12041 <= not w12037 and not w12040;
w12042 <= not w3102 and not w10443;
w12043 <= not w10440 and w12042;
w12044 <= w10445 and not w12043;
w12045 <= not w10441 and w10443;
w12046 <= not w12044 and not w12045;
w12047 <= not w3130 and not w10429;
w12048 <= not w10426 and w12047;
w12049 <= w10431 and not w12048;
w12050 <= not w10427 and w10429;
w12051 <= not w12049 and not w12050;
w12052 <= not w12046 and w12051;
w12053 <= w12046 and not w12051;
w12054 <= not w12052 and not w12053;
w12055 <= not w12041 and not w12054;
w12056 <= not w12040 and not w12052;
w12057 <= not w12053 and w12056;
w12058 <= not w12037 and w12057;
w12059 <= not w12055 and not w12058;
w12060 <= not w12035 and w12059;
w12061 <= w12035 and not w12059;
w12062 <= not w12060 and not w12061;
w12063 <= not w12011 and not w12062;
w12064 <= w12011 and w12062;
w12065 <= not w12063 and not w12064;
w12066 <= not w10379 and not w10415;
w12067 <= not w10343 and not w12066;
w12068 <= w10379 and w10415;
w12069 <= not w12067 and not w12068;
w12070 <= not w10395 and not w10409;
w12071 <= not w10381 and not w12070;
w12072 <= not w10394 and not w10408;
w12073 <= not w10405 and w12072;
w12074 <= not w10391 and w12073;
w12075 <= not w12071 and not w12074;
w12076 <= not w3009 and not w10399;
w12077 <= not w10396 and w12076;
w12078 <= w10401 and not w12077;
w12079 <= not w10397 and w10399;
w12080 <= not w12078 and not w12079;
w12081 <= not w2994 and not w10385;
w12082 <= not w10382 and w12081;
w12083 <= w10387 and not w12082;
w12084 <= not w10383 and w10385;
w12085 <= not w12083 and not w12084;
w12086 <= not w12080 and w12085;
w12087 <= w12080 and not w12085;
w12088 <= not w12086 and not w12087;
w12089 <= not w12075 and not w12088;
w12090 <= not w12074 and not w12086;
w12091 <= not w12087 and w12090;
w12092 <= not w12071 and w12091;
w12093 <= not w12089 and not w12092;
w12094 <= not w10359 and not w10373;
w12095 <= not w10345 and not w12094;
w12096 <= not w10358 and not w10372;
w12097 <= not w10369 and w12096;
w12098 <= not w10355 and w12097;
w12099 <= not w12095 and not w12098;
w12100 <= not w3045 and not w10363;
w12101 <= not w10360 and w12100;
w12102 <= w10365 and not w12101;
w12103 <= not w10361 and w10363;
w12104 <= not w12102 and not w12103;
w12105 <= not w3073 and not w10349;
w12106 <= not w10346 and w12105;
w12107 <= w10351 and not w12106;
w12108 <= not w10347 and w10349;
w12109 <= not w12107 and not w12108;
w12110 <= not w12104 and w12109;
w12111 <= w12104 and not w12109;
w12112 <= not w12110 and not w12111;
w12113 <= not w12099 and not w12112;
w12114 <= not w12098 and not w12110;
w12115 <= not w12111 and w12114;
w12116 <= not w12095 and w12115;
w12117 <= not w12113 and not w12116;
w12118 <= not w12093 and w12117;
w12119 <= w12093 and not w12117;
w12120 <= not w12118 and not w12119;
w12121 <= not w12069 and not w12120;
w12122 <= w12069 and w12120;
w12123 <= not w12121 and not w12122;
w12124 <= not w12065 and w12123;
w12125 <= w12065 and not w12123;
w12126 <= not w12124 and not w12125;
w12127 <= not w12007 and not w12126;
w12128 <= w12007 and w12126;
w12129 <= not w12127 and not w12128;
w12130 <= not w10253 and not w10333;
w12131 <= not w10173 and not w12130;
w12132 <= w10253 and w10333;
w12133 <= not w12131 and not w12132;
w12134 <= not w10291 and not w10327;
w12135 <= not w10255 and not w12134;
w12136 <= w10291 and w10327;
w12137 <= not w12135 and not w12136;
w12138 <= not w10307 and not w10321;
w12139 <= not w10293 and not w12138;
w12140 <= not w10306 and not w10320;
w12141 <= not w10317 and w12140;
w12142 <= not w10303 and w12141;
w12143 <= not w12139 and not w12142;
w12144 <= not w3300 and not w10311;
w12145 <= not w10308 and w12144;
w12146 <= w10313 and not w12145;
w12147 <= not w10309 and w10311;
w12148 <= not w12146 and not w12147;
w12149 <= not w3285 and not w10297;
w12150 <= not w10294 and w12149;
w12151 <= w10299 and not w12150;
w12152 <= not w10295 and w10297;
w12153 <= not w12151 and not w12152;
w12154 <= not w12148 and w12153;
w12155 <= w12148 and not w12153;
w12156 <= not w12154 and not w12155;
w12157 <= not w12143 and not w12156;
w12158 <= not w12142 and not w12154;
w12159 <= not w12155 and w12158;
w12160 <= not w12139 and w12159;
w12161 <= not w12157 and not w12160;
w12162 <= not w10271 and not w10285;
w12163 <= not w10257 and not w12162;
w12164 <= not w10270 and not w10284;
w12165 <= not w10281 and w12164;
w12166 <= not w10267 and w12165;
w12167 <= not w12163 and not w12166;
w12168 <= not w3231 and not w10275;
w12169 <= not w10272 and w12168;
w12170 <= w10277 and not w12169;
w12171 <= not w10273 and w10275;
w12172 <= not w12170 and not w12171;
w12173 <= not w3259 and not w10261;
w12174 <= not w10258 and w12173;
w12175 <= w10263 and not w12174;
w12176 <= not w10259 and w10261;
w12177 <= not w12175 and not w12176;
w12178 <= not w12172 and w12177;
w12179 <= w12172 and not w12177;
w12180 <= not w12178 and not w12179;
w12181 <= not w12167 and not w12180;
w12182 <= not w12166 and not w12178;
w12183 <= not w12179 and w12182;
w12184 <= not w12163 and w12183;
w12185 <= not w12181 and not w12184;
w12186 <= not w12161 and w12185;
w12187 <= w12161 and not w12185;
w12188 <= not w12186 and not w12187;
w12189 <= not w12137 and not w12188;
w12190 <= w12137 and w12188;
w12191 <= not w12189 and not w12190;
w12192 <= not w10211 and not w10247;
w12193 <= not w10175 and not w12192;
w12194 <= w10211 and w10247;
w12195 <= not w12193 and not w12194;
w12196 <= not w10227 and not w10241;
w12197 <= not w10213 and not w12196;
w12198 <= not w10226 and not w10240;
w12199 <= not w10237 and w12198;
w12200 <= not w10223 and w12199;
w12201 <= not w12197 and not w12200;
w12202 <= not w3367 and not w10231;
w12203 <= not w10228 and w12202;
w12204 <= w10233 and not w12203;
w12205 <= not w10229 and w10231;
w12206 <= not w12204 and not w12205;
w12207 <= not w3352 and not w10217;
w12208 <= not w10214 and w12207;
w12209 <= w10219 and not w12208;
w12210 <= not w10215 and w10217;
w12211 <= not w12209 and not w12210;
w12212 <= not w12206 and w12211;
w12213 <= w12206 and not w12211;
w12214 <= not w12212 and not w12213;
w12215 <= not w12201 and not w12214;
w12216 <= not w12200 and not w12212;
w12217 <= not w12213 and w12216;
w12218 <= not w12197 and w12217;
w12219 <= not w12215 and not w12218;
w12220 <= not w10191 and not w10205;
w12221 <= not w10177 and not w12220;
w12222 <= not w10190 and not w10204;
w12223 <= not w10201 and w12222;
w12224 <= not w10187 and w12223;
w12225 <= not w12221 and not w12224;
w12226 <= not w3403 and not w10195;
w12227 <= not w10192 and w12226;
w12228 <= w10197 and not w12227;
w12229 <= not w10193 and w10195;
w12230 <= not w12228 and not w12229;
w12231 <= not w3431 and not w10181;
w12232 <= not w10178 and w12231;
w12233 <= w10183 and not w12232;
w12234 <= not w10179 and w10181;
w12235 <= not w12233 and not w12234;
w12236 <= not w12230 and w12235;
w12237 <= w12230 and not w12235;
w12238 <= not w12236 and not w12237;
w12239 <= not w12225 and not w12238;
w12240 <= not w12224 and not w12236;
w12241 <= not w12237 and w12240;
w12242 <= not w12221 and w12241;
w12243 <= not w12239 and not w12242;
w12244 <= not w12219 and w12243;
w12245 <= w12219 and not w12243;
w12246 <= not w12244 and not w12245;
w12247 <= not w12195 and not w12246;
w12248 <= w12195 and w12246;
w12249 <= not w12247 and not w12248;
w12250 <= not w12191 and w12249;
w12251 <= w12191 and not w12249;
w12252 <= not w12250 and not w12251;
w12253 <= not w12133 and not w12252;
w12254 <= w12133 and w12252;
w12255 <= not w12253 and not w12254;
w12256 <= not w12129 and w12255;
w12257 <= w12129 and not w12255;
w12258 <= not w12256 and not w12257;
w12259 <= not w12003 and not w12258;
w12260 <= w12003 and w12258;
w12261 <= not w12259 and not w12260;
w12262 <= not w11999 and w12261;
w12263 <= w11999 and not w12261;
w12264 <= not w12262 and not w12263;
w12265 <= not w11737 and not w12264;
w12266 <= w11737 and w12264;
w12267 <= not w12265 and not w12266;
w12268 <= not w11733 and not w12267;
w12269 <= not w10868 and not w12268;
w12270 <= not w11731 and w12267;
w12271 <= not w11732 and w12270;
w12272 <= not w12269 and not w12271;
w12273 <= not w11406 and not w11727;
w12274 <= not w10872 and not w12273;
w12275 <= w11406 and w11727;
w12276 <= not w12274 and not w12275;
w12277 <= not w11594 and not w11720;
w12278 <= not w11411 and not w12277;
w12279 <= not w11592 and w11720;
w12280 <= not w11593 and w12279;
w12281 <= not w12278 and not w12280;
w12282 <= not w11529 and not w11587;
w12283 <= not w11416 and not w12282;
w12284 <= not w11527 and w11587;
w12285 <= not w11528 and w12284;
w12286 <= not w12283 and not w12285;
w12287 <= not w11478 and not w11523;
w12288 <= not w11420 and not w12287;
w12289 <= w11478 and w11523;
w12290 <= not w12288 and not w12289;
w12291 <= not w11483 and not w11518;
w12292 <= not w11519 and not w12291;
w12293 <= w11504 and w11509;
w12294 <= not w11499 and not w12293;
w12295 <= not w11504 and not w11509;
w12296 <= not w11490 and not w12295;
w12297 <= not w12294 and w12296;
w12298 <= not w12294 and not w12295;
w12299 <= w11490 and not w12298;
w12300 <= not w12297 and not w12299;
w12301 <= not w12292 and w12300;
w12302 <= not w11519 and not w12300;
w12303 <= not w12291 and w12302;
w12304 <= not w12301 and not w12303;
w12305 <= not w11448 and not w11472;
w12306 <= not w11424 and not w12305;
w12307 <= not w11447 and not w11471;
w12308 <= not w11468 and w12307;
w12309 <= not w11444 and w12308;
w12310 <= not w12306 and not w12309;
w12311 <= w11435 and w11440;
w12312 <= not w11430 and not w12311;
w12313 <= not w11435 and not w11440;
w12314 <= not w12312 and not w12313;
w12315 <= w11459 and w11464;
w12316 <= not w11454 and not w12315;
w12317 <= not w11459 and not w11464;
w12318 <= not w12316 and not w12317;
w12319 <= not w12314 and w12318;
w12320 <= w12314 and not w12318;
w12321 <= not w12319 and not w12320;
w12322 <= not w12310 and not w12321;
w12323 <= not w12309 and not w12319;
w12324 <= not w12320 and w12323;
w12325 <= not w12306 and w12324;
w12326 <= not w12322 and not w12325;
w12327 <= not w12304 and w12326;
w12328 <= w12304 and not w12326;
w12329 <= not w12327 and not w12328;
w12330 <= w12290 and w12329;
w12331 <= not w12290 and not w12329;
w12332 <= not w11557 and not w11581;
w12333 <= not w11533 and not w12332;
w12334 <= not w11556 and not w11580;
w12335 <= not w11577 and w12334;
w12336 <= not w11553 and w12335;
w12337 <= not w12333 and not w12336;
w12338 <= w11544 and w11549;
w12339 <= not w11539 and not w12338;
w12340 <= not w11544 and not w11549;
w12341 <= not w12339 and not w12340;
w12342 <= w11568 and w11573;
w12343 <= not w11563 and not w12342;
w12344 <= not w11568 and not w11573;
w12345 <= not w12343 and not w12344;
w12346 <= not w12341 and w12345;
w12347 <= w12341 and not w12345;
w12348 <= not w12346 and not w12347;
w12349 <= not w12337 and not w12348;
w12350 <= not w12336 and not w12346;
w12351 <= not w12347 and w12350;
w12352 <= not w12333 and w12351;
w12353 <= not w12349 and not w12352;
w12354 <= not w12331 and not w12353;
w12355 <= not w12330 and w12354;
w12356 <= not w12330 and not w12331;
w12357 <= w12353 and not w12356;
w12358 <= not w12355 and not w12357;
w12359 <= w12286 and w12358;
w12360 <= not w12286 and not w12358;
w12361 <= not w11656 and not w11714;
w12362 <= not w11598 and not w12361;
w12363 <= w11656 and w11714;
w12364 <= not w12362 and not w12363;
w12365 <= not w11684 and not w11708;
w12366 <= not w11660 and not w12365;
w12367 <= not w11683 and not w11707;
w12368 <= not w11704 and w12367;
w12369 <= not w11680 and w12368;
w12370 <= not w12366 and not w12369;
w12371 <= w11671 and w11676;
w12372 <= not w11666 and not w12371;
w12373 <= not w11671 and not w11676;
w12374 <= not w12372 and not w12373;
w12375 <= w11695 and w11700;
w12376 <= not w11690 and not w12375;
w12377 <= not w11695 and not w11700;
w12378 <= not w12376 and not w12377;
w12379 <= not w12374 and w12378;
w12380 <= w12374 and not w12378;
w12381 <= not w12379 and not w12380;
w12382 <= not w12370 and not w12381;
w12383 <= not w12369 and not w12379;
w12384 <= not w12380 and w12383;
w12385 <= not w12366 and w12384;
w12386 <= not w12382 and not w12385;
w12387 <= not w11626 and not w11650;
w12388 <= not w11602 and not w12387;
w12389 <= not w11625 and not w11649;
w12390 <= not w11646 and w12389;
w12391 <= not w11622 and w12390;
w12392 <= not w12388 and not w12391;
w12393 <= w11613 and w11618;
w12394 <= not w11608 and not w12393;
w12395 <= not w11613 and not w11618;
w12396 <= not w12394 and not w12395;
w12397 <= w11637 and w11642;
w12398 <= not w11632 and not w12397;
w12399 <= not w11637 and not w11642;
w12400 <= not w12398 and not w12399;
w12401 <= not w12396 and w12400;
w12402 <= w12396 and not w12400;
w12403 <= not w12401 and not w12402;
w12404 <= not w12392 and not w12403;
w12405 <= not w12391 and not w12401;
w12406 <= not w12402 and w12405;
w12407 <= not w12388 and w12406;
w12408 <= not w12404 and not w12407;
w12409 <= not w12386 and w12408;
w12410 <= w12386 and not w12408;
w12411 <= not w12409 and not w12410;
w12412 <= not w12364 and not w12411;
w12413 <= w12364 and w12411;
w12414 <= not w12412 and not w12413;
w12415 <= not w12360 and not w12414;
w12416 <= not w12359 and w12415;
w12417 <= not w12359 and not w12360;
w12418 <= w12414 and not w12417;
w12419 <= not w12416 and not w12418;
w12420 <= not w12281 and not w12419;
w12421 <= w12281 and w12419;
w12422 <= not w12420 and not w12421;
w12423 <= not w11138 and not w11400;
w12424 <= not w10876 and not w12423;
w12425 <= w11138 and w11400;
w12426 <= not w12424 and not w12425;
w12427 <= not w11268 and not w11394;
w12428 <= not w11142 and not w12427;
w12429 <= w11268 and w11394;
w12430 <= not w12428 and not w12429;
w12431 <= not w11330 and not w11388;
w12432 <= not w11272 and not w12431;
w12433 <= w11330 and w11388;
w12434 <= not w12432 and not w12433;
w12435 <= not w11358 and not w11382;
w12436 <= not w11334 and not w12435;
w12437 <= not w11357 and not w11381;
w12438 <= not w11378 and w12437;
w12439 <= not w11354 and w12438;
w12440 <= not w12436 and not w12439;
w12441 <= w11345 and w11350;
w12442 <= not w11340 and not w12441;
w12443 <= not w11345 and not w11350;
w12444 <= not w12442 and not w12443;
w12445 <= w11369 and w11374;
w12446 <= not w11364 and not w12445;
w12447 <= not w11369 and not w11374;
w12448 <= not w12446 and not w12447;
w12449 <= not w12444 and w12448;
w12450 <= w12444 and not w12448;
w12451 <= not w12449 and not w12450;
w12452 <= not w12440 and not w12451;
w12453 <= not w12439 and not w12449;
w12454 <= not w12450 and w12453;
w12455 <= not w12436 and w12454;
w12456 <= not w12452 and not w12455;
w12457 <= not w11300 and not w11324;
w12458 <= not w11276 and not w12457;
w12459 <= not w11299 and not w11323;
w12460 <= not w11320 and w12459;
w12461 <= not w11296 and w12460;
w12462 <= not w12458 and not w12461;
w12463 <= w11287 and w11292;
w12464 <= not w11282 and not w12463;
w12465 <= not w11287 and not w11292;
w12466 <= not w12464 and not w12465;
w12467 <= w11311 and w11316;
w12468 <= not w11306 and not w12467;
w12469 <= not w11311 and not w11316;
w12470 <= not w12468 and not w12469;
w12471 <= not w12466 and w12470;
w12472 <= w12466 and not w12470;
w12473 <= not w12471 and not w12472;
w12474 <= not w12462 and not w12473;
w12475 <= not w12461 and not w12471;
w12476 <= not w12472 and w12475;
w12477 <= not w12458 and w12476;
w12478 <= not w12474 and not w12477;
w12479 <= not w12456 and w12478;
w12480 <= w12456 and not w12478;
w12481 <= not w12479 and not w12480;
w12482 <= not w12434 and not w12481;
w12483 <= w12434 and w12481;
w12484 <= not w12482 and not w12483;
w12485 <= not w11204 and not w11262;
w12486 <= not w11146 and not w12485;
w12487 <= w11204 and w11262;
w12488 <= not w12486 and not w12487;
w12489 <= not w11232 and not w11256;
w12490 <= not w11208 and not w12489;
w12491 <= not w11231 and not w11255;
w12492 <= not w11252 and w12491;
w12493 <= not w11228 and w12492;
w12494 <= not w12490 and not w12493;
w12495 <= w11219 and w11224;
w12496 <= not w11214 and not w12495;
w12497 <= not w11219 and not w11224;
w12498 <= not w12496 and not w12497;
w12499 <= w11243 and w11248;
w12500 <= not w11238 and not w12499;
w12501 <= not w11243 and not w11248;
w12502 <= not w12500 and not w12501;
w12503 <= not w12498 and w12502;
w12504 <= w12498 and not w12502;
w12505 <= not w12503 and not w12504;
w12506 <= not w12494 and not w12505;
w12507 <= not w12493 and not w12503;
w12508 <= not w12504 and w12507;
w12509 <= not w12490 and w12508;
w12510 <= not w12506 and not w12509;
w12511 <= not w11174 and not w11198;
w12512 <= not w11150 and not w12511;
w12513 <= not w11173 and not w11197;
w12514 <= not w11194 and w12513;
w12515 <= not w11170 and w12514;
w12516 <= not w12512 and not w12515;
w12517 <= w11161 and w11166;
w12518 <= not w11156 and not w12517;
w12519 <= not w11161 and not w11166;
w12520 <= not w12518 and not w12519;
w12521 <= w11185 and w11190;
w12522 <= not w11180 and not w12521;
w12523 <= not w11185 and not w11190;
w12524 <= not w12522 and not w12523;
w12525 <= not w12520 and w12524;
w12526 <= w12520 and not w12524;
w12527 <= not w12525 and not w12526;
w12528 <= not w12516 and not w12527;
w12529 <= not w12515 and not w12525;
w12530 <= not w12526 and w12529;
w12531 <= not w12512 and w12530;
w12532 <= not w12528 and not w12531;
w12533 <= not w12510 and w12532;
w12534 <= w12510 and not w12532;
w12535 <= not w12533 and not w12534;
w12536 <= not w12488 and not w12535;
w12537 <= w12488 and w12535;
w12538 <= not w12536 and not w12537;
w12539 <= not w12484 and w12538;
w12540 <= w12484 and not w12538;
w12541 <= not w12539 and not w12540;
w12542 <= not w12430 and not w12541;
w12543 <= w12430 and w12541;
w12544 <= not w12542 and not w12543;
w12545 <= not w11006 and not w11132;
w12546 <= not w10880 and not w12545;
w12547 <= w11006 and w11132;
w12548 <= not w12546 and not w12547;
w12549 <= not w11068 and not w11126;
w12550 <= not w11010 and not w12549;
w12551 <= w11068 and w11126;
w12552 <= not w12550 and not w12551;
w12553 <= not w11096 and not w11120;
w12554 <= not w11072 and not w12553;
w12555 <= not w11095 and not w11119;
w12556 <= not w11116 and w12555;
w12557 <= not w11092 and w12556;
w12558 <= not w12554 and not w12557;
w12559 <= w11083 and w11088;
w12560 <= not w11078 and not w12559;
w12561 <= not w11083 and not w11088;
w12562 <= not w12560 and not w12561;
w12563 <= w11107 and w11112;
w12564 <= not w11102 and not w12563;
w12565 <= not w11107 and not w11112;
w12566 <= not w12564 and not w12565;
w12567 <= not w12562 and w12566;
w12568 <= w12562 and not w12566;
w12569 <= not w12567 and not w12568;
w12570 <= not w12558 and not w12569;
w12571 <= not w12557 and not w12567;
w12572 <= not w12568 and w12571;
w12573 <= not w12554 and w12572;
w12574 <= not w12570 and not w12573;
w12575 <= not w11038 and not w11062;
w12576 <= not w11014 and not w12575;
w12577 <= not w11037 and not w11061;
w12578 <= not w11058 and w12577;
w12579 <= not w11034 and w12578;
w12580 <= not w12576 and not w12579;
w12581 <= w11025 and w11030;
w12582 <= not w11020 and not w12581;
w12583 <= not w11025 and not w11030;
w12584 <= not w12582 and not w12583;
w12585 <= w11049 and w11054;
w12586 <= not w11044 and not w12585;
w12587 <= not w11049 and not w11054;
w12588 <= not w12586 and not w12587;
w12589 <= not w12584 and w12588;
w12590 <= w12584 and not w12588;
w12591 <= not w12589 and not w12590;
w12592 <= not w12580 and not w12591;
w12593 <= not w12579 and not w12589;
w12594 <= not w12590 and w12593;
w12595 <= not w12576 and w12594;
w12596 <= not w12592 and not w12595;
w12597 <= not w12574 and w12596;
w12598 <= w12574 and not w12596;
w12599 <= not w12597 and not w12598;
w12600 <= not w12552 and not w12599;
w12601 <= w12552 and w12599;
w12602 <= not w12600 and not w12601;
w12603 <= not w10942 and not w11000;
w12604 <= not w10884 and not w12603;
w12605 <= w10942 and w11000;
w12606 <= not w12604 and not w12605;
w12607 <= not w10970 and not w10994;
w12608 <= not w10946 and not w12607;
w12609 <= not w10969 and not w10993;
w12610 <= not w10990 and w12609;
w12611 <= not w10966 and w12610;
w12612 <= not w12608 and not w12611;
w12613 <= w10957 and w10962;
w12614 <= not w10952 and not w12613;
w12615 <= not w10957 and not w10962;
w12616 <= not w12614 and not w12615;
w12617 <= w10981 and w10986;
w12618 <= not w10976 and not w12617;
w12619 <= not w10981 and not w10986;
w12620 <= not w12618 and not w12619;
w12621 <= not w12616 and w12620;
w12622 <= w12616 and not w12620;
w12623 <= not w12621 and not w12622;
w12624 <= not w12612 and not w12623;
w12625 <= not w12611 and not w12621;
w12626 <= not w12622 and w12625;
w12627 <= not w12608 and w12626;
w12628 <= not w12624 and not w12627;
w12629 <= not w10912 and not w10936;
w12630 <= not w10888 and not w12629;
w12631 <= not w10911 and not w10935;
w12632 <= not w10932 and w12631;
w12633 <= not w10908 and w12632;
w12634 <= not w12630 and not w12633;
w12635 <= w10899 and w10904;
w12636 <= not w10894 and not w12635;
w12637 <= not w10899 and not w10904;
w12638 <= not w12636 and not w12637;
w12639 <= w10923 and w10928;
w12640 <= not w10918 and not w12639;
w12641 <= not w10923 and not w10928;
w12642 <= not w12640 and not w12641;
w12643 <= not w12638 and w12642;
w12644 <= w12638 and not w12642;
w12645 <= not w12643 and not w12644;
w12646 <= not w12634 and not w12645;
w12647 <= not w12633 and not w12643;
w12648 <= not w12644 and w12647;
w12649 <= not w12630 and w12648;
w12650 <= not w12646 and not w12649;
w12651 <= not w12628 and w12650;
w12652 <= w12628 and not w12650;
w12653 <= not w12651 and not w12652;
w12654 <= not w12606 and not w12653;
w12655 <= w12606 and w12653;
w12656 <= not w12654 and not w12655;
w12657 <= not w12602 and w12656;
w12658 <= w12602 and not w12656;
w12659 <= not w12657 and not w12658;
w12660 <= not w12548 and not w12659;
w12661 <= w12548 and w12659;
w12662 <= not w12660 and not w12661;
w12663 <= not w12544 and w12662;
w12664 <= w12544 and not w12662;
w12665 <= not w12663 and not w12664;
w12666 <= not w12426 and not w12665;
w12667 <= w12426 and w12665;
w12668 <= not w12666 and not w12667;
w12669 <= not w12422 and w12668;
w12670 <= w12422 and not w12668;
w12671 <= not w12669 and not w12670;
w12672 <= not w12276 and not w12671;
w12673 <= w12276 and w12671;
w12674 <= not w12672 and not w12673;
w12675 <= not w11999 and not w12261;
w12676 <= not w11737 and not w12675;
w12677 <= w11999 and w12261;
w12678 <= not w12676 and not w12677;
w12679 <= not w12129 and not w12255;
w12680 <= not w12003 and not w12679;
w12681 <= w12129 and w12255;
w12682 <= not w12680 and not w12681;
w12683 <= not w12191 and not w12249;
w12684 <= not w12133 and not w12683;
w12685 <= w12191 and w12249;
w12686 <= not w12684 and not w12685;
w12687 <= not w12219 and not w12243;
w12688 <= not w12195 and not w12687;
w12689 <= not w12218 and not w12242;
w12690 <= not w12239 and w12689;
w12691 <= not w12215 and w12690;
w12692 <= not w12688 and not w12691;
w12693 <= w12206 and w12211;
w12694 <= not w12201 and not w12693;
w12695 <= not w12206 and not w12211;
w12696 <= not w12694 and not w12695;
w12697 <= w12230 and w12235;
w12698 <= not w12225 and not w12697;
w12699 <= not w12230 and not w12235;
w12700 <= not w12698 and not w12699;
w12701 <= not w12696 and w12700;
w12702 <= w12696 and not w12700;
w12703 <= not w12701 and not w12702;
w12704 <= not w12692 and not w12703;
w12705 <= not w12691 and not w12701;
w12706 <= not w12702 and w12705;
w12707 <= not w12688 and w12706;
w12708 <= not w12704 and not w12707;
w12709 <= not w12161 and not w12185;
w12710 <= not w12137 and not w12709;
w12711 <= not w12160 and not w12184;
w12712 <= not w12181 and w12711;
w12713 <= not w12157 and w12712;
w12714 <= not w12710 and not w12713;
w12715 <= w12148 and w12153;
w12716 <= not w12143 and not w12715;
w12717 <= not w12148 and not w12153;
w12718 <= not w12716 and not w12717;
w12719 <= w12172 and w12177;
w12720 <= not w12167 and not w12719;
w12721 <= not w12172 and not w12177;
w12722 <= not w12720 and not w12721;
w12723 <= not w12718 and w12722;
w12724 <= w12718 and not w12722;
w12725 <= not w12723 and not w12724;
w12726 <= not w12714 and not w12725;
w12727 <= not w12713 and not w12723;
w12728 <= not w12724 and w12727;
w12729 <= not w12710 and w12728;
w12730 <= not w12726 and not w12729;
w12731 <= not w12708 and w12730;
w12732 <= w12708 and not w12730;
w12733 <= not w12731 and not w12732;
w12734 <= not w12686 and not w12733;
w12735 <= w12686 and w12733;
w12736 <= not w12734 and not w12735;
w12737 <= not w12065 and not w12123;
w12738 <= not w12007 and not w12737;
w12739 <= w12065 and w12123;
w12740 <= not w12738 and not w12739;
w12741 <= not w12093 and not w12117;
w12742 <= not w12069 and not w12741;
w12743 <= not w12092 and not w12116;
w12744 <= not w12113 and w12743;
w12745 <= not w12089 and w12744;
w12746 <= not w12742 and not w12745;
w12747 <= w12080 and w12085;
w12748 <= not w12075 and not w12747;
w12749 <= not w12080 and not w12085;
w12750 <= not w12748 and not w12749;
w12751 <= w12104 and w12109;
w12752 <= not w12099 and not w12751;
w12753 <= not w12104 and not w12109;
w12754 <= not w12752 and not w12753;
w12755 <= not w12750 and w12754;
w12756 <= w12750 and not w12754;
w12757 <= not w12755 and not w12756;
w12758 <= not w12746 and not w12757;
w12759 <= not w12745 and not w12755;
w12760 <= not w12756 and w12759;
w12761 <= not w12742 and w12760;
w12762 <= not w12758 and not w12761;
w12763 <= not w12035 and not w12059;
w12764 <= not w12011 and not w12763;
w12765 <= not w12034 and not w12058;
w12766 <= not w12055 and w12765;
w12767 <= not w12031 and w12766;
w12768 <= not w12764 and not w12767;
w12769 <= w12022 and w12027;
w12770 <= not w12017 and not w12769;
w12771 <= not w12022 and not w12027;
w12772 <= not w12770 and not w12771;
w12773 <= w12046 and w12051;
w12774 <= not w12041 and not w12773;
w12775 <= not w12046 and not w12051;
w12776 <= not w12774 and not w12775;
w12777 <= not w12772 and w12776;
w12778 <= w12772 and not w12776;
w12779 <= not w12777 and not w12778;
w12780 <= not w12768 and not w12779;
w12781 <= not w12767 and not w12777;
w12782 <= not w12778 and w12781;
w12783 <= not w12764 and w12782;
w12784 <= not w12780 and not w12783;
w12785 <= not w12762 and w12784;
w12786 <= w12762 and not w12784;
w12787 <= not w12785 and not w12786;
w12788 <= not w12740 and not w12787;
w12789 <= w12740 and w12787;
w12790 <= not w12788 and not w12789;
w12791 <= not w12736 and w12790;
w12792 <= w12736 and not w12790;
w12793 <= not w12791 and not w12792;
w12794 <= not w12682 and not w12793;
w12795 <= w12682 and w12793;
w12796 <= not w12794 and not w12795;
w12797 <= not w11867 and not w11993;
w12798 <= not w11741 and not w12797;
w12799 <= w11867 and w11993;
w12800 <= not w12798 and not w12799;
w12801 <= not w11929 and not w11987;
w12802 <= not w11871 and not w12801;
w12803 <= w11929 and w11987;
w12804 <= not w12802 and not w12803;
w12805 <= not w11957 and not w11981;
w12806 <= not w11933 and not w12805;
w12807 <= not w11956 and not w11980;
w12808 <= not w11977 and w12807;
w12809 <= not w11953 and w12808;
w12810 <= not w12806 and not w12809;
w12811 <= w11944 and w11949;
w12812 <= not w11939 and not w12811;
w12813 <= not w11944 and not w11949;
w12814 <= not w12812 and not w12813;
w12815 <= w11968 and w11973;
w12816 <= not w11963 and not w12815;
w12817 <= not w11968 and not w11973;
w12818 <= not w12816 and not w12817;
w12819 <= not w12814 and w12818;
w12820 <= w12814 and not w12818;
w12821 <= not w12819 and not w12820;
w12822 <= not w12810 and not w12821;
w12823 <= not w12809 and not w12819;
w12824 <= not w12820 and w12823;
w12825 <= not w12806 and w12824;
w12826 <= not w12822 and not w12825;
w12827 <= not w11899 and not w11923;
w12828 <= not w11875 and not w12827;
w12829 <= not w11898 and not w11922;
w12830 <= not w11919 and w12829;
w12831 <= not w11895 and w12830;
w12832 <= not w12828 and not w12831;
w12833 <= w11886 and w11891;
w12834 <= not w11881 and not w12833;
w12835 <= not w11886 and not w11891;
w12836 <= not w12834 and not w12835;
w12837 <= w11910 and w11915;
w12838 <= not w11905 and not w12837;
w12839 <= not w11910 and not w11915;
w12840 <= not w12838 and not w12839;
w12841 <= not w12836 and w12840;
w12842 <= w12836 and not w12840;
w12843 <= not w12841 and not w12842;
w12844 <= not w12832 and not w12843;
w12845 <= not w12831 and not w12841;
w12846 <= not w12842 and w12845;
w12847 <= not w12828 and w12846;
w12848 <= not w12844 and not w12847;
w12849 <= not w12826 and w12848;
w12850 <= w12826 and not w12848;
w12851 <= not w12849 and not w12850;
w12852 <= not w12804 and not w12851;
w12853 <= w12804 and w12851;
w12854 <= not w12852 and not w12853;
w12855 <= not w11803 and not w11861;
w12856 <= not w11745 and not w12855;
w12857 <= w11803 and w11861;
w12858 <= not w12856 and not w12857;
w12859 <= not w11831 and not w11855;
w12860 <= not w11807 and not w12859;
w12861 <= not w11830 and not w11854;
w12862 <= not w11851 and w12861;
w12863 <= not w11827 and w12862;
w12864 <= not w12860 and not w12863;
w12865 <= w11818 and w11823;
w12866 <= not w11813 and not w12865;
w12867 <= not w11818 and not w11823;
w12868 <= not w12866 and not w12867;
w12869 <= w11842 and w11847;
w12870 <= not w11837 and not w12869;
w12871 <= not w11842 and not w11847;
w12872 <= not w12870 and not w12871;
w12873 <= not w12868 and w12872;
w12874 <= w12868 and not w12872;
w12875 <= not w12873 and not w12874;
w12876 <= not w12864 and not w12875;
w12877 <= not w12863 and not w12873;
w12878 <= not w12874 and w12877;
w12879 <= not w12860 and w12878;
w12880 <= not w12876 and not w12879;
w12881 <= not w11773 and not w11797;
w12882 <= not w11749 and not w12881;
w12883 <= not w11772 and not w11796;
w12884 <= not w11793 and w12883;
w12885 <= not w11769 and w12884;
w12886 <= not w12882 and not w12885;
w12887 <= w11760 and w11765;
w12888 <= not w11755 and not w12887;
w12889 <= not w11760 and not w11765;
w12890 <= not w12888 and not w12889;
w12891 <= w11784 and w11789;
w12892 <= not w11779 and not w12891;
w12893 <= not w11784 and not w11789;
w12894 <= not w12892 and not w12893;
w12895 <= not w12890 and w12894;
w12896 <= w12890 and not w12894;
w12897 <= not w12895 and not w12896;
w12898 <= not w12886 and not w12897;
w12899 <= not w12885 and not w12895;
w12900 <= not w12896 and w12899;
w12901 <= not w12882 and w12900;
w12902 <= not w12898 and not w12901;
w12903 <= not w12880 and w12902;
w12904 <= w12880 and not w12902;
w12905 <= not w12903 and not w12904;
w12906 <= not w12858 and not w12905;
w12907 <= w12858 and w12905;
w12908 <= not w12906 and not w12907;
w12909 <= not w12854 and w12908;
w12910 <= w12854 and not w12908;
w12911 <= not w12909 and not w12910;
w12912 <= not w12800 and not w12911;
w12913 <= w12800 and w12911;
w12914 <= not w12912 and not w12913;
w12915 <= not w12796 and w12914;
w12916 <= w12796 and not w12914;
w12917 <= not w12915 and not w12916;
w12918 <= not w12678 and not w12917;
w12919 <= w12678 and w12917;
w12920 <= not w12918 and not w12919;
w12921 <= not w12674 and not w12920;
w12922 <= not w12272 and not w12921;
w12923 <= not w12672 and w12920;
w12924 <= not w12673 and w12923;
w12925 <= not w12922 and not w12924;
w12926 <= not w12422 and not w12668;
w12927 <= not w12276 and not w12926;
w12928 <= w12422 and w12668;
w12929 <= not w12927 and not w12928;
w12930 <= not w12544 and not w12662;
w12931 <= not w12426 and not w12930;
w12932 <= w12544 and w12662;
w12933 <= not w12931 and not w12932;
w12934 <= not w12602 and not w12656;
w12935 <= not w12548 and not w12934;
w12936 <= w12602 and w12656;
w12937 <= not w12935 and not w12936;
w12938 <= not w12628 and not w12650;
w12939 <= not w12606 and not w12938;
w12940 <= not w12627 and not w12649;
w12941 <= not w12646 and w12940;
w12942 <= not w12624 and w12941;
w12943 <= not w12939 and not w12942;
w12944 <= not w12637 and not w12641;
w12945 <= not w12640 and w12944;
w12946 <= not w12636 and w12945;
w12947 <= not w12634 and not w12946;
w12948 <= not w12638 and not w12642;
w12949 <= not w12947 and not w12948;
w12950 <= not w12615 and not w12619;
w12951 <= not w12618 and w12950;
w12952 <= not w12614 and w12951;
w12953 <= not w12612 and not w12952;
w12954 <= not w12616 and not w12620;
w12955 <= not w12953 and not w12954;
w12956 <= not w12949 and w12955;
w12957 <= w12949 and not w12955;
w12958 <= not w12956 and not w12957;
w12959 <= not w12943 and not w12958;
w12960 <= not w12942 and not w12956;
w12961 <= not w12957 and w12960;
w12962 <= not w12939 and w12961;
w12963 <= not w12959 and not w12962;
w12964 <= not w12574 and not w12596;
w12965 <= not w12552 and not w12964;
w12966 <= not w12573 and not w12595;
w12967 <= not w12592 and w12966;
w12968 <= not w12570 and w12967;
w12969 <= not w12965 and not w12968;
w12970 <= not w12583 and not w12587;
w12971 <= not w12586 and w12970;
w12972 <= not w12582 and w12971;
w12973 <= not w12580 and not w12972;
w12974 <= not w12584 and not w12588;
w12975 <= not w12973 and not w12974;
w12976 <= not w12561 and not w12565;
w12977 <= not w12564 and w12976;
w12978 <= not w12560 and w12977;
w12979 <= not w12558 and not w12978;
w12980 <= not w12562 and not w12566;
w12981 <= not w12979 and not w12980;
w12982 <= not w12975 and w12981;
w12983 <= w12975 and not w12981;
w12984 <= not w12982 and not w12983;
w12985 <= not w12969 and not w12984;
w12986 <= not w12968 and not w12982;
w12987 <= not w12983 and w12986;
w12988 <= not w12965 and w12987;
w12989 <= not w12985 and not w12988;
w12990 <= not w12963 and w12989;
w12991 <= w12963 and not w12989;
w12992 <= not w12990 and not w12991;
w12993 <= not w12937 and not w12992;
w12994 <= w12937 and w12992;
w12995 <= not w12993 and not w12994;
w12996 <= not w12484 and not w12538;
w12997 <= not w12430 and not w12996;
w12998 <= w12484 and w12538;
w12999 <= not w12997 and not w12998;
w13000 <= not w12510 and not w12532;
w13001 <= not w12488 and not w13000;
w13002 <= not w12509 and not w12531;
w13003 <= not w12528 and w13002;
w13004 <= not w12506 and w13003;
w13005 <= not w13001 and not w13004;
w13006 <= not w12519 and not w12523;
w13007 <= not w12522 and w13006;
w13008 <= not w12518 and w13007;
w13009 <= not w12516 and not w13008;
w13010 <= not w12520 and not w12524;
w13011 <= not w13009 and not w13010;
w13012 <= not w12497 and not w12501;
w13013 <= not w12500 and w13012;
w13014 <= not w12496 and w13013;
w13015 <= not w12494 and not w13014;
w13016 <= not w12498 and not w12502;
w13017 <= not w13015 and not w13016;
w13018 <= not w13011 and w13017;
w13019 <= w13011 and not w13017;
w13020 <= not w13018 and not w13019;
w13021 <= not w13005 and not w13020;
w13022 <= not w13004 and not w13018;
w13023 <= not w13019 and w13022;
w13024 <= not w13001 and w13023;
w13025 <= not w13021 and not w13024;
w13026 <= not w12456 and not w12478;
w13027 <= not w12434 and not w13026;
w13028 <= not w12455 and not w12477;
w13029 <= not w12474 and w13028;
w13030 <= not w12452 and w13029;
w13031 <= not w13027 and not w13030;
w13032 <= not w12465 and not w12469;
w13033 <= not w12468 and w13032;
w13034 <= not w12464 and w13033;
w13035 <= not w12462 and not w13034;
w13036 <= not w12466 and not w12470;
w13037 <= not w13035 and not w13036;
w13038 <= not w12443 and not w12447;
w13039 <= not w12446 and w13038;
w13040 <= not w12442 and w13039;
w13041 <= not w12440 and not w13040;
w13042 <= not w12444 and not w12448;
w13043 <= not w13041 and not w13042;
w13044 <= not w13037 and w13043;
w13045 <= w13037 and not w13043;
w13046 <= not w13044 and not w13045;
w13047 <= not w13031 and not w13046;
w13048 <= not w13030 and not w13044;
w13049 <= not w13045 and w13048;
w13050 <= not w13027 and w13049;
w13051 <= not w13047 and not w13050;
w13052 <= not w13025 and w13051;
w13053 <= w13025 and not w13051;
w13054 <= not w13052 and not w13053;
w13055 <= not w12999 and not w13054;
w13056 <= w12999 and w13054;
w13057 <= not w13055 and not w13056;
w13058 <= not w12995 and w13057;
w13059 <= w12995 and not w13057;
w13060 <= not w13058 and not w13059;
w13061 <= not w12933 and not w13060;
w13062 <= w12933 and w13060;
w13063 <= not w13061 and not w13062;
w13064 <= not w12414 and not w12417;
w13065 <= not w12281 and not w13064;
w13066 <= not w12360 and w12414;
w13067 <= not w12359 and w13066;
w13068 <= not w13065 and not w13067;
w13069 <= not w12353 and not w12356;
w13070 <= not w12286 and not w13069;
w13071 <= not w12331 and w12353;
w13072 <= not w12330 and w13071;
w13073 <= not w13070 and not w13072;
w13074 <= not w12304 and not w12326;
w13075 <= not w12290 and not w13074;
w13076 <= not w12303 and not w12325;
w13077 <= not w12322 and w13076;
w13078 <= not w12301 and w13077;
w13079 <= not w13075 and not w13078;
w13080 <= not w12313 and not w12317;
w13081 <= not w12316 and w13080;
w13082 <= not w12312 and w13081;
w13083 <= not w12310 and not w13082;
w13084 <= not w12314 and not w12318;
w13085 <= not w13083 and not w13084;
w13086 <= not w12292 and not w12297;
w13087 <= not w12299 and not w13086;
w13088 <= not w13085 and w13087;
w13089 <= w13085 and not w13087;
w13090 <= not w13088 and not w13089;
w13091 <= not w13079 and not w13090;
w13092 <= not w13078 and not w13088;
w13093 <= not w13089 and w13092;
w13094 <= not w13075 and w13093;
w13095 <= not w12340 and not w12344;
w13096 <= not w12343 and w13095;
w13097 <= not w12339 and w13096;
w13098 <= not w12337 and not w13097;
w13099 <= not w12341 and not w12345;
w13100 <= not w13098 and not w13099;
w13101 <= not w13094 and w13100;
w13102 <= not w13091 and w13101;
w13103 <= not w13091 and not w13094;
w13104 <= not w13100 and not w13103;
w13105 <= not w13102 and not w13104;
w13106 <= not w13073 and not w13105;
w13107 <= not w13072 and not w13102;
w13108 <= not w13070 and w13107;
w13109 <= not w13104 and w13108;
w13110 <= not w13106 and not w13109;
w13111 <= not w12386 and not w12408;
w13112 <= not w12364 and not w13111;
w13113 <= not w12385 and not w12407;
w13114 <= not w12404 and w13113;
w13115 <= not w12382 and w13114;
w13116 <= not w13112 and not w13115;
w13117 <= not w12395 and not w12399;
w13118 <= not w12398 and w13117;
w13119 <= not w12394 and w13118;
w13120 <= not w12392 and not w13119;
w13121 <= not w12396 and not w12400;
w13122 <= not w13120 and not w13121;
w13123 <= not w12373 and not w12377;
w13124 <= not w12376 and w13123;
w13125 <= not w12372 and w13124;
w13126 <= not w12370 and not w13125;
w13127 <= not w12374 and not w12378;
w13128 <= not w13126 and not w13127;
w13129 <= not w13122 and w13128;
w13130 <= w13122 and not w13128;
w13131 <= not w13129 and not w13130;
w13132 <= not w13116 and not w13131;
w13133 <= not w13115 and not w13129;
w13134 <= not w13130 and w13133;
w13135 <= not w13112 and w13134;
w13136 <= not w13132 and not w13135;
w13137 <= not w13110 and w13136;
w13138 <= not w13106 and not w13136;
w13139 <= not w13109 and w13138;
w13140 <= not w13137 and not w13139;
w13141 <= not w13068 and not w13140;
w13142 <= w13068 and w13140;
w13143 <= not w13141 and not w13142;
w13144 <= not w13063 and w13143;
w13145 <= w13063 and not w13143;
w13146 <= not w13144 and not w13145;
w13147 <= not w12929 and not w13146;
w13148 <= w12929 and w13146;
w13149 <= not w13147 and not w13148;
w13150 <= not w12796 and not w12914;
w13151 <= not w12678 and not w13150;
w13152 <= w12796 and w12914;
w13153 <= not w13151 and not w13152;
w13154 <= not w12854 and not w12908;
w13155 <= not w12800 and not w13154;
w13156 <= w12854 and w12908;
w13157 <= not w13155 and not w13156;
w13158 <= not w12880 and not w12902;
w13159 <= not w12858 and not w13158;
w13160 <= not w12879 and not w12901;
w13161 <= not w12898 and w13160;
w13162 <= not w12876 and w13161;
w13163 <= not w13159 and not w13162;
w13164 <= not w12889 and not w12893;
w13165 <= not w12892 and w13164;
w13166 <= not w12888 and w13165;
w13167 <= not w12886 and not w13166;
w13168 <= not w12890 and not w12894;
w13169 <= not w13167 and not w13168;
w13170 <= not w12867 and not w12871;
w13171 <= not w12870 and w13170;
w13172 <= not w12866 and w13171;
w13173 <= not w12864 and not w13172;
w13174 <= not w12868 and not w12872;
w13175 <= not w13173 and not w13174;
w13176 <= not w13169 and w13175;
w13177 <= w13169 and not w13175;
w13178 <= not w13176 and not w13177;
w13179 <= not w13163 and not w13178;
w13180 <= not w13162 and not w13176;
w13181 <= not w13177 and w13180;
w13182 <= not w13159 and w13181;
w13183 <= not w13179 and not w13182;
w13184 <= not w12826 and not w12848;
w13185 <= not w12804 and not w13184;
w13186 <= not w12825 and not w12847;
w13187 <= not w12844 and w13186;
w13188 <= not w12822 and w13187;
w13189 <= not w13185 and not w13188;
w13190 <= not w12835 and not w12839;
w13191 <= not w12838 and w13190;
w13192 <= not w12834 and w13191;
w13193 <= not w12832 and not w13192;
w13194 <= not w12836 and not w12840;
w13195 <= not w13193 and not w13194;
w13196 <= not w12813 and not w12817;
w13197 <= not w12816 and w13196;
w13198 <= not w12812 and w13197;
w13199 <= not w12810 and not w13198;
w13200 <= not w12814 and not w12818;
w13201 <= not w13199 and not w13200;
w13202 <= not w13195 and w13201;
w13203 <= w13195 and not w13201;
w13204 <= not w13202 and not w13203;
w13205 <= not w13189 and not w13204;
w13206 <= not w13188 and not w13202;
w13207 <= not w13203 and w13206;
w13208 <= not w13185 and w13207;
w13209 <= not w13205 and not w13208;
w13210 <= not w13183 and w13209;
w13211 <= w13183 and not w13209;
w13212 <= not w13210 and not w13211;
w13213 <= not w13157 and not w13212;
w13214 <= w13157 and w13212;
w13215 <= not w13213 and not w13214;
w13216 <= not w12736 and not w12790;
w13217 <= not w12682 and not w13216;
w13218 <= w12736 and w12790;
w13219 <= not w13217 and not w13218;
w13220 <= not w12762 and not w12784;
w13221 <= not w12740 and not w13220;
w13222 <= not w12761 and not w12783;
w13223 <= not w12780 and w13222;
w13224 <= not w12758 and w13223;
w13225 <= not w13221 and not w13224;
w13226 <= not w12771 and not w12775;
w13227 <= not w12774 and w13226;
w13228 <= not w12770 and w13227;
w13229 <= not w12768 and not w13228;
w13230 <= not w12772 and not w12776;
w13231 <= not w13229 and not w13230;
w13232 <= not w12749 and not w12753;
w13233 <= not w12752 and w13232;
w13234 <= not w12748 and w13233;
w13235 <= not w12746 and not w13234;
w13236 <= not w12750 and not w12754;
w13237 <= not w13235 and not w13236;
w13238 <= not w13231 and w13237;
w13239 <= w13231 and not w13237;
w13240 <= not w13238 and not w13239;
w13241 <= not w13225 and not w13240;
w13242 <= not w13224 and not w13238;
w13243 <= not w13239 and w13242;
w13244 <= not w13221 and w13243;
w13245 <= not w13241 and not w13244;
w13246 <= not w12708 and not w12730;
w13247 <= not w12686 and not w13246;
w13248 <= not w12707 and not w12729;
w13249 <= not w12726 and w13248;
w13250 <= not w12704 and w13249;
w13251 <= not w13247 and not w13250;
w13252 <= not w12717 and not w12721;
w13253 <= not w12720 and w13252;
w13254 <= not w12716 and w13253;
w13255 <= not w12714 and not w13254;
w13256 <= not w12718 and not w12722;
w13257 <= not w13255 and not w13256;
w13258 <= not w12695 and not w12699;
w13259 <= not w12698 and w13258;
w13260 <= not w12694 and w13259;
w13261 <= not w12692 and not w13260;
w13262 <= not w12696 and not w12700;
w13263 <= not w13261 and not w13262;
w13264 <= not w13257 and w13263;
w13265 <= w13257 and not w13263;
w13266 <= not w13264 and not w13265;
w13267 <= not w13251 and not w13266;
w13268 <= not w13250 and not w13264;
w13269 <= not w13265 and w13268;
w13270 <= not w13247 and w13269;
w13271 <= not w13267 and not w13270;
w13272 <= not w13245 and w13271;
w13273 <= w13245 and not w13271;
w13274 <= not w13272 and not w13273;
w13275 <= not w13219 and not w13274;
w13276 <= w13219 and w13274;
w13277 <= not w13275 and not w13276;
w13278 <= not w13215 and w13277;
w13279 <= w13215 and not w13277;
w13280 <= not w13278 and not w13279;
w13281 <= not w13153 and not w13280;
w13282 <= w13153 and w13280;
w13283 <= not w13281 and not w13282;
w13284 <= not w13149 and not w13283;
w13285 <= not w12925 and not w13284;
w13286 <= not w13147 and w13283;
w13287 <= not w13148 and w13286;
w13288 <= not w13285 and not w13287;
w13289 <= not w13063 and not w13143;
w13290 <= not w12929 and not w13289;
w13291 <= w13063 and w13143;
w13292 <= not w13290 and not w13291;
w13293 <= not w13110 and not w13136;
w13294 <= not w13068 and not w13293;
w13295 <= not w13106 and w13136;
w13296 <= not w13109 and w13295;
w13297 <= not w13294 and not w13296;
w13298 <= not w13121 and not w13127;
w13299 <= not w13126 and w13298;
w13300 <= not w13120 and w13299;
w13301 <= not w13116 and not w13300;
w13302 <= not w13122 and not w13128;
w13303 <= not w13301 and not w13302;
w13304 <= w13100 and not w13103;
w13305 <= not w13073 and not w13304;
w13306 <= not w13094 and not w13100;
w13307 <= not w13091 and w13306;
w13308 <= not w13305 and not w13307;
w13309 <= not w12299 and not w13084;
w13310 <= not w13086 and w13309;
w13311 <= not w13083 and w13310;
w13312 <= not w13079 and not w13311;
w13313 <= not w13085 and not w13087;
w13314 <= not w13312 and not w13313;
w13315 <= not w13308 and w13314;
w13316 <= not w13307 and not w13314;
w13317 <= not w13305 and w13316;
w13318 <= not w13315 and not w13317;
w13319 <= not w13303 and not w13318;
w13320 <= w13303 and not w13317;
w13321 <= not w13315 and w13320;
w13322 <= not w13319 and not w13321;
w13323 <= not w13297 and w13322;
w13324 <= w13297 and not w13322;
w13325 <= not w13323 and not w13324;
w13326 <= not w12995 and not w13057;
w13327 <= not w12933 and not w13326;
w13328 <= w12995 and w13057;
w13329 <= not w13327 and not w13328;
w13330 <= not w13025 and not w13051;
w13331 <= not w12999 and not w13330;
w13332 <= not w13024 and not w13050;
w13333 <= not w13047 and w13332;
w13334 <= not w13021 and w13333;
w13335 <= not w13331 and not w13334;
w13336 <= not w13010 and not w13016;
w13337 <= not w13015 and w13336;
w13338 <= not w13009 and w13337;
w13339 <= not w13005 and not w13338;
w13340 <= not w13011 and not w13017;
w13341 <= not w13339 and not w13340;
w13342 <= not w13036 and not w13042;
w13343 <= not w13041 and w13342;
w13344 <= not w13035 and w13343;
w13345 <= not w13031 and not w13344;
w13346 <= not w13037 and not w13043;
w13347 <= not w13345 and not w13346;
w13348 <= not w13341 and w13347;
w13349 <= w13341 and not w13347;
w13350 <= not w13348 and not w13349;
w13351 <= not w13335 and not w13350;
w13352 <= not w13334 and not w13348;
w13353 <= not w13349 and w13352;
w13354 <= not w13331 and w13353;
w13355 <= not w13351 and not w13354;
w13356 <= not w12963 and not w12989;
w13357 <= not w12937 and not w13356;
w13358 <= not w12962 and not w12988;
w13359 <= not w12985 and w13358;
w13360 <= not w12959 and w13359;
w13361 <= not w13357 and not w13360;
w13362 <= not w12948 and not w12954;
w13363 <= not w12953 and w13362;
w13364 <= not w12947 and w13363;
w13365 <= not w12943 and not w13364;
w13366 <= not w12949 and not w12955;
w13367 <= not w13365 and not w13366;
w13368 <= not w12974 and not w12980;
w13369 <= not w12979 and w13368;
w13370 <= not w12973 and w13369;
w13371 <= not w12969 and not w13370;
w13372 <= not w12975 and not w12981;
w13373 <= not w13371 and not w13372;
w13374 <= not w13367 and w13373;
w13375 <= w13367 and not w13373;
w13376 <= not w13374 and not w13375;
w13377 <= not w13361 and not w13376;
w13378 <= not w13360 and not w13374;
w13379 <= not w13375 and w13378;
w13380 <= not w13357 and w13379;
w13381 <= not w13377 and not w13380;
w13382 <= not w13355 and w13381;
w13383 <= w13355 and not w13381;
w13384 <= not w13382 and not w13383;
w13385 <= not w13329 and not w13384;
w13386 <= w13329 and w13384;
w13387 <= not w13385 and not w13386;
w13388 <= not w13325 and w13387;
w13389 <= w13325 and not w13387;
w13390 <= not w13388 and not w13389;
w13391 <= not w13292 and not w13390;
w13392 <= w13292 and w13390;
w13393 <= not w13391 and not w13392;
w13394 <= not w13215 and not w13277;
w13395 <= not w13153 and not w13394;
w13396 <= w13215 and w13277;
w13397 <= not w13395 and not w13396;
w13398 <= not w13245 and not w13271;
w13399 <= not w13219 and not w13398;
w13400 <= not w13244 and not w13270;
w13401 <= not w13267 and w13400;
w13402 <= not w13241 and w13401;
w13403 <= not w13399 and not w13402;
w13404 <= not w13230 and not w13236;
w13405 <= not w13235 and w13404;
w13406 <= not w13229 and w13405;
w13407 <= not w13225 and not w13406;
w13408 <= not w13231 and not w13237;
w13409 <= not w13407 and not w13408;
w13410 <= not w13256 and not w13262;
w13411 <= not w13261 and w13410;
w13412 <= not w13255 and w13411;
w13413 <= not w13251 and not w13412;
w13414 <= not w13257 and not w13263;
w13415 <= not w13413 and not w13414;
w13416 <= not w13409 and w13415;
w13417 <= w13409 and not w13415;
w13418 <= not w13416 and not w13417;
w13419 <= not w13403 and not w13418;
w13420 <= not w13402 and not w13416;
w13421 <= not w13417 and w13420;
w13422 <= not w13399 and w13421;
w13423 <= not w13419 and not w13422;
w13424 <= not w13183 and not w13209;
w13425 <= not w13157 and not w13424;
w13426 <= not w13182 and not w13208;
w13427 <= not w13205 and w13426;
w13428 <= not w13179 and w13427;
w13429 <= not w13425 and not w13428;
w13430 <= not w13168 and not w13174;
w13431 <= not w13173 and w13430;
w13432 <= not w13167 and w13431;
w13433 <= not w13163 and not w13432;
w13434 <= not w13169 and not w13175;
w13435 <= not w13433 and not w13434;
w13436 <= not w13194 and not w13200;
w13437 <= not w13199 and w13436;
w13438 <= not w13193 and w13437;
w13439 <= not w13189 and not w13438;
w13440 <= not w13195 and not w13201;
w13441 <= not w13439 and not w13440;
w13442 <= not w13435 and w13441;
w13443 <= w13435 and not w13441;
w13444 <= not w13442 and not w13443;
w13445 <= not w13429 and not w13444;
w13446 <= not w13428 and not w13442;
w13447 <= not w13443 and w13446;
w13448 <= not w13425 and w13447;
w13449 <= not w13445 and not w13448;
w13450 <= not w13423 and w13449;
w13451 <= w13423 and not w13449;
w13452 <= not w13450 and not w13451;
w13453 <= not w13397 and not w13452;
w13454 <= w13397 and w13452;
w13455 <= not w13453 and not w13454;
w13456 <= not w13393 and not w13455;
w13457 <= not w13288 and not w13456;
w13458 <= not w13391 and w13455;
w13459 <= not w13392 and w13458;
w13460 <= not w13457 and not w13459;
w13461 <= not w13325 and not w13387;
w13462 <= not w13292 and not w13461;
w13463 <= w13325 and w13387;
w13464 <= not w13462 and not w13463;
w13465 <= not w13297 and not w13321;
w13466 <= not w13319 and not w13465;
w13467 <= not w13308 and not w13314;
w13468 <= not w13466 and w13467;
w13469 <= not w13319 and not w13467;
w13470 <= not w13465 and w13469;
w13471 <= not w13468 and not w13470;
w13472 <= not w13355 and not w13381;
w13473 <= not w13329 and not w13472;
w13474 <= not w13354 and not w13380;
w13475 <= not w13377 and w13474;
w13476 <= not w13351 and w13475;
w13477 <= not w13473 and not w13476;
w13478 <= not w13366 and not w13372;
w13479 <= not w13371 and w13478;
w13480 <= not w13365 and w13479;
w13481 <= not w13361 and not w13480;
w13482 <= not w13367 and not w13373;
w13483 <= not w13481 and not w13482;
w13484 <= not w13340 and not w13346;
w13485 <= not w13345 and w13484;
w13486 <= not w13339 and w13485;
w13487 <= not w13335 and not w13486;
w13488 <= not w13341 and not w13347;
w13489 <= not w13487 and not w13488;
w13490 <= not w13483 and w13489;
w13491 <= w13483 and not w13489;
w13492 <= not w13490 and not w13491;
w13493 <= not w13477 and not w13492;
w13494 <= not w13476 and not w13490;
w13495 <= not w13491 and w13494;
w13496 <= not w13473 and w13495;
w13497 <= not w13493 and not w13496;
w13498 <= not w13471 and not w13497;
w13499 <= not w13470 and not w13496;
w13500 <= not w13468 and w13499;
w13501 <= not w13493 and w13500;
w13502 <= not w13498 and not w13501;
w13503 <= not w13464 and w13502;
w13504 <= w13464 and not w13502;
w13505 <= not w13503 and not w13504;
w13506 <= not w13423 and not w13449;
w13507 <= not w13397 and not w13506;
w13508 <= not w13422 and not w13448;
w13509 <= not w13445 and w13508;
w13510 <= not w13419 and w13509;
w13511 <= not w13507 and not w13510;
w13512 <= not w13434 and not w13440;
w13513 <= not w13439 and w13512;
w13514 <= not w13433 and w13513;
w13515 <= not w13429 and not w13514;
w13516 <= not w13435 and not w13441;
w13517 <= not w13515 and not w13516;
w13518 <= not w13408 and not w13414;
w13519 <= not w13413 and w13518;
w13520 <= not w13407 and w13519;
w13521 <= not w13403 and not w13520;
w13522 <= not w13409 and not w13415;
w13523 <= not w13521 and not w13522;
w13524 <= not w13517 and w13523;
w13525 <= w13517 and not w13523;
w13526 <= not w13524 and not w13525;
w13527 <= not w13511 and not w13526;
w13528 <= not w13510 and not w13524;
w13529 <= not w13525 and w13528;
w13530 <= not w13507 and w13529;
w13531 <= not w13527 and not w13530;
w13532 <= not w13505 and not w13531;
w13533 <= not w13460 and not w13532;
w13534 <= not w13503 and w13531;
w13535 <= not w13504 and w13534;
w13536 <= not w13533 and not w13535;
w13537 <= not w13464 and not w13498;
w13538 <= not w13501 and not w13537;
w13539 <= not w13482 and not w13488;
w13540 <= not w13487 and w13539;
w13541 <= not w13481 and w13540;
w13542 <= not w13477 and not w13541;
w13543 <= not w13483 and not w13489;
w13544 <= not w13468 and not w13543;
w13545 <= not w13542 and w13544;
w13546 <= not w13542 and not w13543;
w13547 <= w13468 and not w13546;
w13548 <= not w13545 and not w13547;
w13549 <= not w13538 and w13548;
w13550 <= not w13501 and not w13548;
w13551 <= not w13537 and w13550;
w13552 <= not w13549 and not w13551;
w13553 <= not w13516 and not w13522;
w13554 <= not w13521 and w13553;
w13555 <= not w13515 and w13554;
w13556 <= not w13511 and not w13555;
w13557 <= not w13517 and not w13523;
w13558 <= not w13556 and not w13557;
w13559 <= not w13552 and w13558;
w13560 <= not w13536 and not w13559;
w13561 <= not w13551 and not w13558;
w13562 <= not w13549 and w13561;
w13563 <= not w13560 and not w13562;
w13564 <= not w13538 and not w13545;
w13565 <= not w13547 and not w13564;
w13566 <= not w13563 and w13565;
w13567 <= not w13562 and not w13565;
w13568 <= not w13560 and w13567;
w13569 <= not w13566 and not w13568;
w13570 <= not w13552 and not w13558;
w13571 <= not w13551 and w13558;
w13572 <= not w13549 and w13571;
w13573 <= not w13535 and not w13572;
w13574 <= not w13533 and w13573;
w13575 <= not w13570 and w13574;
w13576 <= not w13570 and not w13572;
w13577 <= not w13536 and not w13576;
w13578 <= not w13505 and w13531;
w13579 <= not w13503 and not w13531;
w13580 <= not w13504 and w13579;
w13581 <= not w13578 and not w13580;
w13582 <= w13460 and w13581;
w13583 <= not w13460 and not w13581;
w13584 <= not w13391 and not w13455;
w13585 <= not w13392 and w13584;
w13586 <= not w13393 and w13455;
w13587 <= not w13585 and not w13586;
w13588 <= w13288 and w13587;
w13589 <= not w13288 and not w13587;
w13590 <= not w13149 and w13283;
w13591 <= not w13147 and not w13283;
w13592 <= not w13148 and w13591;
w13593 <= not w13590 and not w13592;
w13594 <= w12925 and w13593;
w13595 <= not w12925 and not w13593;
w13596 <= not w12672 and not w12920;
w13597 <= not w12673 and w13596;
w13598 <= not w12674 and w12920;
w13599 <= not w13597 and not w13598;
w13600 <= w12272 and w13599;
w13601 <= not w12272 and not w13599;
w13602 <= not w11733 and w12267;
w13603 <= not w11731 and not w12267;
w13604 <= not w11732 and w13603;
w13605 <= not w13602 and not w13604;
w13606 <= w10868 and w13605;
w13607 <= not w10868 and not w13605;
w13608 <= not w10165 and not w10863;
w13609 <= not w10166 and w13608;
w13610 <= not w10167 and w10863;
w13611 <= not w13609 and not w13610;
w13612 <= not w9044 and not w13611;
w13613 <= not w9029 and not w9030;
w13614 <= not w9031 and w13613;
w13615 <= w9029 and not w9032;
w13616 <= not w13614 and not w13615;
w13617 <= A(1000) and not w13616;
w13618 <= not w13612 and w13617;
w13619 <= w9044 and w13611;
w13620 <= w9033 and not w9038;
w13621 <= not w9026 and w13620;
w13622 <= not w9033 and not w9042;
w13623 <= not w13621 and not w13622;
w13624 <= w3469 and not w13623;
w13625 <= not w9040 and not w9043;
w13626 <= not w3469 and not w13625;
w13627 <= not w13624 and not w13626;
w13628 <= not w13619 and not w13627;
w13629 <= w13618 and w13628;
w13630 <= not w13607 and w13629;
w13631 <= not w13606 and w13630;
w13632 <= not w13601 and w13631;
w13633 <= not w13600 and w13632;
w13634 <= not w13595 and w13633;
w13635 <= not w13594 and w13634;
w13636 <= not w13589 and w13635;
w13637 <= not w13588 and w13636;
w13638 <= not w13583 and w13637;
w13639 <= not w13582 and w13638;
w13640 <= not w13577 and w13639;
w13641 <= not w13575 and w13640;
w13642 <= w13569 and w13641;
w13643 <= not w13569 and not w13641;
w13644 <= not w13642 and not w13643;
w13645 <= not w13575 and not w13577;
w13646 <= not w13639 and not w13645;
w13647 <= not w13582 and not w13583;
w13648 <= not w13637 and not w13647;
w13649 <= not w13588 and not w13589;
w13650 <= not w13635 and not w13649;
w13651 <= not w13606 and not w13607;
w13652 <= not w13629 and not w13651;
w13653 <= not w13612 and not w13619;
w13654 <= w13617 and not w13627;
w13655 <= not w13653 and not w13654;
w13656 <= not w13629 and not w13655;
w13657 <= w13617 and not w13624;
w13658 <= not w13626 and w13657;
w13659 <= not w13617 and not w13627;
w13660 <= not w13658 and not w13659;
w13661 <= not w13656 and w13660;
w13662 <= not w13631 and not w13661;
w13663 <= not w13652 and w13662;
w13664 <= not w13600 and not w13601;
w13665 <= not w13631 and not w13664;
w13666 <= not w13633 and not w13665;
w13667 <= not w13663 and not w13666;
w13668 <= not w13594 and not w13595;
w13669 <= not w13633 and not w13668;
w13670 <= not w13635 and not w13669;
w13671 <= not w13667 and w13670;
w13672 <= not w13637 and w13671;
w13673 <= not w13650 and w13672;
w13674 <= not w13639 and w13673;
w13675 <= not w13648 and w13674;
w13676 <= not w13641 and w13675;
w13677 <= not w13646 and w13676;
w13678 <= not w13644 and w13677;
w13679 <= not w13569 and w13641;
w13680 <= not w13563 and not w13565;
w13681 <= not w13679 and w13680;
w13682 <= w13641 and not w13680;
w13683 <= not w13569 and w13682;
w13684 <= not w13565 and w13637;
w13685 <= w13647 and w13684;
w13686 <= not w13577 and w13685;
w13687 <= not w13575 and w13686;
w13688 <= not w13563 and w13687;
w13689 <= not w13569 and w13688;
w13690 <= not w13683 and not w13689;
w13691 <= not w13681 and w13690;
w13692 <= not w13678 and w13691;
w13693 <= not w13639 and not w13648;
w13694 <= not w13631 and not w13652;
w13695 <= w13661 and not w13694;
w13696 <= not w13663 and not w13695;
w13697 <= w13656 and not w13660;
w13698 <= A(1000) and not w13614;
w13699 <= not w13615 and w13698;
w13700 <= not A(1000) and not w13616;
w13701 <= not w13699 and not w13700;
w13702 <= not w13661 and w13701;
w13703 <= not w13697 and w13702;
w13704 <= w13656 and not w13703;
w13705 <= not w13661 and not w13697;
w13706 <= not w13701 and not w13705;
w13707 <= not w13704 and not w13706;
w13708 <= not w13696 and w13707;
w13709 <= w13694 and not w13708;
w13710 <= w13696 and not w13707;
w13711 <= not w13709 and not w13710;
w13712 <= not w13663 and not w13711;
w13713 <= not w13633 and w13663;
w13714 <= not w13665 and w13713;
w13715 <= w13667 and not w13670;
w13716 <= not w13671 and not w13715;
w13717 <= not w13714 and not w13716;
w13718 <= not w13712 and w13717;
w13719 <= w13670 and not w13718;
w13720 <= not w13712 and not w13714;
w13721 <= w13716 and not w13720;
w13722 <= not w13719 and not w13721;
w13723 <= w13671 and not w13722;
w13724 <= not w13637 and not w13650;
w13725 <= not w13671 and w13724;
w13726 <= not w13673 and not w13693;
w13727 <= not w13675 and not w13726;
w13728 <= not w13725 and not w13727;
w13729 <= not w13723 and w13728;
w13730 <= w13693 and not w13729;
w13731 <= not w13723 and not w13725;
w13732 <= w13727 and not w13731;
w13733 <= not w13730 and not w13732;
w13734 <= w13675 and not w13677;
w13735 <= not w13733 and w13734;
w13736 <= w13677 and not w13730;
w13737 <= not w13732 and w13736;
w13738 <= not w13641 and not w13646;
w13739 <= not w13737 and w13738;
w13740 <= not w13735 and not w13739;
w13741 <= w13677 and not w13678;
w13742 <= not w13740 and w13741;
w13743 <= w13678 and not w13735;
w13744 <= not w13739 and w13743;
w13745 <= not w13644 and not w13744;
w13746 <= not w13678 and not w13745;
w13747 <= not w13742 and w13746;
w13748 <= w13677 and not w13683;
w13749 <= not w13681 and w13748;
w13750 <= not w13644 and w13749;
w13751 <= not w13681 and not w13683;
w13752 <= not w13678 and w13751;
w13753 <= w13689 and not w13752;
w13754 <= not w13692 and not w13753;
w13755 <= not w13750 and not w13754;
w13756 <= not w13747 and w13755;
w13757 <= w13692 and not w13756;
one <= '1';
maj <= not w13757;-- level 70
end Behavioral;
