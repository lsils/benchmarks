library ieee;
use ieee.std_logic_1164.all;

entity top is
 port(pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203: in std_logic;
po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230: out std_logic);
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200, w19201, w19202, w19203, w19204, w19205, w19206, w19207, w19208, w19209, w19210, w19211, w19212, w19213, w19214, w19215, w19216, w19217, w19218, w19219, w19220, w19221, w19222, w19223, w19224, w19225, w19226, w19227, w19228, w19229, w19230, w19231, w19232, w19233, w19234, w19235, w19236, w19237, w19238, w19239, w19240, w19241, w19242, w19243, w19244, w19245, w19246, w19247, w19248, w19249, w19250, w19251, w19252, w19253, w19254, w19255, w19256, w19257, w19258, w19259, w19260, w19261, w19262, w19263, w19264, w19265, w19266, w19267, w19268, w19269, w19270, w19271, w19272, w19273, w19274, w19275, w19276, w19277, w19278, w19279, w19280, w19281, w19282, w19283, w19284, w19285, w19286, w19287, w19288, w19289, w19290, w19291, w19292, w19293, w19294, w19295, w19296, w19297, w19298, w19299, w19300, w19301, w19302, w19303, w19304, w19305, w19306, w19307, w19308, w19309, w19310, w19311, w19312, w19313, w19314, w19315, w19316, w19317, w19318, w19319, w19320, w19321, w19322, w19323, w19324, w19325, w19326, w19327, w19328, w19329, w19330, w19331, w19332, w19333, w19334, w19335, w19336, w19337, w19338, w19339, w19340, w19341, w19342, w19343, w19344, w19345, w19346, w19347, w19348, w19349, w19350, w19351, w19352, w19353, w19354, w19355, w19356, w19357, w19358, w19359, w19360, w19361, w19362, w19363, w19364, w19365, w19366, w19367, w19368, w19369, w19370, w19371, w19372, w19373, w19374, w19375, w19376, w19377, w19378, w19379, w19380, w19381, w19382, w19383, w19384, w19385, w19386, w19387, w19388, w19389, w19390, w19391, w19392, w19393, w19394, w19395, w19396, w19397, w19398, w19399, w19400, w19401, w19402, w19403, w19404, w19405, w19406, w19407, w19408, w19409, w19410, w19411, w19412, w19413, w19414, w19415, w19416, w19417, w19418, w19419, w19420, w19421, w19422, w19423, w19424, w19425, w19426, w19427, w19428, w19429, w19430, w19431, w19432, w19433, w19434, w19435, w19436, w19437, w19438, w19439, w19440, w19441, w19442, w19443, w19444, w19445, w19446, w19447, w19448, w19449, w19450, w19451, w19452, w19453, w19454, w19455, w19456, w19457, w19458, w19459, w19460, w19461, w19462, w19463, w19464, w19465, w19466, w19467, w19468, w19469, w19470, w19471, w19472, w19473, w19474, w19475, w19476, w19477, w19478, w19479, w19480, w19481, w19482, w19483, w19484, w19485, w19486, w19487, w19488, w19489, w19490, w19491, w19492, w19493, w19494, w19495, w19496, w19497, w19498, w19499, w19500, w19501, w19502, w19503, w19504, w19505, w19506, w19507, w19508, w19509, w19510, w19511, w19512, w19513, w19514, w19515, w19516, w19517, w19518, w19519, w19520, w19521, w19522, w19523, w19524, w19525, w19526, w19527, w19528, w19529, w19530, w19531, w19532, w19533, w19534, w19535, w19536, w19537, w19538, w19539, w19540, w19541, w19542, w19543, w19544, w19545, w19546, w19547, w19548, w19549, w19550, w19551, w19552, w19553, w19554, w19555, w19556, w19557, w19558, w19559, w19560, w19561, w19562, w19563, w19564, w19565, w19566, w19567, w19568, w19569, w19570, w19571, w19572, w19573, w19574, w19575, w19576, w19577, w19578, w19579, w19580, w19581, w19582, w19583, w19584, w19585, w19586, w19587, w19588, w19589, w19590, w19591, w19592, w19593, w19594, w19595, w19596, w19597, w19598, w19599, w19600, w19601, w19602, w19603, w19604, w19605, w19606, w19607, w19608, w19609, w19610, w19611, w19612, w19613, w19614, w19615, w19616, w19617, w19618, w19619, w19620, w19621, w19622, w19623, w19624, w19625, w19626, w19627, w19628, w19629, w19630, w19631, w19632, w19633, w19634, w19635, w19636, w19637, w19638, w19639, w19640, w19641, w19642, w19643, w19644, w19645, w19646, w19647, w19648, w19649, w19650, w19651, w19652, w19653, w19654, w19655, w19656, w19657, w19658, w19659, w19660, w19661, w19662, w19663, w19664, w19665, w19666, w19667, w19668, w19669, w19670, w19671, w19672, w19673, w19674, w19675, w19676, w19677, w19678, w19679, w19680, w19681, w19682, w19683, w19684, w19685, w19686, w19687, w19688, w19689, w19690, w19691, w19692, w19693, w19694, w19695, w19696, w19697, w19698, w19699, w19700, w19701, w19702, w19703, w19704, w19705, w19706, w19707, w19708, w19709, w19710, w19711, w19712, w19713, w19714, w19715, w19716, w19717, w19718, w19719, w19720, w19721, w19722, w19723, w19724, w19725, w19726, w19727, w19728, w19729, w19730, w19731, w19732, w19733, w19734, w19735, w19736, w19737, w19738, w19739, w19740, w19741, w19742, w19743, w19744, w19745, w19746, w19747, w19748, w19749, w19750, w19751, w19752, w19753, w19754, w19755, w19756, w19757, w19758, w19759, w19760, w19761, w19762, w19763, w19764, w19765, w19766, w19767, w19768, w19769, w19770, w19771, w19772, w19773, w19774, w19775, w19776, w19777, w19778, w19779, w19780, w19781, w19782, w19783, w19784, w19785, w19786, w19787, w19788, w19789, w19790, w19791, w19792, w19793, w19794, w19795, w19796, w19797, w19798, w19799, w19800, w19801, w19802, w19803, w19804, w19805, w19806, w19807, w19808, w19809, w19810, w19811, w19812, w19813, w19814, w19815, w19816, w19817, w19818, w19819, w19820, w19821, w19822, w19823, w19824, w19825, w19826, w19827, w19828, w19829, w19830, w19831, w19832, w19833, w19834, w19835, w19836, w19837, w19838, w19839, w19840, w19841, w19842, w19843, w19844, w19845, w19846, w19847, w19848, w19849, w19850, w19851, w19852, w19853, w19854, w19855, w19856, w19857, w19858, w19859, w19860, w19861, w19862, w19863, w19864, w19865, w19866, w19867, w19868, w19869, w19870, w19871, w19872, w19873, w19874, w19875, w19876, w19877, w19878, w19879, w19880, w19881, w19882, w19883, w19884, w19885, w19886, w19887, w19888, w19889, w19890, w19891, w19892, w19893, w19894, w19895, w19896, w19897, w19898, w19899, w19900, w19901, w19902, w19903, w19904, w19905, w19906, w19907, w19908, w19909, w19910, w19911, w19912, w19913, w19914, w19915, w19916, w19917, w19918, w19919, w19920, w19921, w19922, w19923, w19924, w19925, w19926, w19927, w19928, w19929, w19930, w19931, w19932, w19933, w19934, w19935, w19936, w19937, w19938, w19939, w19940, w19941, w19942, w19943, w19944, w19945, w19946, w19947, w19948, w19949, w19950, w19951, w19952, w19953, w19954, w19955, w19956, w19957, w19958, w19959, w19960, w19961, w19962, w19963, w19964, w19965, w19966, w19967, w19968, w19969, w19970, w19971, w19972, w19973, w19974, w19975, w19976, w19977, w19978, w19979, w19980, w19981, w19982, w19983, w19984, w19985, w19986, w19987, w19988, w19989, w19990, w19991, w19992, w19993, w19994, w19995, w19996, w19997, w19998, w19999, w20000, w20001, w20002, w20003, w20004, w20005, w20006, w20007, w20008, w20009, w20010, w20011, w20012, w20013, w20014, w20015, w20016, w20017, w20018, w20019, w20020, w20021, w20022, w20023, w20024, w20025, w20026, w20027, w20028, w20029, w20030, w20031, w20032, w20033, w20034, w20035, w20036, w20037, w20038, w20039, w20040, w20041, w20042, w20043, w20044, w20045, w20046, w20047, w20048, w20049, w20050, w20051, w20052, w20053, w20054, w20055, w20056, w20057, w20058, w20059, w20060, w20061, w20062, w20063, w20064, w20065, w20066, w20067, w20068, w20069, w20070, w20071, w20072, w20073, w20074, w20075, w20076, w20077, w20078, w20079, w20080, w20081, w20082, w20083, w20084, w20085, w20086, w20087, w20088, w20089, w20090, w20091, w20092, w20093, w20094, w20095, w20096, w20097, w20098, w20099, w20100, w20101, w20102, w20103, w20104, w20105, w20106, w20107, w20108, w20109, w20110, w20111, w20112, w20113, w20114, w20115, w20116, w20117, w20118, w20119, w20120, w20121, w20122, w20123, w20124, w20125, w20126, w20127, w20128, w20129, w20130, w20131, w20132, w20133, w20134, w20135, w20136, w20137, w20138, w20139, w20140, w20141, w20142, w20143, w20144, w20145, w20146, w20147, w20148, w20149, w20150, w20151, w20152, w20153, w20154, w20155, w20156, w20157, w20158, w20159, w20160, w20161, w20162, w20163, w20164, w20165, w20166, w20167, w20168, w20169, w20170, w20171, w20172, w20173, w20174, w20175, w20176, w20177, w20178, w20179, w20180, w20181, w20182, w20183, w20184, w20185, w20186, w20187, w20188, w20189, w20190, w20191, w20192, w20193, w20194, w20195, w20196, w20197, w20198, w20199, w20200, w20201, w20202, w20203, w20204, w20205, w20206, w20207, w20208, w20209, w20210, w20211, w20212, w20213, w20214, w20215, w20216, w20217, w20218, w20219, w20220, w20221, w20222, w20223, w20224, w20225, w20226, w20227, w20228, w20229, w20230, w20231, w20232, w20233, w20234, w20235, w20236, w20237, w20238, w20239, w20240, w20241, w20242, w20243, w20244, w20245, w20246, w20247, w20248, w20249, w20250, w20251, w20252, w20253, w20254, w20255, w20256, w20257, w20258, w20259, w20260, w20261, w20262, w20263, w20264, w20265, w20266, w20267, w20268, w20269, w20270, w20271, w20272, w20273, w20274, w20275, w20276, w20277, w20278, w20279, w20280, w20281, w20282, w20283, w20284, w20285, w20286, w20287, w20288, w20289, w20290, w20291, w20292, w20293, w20294, w20295, w20296, w20297, w20298, w20299, w20300, w20301, w20302, w20303, w20304, w20305, w20306, w20307, w20308, w20309, w20310, w20311, w20312, w20313, w20314, w20315, w20316, w20317, w20318, w20319, w20320, w20321, w20322, w20323, w20324, w20325, w20326, w20327, w20328, w20329, w20330, w20331, w20332, w20333, w20334, w20335, w20336, w20337, w20338, w20339, w20340, w20341, w20342, w20343, w20344, w20345, w20346, w20347, w20348, w20349, w20350, w20351, w20352, w20353, w20354, w20355, w20356, w20357, w20358, w20359, w20360, w20361, w20362, w20363, w20364, w20365, w20366, w20367, w20368, w20369, w20370, w20371, w20372, w20373, w20374, w20375, w20376, w20377, w20378, w20379, w20380, w20381, w20382, w20383, w20384, w20385, w20386, w20387, w20388, w20389, w20390, w20391, w20392, w20393, w20394, w20395, w20396, w20397, w20398, w20399, w20400, w20401, w20402, w20403, w20404, w20405, w20406, w20407, w20408, w20409, w20410, w20411, w20412, w20413, w20414, w20415, w20416, w20417, w20418, w20419, w20420, w20421, w20422, w20423, w20424, w20425, w20426, w20427, w20428, w20429, w20430, w20431, w20432, w20433, w20434, w20435, w20436, w20437, w20438, w20439, w20440, w20441, w20442, w20443, w20444, w20445, w20446, w20447, w20448, w20449, w20450, w20451, w20452, w20453, w20454, w20455, w20456, w20457, w20458, w20459, w20460, w20461, w20462, w20463, w20464, w20465, w20466, w20467, w20468, w20469, w20470, w20471, w20472, w20473, w20474, w20475, w20476, w20477, w20478, w20479, w20480, w20481, w20482, w20483, w20484, w20485, w20486, w20487, w20488, w20489, w20490, w20491, w20492, w20493, w20494, w20495, w20496, w20497, w20498, w20499, w20500, w20501, w20502, w20503, w20504, w20505, w20506, w20507, w20508, w20509, w20510, w20511, w20512, w20513, w20514, w20515, w20516, w20517, w20518, w20519, w20520, w20521, w20522, w20523, w20524, w20525, w20526, w20527, w20528, w20529, w20530, w20531, w20532, w20533, w20534, w20535, w20536, w20537, w20538, w20539, w20540, w20541, w20542, w20543, w20544, w20545, w20546, w20547, w20548, w20549, w20550, w20551, w20552, w20553, w20554, w20555, w20556, w20557, w20558, w20559, w20560, w20561, w20562, w20563, w20564, w20565, w20566, w20567, w20568, w20569, w20570, w20571, w20572, w20573, w20574, w20575, w20576, w20577, w20578, w20579, w20580, w20581, w20582, w20583, w20584, w20585, w20586, w20587, w20588, w20589, w20590, w20591, w20592, w20593, w20594, w20595, w20596, w20597, w20598, w20599, w20600, w20601, w20602, w20603, w20604, w20605, w20606, w20607, w20608, w20609, w20610, w20611, w20612, w20613, w20614, w20615, w20616, w20617, w20618, w20619, w20620, w20621, w20622, w20623, w20624, w20625, w20626, w20627, w20628, w20629, w20630, w20631, w20632, w20633, w20634, w20635, w20636, w20637, w20638, w20639, w20640, w20641, w20642, w20643, w20644, w20645, w20646, w20647, w20648, w20649, w20650, w20651, w20652, w20653, w20654, w20655, w20656, w20657, w20658, w20659, w20660, w20661, w20662, w20663, w20664, w20665, w20666, w20667, w20668, w20669, w20670, w20671, w20672, w20673, w20674, w20675, w20676, w20677, w20678, w20679, w20680, w20681, w20682, w20683, w20684, w20685, w20686, w20687, w20688, w20689, w20690, w20691, w20692, w20693, w20694, w20695, w20696, w20697, w20698, w20699, w20700, w20701, w20702, w20703, w20704, w20705, w20706, w20707, w20708, w20709, w20710, w20711, w20712, w20713, w20714, w20715, w20716, w20717, w20718, w20719, w20720, w20721, w20722, w20723, w20724, w20725, w20726, w20727, w20728, w20729, w20730, w20731, w20732, w20733, w20734, w20735, w20736, w20737, w20738, w20739, w20740, w20741, w20742, w20743, w20744, w20745, w20746, w20747, w20748, w20749, w20750, w20751, w20752, w20753, w20754, w20755, w20756, w20757, w20758, w20759, w20760, w20761, w20762, w20763, w20764, w20765, w20766, w20767, w20768, w20769, w20770, w20771, w20772, w20773, w20774, w20775, w20776, w20777, w20778, w20779, w20780, w20781, w20782, w20783, w20784, w20785, w20786, w20787, w20788, w20789, w20790, w20791, w20792, w20793, w20794, w20795, w20796, w20797, w20798, w20799, w20800, w20801, w20802, w20803, w20804, w20805, w20806, w20807, w20808, w20809, w20810, w20811, w20812, w20813, w20814, w20815, w20816, w20817, w20818, w20819, w20820, w20821, w20822, w20823, w20824, w20825, w20826, w20827, w20828, w20829, w20830, w20831, w20832, w20833, w20834, w20835, w20836, w20837, w20838, w20839, w20840, w20841, w20842, w20843, w20844, w20845, w20846, w20847, w20848, w20849, w20850, w20851, w20852, w20853, w20854, w20855, w20856, w20857, w20858, w20859, w20860, w20861, w20862, w20863, w20864, w20865, w20866, w20867, w20868, w20869, w20870, w20871, w20872, w20873, w20874, w20875, w20876, w20877, w20878, w20879, w20880, w20881, w20882, w20883, w20884, w20885, w20886, w20887, w20888, w20889, w20890, w20891, w20892, w20893, w20894, w20895, w20896, w20897, w20898, w20899, w20900, w20901, w20902, w20903, w20904, w20905, w20906, w20907, w20908, w20909, w20910, w20911, w20912, w20913, w20914, w20915, w20916, w20917, w20918, w20919, w20920, w20921, w20922, w20923, w20924, w20925, w20926, w20927, w20928, w20929, w20930, w20931, w20932, w20933, w20934, w20935, w20936, w20937, w20938, w20939, w20940, w20941, w20942, w20943, w20944, w20945, w20946, w20947, w20948, w20949, w20950, w20951, w20952, w20953, w20954, w20955, w20956, w20957, w20958, w20959, w20960, w20961, w20962, w20963, w20964, w20965, w20966, w20967, w20968, w20969, w20970, w20971, w20972, w20973, w20974, w20975, w20976, w20977, w20978, w20979, w20980, w20981, w20982, w20983, w20984, w20985, w20986, w20987, w20988, w20989, w20990, w20991, w20992, w20993, w20994, w20995, w20996, w20997, w20998, w20999, w21000, w21001, w21002, w21003, w21004, w21005, w21006, w21007, w21008, w21009, w21010, w21011, w21012, w21013, w21014, w21015, w21016, w21017, w21018, w21019, w21020, w21021, w21022, w21023, w21024, w21025, w21026, w21027, w21028, w21029, w21030, w21031, w21032, w21033, w21034, w21035, w21036, w21037, w21038, w21039, w21040, w21041, w21042, w21043, w21044, w21045, w21046, w21047, w21048, w21049, w21050, w21051, w21052, w21053, w21054, w21055, w21056, w21057, w21058, w21059, w21060, w21061, w21062, w21063, w21064, w21065, w21066, w21067, w21068, w21069, w21070, w21071, w21072, w21073, w21074, w21075, w21076, w21077, w21078, w21079, w21080, w21081, w21082, w21083, w21084, w21085, w21086, w21087, w21088, w21089, w21090, w21091, w21092, w21093, w21094, w21095, w21096, w21097, w21098, w21099, w21100, w21101, w21102, w21103, w21104, w21105, w21106, w21107, w21108, w21109, w21110, w21111, w21112, w21113, w21114, w21115, w21116, w21117, w21118, w21119, w21120, w21121, w21122, w21123, w21124, w21125, w21126, w21127, w21128, w21129, w21130, w21131, w21132, w21133, w21134, w21135, w21136, w21137, w21138, w21139, w21140, w21141, w21142, w21143, w21144, w21145, w21146, w21147, w21148, w21149, w21150, w21151, w21152, w21153, w21154, w21155, w21156, w21157, w21158, w21159, w21160, w21161, w21162, w21163, w21164, w21165, w21166, w21167, w21168, w21169, w21170, w21171, w21172, w21173, w21174, w21175, w21176, w21177, w21178, w21179, w21180, w21181, w21182, w21183, w21184, w21185, w21186, w21187, w21188, w21189, w21190, w21191, w21192, w21193, w21194, w21195, w21196, w21197, w21198, w21199, w21200, w21201, w21202, w21203, w21204, w21205, w21206, w21207, w21208, w21209, w21210, w21211, w21212, w21213, w21214, w21215, w21216, w21217, w21218, w21219, w21220, w21221, w21222, w21223, w21224, w21225, w21226, w21227, w21228, w21229, w21230, w21231, w21232, w21233, w21234, w21235, w21236, w21237, w21238, w21239, w21240, w21241, w21242, w21243, w21244, w21245, w21246, w21247, w21248, w21249, w21250, w21251, w21252, w21253, w21254, w21255, w21256, w21257, w21258, w21259, w21260, w21261, w21262, w21263, w21264, w21265, w21266, w21267, w21268, w21269, w21270, w21271, w21272, w21273, w21274, w21275, w21276, w21277, w21278, w21279, w21280, w21281, w21282, w21283, w21284, w21285, w21286, w21287, w21288, w21289, w21290, w21291, w21292, w21293, w21294, w21295, w21296, w21297, w21298, w21299, w21300, w21301, w21302, w21303, w21304, w21305, w21306, w21307, w21308, w21309, w21310, w21311, w21312, w21313, w21314, w21315, w21316, w21317, w21318, w21319, w21320, w21321, w21322, w21323, w21324, w21325, w21326, w21327, w21328, w21329, w21330, w21331, w21332, w21333, w21334, w21335, w21336, w21337, w21338, w21339, w21340, w21341, w21342, w21343, w21344, w21345, w21346, w21347, w21348, w21349, w21350, w21351, w21352, w21353, w21354, w21355, w21356, w21357, w21358, w21359, w21360, w21361, w21362, w21363, w21364, w21365, w21366, w21367, w21368, w21369, w21370, w21371, w21372, w21373, w21374, w21375, w21376, w21377, w21378, w21379, w21380, w21381, w21382, w21383, w21384, w21385, w21386, w21387, w21388, w21389, w21390, w21391, w21392, w21393, w21394, w21395, w21396, w21397, w21398, w21399, w21400, w21401, w21402, w21403, w21404, w21405, w21406, w21407, w21408, w21409, w21410, w21411, w21412, w21413, w21414, w21415, w21416, w21417, w21418, w21419, w21420, w21421, w21422, w21423, w21424, w21425, w21426, w21427, w21428, w21429, w21430, w21431, w21432, w21433, w21434, w21435, w21436, w21437, w21438, w21439, w21440, w21441, w21442, w21443, w21444, w21445, w21446, w21447, w21448, w21449, w21450, w21451, w21452, w21453, w21454, w21455, w21456, w21457, w21458, w21459, w21460, w21461, w21462, w21463, w21464, w21465, w21466, w21467, w21468, w21469, w21470, w21471, w21472, w21473, w21474, w21475, w21476, w21477, w21478, w21479, w21480, w21481, w21482, w21483, w21484, w21485, w21486, w21487, w21488, w21489, w21490, w21491, w21492, w21493, w21494, w21495, w21496, w21497, w21498, w21499, w21500, w21501, w21502, w21503, w21504, w21505, w21506, w21507, w21508, w21509, w21510, w21511, w21512, w21513, w21514, w21515, w21516, w21517, w21518, w21519, w21520, w21521, w21522, w21523, w21524, w21525, w21526, w21527, w21528, w21529, w21530, w21531, w21532, w21533, w21534, w21535, w21536, w21537, w21538, w21539, w21540, w21541, w21542, w21543, w21544, w21545, w21546, w21547, w21548, w21549, w21550, w21551, w21552, w21553, w21554, w21555, w21556, w21557, w21558, w21559, w21560, w21561, w21562, w21563, w21564, w21565, w21566, w21567, w21568, w21569, w21570, w21571, w21572, w21573, w21574, w21575, w21576, w21577, w21578, w21579, w21580, w21581, w21582, w21583, w21584, w21585, w21586, w21587, w21588, w21589, w21590, w21591, w21592, w21593, w21594, w21595, w21596, w21597, w21598, w21599, w21600, w21601, w21602, w21603, w21604, w21605, w21606, w21607, w21608, w21609, w21610, w21611, w21612, w21613, w21614, w21615, w21616, w21617, w21618, w21619, w21620, w21621, w21622, w21623, w21624, w21625, w21626, w21627, w21628, w21629, w21630, w21631, w21632, w21633, w21634, w21635, w21636, w21637, w21638, w21639, w21640, w21641, w21642, w21643, w21644, w21645, w21646, w21647, w21648, w21649, w21650, w21651, w21652, w21653, w21654, w21655, w21656, w21657, w21658, w21659, w21660, w21661, w21662, w21663, w21664, w21665, w21666, w21667, w21668, w21669, w21670, w21671, w21672, w21673, w21674, w21675, w21676, w21677, w21678, w21679, w21680, w21681, w21682, w21683, w21684, w21685, w21686, w21687, w21688, w21689, w21690, w21691, w21692, w21693, w21694, w21695, w21696, w21697, w21698, w21699, w21700, w21701, w21702, w21703, w21704, w21705, w21706, w21707, w21708, w21709, w21710, w21711, w21712, w21713, w21714, w21715, w21716, w21717, w21718, w21719, w21720, w21721, w21722, w21723, w21724, w21725, w21726, w21727, w21728, w21729, w21730, w21731, w21732, w21733, w21734, w21735, w21736, w21737, w21738, w21739, w21740, w21741, w21742, w21743, w21744, w21745, w21746, w21747, w21748, w21749, w21750, w21751, w21752, w21753, w21754, w21755, w21756, w21757, w21758, w21759, w21760, w21761, w21762, w21763, w21764, w21765, w21766, w21767, w21768, w21769, w21770, w21771, w21772, w21773, w21774, w21775, w21776, w21777, w21778, w21779, w21780, w21781, w21782, w21783, w21784, w21785, w21786, w21787, w21788, w21789, w21790, w21791, w21792, w21793, w21794, w21795, w21796, w21797, w21798, w21799, w21800, w21801, w21802, w21803, w21804, w21805, w21806, w21807, w21808, w21809, w21810, w21811, w21812, w21813, w21814, w21815, w21816, w21817, w21818, w21819, w21820, w21821, w21822, w21823, w21824, w21825, w21826, w21827, w21828, w21829, w21830, w21831, w21832, w21833, w21834, w21835, w21836, w21837, w21838, w21839, w21840, w21841, w21842, w21843, w21844, w21845, w21846, w21847, w21848, w21849, w21850, w21851, w21852, w21853, w21854, w21855, w21856, w21857, w21858, w21859, w21860, w21861, w21862, w21863, w21864, w21865, w21866, w21867, w21868, w21869, w21870, w21871, w21872, w21873, w21874, w21875, w21876, w21877, w21878, w21879, w21880, w21881, w21882, w21883, w21884, w21885, w21886, w21887, w21888, w21889, w21890, w21891, w21892, w21893, w21894, w21895, w21896, w21897, w21898, w21899, w21900, w21901, w21902, w21903, w21904, w21905, w21906, w21907, w21908, w21909, w21910, w21911, w21912, w21913, w21914, w21915, w21916, w21917, w21918, w21919, w21920, w21921, w21922, w21923, w21924, w21925, w21926, w21927, w21928, w21929, w21930, w21931, w21932, w21933, w21934, w21935, w21936, w21937, w21938, w21939, w21940, w21941, w21942, w21943, w21944, w21945, w21946, w21947, w21948, w21949, w21950, w21951, w21952, w21953, w21954, w21955, w21956, w21957, w21958, w21959, w21960, w21961, w21962, w21963, w21964, w21965, w21966, w21967, w21968, w21969, w21970, w21971, w21972, w21973, w21974, w21975, w21976, w21977, w21978, w21979, w21980, w21981, w21982, w21983, w21984, w21985, w21986, w21987, w21988, w21989, w21990, w21991, w21992, w21993, w21994, w21995, w21996, w21997, w21998, w21999, w22000, w22001, w22002, w22003, w22004, w22005, w22006, w22007, w22008, w22009, w22010, w22011, w22012, w22013, w22014, w22015, w22016, w22017, w22018, w22019, w22020, w22021, w22022, w22023, w22024, w22025, w22026, w22027, w22028, w22029, w22030, w22031, w22032, w22033, w22034, w22035, w22036, w22037, w22038, w22039, w22040, w22041, w22042, w22043, w22044, w22045, w22046, w22047, w22048, w22049, w22050, w22051, w22052, w22053, w22054, w22055, w22056, w22057, w22058, w22059, w22060, w22061, w22062, w22063, w22064, w22065, w22066, w22067, w22068, w22069, w22070, w22071, w22072, w22073, w22074, w22075, w22076, w22077, w22078, w22079, w22080, w22081, w22082, w22083, w22084, w22085, w22086, w22087, w22088, w22089, w22090, w22091, w22092, w22093, w22094, w22095, w22096, w22097, w22098, w22099, w22100, w22101, w22102, w22103, w22104, w22105, w22106, w22107, w22108, w22109, w22110, w22111, w22112, w22113, w22114, w22115, w22116, w22117, w22118, w22119, w22120, w22121, w22122, w22123, w22124, w22125, w22126, w22127, w22128, w22129, w22130, w22131, w22132, w22133, w22134, w22135, w22136, w22137, w22138, w22139, w22140, w22141, w22142, w22143, w22144, w22145, w22146, w22147, w22148, w22149, w22150, w22151, w22152, w22153, w22154, w22155, w22156, w22157, w22158, w22159, w22160, w22161, w22162, w22163, w22164, w22165, w22166, w22167, w22168, w22169, w22170, w22171, w22172, w22173, w22174, w22175, w22176, w22177, w22178, w22179, w22180, w22181, w22182, w22183, w22184, w22185, w22186, w22187, w22188, w22189, w22190, w22191, w22192, w22193, w22194, w22195, w22196, w22197, w22198, w22199, w22200, w22201, w22202, w22203, w22204, w22205, w22206, w22207, w22208, w22209, w22210, w22211, w22212, w22213, w22214, w22215, w22216, w22217, w22218, w22219, w22220, w22221, w22222, w22223, w22224, w22225, w22226, w22227, w22228, w22229, w22230, w22231, w22232, w22233, w22234, w22235, w22236, w22237, w22238, w22239, w22240, w22241, w22242, w22243, w22244, w22245, w22246, w22247, w22248, w22249, w22250, w22251, w22252, w22253, w22254, w22255, w22256, w22257, w22258, w22259, w22260, w22261, w22262, w22263, w22264, w22265, w22266, w22267, w22268, w22269, w22270, w22271, w22272, w22273, w22274, w22275, w22276, w22277, w22278, w22279, w22280, w22281, w22282, w22283, w22284, w22285, w22286, w22287, w22288, w22289, w22290, w22291, w22292, w22293, w22294, w22295, w22296, w22297, w22298, w22299, w22300, w22301, w22302, w22303, w22304, w22305, w22306, w22307, w22308, w22309, w22310, w22311, w22312, w22313, w22314, w22315, w22316, w22317, w22318, w22319, w22320, w22321, w22322, w22323, w22324, w22325, w22326, w22327, w22328, w22329, w22330, w22331, w22332, w22333, w22334, w22335, w22336, w22337, w22338, w22339, w22340, w22341, w22342, w22343, w22344, w22345, w22346, w22347, w22348, w22349, w22350, w22351, w22352, w22353, w22354, w22355, w22356, w22357, w22358, w22359, w22360, w22361, w22362, w22363, w22364, w22365, w22366, w22367, w22368, w22369, w22370, w22371, w22372, w22373, w22374, w22375, w22376, w22377, w22378, w22379, w22380, w22381, w22382, w22383, w22384, w22385, w22386, w22387, w22388, w22389, w22390, w22391, w22392, w22393, w22394, w22395, w22396, w22397, w22398, w22399, w22400, w22401, w22402, w22403, w22404, w22405, w22406, w22407, w22408, w22409, w22410, w22411, w22412, w22413, w22414, w22415, w22416, w22417, w22418, w22419, w22420, w22421, w22422, w22423, w22424, w22425, w22426, w22427, w22428, w22429, w22430, w22431, w22432, w22433, w22434, w22435, w22436, w22437, w22438, w22439, w22440, w22441, w22442, w22443, w22444, w22445, w22446, w22447, w22448, w22449, w22450, w22451, w22452, w22453, w22454, w22455, w22456, w22457, w22458, w22459, w22460, w22461, w22462, w22463, w22464, w22465, w22466, w22467, w22468, w22469, w22470, w22471, w22472, w22473, w22474, w22475, w22476, w22477, w22478, w22479, w22480, w22481, w22482, w22483, w22484, w22485, w22486, w22487, w22488, w22489, w22490, w22491, w22492, w22493, w22494, w22495, w22496, w22497, w22498, w22499, w22500, w22501, w22502, w22503, w22504, w22505, w22506, w22507, w22508, w22509, w22510, w22511, w22512, w22513, w22514, w22515, w22516, w22517, w22518, w22519, w22520, w22521, w22522, w22523, w22524, w22525, w22526, w22527, w22528, w22529, w22530, w22531, w22532, w22533, w22534, w22535, w22536, w22537, w22538, w22539, w22540, w22541, w22542, w22543, w22544, w22545, w22546, w22547, w22548, w22549, w22550, w22551, w22552, w22553, w22554, w22555, w22556, w22557, w22558, w22559, w22560, w22561, w22562, w22563, w22564, w22565, w22566, w22567, w22568, w22569, w22570, w22571, w22572, w22573, w22574, w22575, w22576, w22577, w22578, w22579, w22580, w22581, w22582, w22583, w22584, w22585, w22586, w22587, w22588, w22589, w22590, w22591, w22592, w22593, w22594, w22595, w22596, w22597, w22598, w22599, w22600, w22601, w22602, w22603, w22604, w22605, w22606, w22607, w22608, w22609, w22610, w22611, w22612, w22613, w22614, w22615, w22616, w22617, w22618, w22619, w22620, w22621, w22622, w22623, w22624, w22625, w22626, w22627, w22628, w22629, w22630, w22631, w22632, w22633, w22634, w22635, w22636, w22637, w22638, w22639, w22640, w22641, w22642, w22643, w22644, w22645, w22646, w22647, w22648, w22649, w22650, w22651, w22652, w22653, w22654, w22655, w22656, w22657, w22658, w22659, w22660, w22661, w22662, w22663, w22664, w22665, w22666, w22667, w22668, w22669, w22670, w22671, w22672, w22673, w22674, w22675, w22676, w22677, w22678, w22679, w22680, w22681, w22682, w22683, w22684, w22685, w22686, w22687, w22688, w22689, w22690, w22691, w22692, w22693, w22694, w22695, w22696, w22697, w22698, w22699, w22700, w22701, w22702, w22703, w22704, w22705, w22706, w22707, w22708, w22709, w22710, w22711, w22712, w22713, w22714, w22715, w22716, w22717, w22718, w22719, w22720, w22721, w22722, w22723, w22724, w22725, w22726, w22727, w22728, w22729, w22730, w22731, w22732, w22733, w22734, w22735, w22736, w22737, w22738, w22739, w22740, w22741, w22742, w22743, w22744, w22745, w22746, w22747, w22748, w22749, w22750, w22751, w22752, w22753, w22754, w22755, w22756, w22757, w22758, w22759, w22760, w22761, w22762, w22763, w22764, w22765, w22766, w22767, w22768, w22769, w22770, w22771, w22772, w22773, w22774, w22775, w22776, w22777, w22778, w22779, w22780, w22781, w22782, w22783, w22784, w22785, w22786, w22787, w22788, w22789, w22790, w22791, w22792, w22793, w22794, w22795, w22796, w22797, w22798, w22799, w22800, w22801, w22802, w22803, w22804, w22805, w22806, w22807, w22808, w22809, w22810, w22811, w22812, w22813, w22814, w22815, w22816, w22817, w22818, w22819, w22820, w22821, w22822, w22823, w22824, w22825, w22826, w22827, w22828, w22829, w22830, w22831, w22832, w22833, w22834, w22835, w22836, w22837, w22838, w22839, w22840, w22841, w22842, w22843, w22844, w22845, w22846, w22847, w22848, w22849, w22850, w22851, w22852, w22853, w22854, w22855, w22856, w22857, w22858, w22859, w22860, w22861, w22862, w22863, w22864, w22865, w22866, w22867, w22868, w22869, w22870, w22871, w22872, w22873, w22874, w22875, w22876, w22877, w22878, w22879, w22880, w22881, w22882, w22883, w22884, w22885, w22886, w22887, w22888, w22889, w22890, w22891, w22892, w22893, w22894, w22895, w22896, w22897, w22898, w22899, w22900, w22901, w22902, w22903, w22904, w22905, w22906, w22907, w22908, w22909, w22910, w22911, w22912, w22913, w22914, w22915, w22916, w22917, w22918, w22919, w22920, w22921, w22922, w22923, w22924, w22925, w22926, w22927, w22928, w22929, w22930, w22931, w22932, w22933, w22934, w22935, w22936, w22937, w22938, w22939, w22940, w22941, w22942, w22943, w22944, w22945, w22946, w22947, w22948, w22949, w22950, w22951, w22952, w22953, w22954, w22955, w22956, w22957, w22958, w22959, w22960, w22961, w22962, w22963, w22964, w22965, w22966, w22967, w22968, w22969, w22970, w22971, w22972, w22973, w22974, w22975, w22976, w22977, w22978, w22979, w22980, w22981, w22982, w22983, w22984, w22985, w22986, w22987, w22988, w22989, w22990, w22991, w22992, w22993, w22994, w22995, w22996, w22997, w22998, w22999, w23000, w23001, w23002, w23003, w23004, w23005, w23006, w23007, w23008, w23009, w23010, w23011, w23012, w23013, w23014, w23015, w23016, w23017, w23018, w23019, w23020, w23021, w23022, w23023, w23024, w23025, w23026, w23027, w23028, w23029, w23030, w23031, w23032, w23033, w23034, w23035, w23036, w23037, w23038, w23039, w23040, w23041, w23042, w23043, w23044, w23045, w23046, w23047, w23048, w23049, w23050, w23051, w23052, w23053, w23054, w23055, w23056, w23057, w23058, w23059, w23060, w23061, w23062, w23063, w23064, w23065, w23066, w23067, w23068, w23069, w23070, w23071, w23072, w23073, w23074, w23075, w23076, w23077, w23078, w23079, w23080, w23081, w23082, w23083, w23084, w23085, w23086, w23087, w23088, w23089, w23090, w23091, w23092, w23093, w23094, w23095, w23096, w23097, w23098, w23099, w23100, w23101, w23102, w23103, w23104, w23105, w23106, w23107, w23108, w23109, w23110, w23111, w23112, w23113, w23114, w23115, w23116, w23117, w23118, w23119, w23120, w23121, w23122, w23123, w23124, w23125, w23126, w23127, w23128, w23129, w23130, w23131, w23132, w23133, w23134, w23135, w23136, w23137, w23138, w23139, w23140, w23141, w23142, w23143, w23144, w23145, w23146, w23147, w23148, w23149, w23150, w23151, w23152, w23153, w23154, w23155, w23156, w23157, w23158, w23159, w23160, w23161, w23162, w23163, w23164, w23165, w23166, w23167, w23168, w23169, w23170, w23171, w23172, w23173, w23174, w23175, w23176, w23177, w23178, w23179, w23180, w23181, w23182, w23183, w23184, w23185, w23186, w23187, w23188, w23189, w23190, w23191, w23192, w23193, w23194, w23195, w23196, w23197, w23198, w23199, w23200, w23201, w23202, w23203, w23204, w23205, w23206, w23207, w23208, w23209, w23210, w23211, w23212, w23213, w23214, w23215, w23216, w23217, w23218, w23219, w23220, w23221, w23222, w23223, w23224, w23225, w23226, w23227, w23228, w23229, w23230, w23231, w23232, w23233, w23234, w23235, w23236, w23237, w23238, w23239, w23240, w23241, w23242, w23243, w23244, w23245, w23246, w23247, w23248, w23249, w23250, w23251, w23252, w23253, w23254, w23255, w23256, w23257, w23258, w23259, w23260, w23261, w23262, w23263, w23264, w23265, w23266, w23267, w23268, w23269, w23270, w23271, w23272, w23273, w23274, w23275, w23276, w23277, w23278, w23279, w23280, w23281, w23282, w23283, w23284, w23285, w23286, w23287, w23288, w23289, w23290, w23291, w23292, w23293, w23294, w23295, w23296, w23297, w23298, w23299, w23300, w23301, w23302, w23303, w23304, w23305, w23306, w23307, w23308, w23309, w23310, w23311, w23312, w23313, w23314, w23315, w23316, w23317, w23318, w23319, w23320, w23321, w23322, w23323, w23324, w23325, w23326, w23327, w23328, w23329, w23330, w23331, w23332, w23333, w23334, w23335, w23336, w23337, w23338, w23339, w23340, w23341, w23342, w23343, w23344, w23345, w23346, w23347, w23348, w23349, w23350, w23351, w23352, w23353, w23354, w23355, w23356, w23357, w23358, w23359, w23360, w23361, w23362, w23363, w23364, w23365, w23366, w23367, w23368, w23369, w23370, w23371, w23372, w23373, w23374, w23375, w23376, w23377, w23378, w23379, w23380, w23381, w23382, w23383, w23384, w23385, w23386, w23387, w23388, w23389, w23390, w23391, w23392, w23393, w23394, w23395, w23396, w23397, w23398, w23399, w23400, w23401, w23402, w23403, w23404, w23405, w23406, w23407, w23408, w23409, w23410, w23411, w23412, w23413, w23414, w23415, w23416, w23417, w23418, w23419, w23420, w23421, w23422, w23423, w23424, w23425, w23426, w23427, w23428, w23429, w23430, w23431, w23432, w23433, w23434, w23435, w23436, w23437, w23438, w23439, w23440, w23441, w23442, w23443, w23444, w23445, w23446, w23447, w23448, w23449, w23450, w23451, w23452, w23453, w23454, w23455, w23456, w23457, w23458, w23459, w23460, w23461, w23462, w23463, w23464, w23465, w23466, w23467, w23468, w23469, w23470, w23471, w23472, w23473, w23474, w23475, w23476, w23477, w23478, w23479, w23480, w23481, w23482, w23483, w23484, w23485, w23486, w23487, w23488, w23489, w23490, w23491, w23492, w23493, w23494, w23495, w23496, w23497, w23498, w23499, w23500, w23501, w23502, w23503, w23504, w23505, w23506, w23507, w23508, w23509, w23510, w23511, w23512, w23513, w23514, w23515, w23516, w23517, w23518, w23519, w23520, w23521, w23522, w23523, w23524, w23525, w23526, w23527, w23528, w23529, w23530, w23531, w23532, w23533, w23534, w23535, w23536, w23537, w23538, w23539, w23540, w23541, w23542, w23543, w23544, w23545, w23546, w23547, w23548, w23549, w23550, w23551, w23552, w23553, w23554, w23555, w23556, w23557, w23558, w23559, w23560, w23561, w23562, w23563, w23564, w23565, w23566, w23567, w23568, w23569, w23570, w23571, w23572, w23573, w23574, w23575, w23576, w23577, w23578, w23579, w23580, w23581, w23582, w23583, w23584, w23585, w23586, w23587, w23588, w23589, w23590, w23591, w23592, w23593, w23594, w23595, w23596, w23597, w23598, w23599, w23600, w23601, w23602, w23603, w23604, w23605, w23606, w23607, w23608, w23609, w23610, w23611, w23612, w23613, w23614, w23615, w23616, w23617, w23618, w23619, w23620, w23621, w23622, w23623, w23624, w23625, w23626, w23627, w23628, w23629, w23630, w23631, w23632, w23633, w23634, w23635, w23636, w23637, w23638, w23639, w23640, w23641, w23642, w23643, w23644, w23645, w23646, w23647, w23648, w23649, w23650, w23651, w23652, w23653, w23654, w23655, w23656, w23657, w23658, w23659, w23660, w23661, w23662, w23663, w23664, w23665, w23666, w23667, w23668, w23669, w23670, w23671, w23672, w23673, w23674, w23675, w23676, w23677, w23678, w23679, w23680, w23681, w23682, w23683, w23684, w23685, w23686, w23687, w23688, w23689, w23690, w23691, w23692, w23693, w23694, w23695, w23696, w23697, w23698, w23699, w23700, w23701, w23702, w23703, w23704, w23705, w23706, w23707, w23708, w23709, w23710, w23711, w23712, w23713, w23714, w23715, w23716, w23717, w23718, w23719, w23720, w23721, w23722, w23723, w23724, w23725, w23726, w23727, w23728, w23729, w23730, w23731, w23732, w23733, w23734, w23735, w23736, w23737, w23738, w23739, w23740, w23741, w23742, w23743, w23744, w23745, w23746, w23747, w23748, w23749, w23750, w23751, w23752, w23753, w23754, w23755, w23756, w23757, w23758, w23759, w23760, w23761, w23762, w23763, w23764, w23765, w23766, w23767, w23768, w23769, w23770, w23771, w23772, w23773, w23774, w23775, w23776, w23777, w23778, w23779, w23780, w23781, w23782, w23783, w23784, w23785, w23786, w23787, w23788, w23789, w23790, w23791, w23792, w23793, w23794, w23795, w23796, w23797, w23798, w23799, w23800, w23801, w23802, w23803, w23804, w23805, w23806, w23807, w23808, w23809, w23810, w23811, w23812, w23813, w23814, w23815, w23816, w23817, w23818, w23819, w23820, w23821, w23822, w23823, w23824, w23825, w23826, w23827, w23828, w23829, w23830, w23831, w23832, w23833, w23834, w23835, w23836, w23837, w23838, w23839, w23840, w23841, w23842, w23843, w23844, w23845, w23846, w23847, w23848, w23849, w23850, w23851, w23852, w23853, w23854, w23855, w23856, w23857, w23858, w23859, w23860, w23861, w23862, w23863, w23864, w23865, w23866, w23867, w23868, w23869, w23870, w23871, w23872, w23873, w23874, w23875, w23876, w23877, w23878, w23879, w23880, w23881, w23882, w23883, w23884, w23885, w23886, w23887, w23888, w23889, w23890, w23891, w23892, w23893, w23894, w23895, w23896, w23897, w23898, w23899, w23900, w23901, w23902, w23903, w23904, w23905, w23906, w23907, w23908, w23909, w23910, w23911, w23912, w23913, w23914, w23915, w23916, w23917, w23918, w23919, w23920, w23921, w23922, w23923, w23924, w23925, w23926, w23927, w23928, w23929, w23930, w23931, w23932, w23933, w23934, w23935, w23936, w23937, w23938, w23939, w23940, w23941, w23942, w23943, w23944, w23945, w23946, w23947, w23948, w23949, w23950, w23951, w23952, w23953, w23954, w23955, w23956, w23957, w23958, w23959, w23960, w23961, w23962, w23963, w23964, w23965, w23966, w23967, w23968, w23969, w23970, w23971, w23972, w23973, w23974, w23975, w23976, w23977, w23978, w23979, w23980, w23981, w23982, w23983, w23984, w23985, w23986, w23987, w23988, w23989, w23990, w23991, w23992, w23993, w23994, w23995, w23996, w23997, w23998, w23999, w24000, w24001, w24002, w24003, w24004, w24005, w24006, w24007, w24008, w24009, w24010, w24011, w24012, w24013, w24014, w24015, w24016, w24017, w24018, w24019, w24020, w24021, w24022, w24023, w24024, w24025, w24026, w24027, w24028, w24029, w24030, w24031, w24032, w24033, w24034, w24035, w24036, w24037, w24038, w24039, w24040, w24041, w24042, w24043, w24044, w24045, w24046, w24047, w24048, w24049, w24050, w24051, w24052, w24053, w24054, w24055, w24056, w24057, w24058, w24059, w24060, w24061, w24062, w24063, w24064, w24065, w24066, w24067, w24068, w24069, w24070, w24071, w24072, w24073, w24074, w24075, w24076, w24077, w24078, w24079, w24080, w24081, w24082, w24083, w24084, w24085, w24086, w24087, w24088, w24089, w24090, w24091, w24092, w24093, w24094, w24095, w24096, w24097, w24098, w24099, w24100, w24101, w24102, w24103, w24104, w24105, w24106, w24107, w24108, w24109, w24110, w24111, w24112, w24113, w24114, w24115, w24116, w24117, w24118, w24119, w24120, w24121, w24122, w24123, w24124, w24125, w24126, w24127, w24128, w24129, w24130, w24131, w24132, w24133, w24134, w24135, w24136, w24137, w24138, w24139, w24140, w24141, w24142, w24143, w24144, w24145, w24146, w24147, w24148, w24149, w24150, w24151, w24152, w24153, w24154, w24155, w24156, w24157, w24158, w24159, w24160, w24161, w24162, w24163, w24164, w24165, w24166, w24167, w24168, w24169, w24170, w24171, w24172, w24173, w24174, w24175, w24176, w24177, w24178, w24179, w24180, w24181, w24182, w24183, w24184, w24185, w24186, w24187, w24188, w24189, w24190, w24191, w24192, w24193, w24194, w24195, w24196, w24197, w24198, w24199, w24200, w24201, w24202, w24203, w24204, w24205, w24206, w24207, w24208, w24209, w24210, w24211, w24212, w24213, w24214, w24215, w24216, w24217, w24218, w24219, w24220, w24221, w24222, w24223, w24224, w24225, w24226, w24227, w24228, w24229, w24230, w24231, w24232, w24233, w24234, w24235, w24236, w24237, w24238, w24239, w24240, w24241, w24242, w24243, w24244, w24245, w24246, w24247, w24248, w24249, w24250, w24251, w24252, w24253, w24254, w24255, w24256, w24257, w24258, w24259, w24260, w24261, w24262, w24263, w24264, w24265, w24266, w24267, w24268, w24269, w24270, w24271, w24272, w24273, w24274, w24275, w24276, w24277, w24278, w24279, w24280, w24281, w24282, w24283, w24284, w24285, w24286, w24287, w24288, w24289, w24290, w24291, w24292, w24293, w24294, w24295, w24296, w24297, w24298, w24299, w24300, w24301, w24302, w24303, w24304, w24305, w24306, w24307, w24308, w24309, w24310, w24311, w24312, w24313, w24314, w24315, w24316, w24317, w24318, w24319, w24320, w24321, w24322, w24323, w24324, w24325, w24326, w24327, w24328, w24329, w24330, w24331, w24332, w24333, w24334, w24335, w24336, w24337, w24338, w24339, w24340, w24341, w24342, w24343, w24344, w24345, w24346, w24347, w24348, w24349, w24350, w24351, w24352, w24353, w24354, w24355, w24356, w24357, w24358, w24359, w24360, w24361, w24362, w24363, w24364, w24365, w24366, w24367, w24368, w24369, w24370, w24371, w24372, w24373, w24374, w24375, w24376, w24377, w24378, w24379, w24380, w24381, w24382, w24383, w24384, w24385, w24386, w24387, w24388, w24389, w24390, w24391, w24392, w24393, w24394, w24395, w24396, w24397, w24398, w24399, w24400, w24401, w24402, w24403, w24404, w24405, w24406, w24407, w24408, w24409, w24410, w24411, w24412, w24413, w24414, w24415, w24416, w24417, w24418, w24419, w24420, w24421, w24422, w24423, w24424, w24425, w24426, w24427, w24428, w24429, w24430, w24431, w24432, w24433, w24434, w24435, w24436, w24437, w24438, w24439, w24440, w24441, w24442, w24443, w24444, w24445, w24446, w24447, w24448, w24449, w24450, w24451, w24452, w24453, w24454, w24455, w24456, w24457, w24458, w24459, w24460, w24461, w24462, w24463, w24464, w24465, w24466, w24467, w24468, w24469, w24470, w24471, w24472, w24473, w24474, w24475, w24476, w24477, w24478, w24479, w24480, w24481, w24482, w24483, w24484, w24485, w24486, w24487, w24488, w24489, w24490, w24491, w24492, w24493, w24494, w24495, w24496, w24497, w24498, w24499, w24500, w24501, w24502, w24503, w24504, w24505, w24506, w24507, w24508, w24509, w24510, w24511, w24512, w24513, w24514, w24515, w24516, w24517, w24518, w24519, w24520, w24521, w24522, w24523, w24524, w24525, w24526, w24527, w24528, w24529, w24530, w24531, w24532, w24533, w24534, w24535, w24536, w24537, w24538, w24539, w24540, w24541, w24542, w24543, w24544, w24545, w24546, w24547, w24548, w24549, w24550, w24551, w24552, w24553, w24554, w24555, w24556, w24557, w24558, w24559, w24560, w24561, w24562, w24563, w24564, w24565, w24566, w24567, w24568, w24569, w24570, w24571, w24572, w24573, w24574, w24575, w24576, w24577, w24578, w24579, w24580, w24581, w24582, w24583, w24584, w24585, w24586, w24587, w24588, w24589, w24590, w24591, w24592, w24593, w24594, w24595, w24596, w24597, w24598, w24599, w24600, w24601, w24602, w24603, w24604, w24605, w24606, w24607, w24608, w24609, w24610, w24611, w24612, w24613, w24614, w24615, w24616, w24617, w24618, w24619, w24620, w24621, w24622, w24623, w24624, w24625, w24626, w24627, w24628, w24629, w24630, w24631, w24632, w24633, w24634, w24635, w24636, w24637, w24638, w24639, w24640, w24641, w24642, w24643, w24644, w24645, w24646, w24647, w24648, w24649, w24650, w24651, w24652, w24653, w24654, w24655, w24656, w24657, w24658, w24659, w24660, w24661, w24662, w24663, w24664, w24665, w24666, w24667, w24668, w24669, w24670, w24671, w24672, w24673, w24674, w24675, w24676, w24677, w24678, w24679, w24680, w24681, w24682, w24683, w24684, w24685, w24686, w24687, w24688, w24689, w24690, w24691, w24692, w24693, w24694, w24695, w24696, w24697, w24698, w24699, w24700, w24701, w24702, w24703, w24704, w24705, w24706, w24707, w24708, w24709, w24710, w24711, w24712, w24713, w24714, w24715, w24716, w24717, w24718, w24719, w24720, w24721, w24722, w24723, w24724, w24725, w24726, w24727, w24728, w24729, w24730, w24731, w24732, w24733, w24734, w24735, w24736, w24737, w24738, w24739, w24740, w24741, w24742, w24743, w24744, w24745, w24746, w24747, w24748, w24749, w24750, w24751, w24752, w24753, w24754, w24755, w24756, w24757, w24758, w24759, w24760, w24761, w24762, w24763, w24764, w24765, w24766, w24767, w24768, w24769, w24770, w24771, w24772, w24773, w24774, w24775, w24776, w24777, w24778, w24779, w24780, w24781, w24782, w24783, w24784, w24785, w24786, w24787, w24788, w24789, w24790, w24791, w24792, w24793, w24794, w24795, w24796, w24797, w24798, w24799, w24800, w24801, w24802, w24803, w24804, w24805, w24806, w24807, w24808, w24809, w24810, w24811, w24812, w24813, w24814, w24815, w24816, w24817, w24818, w24819, w24820, w24821, w24822, w24823, w24824, w24825, w24826, w24827, w24828, w24829, w24830, w24831, w24832, w24833, w24834, w24835, w24836, w24837, w24838, w24839, w24840, w24841, w24842, w24843, w24844, w24845, w24846, w24847, w24848, w24849, w24850, w24851, w24852, w24853, w24854, w24855, w24856, w24857, w24858, w24859, w24860, w24861, w24862, w24863, w24864, w24865, w24866, w24867, w24868, w24869, w24870, w24871, w24872, w24873, w24874, w24875, w24876, w24877, w24878, w24879, w24880, w24881, w24882, w24883, w24884, w24885, w24886, w24887, w24888, w24889, w24890, w24891, w24892, w24893, w24894, w24895, w24896, w24897, w24898, w24899, w24900, w24901, w24902, w24903, w24904, w24905, w24906, w24907, w24908, w24909, w24910, w24911, w24912, w24913, w24914, w24915, w24916, w24917, w24918, w24919, w24920, w24921, w24922, w24923, w24924, w24925, w24926, w24927, w24928, w24929, w24930, w24931, w24932, w24933, w24934, w24935, w24936, w24937, w24938, w24939, w24940, w24941, w24942, w24943, w24944, w24945, w24946, w24947, w24948, w24949, w24950, w24951, w24952, w24953, w24954, w24955, w24956, w24957, w24958, w24959, w24960, w24961, w24962, w24963, w24964, w24965, w24966, w24967, w24968, w24969, w24970, w24971, w24972, w24973, w24974, w24975, w24976, w24977, w24978, w24979, w24980, w24981, w24982, w24983, w24984, w24985, w24986, w24987, w24988, w24989, w24990, w24991, w24992, w24993, w24994, w24995, w24996, w24997, w24998, w24999, w25000, w25001, w25002, w25003, w25004, w25005, w25006, w25007, w25008, w25009, w25010, w25011, w25012, w25013, w25014, w25015, w25016, w25017, w25018, w25019, w25020, w25021, w25022, w25023, w25024, w25025, w25026, w25027, w25028, w25029, w25030, w25031, w25032, w25033, w25034, w25035, w25036, w25037, w25038, w25039, w25040, w25041, w25042, w25043, w25044, w25045, w25046, w25047, w25048, w25049, w25050, w25051, w25052, w25053, w25054, w25055, w25056, w25057, w25058, w25059, w25060, w25061, w25062, w25063, w25064, w25065, w25066, w25067, w25068, w25069, w25070, w25071, w25072, w25073, w25074, w25075, w25076, w25077, w25078, w25079, w25080, w25081, w25082, w25083, w25084, w25085, w25086, w25087, w25088, w25089, w25090, w25091, w25092, w25093, w25094, w25095, w25096, w25097, w25098, w25099, w25100, w25101, w25102, w25103, w25104, w25105, w25106, w25107, w25108, w25109, w25110, w25111, w25112, w25113, w25114, w25115, w25116, w25117, w25118, w25119, w25120, w25121, w25122, w25123, w25124, w25125, w25126, w25127, w25128, w25129, w25130, w25131, w25132, w25133, w25134, w25135, w25136, w25137, w25138, w25139, w25140, w25141, w25142, w25143, w25144, w25145, w25146, w25147, w25148, w25149, w25150, w25151, w25152, w25153, w25154, w25155, w25156, w25157, w25158, w25159, w25160, w25161, w25162, w25163, w25164, w25165, w25166, w25167, w25168, w25169, w25170, w25171, w25172, w25173, w25174, w25175, w25176, w25177, w25178, w25179, w25180, w25181, w25182, w25183, w25184, w25185, w25186, w25187, w25188, w25189, w25190, w25191, w25192, w25193, w25194, w25195, w25196, w25197, w25198, w25199, w25200, w25201, w25202, w25203, w25204, w25205, w25206, w25207, w25208, w25209, w25210, w25211, w25212, w25213, w25214, w25215, w25216, w25217, w25218, w25219, w25220, w25221, w25222, w25223, w25224, w25225, w25226, w25227, w25228, w25229, w25230, w25231, w25232, w25233, w25234, w25235, w25236, w25237, w25238, w25239, w25240, w25241, w25242, w25243, w25244, w25245, w25246, w25247, w25248, w25249, w25250, w25251, w25252, w25253, w25254, w25255, w25256, w25257, w25258, w25259, w25260, w25261, w25262, w25263, w25264, w25265, w25266, w25267, w25268, w25269, w25270, w25271, w25272, w25273, w25274, w25275, w25276, w25277, w25278, w25279, w25280, w25281, w25282, w25283, w25284, w25285, w25286, w25287, w25288, w25289, w25290, w25291, w25292, w25293, w25294, w25295, w25296, w25297, w25298, w25299, w25300, w25301, w25302, w25303, w25304, w25305, w25306, w25307, w25308, w25309, w25310, w25311, w25312, w25313, w25314, w25315, w25316, w25317, w25318, w25319, w25320, w25321, w25322, w25323, w25324, w25325, w25326, w25327, w25328, w25329, w25330, w25331, w25332, w25333, w25334, w25335, w25336, w25337, w25338, w25339, w25340, w25341, w25342, w25343, w25344, w25345, w25346, w25347, w25348, w25349, w25350, w25351, w25352, w25353, w25354, w25355, w25356, w25357, w25358, w25359, w25360, w25361, w25362, w25363, w25364, w25365, w25366, w25367, w25368, w25369, w25370, w25371, w25372, w25373, w25374, w25375, w25376, w25377, w25378, w25379, w25380, w25381, w25382, w25383, w25384, w25385, w25386, w25387, w25388, w25389, w25390, w25391, w25392, w25393, w25394, w25395, w25396, w25397, w25398, w25399, w25400, w25401, w25402, w25403, w25404, w25405, w25406, w25407, w25408, w25409, w25410, w25411, w25412, w25413, w25414, w25415, w25416, w25417, w25418, w25419, w25420, w25421, w25422, w25423, w25424, w25425, w25426, w25427, w25428, w25429, w25430, w25431, w25432, w25433, w25434, w25435, w25436, w25437, w25438, w25439, w25440, w25441, w25442, w25443, w25444, w25445, w25446, w25447, w25448, w25449, w25450, w25451, w25452, w25453, w25454, w25455, w25456, w25457, w25458, w25459, w25460, w25461, w25462, w25463, w25464, w25465, w25466, w25467, w25468, w25469, w25470, w25471, w25472, w25473, w25474, w25475, w25476, w25477, w25478, w25479, w25480, w25481, w25482, w25483, w25484, w25485, w25486, w25487, w25488, w25489, w25490, w25491, w25492, w25493, w25494, w25495, w25496, w25497, w25498, w25499, w25500, w25501, w25502, w25503, w25504, w25505, w25506, w25507, w25508, w25509, w25510, w25511, w25512, w25513, w25514, w25515, w25516, w25517, w25518, w25519, w25520, w25521, w25522, w25523, w25524, w25525, w25526, w25527, w25528, w25529, w25530, w25531, w25532, w25533, w25534, w25535, w25536, w25537, w25538, w25539, w25540, w25541, w25542, w25543, w25544, w25545, w25546, w25547, w25548, w25549, w25550, w25551, w25552, w25553, w25554, w25555, w25556, w25557, w25558, w25559, w25560, w25561, w25562, w25563, w25564, w25565, w25566, w25567, w25568, w25569, w25570, w25571, w25572, w25573, w25574, w25575, w25576, w25577, w25578, w25579, w25580, w25581, w25582, w25583, w25584, w25585, w25586, w25587, w25588, w25589, w25590, w25591, w25592, w25593, w25594, w25595, w25596, w25597, w25598, w25599, w25600, w25601, w25602, w25603, w25604, w25605, w25606, w25607, w25608, w25609, w25610, w25611, w25612, w25613, w25614, w25615, w25616, w25617, w25618, w25619, w25620, w25621, w25622, w25623, w25624, w25625, w25626, w25627, w25628, w25629, w25630, w25631, w25632, w25633, w25634, w25635, w25636, w25637, w25638, w25639, w25640, w25641, w25642, w25643, w25644, w25645, w25646, w25647, w25648, w25649, w25650, w25651, w25652, w25653, w25654, w25655, w25656, w25657, w25658, w25659, w25660, w25661, w25662, w25663, w25664, w25665, w25666, w25667, w25668, w25669, w25670, w25671, w25672, w25673, w25674, w25675, w25676, w25677, w25678, w25679, w25680, w25681, w25682, w25683, w25684, w25685, w25686, w25687, w25688, w25689, w25690, w25691, w25692, w25693, w25694, w25695, w25696, w25697, w25698, w25699, w25700, w25701, w25702, w25703, w25704, w25705, w25706, w25707, w25708, w25709, w25710, w25711, w25712, w25713, w25714, w25715, w25716, w25717, w25718, w25719, w25720, w25721, w25722, w25723, w25724, w25725, w25726, w25727, w25728, w25729, w25730, w25731, w25732, w25733, w25734, w25735, w25736, w25737, w25738, w25739, w25740, w25741, w25742, w25743, w25744, w25745, w25746, w25747, w25748, w25749, w25750, w25751, w25752, w25753, w25754, w25755, w25756, w25757, w25758, w25759, w25760, w25761, w25762, w25763, w25764, w25765, w25766, w25767, w25768, w25769, w25770, w25771, w25772, w25773, w25774, w25775, w25776, w25777, w25778, w25779, w25780, w25781, w25782, w25783, w25784, w25785, w25786, w25787, w25788, w25789, w25790, w25791, w25792, w25793, w25794, w25795, w25796, w25797, w25798, w25799, w25800, w25801, w25802, w25803, w25804, w25805, w25806, w25807, w25808, w25809, w25810, w25811, w25812, w25813, w25814, w25815, w25816, w25817, w25818, w25819, w25820, w25821, w25822, w25823, w25824, w25825, w25826, w25827, w25828, w25829, w25830, w25831, w25832, w25833, w25834, w25835, w25836, w25837, w25838, w25839, w25840, w25841, w25842, w25843, w25844, w25845, w25846, w25847, w25848, w25849, w25850, w25851, w25852, w25853, w25854, w25855, w25856, w25857, w25858, w25859, w25860, w25861, w25862, w25863, w25864, w25865, w25866, w25867, w25868, w25869, w25870, w25871, w25872, w25873, w25874, w25875, w25876, w25877, w25878, w25879, w25880, w25881, w25882, w25883, w25884, w25885, w25886, w25887, w25888, w25889, w25890, w25891, w25892, w25893, w25894, w25895, w25896, w25897, w25898, w25899, w25900, w25901, w25902, w25903, w25904, w25905, w25906, w25907, w25908, w25909, w25910, w25911, w25912, w25913, w25914, w25915, w25916, w25917, w25918, w25919, w25920, w25921, w25922, w25923, w25924, w25925, w25926, w25927, w25928, w25929, w25930, w25931, w25932, w25933, w25934, w25935, w25936, w25937, w25938, w25939, w25940, w25941, w25942, w25943, w25944, w25945, w25946, w25947, w25948, w25949, w25950, w25951, w25952, w25953, w25954, w25955, w25956, w25957, w25958, w25959, w25960, w25961, w25962, w25963, w25964, w25965, w25966, w25967, w25968, w25969, w25970, w25971, w25972, w25973, w25974, w25975, w25976, w25977, w25978, w25979, w25980, w25981, w25982, w25983, w25984, w25985, w25986, w25987, w25988, w25989, w25990, w25991, w25992, w25993, w25994, w25995, w25996, w25997, w25998, w25999, w26000, w26001, w26002, w26003, w26004, w26005, w26006, w26007, w26008, w26009, w26010, w26011, w26012, w26013, w26014, w26015, w26016, w26017, w26018, w26019, w26020, w26021, w26022, w26023, w26024, w26025, w26026, w26027, w26028, w26029, w26030, w26031, w26032, w26033, w26034, w26035, w26036, w26037, w26038, w26039, w26040, w26041, w26042, w26043, w26044, w26045, w26046, w26047, w26048, w26049, w26050, w26051, w26052, w26053, w26054, w26055, w26056, w26057, w26058, w26059, w26060, w26061, w26062, w26063, w26064, w26065, w26066, w26067, w26068, w26069, w26070, w26071, w26072, w26073, w26074, w26075, w26076, w26077, w26078, w26079, w26080, w26081, w26082, w26083, w26084, w26085, w26086, w26087, w26088, w26089, w26090, w26091, w26092, w26093, w26094, w26095, w26096, w26097, w26098, w26099, w26100, w26101, w26102, w26103, w26104, w26105, w26106, w26107, w26108, w26109, w26110, w26111, w26112, w26113, w26114, w26115, w26116, w26117, w26118, w26119, w26120, w26121, w26122, w26123, w26124, w26125, w26126, w26127, w26128, w26129, w26130, w26131, w26132, w26133, w26134, w26135, w26136, w26137, w26138, w26139, w26140, w26141, w26142, w26143, w26144, w26145, w26146, w26147, w26148, w26149, w26150, w26151, w26152, w26153, w26154, w26155, w26156, w26157, w26158, w26159, w26160, w26161, w26162, w26163, w26164, w26165, w26166, w26167, w26168, w26169, w26170, w26171, w26172, w26173, w26174, w26175, w26176, w26177, w26178, w26179, w26180, w26181, w26182, w26183, w26184, w26185, w26186, w26187, w26188, w26189, w26190, w26191, w26192, w26193, w26194, w26195, w26196, w26197, w26198, w26199, w26200, w26201, w26202, w26203, w26204, w26205, w26206, w26207, w26208, w26209, w26210, w26211, w26212, w26213, w26214, w26215, w26216, w26217, w26218, w26219, w26220, w26221, w26222, w26223, w26224, w26225, w26226, w26227, w26228, w26229, w26230, w26231, w26232, w26233, w26234, w26235, w26236, w26237, w26238, w26239, w26240, w26241, w26242, w26243, w26244, w26245, w26246, w26247, w26248, w26249, w26250, w26251, w26252, w26253, w26254, w26255, w26256, w26257, w26258, w26259, w26260, w26261, w26262, w26263, w26264, w26265, w26266, w26267, w26268, w26269, w26270, w26271, w26272, w26273, w26274, w26275, w26276, w26277, w26278, w26279, w26280, w26281, w26282, w26283, w26284, w26285, w26286, w26287, w26288, w26289, w26290, w26291, w26292, w26293, w26294, w26295, w26296, w26297, w26298, w26299, w26300, w26301, w26302, w26303, w26304, w26305, w26306, w26307, w26308, w26309, w26310, w26311, w26312, w26313, w26314, w26315, w26316, w26317, w26318, w26319, w26320, w26321, w26322, w26323, w26324, w26325, w26326, w26327, w26328, w26329, w26330, w26331, w26332, w26333, w26334, w26335, w26336, w26337, w26338, w26339, w26340, w26341, w26342, w26343, w26344, w26345, w26346, w26347, w26348, w26349, w26350, w26351, w26352, w26353, w26354, w26355, w26356, w26357, w26358, w26359, w26360, w26361, w26362, w26363, w26364, w26365, w26366, w26367, w26368, w26369, w26370, w26371, w26372, w26373, w26374, w26375, w26376, w26377, w26378, w26379, w26380, w26381, w26382, w26383, w26384, w26385, w26386, w26387, w26388, w26389, w26390, w26391, w26392, w26393, w26394, w26395, w26396, w26397, w26398, w26399, w26400, w26401, w26402, w26403, w26404, w26405, w26406, w26407, w26408, w26409, w26410, w26411, w26412, w26413, w26414, w26415, w26416, w26417, w26418, w26419, w26420, w26421, w26422, w26423, w26424, w26425, w26426, w26427, w26428, w26429, w26430, w26431, w26432, w26433, w26434, w26435, w26436, w26437, w26438, w26439, w26440, w26441, w26442, w26443, w26444, w26445, w26446, w26447, w26448, w26449, w26450, w26451, w26452, w26453, w26454, w26455, w26456, w26457, w26458, w26459, w26460, w26461, w26462, w26463, w26464, w26465, w26466, w26467, w26468, w26469, w26470, w26471, w26472, w26473, w26474, w26475, w26476, w26477, w26478, w26479, w26480, w26481, w26482, w26483, w26484, w26485, w26486, w26487, w26488, w26489, w26490, w26491, w26492, w26493, w26494, w26495, w26496, w26497, w26498, w26499, w26500, w26501, w26502, w26503, w26504, w26505, w26506, w26507, w26508, w26509, w26510, w26511, w26512, w26513, w26514, w26515, w26516, w26517, w26518, w26519, w26520, w26521, w26522, w26523, w26524, w26525, w26526, w26527, w26528, w26529, w26530, w26531, w26532, w26533, w26534, w26535, w26536, w26537, w26538, w26539, w26540, w26541, w26542, w26543, w26544, w26545, w26546, w26547, w26548, w26549, w26550, w26551, w26552, w26553, w26554, w26555, w26556, w26557, w26558, w26559, w26560, w26561, w26562, w26563, w26564, w26565, w26566, w26567, w26568, w26569, w26570, w26571, w26572, w26573, w26574, w26575, w26576, w26577, w26578, w26579, w26580, w26581, w26582, w26583, w26584, w26585, w26586, w26587, w26588, w26589, w26590, w26591, w26592, w26593, w26594, w26595, w26596, w26597, w26598, w26599, w26600, w26601, w26602, w26603, w26604, w26605, w26606, w26607, w26608, w26609, w26610, w26611, w26612, w26613, w26614, w26615, w26616, w26617, w26618, w26619, w26620, w26621, w26622, w26623, w26624, w26625, w26626, w26627, w26628, w26629, w26630, w26631, w26632, w26633, w26634, w26635, w26636, w26637, w26638, w26639, w26640, w26641, w26642, w26643, w26644, w26645, w26646, w26647, w26648, w26649, w26650, w26651, w26652, w26653, w26654, w26655, w26656, w26657, w26658, w26659, w26660, w26661, w26662, w26663, w26664, w26665, w26666, w26667, w26668, w26669, w26670, w26671, w26672, w26673, w26674, w26675, w26676, w26677, w26678, w26679, w26680, w26681, w26682, w26683, w26684, w26685, w26686, w26687, w26688, w26689, w26690, w26691, w26692, w26693, w26694, w26695, w26696, w26697, w26698, w26699, w26700, w26701, w26702, w26703, w26704, w26705, w26706, w26707, w26708, w26709, w26710, w26711, w26712, w26713, w26714, w26715, w26716, w26717, w26718, w26719, w26720, w26721, w26722, w26723, w26724, w26725, w26726, w26727, w26728, w26729, w26730, w26731, w26732, w26733, w26734, w26735, w26736, w26737, w26738, w26739, w26740, w26741, w26742, w26743, w26744, w26745, w26746, w26747, w26748, w26749, w26750, w26751, w26752, w26753, w26754, w26755, w26756, w26757, w26758, w26759, w26760, w26761, w26762, w26763, w26764, w26765, w26766, w26767, w26768, w26769, w26770, w26771, w26772, w26773, w26774, w26775, w26776, w26777, w26778, w26779, w26780, w26781, w26782, w26783, w26784, w26785, w26786, w26787, w26788, w26789, w26790, w26791, w26792, w26793, w26794, w26795, w26796, w26797, w26798, w26799, w26800, w26801, w26802, w26803, w26804, w26805, w26806, w26807, w26808, w26809, w26810, w26811, w26812, w26813, w26814, w26815, w26816, w26817, w26818, w26819, w26820, w26821, w26822, w26823, w26824, w26825, w26826, w26827, w26828, w26829, w26830, w26831, w26832, w26833, w26834, w26835, w26836, w26837, w26838, w26839, w26840, w26841, w26842, w26843, w26844, w26845, w26846, w26847, w26848, w26849, w26850, w26851, w26852, w26853, w26854, w26855, w26856, w26857, w26858, w26859, w26860, w26861, w26862, w26863, w26864, w26865, w26866, w26867, w26868, w26869, w26870, w26871, w26872, w26873, w26874, w26875, w26876, w26877, w26878, w26879, w26880, w26881, w26882, w26883, w26884, w26885, w26886, w26887, w26888, w26889, w26890, w26891, w26892, w26893, w26894, w26895, w26896, w26897, w26898, w26899, w26900, w26901, w26902, w26903, w26904, w26905, w26906, w26907, w26908, w26909, w26910, w26911, w26912, w26913, w26914, w26915, w26916, w26917, w26918, w26919, w26920, w26921, w26922, w26923, w26924, w26925, w26926, w26927, w26928, w26929, w26930, w26931, w26932, w26933, w26934, w26935, w26936, w26937, w26938, w26939, w26940, w26941, w26942, w26943, w26944, w26945, w26946, w26947, w26948, w26949, w26950, w26951, w26952, w26953, w26954, w26955, w26956, w26957, w26958, w26959, w26960, w26961, w26962, w26963, w26964, w26965, w26966, w26967, w26968, w26969, w26970, w26971, w26972, w26973, w26974, w26975, w26976, w26977, w26978, w26979, w26980, w26981, w26982, w26983, w26984, w26985, w26986, w26987, w26988, w26989, w26990, w26991, w26992, w26993, w26994, w26995, w26996, w26997, w26998, w26999, w27000, w27001, w27002, w27003, w27004, w27005, w27006, w27007, w27008, w27009, w27010, w27011, w27012, w27013, w27014, w27015, w27016, w27017, w27018, w27019, w27020, w27021, w27022, w27023, w27024, w27025, w27026, w27027, w27028, w27029, w27030, w27031, w27032, w27033, w27034, w27035, w27036, w27037, w27038, w27039, w27040, w27041, w27042, w27043, w27044, w27045, w27046, w27047, w27048, w27049, w27050, w27051, w27052, w27053, w27054, w27055, w27056, w27057, w27058, w27059, w27060, w27061, w27062, w27063, w27064, w27065, w27066, w27067, w27068, w27069, w27070, w27071, w27072, w27073, w27074, w27075, w27076, w27077, w27078, w27079, w27080, w27081, w27082, w27083, w27084, w27085, w27086, w27087, w27088, w27089, w27090, w27091, w27092, w27093, w27094, w27095, w27096, w27097, w27098, w27099, w27100, w27101, w27102, w27103, w27104, w27105, w27106, w27107, w27108, w27109, w27110, w27111, w27112, w27113, w27114, w27115, w27116, w27117, w27118, w27119, w27120, w27121, w27122, w27123, w27124, w27125, w27126, w27127, w27128, w27129, w27130, w27131, w27132, w27133, w27134, w27135, w27136, w27137, w27138, w27139, w27140, w27141, w27142, w27143, w27144, w27145, w27146, w27147, w27148, w27149, w27150, w27151, w27152, w27153, w27154, w27155, w27156, w27157, w27158, w27159, w27160, w27161, w27162, w27163, w27164, w27165, w27166, w27167, w27168, w27169, w27170, w27171, w27172, w27173, w27174, w27175, w27176, w27177, w27178, w27179, w27180, w27181, w27182, w27183, w27184, w27185, w27186, w27187, w27188, w27189, w27190, w27191, w27192, w27193, w27194, w27195, w27196, w27197, w27198, w27199, w27200, w27201, w27202, w27203, w27204, w27205, w27206, w27207, w27208, w27209, w27210, w27211, w27212, w27213, w27214, w27215, w27216, w27217, w27218, w27219, w27220, w27221, w27222, w27223, w27224, w27225, w27226, w27227, w27228, w27229, w27230, w27231, w27232, w27233, w27234, w27235, w27236, w27237, w27238, w27239, w27240, w27241, w27242, w27243, w27244, w27245, w27246, w27247, w27248, w27249, w27250, w27251, w27252, w27253, w27254, w27255, w27256, w27257, w27258, w27259, w27260, w27261, w27262, w27263, w27264, w27265, w27266, w27267, w27268, w27269, w27270, w27271, w27272, w27273, w27274, w27275, w27276, w27277, w27278, w27279, w27280, w27281, w27282, w27283, w27284, w27285, w27286, w27287, w27288, w27289, w27290, w27291, w27292, w27293, w27294, w27295, w27296, w27297, w27298, w27299, w27300, w27301, w27302, w27303, w27304, w27305, w27306, w27307, w27308, w27309, w27310, w27311, w27312, w27313, w27314, w27315, w27316, w27317, w27318, w27319, w27320, w27321, w27322, w27323, w27324, w27325, w27326, w27327, w27328, w27329, w27330, w27331, w27332, w27333, w27334, w27335, w27336, w27337, w27338, w27339, w27340, w27341, w27342, w27343, w27344, w27345, w27346, w27347, w27348, w27349, w27350, w27351, w27352, w27353, w27354, w27355, w27356, w27357, w27358, w27359, w27360, w27361, w27362, w27363, w27364, w27365, w27366, w27367, w27368, w27369, w27370, w27371, w27372, w27373, w27374, w27375, w27376, w27377, w27378, w27379, w27380, w27381, w27382, w27383, w27384, w27385, w27386, w27387, w27388, w27389, w27390, w27391, w27392, w27393, w27394, w27395, w27396, w27397, w27398, w27399, w27400, w27401, w27402, w27403, w27404, w27405, w27406, w27407, w27408, w27409, w27410, w27411, w27412, w27413, w27414, w27415, w27416, w27417, w27418, w27419, w27420, w27421, w27422, w27423, w27424, w27425, w27426, w27427, w27428, w27429, w27430, w27431, w27432, w27433, w27434, w27435, w27436, w27437, w27438, w27439, w27440, w27441, w27442, w27443, w27444, w27445, w27446, w27447, w27448, w27449, w27450, w27451, w27452, w27453, w27454, w27455, w27456, w27457, w27458, w27459, w27460, w27461, w27462, w27463, w27464, w27465, w27466, w27467, w27468, w27469, w27470, w27471, w27472, w27473, w27474, w27475, w27476, w27477, w27478, w27479, w27480, w27481, w27482, w27483, w27484, w27485, w27486, w27487, w27488, w27489, w27490, w27491, w27492, w27493, w27494, w27495, w27496, w27497, w27498, w27499, w27500, w27501, w27502, w27503, w27504, w27505, w27506, w27507, w27508, w27509, w27510, w27511, w27512, w27513, w27514, w27515, w27516, w27517, w27518, w27519, w27520, w27521, w27522, w27523, w27524, w27525, w27526, w27527, w27528, w27529, w27530, w27531, w27532, w27533, w27534, w27535, w27536, w27537, w27538, w27539, w27540, w27541, w27542, w27543, w27544, w27545, w27546, w27547, w27548, w27549, w27550, w27551, w27552, w27553, w27554, w27555, w27556, w27557, w27558, w27559, w27560, w27561, w27562, w27563, w27564, w27565, w27566, w27567, w27568, w27569, w27570, w27571, w27572, w27573, w27574, w27575, w27576, w27577, w27578, w27579, w27580, w27581, w27582, w27583, w27584, w27585, w27586, w27587, w27588, w27589, w27590, w27591, w27592, w27593, w27594, w27595, w27596, w27597, w27598, w27599, w27600, w27601, w27602, w27603, w27604, w27605, w27606, w27607, w27608, w27609, w27610, w27611, w27612, w27613, w27614, w27615, w27616, w27617, w27618, w27619, w27620, w27621, w27622, w27623, w27624, w27625, w27626, w27627, w27628, w27629, w27630, w27631, w27632, w27633, w27634, w27635, w27636, w27637, w27638, w27639, w27640, w27641, w27642, w27643, w27644, w27645, w27646, w27647, w27648, w27649, w27650, w27651, w27652, w27653, w27654, w27655, w27656, w27657, w27658, w27659, w27660, w27661, w27662, w27663, w27664, w27665, w27666, w27667, w27668, w27669, w27670, w27671, w27672, w27673, w27674, w27675, w27676, w27677, w27678, w27679, w27680, w27681, w27682, w27683, w27684, w27685, w27686, w27687, w27688, w27689, w27690, w27691, w27692, w27693, w27694, w27695, w27696, w27697, w27698, w27699, w27700, w27701, w27702, w27703, w27704, w27705, w27706, w27707, w27708, w27709, w27710, w27711, w27712, w27713, w27714, w27715, w27716, w27717, w27718, w27719, w27720, w27721, w27722, w27723, w27724, w27725, w27726, w27727, w27728, w27729, w27730, w27731, w27732, w27733, w27734, w27735, w27736, w27737, w27738, w27739, w27740, w27741, w27742, w27743, w27744, w27745, w27746, w27747, w27748, w27749, w27750, w27751, w27752, w27753, w27754, w27755, w27756, w27757, w27758, w27759, w27760, w27761, w27762, w27763, w27764, w27765, w27766, w27767, w27768, w27769, w27770, w27771, w27772, w27773, w27774, w27775, w27776, w27777, w27778, w27779, w27780, w27781, w27782, w27783, w27784, w27785, w27786, w27787, w27788, w27789, w27790, w27791, w27792, w27793, w27794, w27795, w27796, w27797, w27798, w27799, w27800, w27801, w27802, w27803, w27804, w27805, w27806, w27807, w27808, w27809, w27810, w27811, w27812, w27813, w27814, w27815, w27816, w27817, w27818, w27819, w27820, w27821, w27822, w27823, w27824, w27825, w27826, w27827, w27828, w27829, w27830, w27831, w27832, w27833, w27834, w27835, w27836, w27837, w27838, w27839, w27840, w27841, w27842, w27843, w27844, w27845, w27846, w27847, w27848, w27849, w27850, w27851, w27852, w27853, w27854, w27855, w27856, w27857, w27858, w27859, w27860, w27861, w27862, w27863, w27864, w27865, w27866, w27867, w27868, w27869, w27870, w27871, w27872, w27873, w27874, w27875, w27876, w27877, w27878, w27879, w27880, w27881, w27882, w27883, w27884, w27885, w27886, w27887, w27888, w27889, w27890, w27891, w27892, w27893, w27894, w27895, w27896, w27897, w27898, w27899, w27900, w27901, w27902, w27903, w27904, w27905, w27906, w27907, w27908, w27909, w27910, w27911, w27912, w27913, w27914, w27915, w27916, w27917, w27918, w27919, w27920, w27921, w27922, w27923, w27924, w27925, w27926, w27927, w27928, w27929, w27930, w27931, w27932, w27933, w27934, w27935, w27936, w27937, w27938, w27939, w27940, w27941, w27942, w27943, w27944, w27945, w27946, w27947, w27948, w27949, w27950, w27951, w27952, w27953, w27954, w27955, w27956, w27957, w27958, w27959, w27960, w27961, w27962, w27963, w27964, w27965, w27966, w27967, w27968, w27969, w27970, w27971, w27972, w27973, w27974, w27975, w27976, w27977, w27978, w27979, w27980, w27981, w27982, w27983, w27984, w27985, w27986, w27987, w27988, w27989, w27990, w27991, w27992, w27993, w27994, w27995, w27996, w27997, w27998, w27999, w28000, w28001, w28002, w28003, w28004, w28005, w28006, w28007, w28008, w28009, w28010, w28011, w28012, w28013, w28014, w28015, w28016, w28017, w28018, w28019, w28020, w28021, w28022, w28023, w28024, w28025, w28026, w28027, w28028, w28029, w28030, w28031, w28032, w28033, w28034, w28035, w28036, w28037, w28038, w28039, w28040, w28041, w28042, w28043, w28044, w28045, w28046, w28047, w28048, w28049, w28050, w28051, w28052, w28053, w28054, w28055, w28056, w28057, w28058, w28059, w28060, w28061, w28062, w28063, w28064, w28065, w28066, w28067, w28068, w28069, w28070, w28071, w28072, w28073, w28074, w28075, w28076, w28077, w28078, w28079, w28080, w28081, w28082, w28083, w28084, w28085, w28086, w28087, w28088, w28089, w28090, w28091, w28092, w28093, w28094, w28095, w28096, w28097, w28098, w28099, w28100, w28101, w28102, w28103, w28104, w28105, w28106, w28107, w28108, w28109, w28110, w28111, w28112, w28113, w28114, w28115, w28116, w28117, w28118, w28119, w28120, w28121, w28122, w28123, w28124, w28125, w28126, w28127, w28128, w28129, w28130, w28131, w28132, w28133, w28134, w28135, w28136, w28137, w28138, w28139, w28140, w28141, w28142, w28143, w28144, w28145, w28146, w28147, w28148, w28149, w28150, w28151, w28152, w28153, w28154, w28155, w28156, w28157, w28158, w28159, w28160, w28161, w28162, w28163, w28164, w28165, w28166, w28167, w28168, w28169, w28170, w28171, w28172, w28173, w28174, w28175, w28176, w28177, w28178, w28179, w28180, w28181, w28182, w28183, w28184, w28185, w28186, w28187, w28188, w28189, w28190, w28191, w28192, w28193, w28194, w28195, w28196, w28197, w28198, w28199, w28200, w28201, w28202, w28203, w28204, w28205, w28206, w28207, w28208, w28209, w28210, w28211, w28212, w28213, w28214, w28215, w28216, w28217, w28218, w28219, w28220, w28221, w28222, w28223, w28224, w28225, w28226, w28227, w28228, w28229, w28230, w28231, w28232, w28233, w28234, w28235, w28236, w28237, w28238, w28239, w28240, w28241, w28242, w28243, w28244, w28245, w28246, w28247, w28248, w28249, w28250, w28251, w28252, w28253, w28254, w28255, w28256, w28257, w28258, w28259, w28260, w28261, w28262, w28263, w28264, w28265, w28266, w28267, w28268, w28269, w28270, w28271, w28272, w28273, w28274, w28275, w28276, w28277, w28278, w28279, w28280, w28281, w28282, w28283, w28284, w28285, w28286, w28287, w28288, w28289, w28290, w28291, w28292, w28293, w28294, w28295, w28296, w28297, w28298, w28299, w28300, w28301, w28302, w28303, w28304, w28305, w28306, w28307, w28308, w28309, w28310, w28311, w28312, w28313, w28314, w28315, w28316, w28317, w28318, w28319, w28320, w28321, w28322, w28323, w28324, w28325, w28326, w28327, w28328, w28329, w28330, w28331, w28332, w28333, w28334, w28335, w28336, w28337, w28338, w28339, w28340, w28341, w28342, w28343, w28344, w28345, w28346, w28347, w28348, w28349, w28350, w28351, w28352, w28353, w28354, w28355, w28356, w28357, w28358, w28359, w28360, w28361, w28362, w28363, w28364, w28365, w28366, w28367, w28368, w28369, w28370, w28371, w28372, w28373, w28374, w28375, w28376, w28377, w28378, w28379, w28380, w28381, w28382, w28383, w28384, w28385, w28386, w28387, w28388, w28389, w28390, w28391, w28392, w28393, w28394, w28395, w28396, w28397, w28398, w28399, w28400, w28401, w28402, w28403, w28404, w28405, w28406, w28407, w28408, w28409, w28410, w28411, w28412, w28413, w28414, w28415, w28416, w28417, w28418, w28419, w28420, w28421, w28422, w28423, w28424, w28425, w28426, w28427, w28428, w28429, w28430, w28431, w28432, w28433, w28434, w28435, w28436, w28437, w28438, w28439, w28440, w28441, w28442, w28443, w28444, w28445, w28446, w28447, w28448, w28449, w28450, w28451, w28452, w28453, w28454, w28455, w28456, w28457, w28458, w28459, w28460, w28461, w28462, w28463, w28464, w28465, w28466, w28467, w28468, w28469, w28470, w28471, w28472, w28473, w28474, w28475, w28476, w28477, w28478, w28479, w28480, w28481, w28482, w28483, w28484, w28485, w28486, w28487, w28488, w28489, w28490, w28491, w28492, w28493, w28494, w28495, w28496, w28497, w28498, w28499, w28500, w28501, w28502, w28503, w28504, w28505, w28506, w28507, w28508, w28509, w28510, w28511, w28512, w28513, w28514, w28515, w28516, w28517, w28518, w28519, w28520, w28521, w28522, w28523, w28524, w28525, w28526, w28527, w28528, w28529, w28530, w28531, w28532, w28533, w28534, w28535, w28536, w28537, w28538, w28539, w28540, w28541, w28542, w28543, w28544, w28545, w28546, w28547, w28548, w28549, w28550, w28551, w28552, w28553, w28554, w28555, w28556, w28557, w28558, w28559, w28560, w28561, w28562, w28563, w28564, w28565, w28566, w28567, w28568, w28569, w28570, w28571, w28572, w28573, w28574, w28575, w28576, w28577, w28578, w28579, w28580, w28581, w28582, w28583, w28584, w28585, w28586, w28587, w28588, w28589, w28590, w28591, w28592, w28593, w28594, w28595, w28596, w28597, w28598, w28599, w28600, w28601, w28602, w28603, w28604, w28605, w28606, w28607, w28608, w28609, w28610, w28611, w28612, w28613, w28614, w28615, w28616, w28617, w28618, w28619, w28620, w28621, w28622, w28623, w28624, w28625, w28626, w28627, w28628, w28629, w28630, w28631, w28632, w28633, w28634, w28635, w28636, w28637, w28638, w28639, w28640, w28641, w28642, w28643, w28644, w28645, w28646, w28647, w28648, w28649, w28650, w28651, w28652, w28653, w28654, w28655, w28656, w28657, w28658, w28659, w28660, w28661, w28662, w28663, w28664, w28665, w28666, w28667, w28668, w28669, w28670, w28671, w28672, w28673, w28674, w28675, w28676, w28677, w28678, w28679, w28680, w28681, w28682, w28683, w28684, w28685, w28686, w28687, w28688, w28689, w28690, w28691, w28692, w28693, w28694, w28695, w28696, w28697, w28698, w28699, w28700, w28701, w28702, w28703, w28704, w28705, w28706, w28707, w28708, w28709, w28710, w28711, w28712, w28713, w28714, w28715, w28716, w28717, w28718, w28719, w28720, w28721, w28722, w28723, w28724, w28725, w28726, w28727, w28728, w28729, w28730, w28731, w28732, w28733, w28734, w28735, w28736, w28737, w28738, w28739, w28740, w28741, w28742, w28743, w28744, w28745, w28746, w28747, w28748, w28749, w28750, w28751, w28752, w28753, w28754, w28755, w28756, w28757, w28758, w28759, w28760, w28761, w28762, w28763, w28764, w28765, w28766, w28767, w28768, w28769, w28770, w28771, w28772, w28773, w28774, w28775, w28776, w28777, w28778, w28779, w28780, w28781, w28782, w28783, w28784, w28785, w28786, w28787, w28788, w28789, w28790, w28791, w28792, w28793, w28794, w28795, w28796, w28797, w28798, w28799, w28800, w28801, w28802, w28803, w28804, w28805, w28806, w28807, w28808, w28809, w28810, w28811, w28812, w28813, w28814, w28815, w28816, w28817, w28818, w28819, w28820, w28821, w28822, w28823, w28824, w28825, w28826, w28827, w28828, w28829, w28830, w28831, w28832, w28833, w28834, w28835, w28836, w28837, w28838, w28839, w28840, w28841, w28842, w28843, w28844, w28845, w28846, w28847, w28848, w28849, w28850, w28851, w28852, w28853, w28854, w28855, w28856, w28857, w28858, w28859, w28860, w28861, w28862, w28863, w28864, w28865, w28866, w28867, w28868, w28869, w28870, w28871, w28872, w28873, w28874, w28875, w28876, w28877, w28878, w28879, w28880, w28881, w28882, w28883, w28884, w28885, w28886, w28887, w28888, w28889, w28890, w28891, w28892, w28893, w28894, w28895, w28896, w28897, w28898, w28899, w28900, w28901, w28902, w28903, w28904, w28905, w28906, w28907, w28908, w28909, w28910, w28911, w28912, w28913, w28914, w28915, w28916, w28917, w28918, w28919, w28920, w28921, w28922, w28923, w28924, w28925, w28926, w28927, w28928, w28929, w28930, w28931, w28932, w28933, w28934, w28935, w28936, w28937, w28938, w28939, w28940, w28941, w28942, w28943, w28944, w28945, w28946, w28947, w28948, w28949, w28950, w28951, w28952, w28953, w28954, w28955, w28956, w28957, w28958, w28959, w28960, w28961, w28962, w28963, w28964, w28965, w28966, w28967, w28968, w28969, w28970, w28971, w28972, w28973, w28974, w28975, w28976, w28977, w28978, w28979, w28980, w28981, w28982, w28983, w28984, w28985, w28986, w28987, w28988, w28989, w28990, w28991, w28992, w28993, w28994, w28995, w28996, w28997, w28998, w28999, w29000, w29001, w29002, w29003, w29004, w29005, w29006, w29007, w29008, w29009, w29010, w29011, w29012, w29013, w29014, w29015, w29016, w29017, w29018, w29019, w29020, w29021, w29022, w29023, w29024, w29025, w29026, w29027, w29028, w29029, w29030, w29031, w29032, w29033, w29034, w29035, w29036, w29037, w29038, w29039, w29040, w29041, w29042, w29043, w29044, w29045, w29046, w29047, w29048, w29049, w29050, w29051, w29052, w29053, w29054, w29055, w29056, w29057, w29058, w29059, w29060, w29061, w29062, w29063, w29064, w29065, w29066, w29067, w29068, w29069, w29070, w29071, w29072, w29073, w29074, w29075, w29076, w29077, w29078, w29079, w29080, w29081, w29082, w29083, w29084, w29085, w29086, w29087, w29088, w29089, w29090, w29091, w29092, w29093, w29094, w29095, w29096, w29097, w29098, w29099, w29100, w29101, w29102, w29103, w29104, w29105, w29106, w29107, w29108, w29109, w29110, w29111, w29112, w29113, w29114, w29115, w29116, w29117, w29118, w29119, w29120, w29121, w29122, w29123, w29124, w29125, w29126, w29127, w29128, w29129, w29130, w29131, w29132, w29133, w29134, w29135, w29136, w29137, w29138, w29139, w29140, w29141, w29142, w29143, w29144, w29145, w29146, w29147, w29148, w29149, w29150, w29151, w29152, w29153, w29154, w29155, w29156, w29157, w29158, w29159, w29160, w29161, w29162, w29163, w29164, w29165, w29166, w29167, w29168, w29169, w29170, w29171, w29172, w29173, w29174, w29175, w29176, w29177, w29178, w29179, w29180, w29181, w29182, w29183, w29184, w29185, w29186, w29187, w29188, w29189, w29190, w29191, w29192, w29193, w29194, w29195, w29196, w29197, w29198, w29199, w29200, w29201, w29202, w29203, w29204, w29205, w29206, w29207, w29208, w29209, w29210, w29211, w29212, w29213, w29214, w29215, w29216, w29217, w29218, w29219, w29220, w29221, w29222, w29223, w29224, w29225, w29226, w29227, w29228, w29229, w29230, w29231, w29232, w29233, w29234, w29235, w29236, w29237, w29238, w29239, w29240, w29241, w29242, w29243, w29244, w29245, w29246, w29247, w29248, w29249, w29250, w29251, w29252, w29253, w29254, w29255, w29256, w29257, w29258, w29259, w29260, w29261, w29262, w29263, w29264, w29265, w29266, w29267, w29268, w29269, w29270, w29271, w29272, w29273, w29274, w29275, w29276, w29277, w29278, w29279, w29280, w29281, w29282, w29283, w29284, w29285, w29286, w29287, w29288, w29289, w29290, w29291, w29292, w29293, w29294, w29295, w29296, w29297, w29298, w29299, w29300, w29301, w29302, w29303, w29304, w29305, w29306, w29307, w29308, w29309, w29310, w29311, w29312, w29313, w29314, w29315, w29316, w29317, w29318, w29319, w29320, w29321, w29322, w29323, w29324, w29325, w29326, w29327, w29328, w29329, w29330, w29331, w29332, w29333, w29334, w29335, w29336, w29337, w29338, w29339, w29340, w29341, w29342, w29343, w29344, w29345, w29346, w29347, w29348, w29349, w29350, w29351, w29352, w29353, w29354, w29355, w29356, w29357, w29358, w29359, w29360, w29361, w29362, w29363, w29364, w29365, w29366, w29367, w29368, w29369, w29370, w29371, w29372, w29373, w29374, w29375, w29376, w29377, w29378, w29379, w29380, w29381, w29382, w29383, w29384, w29385, w29386, w29387, w29388, w29389, w29390, w29391, w29392, w29393, w29394, w29395, w29396, w29397, w29398, w29399, w29400, w29401, w29402, w29403, w29404, w29405, w29406, w29407, w29408, w29409, w29410, w29411, w29412, w29413, w29414, w29415, w29416, w29417, w29418, w29419, w29420, w29421, w29422, w29423, w29424, w29425, w29426, w29427, w29428, w29429, w29430, w29431, w29432, w29433, w29434, w29435, w29436, w29437, w29438, w29439, w29440, w29441, w29442, w29443, w29444, w29445, w29446, w29447, w29448, w29449, w29450, w29451, w29452, w29453, w29454, w29455, w29456, w29457, w29458, w29459, w29460, w29461, w29462, w29463, w29464, w29465, w29466, w29467, w29468, w29469, w29470, w29471, w29472, w29473, w29474, w29475, w29476, w29477, w29478, w29479, w29480, w29481, w29482, w29483, w29484, w29485, w29486, w29487, w29488, w29489, w29490, w29491, w29492, w29493, w29494, w29495, w29496, w29497, w29498, w29499, w29500, w29501, w29502, w29503, w29504, w29505, w29506, w29507, w29508, w29509, w29510, w29511, w29512, w29513, w29514, w29515, w29516, w29517, w29518, w29519, w29520, w29521, w29522, w29523, w29524, w29525, w29526, w29527, w29528, w29529, w29530, w29531, w29532, w29533, w29534, w29535, w29536, w29537, w29538, w29539, w29540, w29541, w29542, w29543, w29544, w29545, w29546, w29547, w29548, w29549, w29550, w29551, w29552, w29553, w29554, w29555, w29556, w29557, w29558, w29559, w29560, w29561, w29562, w29563, w29564, w29565, w29566, w29567, w29568, w29569, w29570, w29571, w29572, w29573, w29574, w29575, w29576, w29577, w29578, w29579, w29580, w29581, w29582, w29583, w29584, w29585, w29586, w29587, w29588, w29589, w29590, w29591, w29592, w29593, w29594, w29595, w29596, w29597, w29598, w29599, w29600, w29601, w29602, w29603, w29604, w29605, w29606, w29607, w29608, w29609, w29610, w29611, w29612, w29613, w29614, w29615, w29616, w29617, w29618, w29619, w29620, w29621, w29622, w29623, w29624, w29625, w29626, w29627, w29628, w29629, w29630, w29631, w29632, w29633, w29634, w29635, w29636, w29637, w29638, w29639, w29640, w29641, w29642, w29643, w29644, w29645, w29646, w29647, w29648, w29649, w29650, w29651, w29652, w29653, w29654, w29655, w29656, w29657, w29658, w29659, w29660, w29661, w29662, w29663, w29664, w29665, w29666, w29667, w29668, w29669, w29670, w29671, w29672, w29673, w29674, w29675, w29676, w29677, w29678, w29679, w29680, w29681, w29682, w29683, w29684, w29685, w29686, w29687, w29688, w29689, w29690, w29691, w29692, w29693, w29694, w29695, w29696, w29697, w29698, w29699, w29700, w29701, w29702, w29703, w29704, w29705, w29706, w29707, w29708, w29709, w29710, w29711, w29712, w29713, w29714, w29715, w29716, w29717, w29718, w29719, w29720, w29721, w29722, w29723, w29724, w29725, w29726, w29727, w29728, w29729, w29730, w29731, w29732, w29733, w29734, w29735, w29736, w29737, w29738, w29739, w29740, w29741, w29742, w29743, w29744, w29745, w29746, w29747, w29748, w29749, w29750, w29751, w29752, w29753, w29754, w29755, w29756, w29757, w29758, w29759, w29760, w29761, w29762, w29763, w29764, w29765, w29766, w29767, w29768, w29769, w29770, w29771, w29772, w29773, w29774, w29775, w29776, w29777, w29778, w29779, w29780, w29781, w29782, w29783, w29784, w29785, w29786, w29787, w29788, w29789, w29790, w29791, w29792, w29793, w29794, w29795, w29796, w29797, w29798, w29799, w29800, w29801, w29802, w29803, w29804, w29805, w29806, w29807, w29808, w29809, w29810, w29811, w29812, w29813, w29814, w29815, w29816, w29817, w29818, w29819, w29820, w29821, w29822, w29823, w29824, w29825, w29826, w29827, w29828, w29829, w29830, w29831, w29832, w29833, w29834, w29835, w29836, w29837, w29838, w29839, w29840, w29841, w29842, w29843, w29844, w29845, w29846, w29847, w29848, w29849, w29850, w29851, w29852, w29853, w29854, w29855, w29856, w29857, w29858, w29859, w29860, w29861, w29862, w29863, w29864, w29865, w29866, w29867, w29868, w29869, w29870, w29871, w29872, w29873, w29874, w29875, w29876, w29877, w29878, w29879, w29880, w29881, w29882, w29883, w29884, w29885, w29886, w29887, w29888, w29889, w29890, w29891, w29892, w29893, w29894, w29895, w29896, w29897, w29898, w29899, w29900, w29901, w29902, w29903, w29904, w29905, w29906, w29907, w29908, w29909, w29910, w29911, w29912, w29913, w29914, w29915, w29916, w29917, w29918, w29919, w29920, w29921, w29922, w29923, w29924, w29925, w29926, w29927, w29928, w29929, w29930, w29931, w29932, w29933, w29934, w29935, w29936, w29937, w29938, w29939, w29940, w29941, w29942, w29943, w29944, w29945, w29946, w29947, w29948, w29949, w29950, w29951, w29952, w29953, w29954, w29955, w29956, w29957, w29958, w29959, w29960, w29961, w29962, w29963, w29964, w29965, w29966, w29967, w29968, w29969, w29970, w29971, w29972, w29973, w29974, w29975, w29976, w29977, w29978, w29979, w29980, w29981, w29982, w29983, w29984, w29985, w29986, w29987, w29988, w29989, w29990, w29991, w29992, w29993, w29994, w29995, w29996, w29997, w29998, w29999, w30000, w30001, w30002, w30003, w30004, w30005, w30006, w30007, w30008, w30009, w30010, w30011, w30012, w30013, w30014, w30015, w30016, w30017, w30018, w30019, w30020, w30021, w30022, w30023, w30024, w30025, w30026, w30027, w30028, w30029, w30030, w30031, w30032, w30033, w30034, w30035, w30036, w30037, w30038, w30039, w30040, w30041, w30042, w30043, w30044, w30045, w30046, w30047, w30048, w30049, w30050, w30051, w30052, w30053, w30054, w30055, w30056, w30057, w30058, w30059, w30060, w30061, w30062, w30063, w30064, w30065, w30066, w30067, w30068, w30069, w30070, w30071, w30072, w30073, w30074, w30075, w30076, w30077, w30078, w30079, w30080, w30081, w30082, w30083, w30084, w30085, w30086, w30087, w30088, w30089, w30090, w30091, w30092, w30093, w30094, w30095, w30096, w30097, w30098, w30099, w30100, w30101, w30102, w30103, w30104, w30105, w30106, w30107, w30108, w30109, w30110, w30111, w30112, w30113, w30114, w30115, w30116, w30117, w30118, w30119, w30120, w30121, w30122, w30123, w30124, w30125, w30126, w30127, w30128, w30129, w30130, w30131, w30132, w30133, w30134, w30135, w30136, w30137, w30138, w30139, w30140, w30141, w30142, w30143, w30144, w30145, w30146, w30147, w30148, w30149, w30150, w30151, w30152, w30153, w30154, w30155, w30156, w30157, w30158, w30159, w30160, w30161, w30162, w30163, w30164, w30165, w30166, w30167, w30168, w30169, w30170, w30171, w30172, w30173, w30174, w30175, w30176, w30177, w30178, w30179, w30180, w30181, w30182, w30183, w30184, w30185, w30186, w30187, w30188, w30189, w30190, w30191, w30192, w30193, w30194, w30195, w30196, w30197, w30198, w30199, w30200, w30201, w30202, w30203, w30204, w30205, w30206, w30207, w30208, w30209, w30210, w30211, w30212, w30213, w30214, w30215, w30216, w30217, w30218, w30219, w30220, w30221, w30222, w30223, w30224, w30225, w30226, w30227, w30228, w30229, w30230, w30231, w30232, w30233, w30234, w30235, w30236, w30237, w30238, w30239, w30240, w30241, w30242, w30243, w30244, w30245, w30246, w30247, w30248, w30249, w30250, w30251, w30252, w30253, w30254, w30255, w30256, w30257, w30258, w30259, w30260, w30261, w30262, w30263, w30264, w30265, w30266, w30267, w30268, w30269, w30270, w30271, w30272, w30273, w30274, w30275, w30276, w30277, w30278, w30279, w30280, w30281, w30282, w30283, w30284, w30285, w30286, w30287, w30288, w30289, w30290, w30291, w30292, w30293, w30294, w30295, w30296, w30297, w30298, w30299, w30300, w30301, w30302, w30303, w30304, w30305, w30306, w30307, w30308, w30309, w30310, w30311, w30312, w30313, w30314, w30315, w30316, w30317, w30318, w30319, w30320, w30321, w30322, w30323, w30324, w30325, w30326, w30327, w30328, w30329, w30330, w30331, w30332, w30333, w30334, w30335, w30336, w30337, w30338, w30339, w30340, w30341, w30342, w30343, w30344, w30345, w30346, w30347, w30348, w30349, w30350, w30351, w30352, w30353, w30354, w30355, w30356, w30357, w30358, w30359, w30360, w30361, w30362, w30363, w30364, w30365, w30366, w30367, w30368, w30369, w30370, w30371, w30372, w30373, w30374, w30375, w30376, w30377, w30378, w30379, w30380, w30381, w30382, w30383, w30384, w30385, w30386, w30387, w30388, w30389, w30390, w30391, w30392, w30393, w30394, w30395, w30396, w30397, w30398, w30399, w30400, w30401, w30402, w30403, w30404, w30405, w30406, w30407, w30408, w30409, w30410, w30411, w30412, w30413, w30414, w30415, w30416, w30417, w30418, w30419, w30420, w30421, w30422, w30423, w30424, w30425, w30426, w30427, w30428, w30429, w30430, w30431, w30432, w30433, w30434, w30435, w30436, w30437, w30438, w30439, w30440, w30441, w30442, w30443, w30444, w30445, w30446, w30447, w30448, w30449, w30450, w30451, w30452, w30453, w30454, w30455, w30456, w30457, w30458, w30459, w30460, w30461, w30462, w30463, w30464, w30465, w30466, w30467, w30468, w30469, w30470, w30471, w30472, w30473, w30474, w30475, w30476, w30477, w30478, w30479, w30480, w30481, w30482, w30483, w30484, w30485, w30486, w30487, w30488, w30489, w30490, w30491, w30492, w30493, w30494, w30495, w30496, w30497, w30498, w30499, w30500, w30501, w30502, w30503, w30504, w30505, w30506, w30507, w30508, w30509, w30510, w30511, w30512, w30513, w30514, w30515, w30516, w30517, w30518, w30519, w30520, w30521, w30522, w30523, w30524, w30525, w30526, w30527, w30528, w30529, w30530, w30531, w30532, w30533, w30534, w30535, w30536, w30537, w30538, w30539, w30540, w30541, w30542, w30543, w30544, w30545, w30546, w30547, w30548, w30549, w30550, w30551, w30552, w30553, w30554, w30555, w30556, w30557, w30558, w30559, w30560, w30561, w30562, w30563, w30564, w30565, w30566, w30567, w30568, w30569, w30570, w30571, w30572, w30573, w30574, w30575, w30576, w30577, w30578, w30579, w30580, w30581, w30582, w30583, w30584, w30585, w30586, w30587, w30588, w30589, w30590, w30591, w30592, w30593, w30594, w30595, w30596, w30597, w30598, w30599, w30600, w30601, w30602, w30603, w30604, w30605, w30606, w30607, w30608, w30609, w30610, w30611, w30612, w30613, w30614, w30615, w30616, w30617, w30618, w30619, w30620, w30621, w30622, w30623, w30624, w30625, w30626, w30627, w30628, w30629, w30630, w30631, w30632, w30633, w30634, w30635, w30636, w30637, w30638, w30639, w30640, w30641, w30642, w30643, w30644, w30645, w30646, w30647, w30648, w30649, w30650, w30651, w30652, w30653, w30654, w30655, w30656, w30657, w30658, w30659, w30660, w30661, w30662, w30663, w30664, w30665, w30666, w30667, w30668, w30669, w30670, w30671, w30672, w30673, w30674, w30675, w30676, w30677, w30678, w30679, w30680, w30681, w30682, w30683, w30684, w30685, w30686, w30687, w30688, w30689, w30690, w30691, w30692, w30693, w30694, w30695, w30696, w30697, w30698, w30699, w30700, w30701, w30702, w30703, w30704, w30705, w30706, w30707, w30708, w30709, w30710, w30711, w30712, w30713, w30714, w30715, w30716, w30717, w30718, w30719, w30720, w30721, w30722, w30723, w30724, w30725, w30726, w30727, w30728, w30729, w30730, w30731, w30732, w30733, w30734, w30735, w30736, w30737, w30738, w30739, w30740, w30741, w30742, w30743, w30744, w30745, w30746, w30747, w30748, w30749, w30750, w30751, w30752, w30753, w30754, w30755, w30756, w30757, w30758, w30759, w30760, w30761, w30762, w30763, w30764, w30765, w30766, w30767, w30768, w30769, w30770, w30771, w30772, w30773, w30774, w30775, w30776, w30777, w30778, w30779, w30780, w30781, w30782, w30783, w30784, w30785, w30786, w30787, w30788, w30789, w30790, w30791, w30792, w30793, w30794, w30795, w30796, w30797, w30798, w30799, w30800, w30801, w30802, w30803, w30804, w30805, w30806, w30807, w30808, w30809, w30810, w30811, w30812, w30813, w30814, w30815, w30816, w30817, w30818, w30819, w30820, w30821, w30822, w30823, w30824, w30825, w30826, w30827, w30828, w30829, w30830, w30831, w30832, w30833, w30834, w30835, w30836, w30837, w30838, w30839, w30840, w30841, w30842, w30843, w30844, w30845, w30846, w30847, w30848, w30849, w30850, w30851, w30852, w30853, w30854, w30855, w30856, w30857, w30858, w30859, w30860, w30861, w30862, w30863, w30864, w30865, w30866, w30867, w30868, w30869, w30870, w30871, w30872, w30873, w30874, w30875, w30876, w30877, w30878, w30879, w30880, w30881, w30882, w30883, w30884, w30885, w30886, w30887, w30888, w30889, w30890, w30891, w30892, w30893, w30894, w30895, w30896, w30897, w30898, w30899, w30900, w30901, w30902, w30903, w30904, w30905, w30906, w30907, w30908, w30909, w30910, w30911, w30912, w30913, w30914, w30915, w30916, w30917, w30918, w30919, w30920, w30921, w30922, w30923, w30924, w30925, w30926, w30927, w30928, w30929, w30930, w30931, w30932, w30933, w30934, w30935, w30936, w30937, w30938, w30939, w30940, w30941, w30942, w30943, w30944, w30945, w30946, w30947, w30948, w30949, w30950, w30951, w30952, w30953, w30954, w30955, w30956, w30957, w30958, w30959, w30960, w30961, w30962, w30963, w30964, w30965, w30966, w30967, w30968, w30969, w30970, w30971, w30972, w30973, w30974, w30975, w30976, w30977, w30978, w30979, w30980, w30981, w30982, w30983, w30984, w30985, w30986, w30987, w30988, w30989, w30990, w30991, w30992, w30993, w30994, w30995, w30996, w30997, w30998, w30999, w31000, w31001, w31002, w31003, w31004, w31005, w31006, w31007, w31008, w31009, w31010, w31011, w31012, w31013, w31014, w31015, w31016, w31017, w31018, w31019, w31020, w31021, w31022, w31023, w31024, w31025, w31026, w31027, w31028, w31029, w31030, w31031, w31032, w31033, w31034, w31035, w31036, w31037, w31038, w31039, w31040, w31041, w31042, w31043, w31044, w31045, w31046, w31047, w31048, w31049, w31050, w31051, w31052, w31053, w31054, w31055, w31056, w31057, w31058, w31059, w31060, w31061, w31062, w31063, w31064, w31065, w31066, w31067, w31068, w31069, w31070, w31071, w31072, w31073, w31074, w31075, w31076, w31077, w31078, w31079, w31080, w31081, w31082, w31083, w31084, w31085, w31086, w31087, w31088, w31089, w31090, w31091, w31092, w31093, w31094, w31095, w31096, w31097, w31098, w31099, w31100, w31101, w31102, w31103, w31104, w31105, w31106, w31107, w31108, w31109, w31110, w31111, w31112, w31113, w31114, w31115, w31116, w31117, w31118, w31119, w31120, w31121, w31122, w31123, w31124, w31125, w31126, w31127, w31128, w31129, w31130, w31131, w31132, w31133, w31134, w31135, w31136, w31137, w31138, w31139, w31140, w31141, w31142, w31143, w31144, w31145, w31146, w31147, w31148, w31149, w31150, w31151, w31152, w31153, w31154, w31155, w31156, w31157, w31158, w31159, w31160, w31161, w31162, w31163, w31164, w31165, w31166, w31167, w31168, w31169, w31170, w31171, w31172, w31173, w31174, w31175, w31176, w31177, w31178, w31179, w31180, w31181, w31182, w31183, w31184, w31185, w31186, w31187, w31188, w31189, w31190, w31191, w31192, w31193, w31194, w31195, w31196, w31197, w31198, w31199, w31200, w31201, w31202, w31203, w31204, w31205, w31206, w31207, w31208, w31209, w31210, w31211, w31212, w31213, w31214, w31215, w31216, w31217, w31218, w31219, w31220, w31221, w31222, w31223, w31224, w31225, w31226, w31227, w31228, w31229, w31230, w31231, w31232, w31233, w31234, w31235, w31236, w31237, w31238, w31239, w31240, w31241, w31242, w31243, w31244, w31245, w31246, w31247, w31248, w31249, w31250, w31251, w31252, w31253, w31254, w31255, w31256, w31257, w31258, w31259, w31260, w31261, w31262, w31263, w31264, w31265, w31266, w31267, w31268, w31269, w31270, w31271, w31272, w31273, w31274, w31275, w31276, w31277, w31278, w31279, w31280, w31281, w31282, w31283, w31284, w31285, w31286, w31287, w31288, w31289, w31290, w31291, w31292, w31293, w31294, w31295, w31296, w31297, w31298, w31299, w31300, w31301, w31302, w31303, w31304, w31305, w31306, w31307, w31308, w31309, w31310, w31311, w31312, w31313, w31314, w31315, w31316, w31317, w31318, w31319, w31320, w31321, w31322, w31323, w31324, w31325, w31326, w31327, w31328, w31329, w31330, w31331, w31332, w31333, w31334, w31335, w31336, w31337, w31338, w31339, w31340, w31341, w31342, w31343, w31344, w31345, w31346, w31347, w31348, w31349, w31350, w31351, w31352, w31353, w31354, w31355, w31356, w31357, w31358, w31359, w31360, w31361, w31362, w31363, w31364, w31365, w31366, w31367, w31368, w31369, w31370, w31371, w31372, w31373, w31374, w31375, w31376, w31377, w31378, w31379, w31380, w31381, w31382, w31383, w31384, w31385, w31386, w31387, w31388, w31389, w31390, w31391, w31392, w31393, w31394, w31395, w31396, w31397, w31398, w31399, w31400, w31401, w31402, w31403, w31404, w31405, w31406, w31407, w31408, w31409, w31410, w31411, w31412, w31413, w31414, w31415, w31416, w31417, w31418, w31419, w31420, w31421, w31422, w31423, w31424, w31425, w31426, w31427, w31428, w31429, w31430, w31431, w31432, w31433, w31434, w31435, w31436, w31437, w31438, w31439, w31440, w31441, w31442, w31443, w31444, w31445, w31446, w31447, w31448, w31449, w31450, w31451, w31452, w31453, w31454, w31455, w31456, w31457, w31458, w31459, w31460, w31461, w31462, w31463, w31464, w31465, w31466, w31467, w31468, w31469, w31470, w31471, w31472, w31473, w31474, w31475, w31476, w31477, w31478, w31479, w31480, w31481, w31482, w31483, w31484, w31485, w31486, w31487, w31488, w31489, w31490, w31491, w31492, w31493, w31494, w31495, w31496, w31497, w31498, w31499, w31500, w31501, w31502, w31503, w31504, w31505, w31506, w31507, w31508, w31509, w31510, w31511, w31512, w31513, w31514, w31515, w31516, w31517, w31518, w31519, w31520, w31521, w31522, w31523, w31524, w31525, w31526, w31527, w31528, w31529, w31530, w31531, w31532, w31533, w31534, w31535, w31536, w31537, w31538, w31539, w31540, w31541, w31542, w31543, w31544, w31545, w31546, w31547, w31548, w31549, w31550, w31551, w31552, w31553, w31554, w31555, w31556, w31557, w31558, w31559, w31560, w31561, w31562, w31563, w31564, w31565, w31566, w31567, w31568, w31569, w31570, w31571, w31572, w31573, w31574, w31575, w31576, w31577, w31578, w31579, w31580, w31581, w31582, w31583, w31584, w31585, w31586, w31587, w31588, w31589, w31590, w31591, w31592, w31593, w31594, w31595, w31596, w31597, w31598, w31599, w31600, w31601, w31602, w31603, w31604, w31605, w31606, w31607, w31608, w31609, w31610, w31611, w31612, w31613, w31614, w31615, w31616, w31617, w31618, w31619, w31620, w31621, w31622, w31623, w31624, w31625, w31626, w31627, w31628, w31629, w31630, w31631, w31632, w31633, w31634, w31635, w31636, w31637, w31638, w31639, w31640, w31641, w31642, w31643, w31644, w31645, w31646, w31647, w31648, w31649, w31650, w31651, w31652, w31653, w31654, w31655, w31656, w31657, w31658, w31659, w31660, w31661, w31662, w31663, w31664, w31665, w31666, w31667, w31668, w31669, w31670, w31671, w31672, w31673, w31674, w31675, w31676, w31677, w31678, w31679, w31680, w31681, w31682, w31683, w31684, w31685, w31686, w31687, w31688, w31689, w31690, w31691, w31692, w31693, w31694, w31695, w31696, w31697, w31698, w31699, w31700, w31701, w31702, w31703, w31704, w31705, w31706, w31707, w31708, w31709, w31710, w31711, w31712, w31713, w31714, w31715, w31716, w31717, w31718, w31719, w31720, w31721, w31722, w31723, w31724, w31725, w31726, w31727, w31728, w31729, w31730, w31731, w31732, w31733, w31734, w31735, w31736, w31737, w31738, w31739, w31740, w31741, w31742, w31743, w31744, w31745, w31746, w31747, w31748, w31749, w31750, w31751, w31752, w31753, w31754, w31755, w31756, w31757, w31758, w31759, w31760, w31761, w31762, w31763, w31764, w31765, w31766, w31767, w31768, w31769, w31770, w31771, w31772, w31773, w31774, w31775, w31776, w31777, w31778, w31779, w31780, w31781, w31782, w31783, w31784, w31785, w31786, w31787, w31788, w31789, w31790, w31791, w31792, w31793, w31794, w31795, w31796, w31797, w31798, w31799, w31800, w31801, w31802, w31803, w31804, w31805, w31806, w31807, w31808, w31809, w31810, w31811, w31812, w31813, w31814, w31815, w31816, w31817, w31818, w31819, w31820, w31821, w31822, w31823, w31824, w31825, w31826, w31827, w31828, w31829, w31830, w31831, w31832, w31833, w31834, w31835, w31836, w31837, w31838, w31839, w31840, w31841, w31842, w31843, w31844, w31845, w31846, w31847, w31848, w31849, w31850, w31851, w31852, w31853, w31854, w31855, w31856, w31857, w31858, w31859, w31860, w31861, w31862, w31863, w31864, w31865, w31866, w31867, w31868, w31869, w31870, w31871, w31872, w31873, w31874, w31875, w31876, w31877, w31878, w31879, w31880, w31881, w31882, w31883, w31884, w31885, w31886, w31887, w31888, w31889, w31890, w31891, w31892, w31893, w31894, w31895, w31896, w31897, w31898, w31899, w31900, w31901, w31902, w31903, w31904, w31905, w31906, w31907, w31908, w31909, w31910, w31911, w31912, w31913, w31914, w31915, w31916, w31917, w31918, w31919, w31920, w31921, w31922, w31923, w31924, w31925, w31926, w31927, w31928, w31929, w31930, w31931, w31932, w31933, w31934, w31935, w31936, w31937, w31938, w31939, w31940, w31941, w31942, w31943, w31944, w31945, w31946, w31947, w31948, w31949, w31950, w31951, w31952, w31953, w31954, w31955, w31956, w31957, w31958, w31959, w31960, w31961, w31962, w31963, w31964, w31965, w31966, w31967, w31968, w31969, w31970, w31971, w31972, w31973, w31974, w31975, w31976, w31977, w31978, w31979, w31980, w31981, w31982, w31983, w31984, w31985, w31986, w31987, w31988, w31989, w31990, w31991, w31992, w31993, w31994, w31995, w31996, w31997, w31998, w31999, w32000, w32001, w32002, w32003, w32004, w32005, w32006, w32007, w32008, w32009, w32010, w32011, w32012, w32013, w32014, w32015, w32016, w32017, w32018, w32019, w32020, w32021, w32022, w32023, w32024, w32025, w32026, w32027, w32028, w32029, w32030, w32031, w32032, w32033, w32034, w32035, w32036, w32037, w32038, w32039, w32040, w32041, w32042, w32043, w32044, w32045, w32046, w32047, w32048, w32049, w32050, w32051, w32052, w32053, w32054, w32055, w32056, w32057, w32058, w32059, w32060, w32061, w32062, w32063, w32064, w32065, w32066, w32067, w32068, w32069, w32070, w32071, w32072, w32073, w32074, w32075, w32076, w32077, w32078, w32079, w32080, w32081, w32082, w32083, w32084, w32085, w32086, w32087, w32088, w32089, w32090, w32091, w32092, w32093, w32094, w32095, w32096, w32097, w32098, w32099, w32100, w32101, w32102, w32103, w32104, w32105, w32106, w32107, w32108, w32109, w32110, w32111, w32112, w32113, w32114, w32115, w32116, w32117, w32118, w32119, w32120, w32121, w32122, w32123, w32124, w32125, w32126, w32127, w32128, w32129, w32130, w32131, w32132, w32133, w32134, w32135, w32136, w32137, w32138, w32139, w32140, w32141, w32142, w32143, w32144, w32145, w32146, w32147, w32148, w32149, w32150, w32151, w32152, w32153, w32154, w32155, w32156, w32157, w32158, w32159, w32160, w32161, w32162, w32163, w32164, w32165, w32166, w32167, w32168, w32169, w32170, w32171, w32172, w32173, w32174, w32175, w32176, w32177, w32178, w32179, w32180, w32181, w32182, w32183, w32184, w32185, w32186, w32187, w32188, w32189, w32190, w32191, w32192, w32193, w32194, w32195, w32196, w32197, w32198, w32199, w32200, w32201, w32202, w32203, w32204, w32205, w32206, w32207, w32208, w32209, w32210, w32211, w32212, w32213, w32214, w32215, w32216, w32217, w32218, w32219, w32220, w32221, w32222, w32223, w32224, w32225, w32226, w32227, w32228, w32229, w32230, w32231, w32232, w32233, w32234, w32235, w32236, w32237, w32238, w32239, w32240, w32241, w32242, w32243, w32244, w32245, w32246, w32247, w32248, w32249, w32250, w32251, w32252, w32253, w32254, w32255, w32256, w32257, w32258, w32259, w32260, w32261, w32262, w32263, w32264, w32265, w32266, w32267, w32268, w32269, w32270, w32271, w32272, w32273, w32274, w32275, w32276, w32277, w32278, w32279, w32280, w32281, w32282, w32283, w32284, w32285, w32286, w32287, w32288, w32289, w32290, w32291, w32292, w32293, w32294, w32295, w32296, w32297, w32298, w32299, w32300, w32301, w32302, w32303, w32304, w32305, w32306, w32307, w32308, w32309, w32310, w32311, w32312, w32313, w32314, w32315, w32316, w32317, w32318, w32319, w32320, w32321, w32322, w32323, w32324, w32325, w32326, w32327, w32328, w32329, w32330, w32331, w32332, w32333, w32334, w32335, w32336, w32337, w32338, w32339, w32340, w32341, w32342, w32343, w32344, w32345, w32346, w32347, w32348, w32349, w32350, w32351, w32352, w32353, w32354, w32355, w32356, w32357, w32358, w32359, w32360, w32361, w32362, w32363, w32364, w32365, w32366, w32367, w32368, w32369, w32370, w32371, w32372, w32373, w32374, w32375, w32376, w32377, w32378, w32379, w32380, w32381, w32382, w32383, w32384, w32385, w32386, w32387, w32388, w32389, w32390, w32391, w32392, w32393, w32394, w32395, w32396, w32397, w32398, w32399, w32400, w32401, w32402, w32403, w32404, w32405, w32406, w32407, w32408, w32409, w32410, w32411, w32412, w32413, w32414, w32415, w32416, w32417, w32418, w32419, w32420, w32421, w32422, w32423, w32424, w32425, w32426, w32427, w32428, w32429, w32430, w32431, w32432, w32433, w32434, w32435, w32436, w32437, w32438, w32439, w32440, w32441, w32442, w32443, w32444, w32445, w32446, w32447, w32448, w32449, w32450, w32451, w32452, w32453, w32454, w32455, w32456, w32457, w32458, w32459, w32460, w32461, w32462, w32463, w32464, w32465, w32466, w32467, w32468, w32469, w32470, w32471, w32472, w32473, w32474, w32475, w32476, w32477, w32478, w32479, w32480, w32481, w32482, w32483, w32484, w32485, w32486, w32487, w32488, w32489, w32490, w32491, w32492, w32493, w32494, w32495, w32496, w32497, w32498, w32499, w32500, w32501, w32502, w32503, w32504, w32505, w32506, w32507, w32508, w32509, w32510, w32511, w32512, w32513, w32514, w32515, w32516, w32517, w32518, w32519, w32520, w32521, w32522, w32523, w32524, w32525, w32526, w32527, w32528, w32529, w32530, w32531, w32532, w32533, w32534, w32535, w32536, w32537, w32538, w32539, w32540, w32541, w32542, w32543, w32544, w32545, w32546, w32547, w32548, w32549, w32550, w32551, w32552, w32553, w32554, w32555, w32556, w32557, w32558, w32559, w32560, w32561, w32562, w32563, w32564, w32565, w32566, w32567, w32568, w32569, w32570, w32571, w32572, w32573, w32574, w32575, w32576, w32577, w32578, w32579, w32580, w32581, w32582, w32583, w32584, w32585, w32586, w32587, w32588, w32589, w32590, w32591, w32592, w32593, w32594, w32595, w32596, w32597, w32598, w32599, w32600, w32601, w32602, w32603, w32604, w32605, w32606, w32607, w32608, w32609, w32610, w32611, w32612, w32613, w32614, w32615, w32616, w32617, w32618, w32619, w32620, w32621, w32622, w32623, w32624, w32625, w32626, w32627, w32628, w32629, w32630, w32631, w32632, w32633, w32634, w32635, w32636, w32637, w32638, w32639, w32640, w32641, w32642, w32643, w32644, w32645, w32646, w32647, w32648, w32649, w32650, w32651, w32652, w32653, w32654, w32655, w32656, w32657, w32658, w32659, w32660, w32661, w32662, w32663, w32664, w32665, w32666, w32667, w32668, w32669, w32670, w32671, w32672, w32673, w32674, w32675, w32676, w32677, w32678, w32679, w32680, w32681, w32682, w32683, w32684, w32685, w32686, w32687, w32688, w32689, w32690, w32691, w32692, w32693, w32694, w32695, w32696, w32697, w32698, w32699, w32700, w32701, w32702, w32703, w32704, w32705, w32706, w32707, w32708, w32709, w32710, w32711, w32712, w32713, w32714, w32715, w32716, w32717, w32718, w32719, w32720, w32721, w32722, w32723, w32724, w32725, w32726, w32727, w32728, w32729, w32730, w32731, w32732, w32733, w32734, w32735, w32736, w32737, w32738, w32739, w32740, w32741, w32742, w32743, w32744, w32745, w32746, w32747, w32748, w32749, w32750, w32751, w32752, w32753, w32754, w32755, w32756, w32757, w32758, w32759, w32760, w32761, w32762, w32763, w32764, w32765, w32766, w32767, w32768, w32769, w32770, w32771, w32772, w32773, w32774, w32775, w32776, w32777, w32778, w32779, w32780, w32781, w32782, w32783, w32784, w32785, w32786, w32787, w32788, w32789, w32790, w32791, w32792, w32793, w32794, w32795, w32796, w32797, w32798, w32799, w32800, w32801, w32802, w32803, w32804, w32805, w32806, w32807, w32808, w32809, w32810, w32811, w32812, w32813, w32814, w32815, w32816, w32817, w32818, w32819, w32820, w32821, w32822, w32823, w32824, w32825, w32826, w32827, w32828, w32829, w32830, w32831, w32832, w32833, w32834, w32835, w32836, w32837, w32838, w32839, w32840, w32841, w32842, w32843, w32844, w32845, w32846, w32847, w32848, w32849, w32850, w32851, w32852, w32853, w32854, w32855, w32856, w32857, w32858, w32859, w32860, w32861, w32862, w32863, w32864, w32865, w32866, w32867, w32868, w32869, w32870, w32871, w32872, w32873, w32874, w32875, w32876, w32877, w32878, w32879, w32880, w32881, w32882, w32883, w32884, w32885, w32886, w32887, w32888, w32889, w32890, w32891, w32892, w32893, w32894, w32895, w32896, w32897, w32898, w32899, w32900, w32901, w32902, w32903, w32904, w32905, w32906, w32907, w32908, w32909, w32910, w32911, w32912, w32913, w32914, w32915, w32916, w32917, w32918, w32919, w32920, w32921, w32922, w32923, w32924, w32925, w32926, w32927, w32928, w32929, w32930, w32931, w32932, w32933, w32934, w32935, w32936, w32937, w32938, w32939, w32940, w32941, w32942, w32943, w32944, w32945, w32946, w32947, w32948, w32949, w32950, w32951, w32952, w32953, w32954, w32955, w32956, w32957, w32958, w32959, w32960, w32961, w32962, w32963, w32964, w32965, w32966, w32967, w32968, w32969, w32970, w32971, w32972, w32973, w32974, w32975, w32976, w32977, w32978, w32979, w32980, w32981, w32982, w32983, w32984, w32985, w32986, w32987, w32988, w32989, w32990, w32991, w32992, w32993, w32994, w32995, w32996, w32997, w32998, w32999, w33000, w33001, w33002, w33003, w33004, w33005, w33006, w33007, w33008, w33009, w33010, w33011, w33012, w33013, w33014, w33015, w33016, w33017, w33018, w33019, w33020, w33021, w33022, w33023, w33024, w33025, w33026, w33027, w33028, w33029, w33030, w33031, w33032, w33033, w33034, w33035, w33036, w33037, w33038, w33039, w33040, w33041, w33042, w33043, w33044, w33045, w33046, w33047, w33048, w33049, w33050, w33051, w33052, w33053, w33054, w33055, w33056, w33057, w33058, w33059, w33060, w33061, w33062, w33063, w33064, w33065, w33066, w33067, w33068, w33069, w33070, w33071, w33072, w33073, w33074, w33075, w33076, w33077, w33078, w33079, w33080, w33081, w33082, w33083, w33084, w33085, w33086, w33087, w33088, w33089, w33090, w33091, w33092, w33093, w33094, w33095, w33096, w33097, w33098, w33099, w33100, w33101, w33102, w33103, w33104, w33105, w33106, w33107, w33108, w33109, w33110, w33111, w33112, w33113, w33114, w33115, w33116, w33117, w33118, w33119, w33120, w33121, w33122, w33123, w33124, w33125, w33126, w33127, w33128, w33129, w33130, w33131, w33132, w33133, w33134, w33135, w33136, w33137, w33138, w33139, w33140, w33141, w33142, w33143, w33144, w33145, w33146, w33147, w33148, w33149, w33150, w33151, w33152, w33153, w33154, w33155, w33156, w33157, w33158, w33159, w33160, w33161, w33162, w33163, w33164, w33165, w33166, w33167, w33168, w33169, w33170, w33171, w33172, w33173, w33174, w33175, w33176, w33177, w33178, w33179, w33180, w33181, w33182, w33183, w33184, w33185, w33186, w33187, w33188, w33189, w33190, w33191, w33192, w33193, w33194, w33195, w33196, w33197, w33198, w33199, w33200, w33201, w33202, w33203, w33204, w33205, w33206, w33207, w33208, w33209, w33210, w33211, w33212, w33213, w33214, w33215, w33216, w33217, w33218, w33219, w33220, w33221, w33222, w33223, w33224, w33225, w33226, w33227, w33228, w33229, w33230, w33231, w33232, w33233, w33234, w33235, w33236, w33237, w33238, w33239, w33240, w33241, w33242, w33243, w33244, w33245, w33246, w33247, w33248, w33249, w33250, w33251, w33252, w33253, w33254, w33255, w33256, w33257, w33258, w33259, w33260, w33261, w33262, w33263, w33264, w33265, w33266, w33267, w33268, w33269, w33270, w33271, w33272, w33273, w33274, w33275, w33276, w33277, w33278, w33279, w33280, w33281, w33282, w33283, w33284, w33285, w33286, w33287, w33288, w33289, w33290, w33291, w33292, w33293, w33294, w33295, w33296, w33297, w33298, w33299, w33300, w33301, w33302, w33303, w33304, w33305, w33306, w33307, w33308, w33309, w33310, w33311, w33312, w33313, w33314, w33315, w33316, w33317, w33318, w33319, w33320, w33321, w33322, w33323, w33324, w33325, w33326, w33327, w33328, w33329, w33330, w33331, w33332, w33333, w33334, w33335, w33336, w33337, w33338, w33339, w33340, w33341, w33342, w33343, w33344, w33345, w33346, w33347, w33348, w33349, w33350, w33351, w33352, w33353, w33354, w33355, w33356, w33357, w33358, w33359, w33360, w33361, w33362, w33363, w33364, w33365, w33366, w33367, w33368, w33369, w33370, w33371, w33372, w33373, w33374, w33375, w33376, w33377, w33378, w33379, w33380, w33381, w33382, w33383, w33384, w33385, w33386, w33387, w33388, w33389, w33390, w33391, w33392, w33393, w33394, w33395, w33396, w33397, w33398, w33399, w33400, w33401, w33402, w33403, w33404, w33405, w33406, w33407, w33408, w33409, w33410, w33411, w33412, w33413, w33414, w33415, w33416, w33417, w33418, w33419, w33420, w33421, w33422, w33423, w33424, w33425, w33426, w33427, w33428, w33429, w33430, w33431, w33432, w33433, w33434, w33435, w33436, w33437, w33438, w33439, w33440, w33441, w33442, w33443, w33444, w33445, w33446, w33447, w33448, w33449, w33450, w33451, w33452, w33453, w33454, w33455, w33456, w33457, w33458, w33459, w33460, w33461, w33462, w33463, w33464, w33465, w33466, w33467, w33468, w33469, w33470, w33471, w33472, w33473, w33474, w33475, w33476, w33477, w33478, w33479, w33480, w33481, w33482, w33483, w33484, w33485, w33486, w33487, w33488, w33489, w33490, w33491, w33492, w33493, w33494, w33495, w33496, w33497, w33498, w33499, w33500, w33501, w33502, w33503, w33504, w33505, w33506, w33507, w33508, w33509, w33510, w33511, w33512, w33513, w33514, w33515, w33516, w33517, w33518, w33519, w33520, w33521, w33522, w33523, w33524, w33525, w33526, w33527, w33528, w33529, w33530, w33531, w33532, w33533, w33534, w33535, w33536, w33537, w33538, w33539, w33540, w33541, w33542, w33543, w33544, w33545, w33546, w33547, w33548, w33549, w33550, w33551, w33552, w33553, w33554, w33555, w33556, w33557, w33558, w33559, w33560, w33561, w33562, w33563, w33564, w33565, w33566, w33567, w33568, w33569, w33570, w33571, w33572, w33573, w33574, w33575, w33576, w33577, w33578, w33579, w33580, w33581, w33582, w33583, w33584, w33585, w33586, w33587, w33588, w33589, w33590, w33591, w33592, w33593, w33594, w33595, w33596, w33597, w33598, w33599, w33600, w33601, w33602, w33603, w33604, w33605, w33606, w33607, w33608, w33609, w33610, w33611, w33612, w33613, w33614, w33615, w33616, w33617, w33618, w33619, w33620, w33621, w33622, w33623, w33624, w33625, w33626, w33627, w33628, w33629, w33630, w33631, w33632, w33633, w33634, w33635, w33636, w33637, w33638, w33639, w33640, w33641, w33642, w33643, w33644, w33645, w33646, w33647, w33648, w33649, w33650, w33651, w33652, w33653, w33654, w33655, w33656, w33657, w33658, w33659, w33660, w33661, w33662, w33663, w33664, w33665, w33666, w33667, w33668, w33669, w33670, w33671, w33672, w33673, w33674, w33675, w33676, w33677, w33678, w33679, w33680, w33681, w33682, w33683, w33684, w33685, w33686, w33687, w33688, w33689, w33690, w33691, w33692, w33693, w33694, w33695, w33696, w33697, w33698, w33699, w33700, w33701, w33702, w33703, w33704, w33705, w33706, w33707, w33708, w33709, w33710, w33711, w33712, w33713, w33714, w33715, w33716, w33717, w33718, w33719, w33720, w33721, w33722, w33723, w33724, w33725, w33726, w33727, w33728, w33729, w33730, w33731, w33732, w33733, w33734, w33735, w33736, w33737, w33738, w33739, w33740, w33741, w33742, w33743, w33744, w33745, w33746, w33747, w33748, w33749, w33750, w33751, w33752, w33753, w33754, w33755, w33756, w33757, w33758, w33759, w33760, w33761, w33762, w33763, w33764, w33765, w33766, w33767, w33768, w33769, w33770, w33771, w33772, w33773, w33774, w33775, w33776, w33777, w33778, w33779, w33780, w33781, w33782, w33783, w33784, w33785, w33786, w33787, w33788, w33789, w33790, w33791, w33792, w33793, w33794, w33795, w33796, w33797, w33798, w33799, w33800, w33801, w33802, w33803, w33804, w33805, w33806, w33807, w33808, w33809, w33810, w33811, w33812, w33813, w33814, w33815, w33816, w33817, w33818, w33819, w33820, w33821, w33822, w33823, w33824, w33825, w33826, w33827, w33828, w33829, w33830, w33831, w33832, w33833, w33834, w33835, w33836, w33837, w33838, w33839, w33840, w33841, w33842, w33843, w33844, w33845, w33846, w33847, w33848, w33849, w33850, w33851, w33852, w33853, w33854, w33855, w33856, w33857, w33858, w33859, w33860, w33861, w33862, w33863, w33864, w33865, w33866, w33867, w33868, w33869, w33870, w33871, w33872, w33873, w33874, w33875, w33876, w33877, w33878, w33879, w33880, w33881, w33882, w33883, w33884, w33885, w33886, w33887, w33888, w33889, w33890, w33891, w33892, w33893, w33894, w33895, w33896, w33897, w33898, w33899, w33900, w33901, w33902, w33903, w33904, w33905, w33906, w33907, w33908, w33909, w33910, w33911, w33912, w33913, w33914, w33915, w33916, w33917, w33918, w33919, w33920, w33921, w33922, w33923, w33924, w33925, w33926, w33927, w33928, w33929, w33930, w33931, w33932, w33933, w33934, w33935, w33936, w33937, w33938, w33939, w33940, w33941, w33942, w33943, w33944, w33945, w33946, w33947, w33948, w33949, w33950, w33951, w33952, w33953, w33954, w33955, w33956, w33957, w33958, w33959, w33960, w33961, w33962, w33963, w33964, w33965, w33966, w33967, w33968, w33969, w33970, w33971, w33972, w33973, w33974, w33975, w33976, w33977, w33978, w33979, w33980, w33981, w33982, w33983, w33984, w33985, w33986, w33987, w33988, w33989, w33990, w33991, w33992, w33993, w33994, w33995, w33996, w33997, w33998, w33999, w34000, w34001, w34002, w34003, w34004, w34005, w34006, w34007, w34008, w34009, w34010, w34011, w34012, w34013, w34014, w34015, w34016, w34017, w34018, w34019, w34020, w34021, w34022, w34023, w34024, w34025, w34026, w34027, w34028, w34029, w34030, w34031, w34032, w34033, w34034, w34035, w34036, w34037, w34038, w34039, w34040, w34041, w34042, w34043, w34044, w34045, w34046, w34047, w34048, w34049, w34050, w34051, w34052, w34053, w34054, w34055, w34056, w34057, w34058, w34059, w34060, w34061, w34062, w34063, w34064, w34065, w34066, w34067, w34068, w34069, w34070, w34071, w34072, w34073, w34074, w34075, w34076, w34077, w34078, w34079, w34080, w34081, w34082, w34083, w34084, w34085, w34086, w34087, w34088, w34089, w34090, w34091, w34092, w34093, w34094, w34095, w34096, w34097, w34098, w34099, w34100, w34101, w34102, w34103, w34104, w34105, w34106, w34107, w34108, w34109, w34110, w34111, w34112, w34113, w34114, w34115, w34116, w34117, w34118, w34119, w34120, w34121, w34122, w34123, w34124, w34125, w34126, w34127, w34128, w34129, w34130, w34131, w34132, w34133, w34134, w34135, w34136, w34137, w34138, w34139, w34140, w34141, w34142, w34143, w34144, w34145, w34146, w34147, w34148, w34149, w34150, w34151, w34152, w34153, w34154, w34155, w34156, w34157, w34158, w34159, w34160, w34161, w34162, w34163, w34164, w34165, w34166, w34167, w34168, w34169, w34170, w34171, w34172, w34173, w34174, w34175, w34176, w34177, w34178, w34179, w34180, w34181, w34182, w34183, w34184, w34185, w34186, w34187, w34188, w34189, w34190, w34191, w34192, w34193, w34194, w34195, w34196, w34197, w34198, w34199, w34200, w34201, w34202, w34203, w34204, w34205, w34206, w34207, w34208, w34209, w34210, w34211, w34212, w34213, w34214, w34215, w34216, w34217, w34218, w34219, w34220, w34221, w34222, w34223, w34224, w34225, w34226, w34227, w34228, w34229, w34230, w34231, w34232, w34233, w34234, w34235, w34236, w34237, w34238, w34239, w34240, w34241, w34242, w34243, w34244, w34245, w34246, w34247, w34248, w34249, w34250, w34251, w34252, w34253, w34254, w34255, w34256, w34257, w34258, w34259, w34260, w34261, w34262, w34263, w34264, w34265, w34266, w34267, w34268, w34269, w34270, w34271, w34272, w34273, w34274, w34275, w34276, w34277, w34278, w34279, w34280, w34281, w34282, w34283, w34284, w34285, w34286, w34287, w34288, w34289, w34290, w34291, w34292, w34293, w34294, w34295, w34296, w34297, w34298, w34299, w34300, w34301, w34302, w34303, w34304, w34305, w34306, w34307, w34308, w34309, w34310, w34311, w34312, w34313, w34314, w34315, w34316, w34317, w34318, w34319, w34320, w34321, w34322, w34323, w34324, w34325, w34326, w34327, w34328, w34329, w34330, w34331, w34332, w34333, w34334, w34335, w34336, w34337, w34338, w34339, w34340, w34341, w34342, w34343, w34344, w34345, w34346, w34347, w34348, w34349, w34350, w34351, w34352, w34353, w34354, w34355, w34356, w34357, w34358, w34359, w34360, w34361, w34362, w34363, w34364, w34365, w34366, w34367, w34368, w34369, w34370, w34371, w34372, w34373, w34374, w34375, w34376, w34377, w34378, w34379, w34380, w34381, w34382, w34383, w34384, w34385, w34386, w34387, w34388, w34389, w34390, w34391, w34392, w34393, w34394, w34395, w34396, w34397, w34398, w34399, w34400, w34401, w34402, w34403, w34404, w34405, w34406, w34407, w34408, w34409, w34410, w34411, w34412, w34413, w34414, w34415, w34416, w34417, w34418, w34419, w34420, w34421, w34422, w34423, w34424, w34425, w34426, w34427, w34428, w34429, w34430, w34431, w34432, w34433, w34434, w34435, w34436, w34437, w34438, w34439, w34440, w34441, w34442, w34443, w34444, w34445, w34446, w34447, w34448, w34449, w34450, w34451, w34452, w34453, w34454, w34455, w34456, w34457, w34458, w34459, w34460, w34461, w34462, w34463, w34464, w34465, w34466, w34467, w34468, w34469, w34470, w34471, w34472, w34473, w34474, w34475, w34476, w34477, w34478, w34479, w34480, w34481, w34482, w34483, w34484, w34485, w34486, w34487, w34488, w34489, w34490, w34491, w34492, w34493, w34494, w34495, w34496, w34497, w34498, w34499, w34500, w34501, w34502, w34503, w34504, w34505, w34506, w34507, w34508, w34509, w34510, w34511, w34512, w34513, w34514, w34515, w34516, w34517, w34518, w34519, w34520, w34521, w34522, w34523, w34524, w34525, w34526, w34527, w34528, w34529, w34530, w34531, w34532, w34533, w34534, w34535, w34536, w34537, w34538, w34539, w34540, w34541, w34542, w34543, w34544, w34545, w34546, w34547, w34548, w34549, w34550, w34551, w34552, w34553, w34554, w34555, w34556, w34557, w34558, w34559, w34560, w34561, w34562, w34563, w34564, w34565, w34566, w34567, w34568, w34569, w34570, w34571, w34572, w34573, w34574, w34575, w34576, w34577, w34578, w34579, w34580, w34581, w34582, w34583, w34584, w34585, w34586, w34587, w34588, w34589, w34590, w34591, w34592, w34593, w34594, w34595, w34596, w34597, w34598, w34599, w34600, w34601, w34602, w34603, w34604, w34605, w34606, w34607, w34608, w34609, w34610, w34611, w34612, w34613, w34614, w34615, w34616, w34617, w34618, w34619, w34620, w34621, w34622, w34623, w34624, w34625, w34626, w34627, w34628, w34629, w34630, w34631, w34632, w34633, w34634, w34635, w34636, w34637, w34638, w34639, w34640, w34641, w34642, w34643, w34644, w34645, w34646, w34647, w34648, w34649, w34650, w34651, w34652, w34653, w34654, w34655, w34656, w34657, w34658, w34659, w34660, w34661, w34662, w34663, w34664, w34665, w34666, w34667, w34668, w34669, w34670, w34671, w34672, w34673, w34674, w34675, w34676, w34677, w34678, w34679, w34680, w34681, w34682, w34683, w34684, w34685, w34686, w34687, w34688, w34689, w34690, w34691, w34692, w34693, w34694, w34695, w34696, w34697, w34698, w34699, w34700, w34701, w34702, w34703, w34704, w34705, w34706, w34707, w34708, w34709, w34710, w34711, w34712, w34713, w34714, w34715, w34716, w34717, w34718, w34719, w34720, w34721, w34722, w34723, w34724, w34725, w34726, w34727, w34728, w34729, w34730, w34731, w34732, w34733, w34734, w34735, w34736, w34737, w34738, w34739, w34740, w34741, w34742, w34743, w34744, w34745, w34746, w34747, w34748, w34749, w34750, w34751, w34752, w34753, w34754, w34755, w34756, w34757, w34758, w34759, w34760, w34761, w34762, w34763, w34764, w34765, w34766, w34767, w34768, w34769, w34770, w34771, w34772, w34773, w34774, w34775, w34776, w34777, w34778, w34779, w34780, w34781, w34782, w34783, w34784, w34785, w34786, w34787, w34788, w34789, w34790, w34791, w34792, w34793, w34794, w34795, w34796, w34797, w34798, w34799, w34800, w34801, w34802, w34803, w34804, w34805, w34806, w34807, w34808, w34809, w34810, w34811, w34812, w34813, w34814, w34815, w34816, w34817, w34818, w34819, w34820, w34821, w34822, w34823, w34824, w34825, w34826, w34827, w34828, w34829, w34830, w34831, w34832, w34833, w34834, w34835, w34836, w34837, w34838, w34839, w34840, w34841, w34842, w34843, w34844, w34845, w34846, w34847, w34848, w34849, w34850, w34851, w34852, w34853, w34854, w34855, w34856, w34857, w34858, w34859, w34860, w34861, w34862, w34863, w34864, w34865, w34866, w34867, w34868, w34869, w34870, w34871, w34872, w34873, w34874, w34875, w34876, w34877, w34878, w34879, w34880, w34881, w34882, w34883, w34884, w34885, w34886, w34887, w34888, w34889, w34890, w34891, w34892, w34893, w34894, w34895, w34896, w34897, w34898, w34899, w34900, w34901, w34902, w34903, w34904, w34905, w34906, w34907, w34908, w34909, w34910, w34911, w34912, w34913, w34914, w34915, w34916, w34917, w34918, w34919, w34920, w34921, w34922, w34923, w34924, w34925, w34926, w34927, w34928, w34929, w34930, w34931, w34932, w34933, w34934, w34935, w34936, w34937, w34938, w34939, w34940, w34941, w34942, w34943, w34944, w34945, w34946, w34947, w34948, w34949, w34950, w34951, w34952, w34953, w34954, w34955, w34956, w34957, w34958, w34959, w34960, w34961, w34962, w34963, w34964, w34965, w34966, w34967, w34968, w34969, w34970, w34971, w34972, w34973, w34974, w34975, w34976, w34977, w34978, w34979, w34980, w34981, w34982, w34983, w34984, w34985, w34986, w34987, w34988, w34989, w34990, w34991, w34992, w34993, w34994, w34995, w34996, w34997, w34998, w34999, w35000, w35001, w35002, w35003, w35004, w35005, w35006, w35007, w35008, w35009, w35010, w35011, w35012, w35013, w35014, w35015, w35016, w35017, w35018, w35019, w35020, w35021, w35022, w35023, w35024, w35025, w35026, w35027, w35028, w35029, w35030, w35031, w35032, w35033, w35034, w35035, w35036, w35037, w35038, w35039, w35040, w35041, w35042, w35043, w35044, w35045, w35046, w35047, w35048, w35049, w35050, w35051, w35052, w35053, w35054, w35055, w35056, w35057, w35058, w35059, w35060, w35061, w35062, w35063, w35064, w35065, w35066, w35067, w35068, w35069, w35070, w35071, w35072, w35073, w35074, w35075, w35076, w35077, w35078, w35079, w35080, w35081, w35082, w35083, w35084, w35085, w35086, w35087, w35088, w35089, w35090, w35091, w35092, w35093, w35094, w35095, w35096, w35097, w35098, w35099, w35100, w35101, w35102, w35103, w35104, w35105, w35106, w35107, w35108, w35109, w35110, w35111, w35112, w35113, w35114, w35115, w35116, w35117, w35118, w35119, w35120, w35121, w35122, w35123, w35124, w35125, w35126, w35127, w35128, w35129, w35130, w35131, w35132, w35133, w35134, w35135, w35136, w35137, w35138, w35139, w35140, w35141, w35142, w35143, w35144, w35145, w35146, w35147, w35148, w35149, w35150, w35151, w35152, w35153, w35154, w35155, w35156, w35157, w35158, w35159, w35160, w35161, w35162, w35163, w35164, w35165, w35166, w35167, w35168, w35169, w35170, w35171, w35172, w35173, w35174, w35175, w35176, w35177, w35178, w35179, w35180, w35181, w35182, w35183, w35184, w35185, w35186, w35187, w35188, w35189, w35190, w35191, w35192, w35193, w35194, w35195, w35196, w35197, w35198, w35199, w35200, w35201, w35202, w35203, w35204, w35205, w35206, w35207, w35208, w35209, w35210, w35211, w35212, w35213, w35214, w35215, w35216, w35217, w35218, w35219, w35220, w35221, w35222, w35223, w35224, w35225, w35226, w35227, w35228, w35229, w35230, w35231, w35232, w35233, w35234, w35235, w35236, w35237, w35238, w35239, w35240, w35241, w35242, w35243, w35244, w35245, w35246, w35247, w35248, w35249, w35250, w35251, w35252, w35253, w35254, w35255, w35256, w35257, w35258, w35259, w35260, w35261, w35262, w35263, w35264, w35265, w35266, w35267, w35268, w35269, w35270, w35271, w35272, w35273, w35274, w35275, w35276, w35277, w35278, w35279, w35280, w35281, w35282, w35283, w35284, w35285, w35286, w35287, w35288, w35289, w35290, w35291, w35292, w35293, w35294, w35295, w35296, w35297, w35298, w35299, w35300, w35301, w35302, w35303, w35304, w35305, w35306, w35307, w35308, w35309, w35310, w35311, w35312, w35313, w35314, w35315, w35316, w35317, w35318, w35319, w35320, w35321, w35322, w35323, w35324, w35325, w35326, w35327, w35328, w35329, w35330, w35331, w35332, w35333, w35334, w35335, w35336, w35337, w35338, w35339, w35340, w35341, w35342, w35343, w35344, w35345, w35346, w35347, w35348, w35349, w35350, w35351, w35352, w35353, w35354, w35355, w35356, w35357, w35358, w35359, w35360, w35361, w35362, w35363, w35364, w35365, w35366, w35367, w35368, w35369, w35370, w35371, w35372, w35373, w35374, w35375, w35376, w35377, w35378, w35379, w35380, w35381, w35382, w35383, w35384, w35385, w35386, w35387, w35388, w35389, w35390, w35391, w35392, w35393, w35394, w35395, w35396, w35397, w35398, w35399, w35400, w35401, w35402, w35403, w35404, w35405, w35406, w35407, w35408, w35409, w35410, w35411, w35412, w35413, w35414, w35415, w35416, w35417, w35418, w35419, w35420, w35421, w35422, w35423, w35424, w35425, w35426, w35427, w35428, w35429, w35430, w35431, w35432, w35433, w35434, w35435, w35436, w35437, w35438, w35439, w35440, w35441, w35442, w35443, w35444, w35445, w35446, w35447, w35448, w35449, w35450, w35451, w35452, w35453, w35454, w35455, w35456, w35457, w35458, w35459, w35460, w35461, w35462, w35463, w35464, w35465, w35466, w35467, w35468, w35469, w35470, w35471, w35472, w35473, w35474, w35475, w35476, w35477, w35478, w35479, w35480, w35481, w35482, w35483, w35484, w35485, w35486, w35487, w35488, w35489, w35490, w35491, w35492, w35493, w35494, w35495, w35496, w35497, w35498, w35499, w35500, w35501, w35502, w35503, w35504, w35505, w35506, w35507, w35508, w35509, w35510, w35511, w35512, w35513, w35514, w35515, w35516, w35517, w35518, w35519, w35520, w35521, w35522, w35523, w35524, w35525, w35526, w35527, w35528, w35529, w35530, w35531, w35532, w35533, w35534, w35535, w35536, w35537, w35538, w35539, w35540, w35541, w35542, w35543, w35544, w35545, w35546, w35547, w35548, w35549, w35550, w35551, w35552, w35553, w35554, w35555, w35556, w35557, w35558, w35559, w35560, w35561, w35562, w35563, w35564, w35565, w35566, w35567, w35568, w35569, w35570, w35571, w35572, w35573, w35574, w35575, w35576, w35577, w35578, w35579, w35580, w35581, w35582, w35583, w35584, w35585, w35586, w35587, w35588, w35589, w35590, w35591, w35592, w35593, w35594, w35595, w35596, w35597, w35598, w35599, w35600, w35601, w35602, w35603, w35604, w35605, w35606, w35607, w35608, w35609, w35610, w35611, w35612, w35613, w35614, w35615, w35616, w35617, w35618, w35619, w35620, w35621, w35622, w35623, w35624, w35625, w35626, w35627, w35628, w35629, w35630, w35631, w35632, w35633, w35634, w35635, w35636, w35637, w35638, w35639, w35640, w35641, w35642, w35643, w35644, w35645, w35646, w35647, w35648, w35649, w35650, w35651, w35652, w35653, w35654, w35655, w35656, w35657, w35658, w35659, w35660, w35661, w35662, w35663, w35664, w35665, w35666, w35667, w35668, w35669, w35670, w35671, w35672, w35673, w35674, w35675, w35676, w35677, w35678, w35679, w35680, w35681, w35682, w35683, w35684, w35685, w35686, w35687, w35688, w35689, w35690, w35691, w35692, w35693, w35694, w35695, w35696, w35697, w35698, w35699, w35700, w35701, w35702, w35703, w35704, w35705, w35706, w35707, w35708, w35709, w35710, w35711, w35712, w35713, w35714, w35715, w35716, w35717, w35718, w35719, w35720, w35721, w35722, w35723, w35724, w35725, w35726, w35727, w35728, w35729, w35730, w35731, w35732, w35733, w35734, w35735, w35736, w35737, w35738, w35739, w35740, w35741, w35742, w35743, w35744, w35745, w35746, w35747, w35748, w35749, w35750, w35751, w35752, w35753, w35754, w35755, w35756, w35757, w35758, w35759, w35760, w35761, w35762, w35763, w35764, w35765, w35766, w35767, w35768, w35769, w35770, w35771, w35772, w35773, w35774, w35775, w35776, w35777, w35778, w35779, w35780, w35781, w35782, w35783, w35784, w35785, w35786, w35787, w35788, w35789, w35790, w35791, w35792, w35793, w35794, w35795, w35796, w35797, w35798, w35799, w35800, w35801, w35802, w35803, w35804, w35805, w35806, w35807, w35808, w35809, w35810, w35811, w35812, w35813, w35814, w35815, w35816, w35817, w35818, w35819, w35820, w35821, w35822, w35823, w35824, w35825, w35826, w35827, w35828, w35829, w35830, w35831, w35832, w35833, w35834, w35835, w35836, w35837, w35838, w35839, w35840, w35841, w35842, w35843, w35844, w35845, w35846, w35847, w35848, w35849, w35850, w35851, w35852, w35853, w35854, w35855, w35856, w35857, w35858, w35859, w35860, w35861, w35862, w35863, w35864, w35865, w35866, w35867, w35868, w35869, w35870, w35871, w35872, w35873, w35874, w35875, w35876, w35877, w35878, w35879, w35880, w35881, w35882, w35883, w35884, w35885, w35886, w35887, w35888, w35889, w35890, w35891, w35892, w35893, w35894, w35895, w35896, w35897, w35898, w35899, w35900, w35901, w35902, w35903, w35904, w35905, w35906, w35907, w35908, w35909, w35910, w35911, w35912, w35913, w35914, w35915, w35916, w35917, w35918, w35919, w35920, w35921, w35922, w35923, w35924, w35925, w35926, w35927, w35928, w35929, w35930, w35931, w35932, w35933, w35934, w35935, w35936, w35937, w35938, w35939, w35940, w35941, w35942, w35943, w35944, w35945, w35946, w35947, w35948, w35949, w35950, w35951, w35952, w35953, w35954, w35955, w35956, w35957, w35958, w35959, w35960, w35961, w35962, w35963, w35964, w35965, w35966, w35967, w35968, w35969, w35970, w35971, w35972, w35973, w35974, w35975, w35976, w35977, w35978, w35979, w35980, w35981, w35982, w35983, w35984, w35985, w35986, w35987, w35988, w35989, w35990, w35991, w35992, w35993, w35994, w35995, w35996, w35997, w35998, w35999, w36000, w36001, w36002, w36003, w36004, w36005, w36006, w36007, w36008, w36009, w36010, w36011, w36012, w36013, w36014, w36015, w36016, w36017, w36018, w36019, w36020, w36021, w36022, w36023, w36024, w36025, w36026, w36027, w36028, w36029, w36030, w36031, w36032, w36033, w36034, w36035, w36036, w36037, w36038, w36039, w36040, w36041, w36042, w36043, w36044, w36045, w36046, w36047, w36048, w36049, w36050, w36051, w36052, w36053, w36054, w36055, w36056, w36057, w36058, w36059, w36060, w36061, w36062, w36063, w36064, w36065, w36066, w36067, w36068, w36069, w36070, w36071, w36072, w36073, w36074, w36075, w36076, w36077, w36078, w36079, w36080, w36081, w36082, w36083, w36084, w36085, w36086, w36087, w36088, w36089, w36090, w36091, w36092, w36093, w36094, w36095, w36096, w36097, w36098, w36099, w36100, w36101, w36102, w36103, w36104, w36105, w36106, w36107, w36108, w36109, w36110, w36111, w36112, w36113, w36114, w36115, w36116, w36117, w36118, w36119, w36120, w36121, w36122, w36123, w36124, w36125, w36126, w36127, w36128, w36129, w36130, w36131, w36132, w36133, w36134, w36135, w36136, w36137, w36138, w36139, w36140, w36141, w36142, w36143, w36144, w36145, w36146, w36147, w36148, w36149, w36150, w36151, w36152, w36153, w36154, w36155, w36156, w36157, w36158, w36159, w36160, w36161, w36162, w36163, w36164, w36165, w36166, w36167, w36168, w36169, w36170, w36171, w36172, w36173, w36174, w36175, w36176, w36177, w36178, w36179, w36180, w36181, w36182, w36183, w36184, w36185, w36186, w36187, w36188, w36189, w36190, w36191, w36192, w36193, w36194, w36195, w36196, w36197, w36198, w36199, w36200, w36201, w36202, w36203, w36204, w36205, w36206, w36207, w36208, w36209, w36210, w36211, w36212, w36213, w36214, w36215, w36216, w36217, w36218, w36219, w36220, w36221, w36222, w36223, w36224, w36225, w36226, w36227, w36228, w36229, w36230, w36231, w36232, w36233, w36234, w36235, w36236, w36237, w36238, w36239, w36240, w36241, w36242, w36243, w36244, w36245, w36246, w36247, w36248, w36249, w36250, w36251, w36252, w36253, w36254, w36255, w36256, w36257, w36258, w36259, w36260, w36261, w36262, w36263, w36264, w36265, w36266, w36267, w36268, w36269, w36270, w36271, w36272, w36273, w36274, w36275, w36276, w36277, w36278, w36279, w36280, w36281, w36282, w36283, w36284, w36285, w36286, w36287, w36288, w36289, w36290, w36291, w36292, w36293, w36294, w36295, w36296, w36297, w36298, w36299, w36300, w36301, w36302, w36303, w36304, w36305, w36306, w36307, w36308, w36309, w36310, w36311, w36312, w36313, w36314, w36315, w36316, w36317, w36318, w36319, w36320, w36321, w36322, w36323, w36324, w36325, w36326, w36327, w36328, w36329, w36330, w36331, w36332, w36333, w36334, w36335, w36336, w36337, w36338, w36339, w36340, w36341, w36342, w36343, w36344, w36345, w36346, w36347, w36348, w36349, w36350, w36351, w36352, w36353, w36354, w36355, w36356, w36357, w36358, w36359, w36360, w36361, w36362, w36363, w36364, w36365, w36366, w36367, w36368, w36369, w36370, w36371, w36372, w36373, w36374, w36375, w36376, w36377, w36378, w36379, w36380, w36381, w36382, w36383, w36384, w36385, w36386, w36387, w36388, w36389, w36390, w36391, w36392, w36393, w36394, w36395, w36396, w36397, w36398, w36399, w36400, w36401, w36402, w36403, w36404, w36405, w36406, w36407, w36408, w36409, w36410, w36411, w36412, w36413, w36414, w36415, w36416, w36417, w36418, w36419, w36420, w36421, w36422, w36423, w36424, w36425, w36426, w36427, w36428, w36429, w36430, w36431, w36432, w36433, w36434, w36435, w36436, w36437, w36438, w36439, w36440, w36441, w36442, w36443, w36444, w36445, w36446, w36447, w36448, w36449, w36450, w36451, w36452, w36453, w36454, w36455, w36456, w36457, w36458, w36459, w36460, w36461, w36462, w36463, w36464, w36465, w36466, w36467, w36468, w36469, w36470, w36471, w36472, w36473, w36474, w36475, w36476, w36477, w36478, w36479, w36480, w36481, w36482, w36483, w36484, w36485, w36486, w36487, w36488, w36489, w36490, w36491, w36492, w36493, w36494, w36495, w36496, w36497, w36498, w36499, w36500, w36501, w36502, w36503, w36504, w36505, w36506, w36507, w36508, w36509, w36510, w36511, w36512, w36513, w36514, w36515, w36516, w36517, w36518, w36519, w36520, w36521, w36522, w36523, w36524, w36525, w36526, w36527, w36528, w36529, w36530, w36531, w36532, w36533, w36534, w36535, w36536, w36537, w36538, w36539, w36540, w36541, w36542, w36543, w36544, w36545, w36546, w36547, w36548, w36549, w36550, w36551, w36552, w36553, w36554, w36555, w36556, w36557, w36558, w36559, w36560, w36561, w36562, w36563, w36564, w36565, w36566, w36567, w36568, w36569, w36570, w36571, w36572, w36573, w36574, w36575, w36576, w36577, w36578, w36579, w36580, w36581, w36582, w36583, w36584, w36585, w36586, w36587, w36588, w36589, w36590, w36591, w36592, w36593, w36594, w36595, w36596, w36597, w36598, w36599, w36600, w36601, w36602, w36603, w36604, w36605, w36606, w36607, w36608, w36609, w36610, w36611, w36612, w36613, w36614, w36615, w36616, w36617, w36618, w36619, w36620, w36621, w36622, w36623, w36624, w36625, w36626, w36627, w36628, w36629, w36630, w36631, w36632, w36633, w36634, w36635, w36636, w36637, w36638, w36639, w36640, w36641, w36642, w36643, w36644, w36645, w36646, w36647, w36648, w36649, w36650, w36651, w36652, w36653, w36654, w36655, w36656, w36657, w36658, w36659, w36660, w36661, w36662, w36663, w36664, w36665, w36666, w36667, w36668, w36669, w36670, w36671, w36672, w36673, w36674, w36675, w36676, w36677, w36678, w36679, w36680, w36681, w36682, w36683, w36684, w36685, w36686, w36687, w36688, w36689, w36690, w36691, w36692, w36693, w36694, w36695, w36696, w36697, w36698, w36699, w36700, w36701, w36702, w36703, w36704, w36705, w36706, w36707, w36708, w36709, w36710, w36711, w36712, w36713, w36714, w36715, w36716, w36717, w36718, w36719, w36720, w36721, w36722, w36723, w36724, w36725, w36726, w36727, w36728, w36729, w36730, w36731, w36732, w36733, w36734, w36735, w36736, w36737, w36738, w36739, w36740, w36741, w36742, w36743, w36744, w36745, w36746, w36747, w36748, w36749, w36750, w36751, w36752, w36753, w36754, w36755, w36756, w36757, w36758, w36759, w36760, w36761, w36762, w36763, w36764, w36765, w36766, w36767, w36768, w36769, w36770, w36771, w36772, w36773, w36774, w36775, w36776, w36777, w36778, w36779, w36780, w36781, w36782, w36783, w36784, w36785, w36786, w36787, w36788, w36789, w36790, w36791, w36792, w36793, w36794, w36795, w36796, w36797, w36798, w36799, w36800, w36801, w36802, w36803, w36804, w36805, w36806, w36807, w36808, w36809, w36810, w36811, w36812, w36813, w36814, w36815, w36816, w36817, w36818, w36819, w36820, w36821, w36822, w36823, w36824, w36825, w36826, w36827, w36828, w36829, w36830, w36831, w36832, w36833, w36834, w36835, w36836, w36837, w36838, w36839, w36840, w36841, w36842, w36843, w36844, w36845, w36846, w36847, w36848, w36849, w36850, w36851, w36852, w36853, w36854, w36855, w36856, w36857, w36858, w36859, w36860, w36861, w36862, w36863, w36864, w36865, w36866, w36867, w36868, w36869, w36870, w36871, w36872, w36873, w36874, w36875, w36876, w36877, w36878, w36879, w36880, w36881, w36882, w36883, w36884, w36885, w36886, w36887, w36888, w36889, w36890, w36891, w36892, w36893, w36894, w36895, w36896, w36897, w36898, w36899, w36900, w36901, w36902, w36903, w36904, w36905, w36906, w36907, w36908, w36909, w36910, w36911, w36912, w36913, w36914, w36915, w36916, w36917, w36918, w36919, w36920, w36921, w36922, w36923, w36924, w36925, w36926, w36927, w36928, w36929, w36930, w36931, w36932, w36933, w36934, w36935, w36936, w36937, w36938, w36939, w36940, w36941, w36942, w36943, w36944, w36945, w36946, w36947, w36948, w36949, w36950, w36951, w36952, w36953, w36954, w36955, w36956, w36957, w36958, w36959, w36960, w36961, w36962, w36963, w36964, w36965, w36966, w36967, w36968, w36969, w36970, w36971, w36972, w36973, w36974, w36975, w36976, w36977, w36978, w36979, w36980, w36981, w36982, w36983, w36984, w36985, w36986, w36987, w36988, w36989, w36990, w36991, w36992, w36993, w36994, w36995, w36996, w36997, w36998, w36999, w37000, w37001, w37002, w37003, w37004, w37005, w37006, w37007, w37008, w37009, w37010, w37011, w37012, w37013, w37014, w37015, w37016, w37017, w37018, w37019, w37020, w37021, w37022, w37023, w37024, w37025, w37026, w37027, w37028, w37029, w37030, w37031, w37032, w37033, w37034, w37035, w37036, w37037, w37038, w37039, w37040, w37041, w37042, w37043, w37044, w37045, w37046, w37047, w37048, w37049, w37050, w37051, w37052, w37053, w37054, w37055, w37056, w37057, w37058, w37059, w37060, w37061, w37062, w37063, w37064, w37065, w37066, w37067, w37068, w37069, w37070, w37071, w37072, w37073, w37074, w37075, w37076, w37077, w37078, w37079, w37080, w37081, w37082, w37083, w37084, w37085, w37086, w37087, w37088, w37089, w37090, w37091, w37092, w37093, w37094, w37095, w37096, w37097, w37098, w37099, w37100, w37101, w37102, w37103, w37104, w37105, w37106, w37107, w37108, w37109, w37110, w37111, w37112, w37113, w37114, w37115, w37116, w37117, w37118, w37119, w37120, w37121, w37122, w37123, w37124, w37125, w37126, w37127, w37128, w37129, w37130, w37131, w37132, w37133, w37134, w37135, w37136, w37137, w37138, w37139, w37140, w37141, w37142, w37143, w37144, w37145, w37146, w37147, w37148, w37149, w37150, w37151, w37152, w37153, w37154, w37155, w37156, w37157, w37158, w37159, w37160, w37161, w37162, w37163, w37164, w37165, w37166, w37167, w37168, w37169, w37170, w37171, w37172, w37173, w37174, w37175, w37176, w37177, w37178, w37179, w37180, w37181, w37182, w37183, w37184, w37185, w37186, w37187, w37188, w37189, w37190, w37191, w37192, w37193, w37194, w37195, w37196, w37197, w37198, w37199, w37200, w37201, w37202, w37203, w37204, w37205, w37206, w37207, w37208, w37209, w37210, w37211, w37212, w37213, w37214, w37215, w37216, w37217, w37218, w37219, w37220, w37221, w37222, w37223, w37224, w37225, w37226, w37227, w37228, w37229, w37230, w37231, w37232, w37233, w37234, w37235, w37236, w37237, w37238, w37239, w37240, w37241, w37242, w37243, w37244, w37245, w37246, w37247, w37248, w37249, w37250, w37251, w37252, w37253, w37254, w37255, w37256, w37257, w37258, w37259, w37260, w37261, w37262, w37263, w37264, w37265, w37266, w37267, w37268, w37269, w37270, w37271, w37272, w37273, w37274, w37275, w37276, w37277, w37278, w37279, w37280, w37281, w37282, w37283, w37284, w37285, w37286, w37287, w37288, w37289, w37290, w37291, w37292, w37293, w37294, w37295, w37296, w37297, w37298, w37299, w37300, w37301, w37302, w37303, w37304, w37305, w37306, w37307, w37308, w37309, w37310, w37311, w37312, w37313, w37314, w37315, w37316, w37317, w37318, w37319, w37320, w37321, w37322, w37323, w37324, w37325, w37326, w37327, w37328, w37329, w37330, w37331, w37332, w37333, w37334, w37335, w37336, w37337, w37338, w37339, w37340, w37341, w37342, w37343, w37344, w37345, w37346, w37347, w37348, w37349, w37350, w37351, w37352, w37353, w37354, w37355, w37356, w37357, w37358, w37359, w37360, w37361, w37362, w37363, w37364, w37365, w37366, w37367, w37368, w37369, w37370, w37371, w37372, w37373, w37374, w37375, w37376, w37377, w37378, w37379, w37380, w37381, w37382, w37383, w37384, w37385, w37386, w37387, w37388, w37389, w37390, w37391, w37392, w37393, w37394, w37395, w37396, w37397, w37398, w37399, w37400, w37401, w37402, w37403, w37404, w37405, w37406, w37407, w37408, w37409, w37410, w37411, w37412, w37413, w37414, w37415, w37416, w37417, w37418, w37419, w37420, w37421, w37422, w37423, w37424, w37425, w37426, w37427, w37428, w37429, w37430, w37431, w37432, w37433, w37434, w37435, w37436, w37437, w37438, w37439, w37440, w37441, w37442, w37443, w37444, w37445, w37446, w37447, w37448, w37449, w37450, w37451, w37452, w37453, w37454, w37455, w37456, w37457, w37458, w37459, w37460, w37461, w37462, w37463, w37464, w37465, w37466, w37467, w37468, w37469, w37470, w37471, w37472, w37473, w37474, w37475, w37476, w37477, w37478, w37479, w37480, w37481, w37482, w37483, w37484, w37485, w37486, w37487, w37488, w37489, w37490, w37491, w37492, w37493, w37494, w37495, w37496, w37497, w37498, w37499, w37500, w37501, w37502, w37503, w37504, w37505, w37506, w37507, w37508, w37509, w37510, w37511, w37512, w37513, w37514, w37515, w37516, w37517, w37518, w37519, w37520, w37521, w37522, w37523, w37524, w37525, w37526, w37527, w37528, w37529, w37530, w37531, w37532, w37533, w37534, w37535, w37536, w37537, w37538, w37539, w37540, w37541, w37542, w37543, w37544, w37545, w37546, w37547, w37548, w37549, w37550, w37551, w37552, w37553, w37554, w37555, w37556, w37557, w37558, w37559, w37560, w37561, w37562, w37563, w37564, w37565, w37566, w37567, w37568, w37569, w37570, w37571, w37572, w37573, w37574, w37575, w37576, w37577, w37578, w37579, w37580, w37581, w37582, w37583, w37584, w37585, w37586, w37587, w37588, w37589, w37590, w37591, w37592, w37593, w37594, w37595, w37596, w37597, w37598, w37599, w37600, w37601, w37602, w37603, w37604, w37605, w37606, w37607, w37608, w37609, w37610, w37611, w37612, w37613, w37614, w37615, w37616, w37617, w37618, w37619, w37620, w37621, w37622, w37623, w37624, w37625, w37626, w37627, w37628, w37629, w37630, w37631, w37632, w37633, w37634, w37635, w37636, w37637, w37638, w37639, w37640, w37641, w37642, w37643, w37644, w37645, w37646, w37647, w37648, w37649, w37650, w37651, w37652, w37653, w37654, w37655, w37656, w37657, w37658, w37659, w37660, w37661, w37662, w37663, w37664, w37665, w37666, w37667, w37668, w37669, w37670, w37671, w37672, w37673, w37674, w37675, w37676, w37677, w37678, w37679, w37680, w37681, w37682, w37683, w37684, w37685, w37686, w37687, w37688, w37689, w37690, w37691, w37692, w37693, w37694, w37695, w37696, w37697, w37698, w37699, w37700, w37701, w37702, w37703, w37704, w37705, w37706, w37707, w37708, w37709, w37710, w37711, w37712, w37713, w37714, w37715, w37716, w37717, w37718, w37719, w37720, w37721, w37722, w37723, w37724, w37725, w37726, w37727, w37728, w37729, w37730, w37731, w37732, w37733, w37734, w37735, w37736, w37737, w37738, w37739, w37740, w37741, w37742, w37743, w37744, w37745, w37746, w37747, w37748, w37749, w37750, w37751, w37752, w37753, w37754, w37755, w37756, w37757, w37758, w37759, w37760, w37761, w37762, w37763, w37764, w37765, w37766, w37767, w37768, w37769, w37770, w37771, w37772, w37773, w37774, w37775, w37776, w37777, w37778, w37779, w37780, w37781, w37782, w37783, w37784, w37785, w37786, w37787, w37788, w37789, w37790, w37791, w37792, w37793, w37794, w37795, w37796, w37797, w37798, w37799, w37800, w37801, w37802, w37803, w37804, w37805, w37806, w37807, w37808, w37809, w37810, w37811, w37812, w37813, w37814, w37815, w37816, w37817, w37818, w37819, w37820, w37821, w37822, w37823, w37824, w37825, w37826, w37827, w37828, w37829, w37830, w37831, w37832, w37833, w37834, w37835, w37836, w37837, w37838, w37839, w37840, w37841, w37842, w37843, w37844, w37845, w37846, w37847, w37848, w37849, w37850, w37851, w37852, w37853, w37854, w37855, w37856, w37857, w37858, w37859, w37860, w37861, w37862, w37863, w37864, w37865, w37866, w37867, w37868, w37869, w37870, w37871, w37872, w37873, w37874, w37875, w37876, w37877, w37878, w37879, w37880, w37881, w37882, w37883, w37884, w37885, w37886, w37887, w37888, w37889, w37890, w37891, w37892, w37893, w37894, w37895, w37896, w37897, w37898, w37899, w37900, w37901, w37902, w37903, w37904, w37905, w37906, w37907, w37908, w37909, w37910, w37911, w37912, w37913, w37914, w37915, w37916, w37917, w37918, w37919, w37920, w37921, w37922, w37923, w37924, w37925, w37926, w37927, w37928, w37929, w37930, w37931, w37932, w37933, w37934, w37935, w37936, w37937, w37938, w37939, w37940, w37941, w37942, w37943, w37944, w37945, w37946, w37947, w37948, w37949, w37950, w37951, w37952, w37953, w37954, w37955, w37956, w37957, w37958, w37959, w37960, w37961, w37962, w37963, w37964, w37965, w37966, w37967, w37968, w37969, w37970, w37971, w37972, w37973, w37974, w37975, w37976, w37977, w37978, w37979, w37980, w37981, w37982, w37983, w37984, w37985, w37986, w37987, w37988, w37989, w37990, w37991, w37992, w37993, w37994, w37995, w37996, w37997, w37998, w37999, w38000, w38001, w38002, w38003, w38004, w38005, w38006, w38007, w38008, w38009, w38010, w38011, w38012, w38013, w38014, w38015, w38016, w38017, w38018, w38019, w38020, w38021, w38022, w38023, w38024, w38025, w38026, w38027, w38028, w38029, w38030, w38031, w38032, w38033, w38034, w38035, w38036, w38037, w38038, w38039, w38040, w38041, w38042, w38043, w38044, w38045, w38046, w38047, w38048, w38049, w38050, w38051, w38052, w38053, w38054, w38055, w38056, w38057, w38058, w38059, w38060, w38061, w38062, w38063, w38064, w38065, w38066, w38067, w38068, w38069, w38070, w38071, w38072, w38073, w38074, w38075, w38076, w38077, w38078, w38079, w38080, w38081, w38082, w38083, w38084, w38085, w38086, w38087, w38088, w38089, w38090, w38091, w38092, w38093, w38094, w38095, w38096, w38097, w38098, w38099, w38100, w38101, w38102, w38103, w38104, w38105, w38106, w38107, w38108, w38109, w38110, w38111, w38112, w38113, w38114, w38115, w38116, w38117, w38118, w38119, w38120, w38121, w38122, w38123, w38124, w38125, w38126, w38127, w38128, w38129, w38130, w38131, w38132, w38133, w38134, w38135, w38136, w38137, w38138, w38139, w38140, w38141, w38142, w38143, w38144, w38145, w38146, w38147, w38148, w38149, w38150, w38151, w38152, w38153, w38154, w38155, w38156, w38157, w38158, w38159, w38160, w38161, w38162, w38163, w38164, w38165, w38166, w38167, w38168, w38169, w38170, w38171, w38172, w38173, w38174, w38175, w38176, w38177, w38178, w38179, w38180, w38181, w38182, w38183, w38184, w38185, w38186, w38187, w38188, w38189, w38190, w38191, w38192, w38193, w38194, w38195, w38196, w38197, w38198, w38199, w38200, w38201, w38202, w38203, w38204, w38205, w38206, w38207, w38208, w38209, w38210, w38211, w38212, w38213, w38214, w38215, w38216, w38217, w38218, w38219, w38220, w38221, w38222, w38223, w38224, w38225, w38226, w38227, w38228, w38229, w38230, w38231, w38232, w38233, w38234, w38235, w38236, w38237, w38238, w38239, w38240, w38241, w38242, w38243, w38244, w38245, w38246, w38247, w38248, w38249, w38250, w38251, w38252, w38253, w38254, w38255, w38256, w38257, w38258, w38259, w38260, w38261, w38262, w38263, w38264, w38265, w38266, w38267, w38268, w38269, w38270, w38271, w38272, w38273, w38274, w38275, w38276, w38277, w38278, w38279, w38280, w38281, w38282, w38283, w38284, w38285, w38286, w38287, w38288, w38289, w38290, w38291, w38292, w38293, w38294, w38295, w38296, w38297, w38298, w38299, w38300, w38301, w38302, w38303, w38304, w38305, w38306, w38307, w38308, w38309, w38310, w38311, w38312, w38313, w38314, w38315, w38316, w38317, w38318, w38319, w38320, w38321, w38322, w38323, w38324, w38325, w38326, w38327, w38328, w38329, w38330, w38331, w38332, w38333, w38334, w38335, w38336, w38337, w38338, w38339, w38340, w38341, w38342, w38343, w38344, w38345, w38346, w38347, w38348, w38349, w38350, w38351, w38352, w38353, w38354, w38355, w38356, w38357, w38358, w38359, w38360, w38361, w38362, w38363, w38364, w38365, w38366, w38367, w38368, w38369, w38370, w38371, w38372, w38373, w38374, w38375, w38376, w38377, w38378, w38379, w38380, w38381, w38382, w38383, w38384, w38385, w38386, w38387, w38388, w38389, w38390, w38391, w38392, w38393, w38394, w38395, w38396, w38397, w38398, w38399, w38400, w38401, w38402, w38403, w38404, w38405, w38406, w38407, w38408, w38409, w38410, w38411, w38412, w38413, w38414, w38415, w38416, w38417, w38418, w38419, w38420, w38421, w38422, w38423, w38424, w38425, w38426, w38427, w38428, w38429, w38430, w38431, w38432, w38433, w38434, w38435, w38436, w38437, w38438, w38439, w38440, w38441, w38442, w38443, w38444, w38445, w38446, w38447, w38448, w38449, w38450, w38451, w38452, w38453, w38454, w38455, w38456, w38457, w38458, w38459, w38460, w38461, w38462, w38463, w38464, w38465, w38466, w38467, w38468, w38469, w38470, w38471, w38472, w38473, w38474, w38475, w38476, w38477, w38478, w38479, w38480, w38481, w38482, w38483, w38484, w38485, w38486, w38487, w38488, w38489, w38490, w38491, w38492, w38493, w38494, w38495, w38496, w38497, w38498, w38499, w38500, w38501, w38502, w38503, w38504, w38505, w38506, w38507, w38508, w38509, w38510, w38511, w38512, w38513, w38514, w38515, w38516, w38517, w38518, w38519, w38520, w38521, w38522, w38523, w38524, w38525, w38526, w38527, w38528, w38529, w38530, w38531, w38532, w38533, w38534, w38535, w38536, w38537, w38538, w38539, w38540, w38541, w38542, w38543, w38544, w38545, w38546, w38547, w38548, w38549, w38550, w38551, w38552, w38553, w38554, w38555, w38556, w38557, w38558, w38559, w38560, w38561, w38562, w38563, w38564, w38565, w38566, w38567, w38568, w38569, w38570, w38571, w38572, w38573, w38574, w38575, w38576, w38577, w38578, w38579, w38580, w38581, w38582, w38583, w38584, w38585, w38586, w38587, w38588, w38589, w38590, w38591, w38592, w38593, w38594, w38595, w38596, w38597, w38598, w38599, w38600, w38601, w38602, w38603, w38604, w38605, w38606, w38607, w38608, w38609, w38610, w38611, w38612, w38613, w38614, w38615, w38616, w38617, w38618, w38619, w38620, w38621, w38622, w38623, w38624, w38625, w38626, w38627, w38628, w38629, w38630, w38631, w38632, w38633, w38634, w38635, w38636, w38637, w38638, w38639, w38640, w38641, w38642, w38643, w38644, w38645, w38646, w38647, w38648, w38649, w38650, w38651, w38652, w38653, w38654, w38655, w38656, w38657, w38658, w38659, w38660, w38661, w38662, w38663, w38664, w38665, w38666, w38667, w38668, w38669, w38670, w38671, w38672, w38673, w38674, w38675, w38676, w38677, w38678, w38679, w38680, w38681, w38682, w38683, w38684, w38685, w38686, w38687, w38688, w38689, w38690, w38691, w38692, w38693, w38694, w38695, w38696, w38697, w38698, w38699, w38700, w38701, w38702, w38703, w38704, w38705, w38706, w38707, w38708, w38709, w38710, w38711, w38712, w38713, w38714, w38715, w38716, w38717, w38718, w38719, w38720, w38721, w38722, w38723, w38724, w38725, w38726, w38727, w38728, w38729, w38730, w38731, w38732, w38733, w38734, w38735, w38736, w38737, w38738, w38739, w38740, w38741, w38742, w38743, w38744, w38745, w38746, w38747, w38748, w38749, w38750, w38751, w38752, w38753, w38754, w38755, w38756, w38757, w38758, w38759, w38760, w38761, w38762, w38763, w38764, w38765, w38766, w38767, w38768, w38769, w38770, w38771, w38772, w38773, w38774, w38775, w38776, w38777, w38778, w38779, w38780, w38781, w38782, w38783, w38784, w38785, w38786, w38787, w38788, w38789, w38790, w38791, w38792, w38793, w38794, w38795, w38796, w38797, w38798, w38799, w38800, w38801, w38802, w38803, w38804, w38805, w38806, w38807, w38808, w38809, w38810, w38811, w38812, w38813, w38814, w38815, w38816, w38817, w38818, w38819, w38820, w38821, w38822, w38823, w38824, w38825, w38826, w38827, w38828, w38829, w38830, w38831, w38832, w38833, w38834, w38835, w38836, w38837, w38838, w38839, w38840, w38841, w38842, w38843, w38844, w38845, w38846, w38847, w38848, w38849, w38850, w38851, w38852, w38853, w38854, w38855, w38856, w38857, w38858, w38859, w38860, w38861, w38862, w38863, w38864, w38865, w38866, w38867, w38868, w38869, w38870, w38871, w38872, w38873, w38874, w38875, w38876, w38877, w38878, w38879, w38880, w38881, w38882, w38883, w38884, w38885, w38886, w38887, w38888, w38889, w38890, w38891, w38892, w38893, w38894, w38895, w38896, w38897, w38898, w38899, w38900, w38901, w38902, w38903, w38904, w38905, w38906, w38907, w38908, w38909, w38910, w38911, w38912, w38913, w38914, w38915, w38916, w38917, w38918, w38919, w38920, w38921, w38922, w38923, w38924, w38925, w38926, w38927, w38928, w38929, w38930, w38931, w38932, w38933, w38934, w38935, w38936, w38937, w38938, w38939, w38940, w38941, w38942, w38943, w38944, w38945, w38946, w38947, w38948, w38949, w38950, w38951, w38952, w38953, w38954, w38955, w38956, w38957, w38958, w38959, w38960, w38961, w38962, w38963, w38964, w38965, w38966, w38967, w38968, w38969, w38970, w38971, w38972, w38973, w38974, w38975, w38976, w38977, w38978, w38979, w38980, w38981, w38982, w38983, w38984, w38985, w38986, w38987, w38988, w38989, w38990, w38991, w38992, w38993, w38994, w38995, w38996, w38997, w38998, w38999, w39000, w39001, w39002, w39003, w39004, w39005, w39006, w39007, w39008, w39009, w39010, w39011, w39012, w39013, w39014, w39015, w39016, w39017, w39018, w39019, w39020, w39021, w39022, w39023, w39024, w39025, w39026, w39027, w39028, w39029, w39030, w39031, w39032, w39033, w39034, w39035, w39036, w39037, w39038, w39039, w39040, w39041, w39042, w39043, w39044, w39045, w39046, w39047, w39048, w39049, w39050, w39051, w39052, w39053, w39054, w39055, w39056, w39057, w39058, w39059, w39060, w39061, w39062, w39063, w39064, w39065, w39066, w39067, w39068, w39069, w39070, w39071, w39072, w39073, w39074, w39075, w39076, w39077, w39078, w39079, w39080, w39081, w39082, w39083, w39084, w39085, w39086, w39087, w39088, w39089, w39090, w39091, w39092, w39093, w39094, w39095, w39096, w39097, w39098, w39099, w39100, w39101, w39102, w39103, w39104, w39105, w39106, w39107, w39108, w39109, w39110, w39111, w39112, w39113, w39114, w39115, w39116, w39117, w39118, w39119, w39120, w39121, w39122, w39123, w39124, w39125, w39126, w39127, w39128, w39129, w39130, w39131, w39132, w39133, w39134, w39135, w39136, w39137, w39138, w39139, w39140, w39141, w39142, w39143, w39144, w39145, w39146, w39147, w39148, w39149, w39150, w39151, w39152, w39153, w39154, w39155, w39156, w39157, w39158, w39159, w39160, w39161, w39162, w39163, w39164, w39165, w39166, w39167, w39168, w39169, w39170, w39171, w39172, w39173, w39174, w39175, w39176, w39177, w39178, w39179, w39180, w39181, w39182, w39183, w39184, w39185, w39186, w39187, w39188, w39189, w39190, w39191, w39192, w39193, w39194, w39195, w39196, w39197, w39198, w39199, w39200, w39201, w39202, w39203, w39204, w39205, w39206, w39207, w39208, w39209, w39210, w39211, w39212, w39213, w39214, w39215, w39216, w39217, w39218, w39219, w39220, w39221, w39222, w39223, w39224, w39225, w39226, w39227, w39228, w39229, w39230, w39231, w39232, w39233, w39234, w39235, w39236, w39237, w39238, w39239, w39240, w39241, w39242, w39243, w39244, w39245, w39246, w39247, w39248, w39249, w39250, w39251, w39252, w39253, w39254, w39255, w39256, w39257, w39258, w39259, w39260, w39261, w39262, w39263, w39264, w39265, w39266, w39267, w39268, w39269, w39270, w39271, w39272, w39273, w39274, w39275, w39276, w39277, w39278, w39279, w39280, w39281, w39282, w39283, w39284, w39285, w39286, w39287, w39288, w39289, w39290, w39291, w39292, w39293, w39294, w39295, w39296, w39297, w39298, w39299, w39300, w39301, w39302, w39303, w39304, w39305, w39306, w39307, w39308, w39309, w39310, w39311, w39312, w39313, w39314, w39315, w39316, w39317, w39318, w39319, w39320, w39321, w39322, w39323, w39324, w39325, w39326, w39327, w39328, w39329, w39330, w39331, w39332, w39333, w39334, w39335, w39336, w39337, w39338, w39339, w39340, w39341, w39342, w39343, w39344, w39345, w39346, w39347, w39348, w39349, w39350, w39351, w39352, w39353, w39354, w39355, w39356, w39357, w39358, w39359, w39360, w39361, w39362, w39363, w39364, w39365, w39366, w39367, w39368, w39369, w39370, w39371, w39372, w39373, w39374, w39375, w39376, w39377, w39378, w39379, w39380, w39381, w39382, w39383, w39384, w39385, w39386, w39387, w39388, w39389, w39390, w39391, w39392, w39393, w39394, w39395, w39396, w39397, w39398, w39399, w39400, w39401, w39402, w39403, w39404, w39405, w39406, w39407, w39408, w39409, w39410, w39411, w39412, w39413, w39414, w39415, w39416, w39417, w39418, w39419, w39420, w39421, w39422, w39423, w39424, w39425, w39426, w39427, w39428, w39429, w39430, w39431, w39432, w39433, w39434, w39435, w39436, w39437, w39438, w39439, w39440, w39441, w39442, w39443, w39444, w39445, w39446, w39447, w39448, w39449, w39450, w39451, w39452, w39453, w39454, w39455, w39456, w39457, w39458, w39459, w39460, w39461, w39462, w39463, w39464, w39465, w39466, w39467, w39468, w39469, w39470, w39471, w39472, w39473, w39474, w39475, w39476, w39477, w39478, w39479, w39480, w39481, w39482, w39483, w39484, w39485, w39486, w39487, w39488, w39489, w39490, w39491, w39492, w39493, w39494, w39495, w39496, w39497, w39498, w39499, w39500, w39501, w39502, w39503, w39504, w39505, w39506, w39507, w39508, w39509, w39510, w39511, w39512, w39513, w39514, w39515, w39516, w39517, w39518, w39519, w39520, w39521, w39522, w39523, w39524, w39525, w39526, w39527, w39528, w39529, w39530, w39531, w39532, w39533, w39534, w39535, w39536, w39537, w39538, w39539, w39540, w39541, w39542, w39543, w39544, w39545, w39546, w39547, w39548, w39549, w39550, w39551, w39552, w39553, w39554, w39555, w39556, w39557, w39558, w39559, w39560, w39561, w39562, w39563, w39564, w39565, w39566, w39567, w39568, w39569, w39570, w39571, w39572, w39573, w39574, w39575, w39576, w39577, w39578, w39579, w39580, w39581, w39582, w39583, w39584, w39585, w39586, w39587, w39588, w39589, w39590, w39591, w39592, w39593, w39594, w39595, w39596, w39597, w39598, w39599, w39600, w39601, w39602, w39603, w39604, w39605, w39606, w39607, w39608, w39609, w39610, w39611, w39612, w39613, w39614, w39615, w39616, w39617, w39618, w39619, w39620, w39621, w39622, w39623, w39624, w39625, w39626, w39627, w39628, w39629, w39630, w39631, w39632, w39633, w39634, w39635, w39636, w39637, w39638, w39639, w39640, w39641, w39642, w39643, w39644, w39645, w39646, w39647, w39648, w39649, w39650, w39651, w39652, w39653, w39654, w39655, w39656, w39657, w39658, w39659, w39660, w39661, w39662, w39663, w39664, w39665, w39666, w39667, w39668, w39669, w39670, w39671, w39672, w39673, w39674, w39675, w39676, w39677, w39678, w39679, w39680, w39681, w39682, w39683, w39684, w39685, w39686, w39687, w39688, w39689, w39690, w39691, w39692, w39693, w39694, w39695, w39696, w39697, w39698, w39699, w39700, w39701, w39702, w39703, w39704, w39705, w39706, w39707, w39708, w39709, w39710, w39711, w39712, w39713, w39714, w39715, w39716, w39717, w39718, w39719, w39720, w39721, w39722, w39723, w39724, w39725, w39726, w39727, w39728, w39729, w39730, w39731, w39732, w39733, w39734, w39735, w39736, w39737, w39738, w39739, w39740, w39741, w39742, w39743, w39744, w39745, w39746, w39747, w39748, w39749, w39750, w39751, w39752, w39753, w39754, w39755, w39756, w39757, w39758, w39759, w39760, w39761, w39762, w39763, w39764, w39765, w39766, w39767, w39768, w39769, w39770, w39771, w39772, w39773, w39774, w39775, w39776, w39777, w39778, w39779, w39780, w39781, w39782, w39783, w39784, w39785, w39786, w39787, w39788, w39789, w39790, w39791, w39792, w39793, w39794, w39795, w39796, w39797, w39798, w39799, w39800, w39801, w39802, w39803, w39804, w39805, w39806, w39807, w39808, w39809, w39810, w39811, w39812, w39813, w39814, w39815, w39816, w39817, w39818, w39819, w39820, w39821, w39822, w39823, w39824, w39825, w39826, w39827, w39828, w39829, w39830, w39831, w39832, w39833, w39834, w39835, w39836, w39837, w39838, w39839, w39840, w39841, w39842, w39843, w39844, w39845, w39846, w39847, w39848, w39849, w39850, w39851, w39852, w39853, w39854, w39855, w39856, w39857, w39858, w39859, w39860, w39861, w39862, w39863, w39864, w39865, w39866, w39867, w39868, w39869, w39870, w39871, w39872, w39873, w39874, w39875, w39876, w39877, w39878, w39879, w39880, w39881, w39882, w39883, w39884, w39885, w39886, w39887, w39888, w39889, w39890, w39891, w39892, w39893, w39894, w39895, w39896, w39897, w39898, w39899, w39900, w39901, w39902, w39903, w39904, w39905, w39906, w39907, w39908, w39909, w39910, w39911, w39912, w39913, w39914, w39915, w39916, w39917, w39918, w39919, w39920, w39921, w39922, w39923, w39924, w39925, w39926, w39927, w39928, w39929, w39930, w39931, w39932, w39933, w39934, w39935, w39936, w39937, w39938, w39939, w39940, w39941, w39942, w39943, w39944, w39945, w39946, w39947, w39948, w39949, w39950, w39951, w39952, w39953, w39954, w39955, w39956, w39957, w39958, w39959, w39960, w39961, w39962, w39963, w39964, w39965, w39966, w39967, w39968, w39969, w39970, w39971, w39972, w39973, w39974, w39975, w39976, w39977, w39978, w39979, w39980, w39981, w39982, w39983, w39984, w39985, w39986, w39987, w39988, w39989, w39990, w39991, w39992, w39993, w39994, w39995, w39996, w39997, w39998, w39999, w40000, w40001, w40002, w40003, w40004, w40005, w40006, w40007, w40008, w40009, w40010, w40011, w40012, w40013, w40014, w40015, w40016, w40017, w40018, w40019, w40020, w40021, w40022, w40023, w40024, w40025, w40026, w40027, w40028, w40029, w40030, w40031, w40032, w40033, w40034, w40035, w40036, w40037, w40038, w40039, w40040, w40041, w40042, w40043, w40044, w40045, w40046, w40047, w40048, w40049, w40050, w40051, w40052, w40053, w40054, w40055, w40056, w40057, w40058, w40059, w40060, w40061, w40062, w40063, w40064, w40065, w40066, w40067, w40068, w40069, w40070, w40071, w40072, w40073, w40074, w40075, w40076, w40077, w40078, w40079, w40080, w40081, w40082, w40083, w40084, w40085, w40086, w40087, w40088, w40089, w40090, w40091, w40092, w40093, w40094, w40095, w40096, w40097, w40098, w40099, w40100, w40101, w40102, w40103, w40104, w40105, w40106, w40107, w40108, w40109, w40110, w40111, w40112, w40113, w40114, w40115, w40116, w40117, w40118, w40119, w40120, w40121, w40122, w40123, w40124, w40125, w40126, w40127, w40128, w40129, w40130, w40131, w40132, w40133, w40134, w40135, w40136, w40137, w40138, w40139, w40140, w40141, w40142, w40143, w40144, w40145, w40146, w40147, w40148, w40149, w40150, w40151, w40152, w40153, w40154, w40155, w40156, w40157, w40158, w40159, w40160, w40161, w40162, w40163, w40164, w40165, w40166, w40167, w40168, w40169, w40170, w40171, w40172, w40173, w40174, w40175, w40176, w40177, w40178, w40179, w40180, w40181, w40182, w40183, w40184, w40185, w40186, w40187, w40188, w40189, w40190, w40191, w40192, w40193, w40194, w40195, w40196, w40197, w40198, w40199, w40200, w40201, w40202, w40203, w40204, w40205, w40206, w40207, w40208, w40209, w40210, w40211, w40212, w40213, w40214, w40215, w40216, w40217, w40218, w40219, w40220, w40221, w40222, w40223, w40224, w40225, w40226, w40227, w40228, w40229, w40230, w40231, w40232, w40233, w40234, w40235, w40236, w40237, w40238, w40239, w40240, w40241, w40242, w40243, w40244, w40245, w40246, w40247, w40248, w40249, w40250, w40251, w40252, w40253, w40254, w40255, w40256, w40257, w40258, w40259, w40260, w40261, w40262, w40263, w40264, w40265, w40266, w40267, w40268, w40269, w40270, w40271, w40272, w40273, w40274, w40275, w40276, w40277, w40278, w40279, w40280, w40281, w40282, w40283, w40284, w40285, w40286, w40287, w40288, w40289, w40290, w40291, w40292, w40293, w40294, w40295, w40296, w40297, w40298, w40299, w40300, w40301, w40302, w40303, w40304, w40305, w40306, w40307, w40308, w40309, w40310, w40311, w40312, w40313, w40314, w40315, w40316, w40317, w40318, w40319, w40320, w40321, w40322, w40323, w40324, w40325, w40326, w40327, w40328, w40329, w40330, w40331, w40332, w40333, w40334, w40335, w40336, w40337, w40338, w40339, w40340, w40341, w40342, w40343, w40344, w40345, w40346, w40347, w40348, w40349, w40350, w40351, w40352, w40353, w40354, w40355, w40356, w40357, w40358, w40359, w40360, w40361, w40362, w40363, w40364, w40365, w40366, w40367, w40368, w40369, w40370, w40371, w40372, w40373, w40374, w40375, w40376, w40377, w40378, w40379, w40380, w40381, w40382, w40383, w40384, w40385, w40386, w40387, w40388, w40389, w40390, w40391, w40392, w40393, w40394, w40395, w40396, w40397, w40398, w40399, w40400, w40401, w40402, w40403, w40404, w40405, w40406, w40407, w40408, w40409, w40410, w40411, w40412, w40413, w40414, w40415, w40416, w40417, w40418, w40419, w40420, w40421, w40422, w40423, w40424, w40425, w40426, w40427, w40428, w40429, w40430, w40431, w40432, w40433, w40434, w40435, w40436, w40437, w40438, w40439, w40440, w40441, w40442, w40443, w40444, w40445, w40446, w40447, w40448, w40449, w40450, w40451, w40452, w40453, w40454, w40455, w40456, w40457, w40458, w40459, w40460, w40461, w40462, w40463, w40464, w40465, w40466, w40467, w40468, w40469, w40470, w40471, w40472, w40473, w40474, w40475, w40476, w40477, w40478, w40479, w40480, w40481, w40482, w40483, w40484, w40485, w40486, w40487, w40488, w40489, w40490, w40491, w40492, w40493, w40494, w40495, w40496, w40497, w40498, w40499, w40500, w40501, w40502, w40503, w40504, w40505, w40506, w40507, w40508, w40509, w40510, w40511, w40512, w40513, w40514, w40515, w40516, w40517, w40518, w40519, w40520, w40521, w40522, w40523, w40524, w40525, w40526, w40527, w40528, w40529, w40530, w40531, w40532, w40533, w40534, w40535, w40536, w40537, w40538, w40539, w40540, w40541, w40542, w40543, w40544, w40545, w40546, w40547, w40548, w40549, w40550, w40551, w40552, w40553, w40554, w40555, w40556, w40557, w40558, w40559, w40560, w40561, w40562, w40563, w40564, w40565, w40566, w40567, w40568, w40569, w40570, w40571, w40572, w40573, w40574, w40575, w40576, w40577, w40578, w40579, w40580, w40581, w40582, w40583, w40584, w40585, w40586, w40587, w40588, w40589, w40590, w40591, w40592, w40593, w40594, w40595, w40596, w40597, w40598, w40599, w40600, w40601, w40602, w40603, w40604, w40605, w40606, w40607, w40608, w40609, w40610, w40611, w40612, w40613, w40614, w40615, w40616, w40617, w40618, w40619, w40620, w40621, w40622, w40623, w40624, w40625, w40626, w40627, w40628, w40629, w40630, w40631, w40632, w40633, w40634, w40635, w40636, w40637, w40638, w40639, w40640, w40641, w40642, w40643, w40644, w40645, w40646, w40647, w40648, w40649, w40650, w40651, w40652, w40653, w40654, w40655, w40656, w40657, w40658, w40659, w40660, w40661, w40662, w40663, w40664, w40665, w40666, w40667, w40668, w40669, w40670, w40671, w40672, w40673, w40674, w40675, w40676, w40677, w40678, w40679, w40680, w40681, w40682, w40683, w40684, w40685, w40686, w40687, w40688, w40689, w40690, w40691, w40692, w40693, w40694, w40695, w40696, w40697, w40698, w40699, w40700, w40701, w40702, w40703, w40704, w40705, w40706, w40707, w40708, w40709, w40710, w40711, w40712, w40713, w40714, w40715, w40716, w40717, w40718, w40719, w40720, w40721, w40722, w40723, w40724, w40725, w40726, w40727, w40728, w40729, w40730, w40731, w40732, w40733, w40734, w40735, w40736, w40737, w40738, w40739, w40740, w40741, w40742, w40743, w40744, w40745, w40746, w40747, w40748, w40749, w40750, w40751, w40752, w40753, w40754, w40755, w40756, w40757, w40758, w40759, w40760, w40761, w40762, w40763, w40764, w40765, w40766, w40767, w40768, w40769, w40770, w40771, w40772, w40773, w40774, w40775, w40776, w40777, w40778, w40779, w40780, w40781, w40782, w40783, w40784, w40785, w40786, w40787, w40788, w40789, w40790, w40791, w40792, w40793, w40794, w40795, w40796, w40797, w40798, w40799, w40800, w40801, w40802, w40803, w40804, w40805, w40806, w40807, w40808, w40809, w40810, w40811, w40812, w40813, w40814, w40815, w40816, w40817, w40818, w40819, w40820, w40821, w40822, w40823, w40824, w40825, w40826, w40827, w40828, w40829, w40830, w40831, w40832, w40833, w40834, w40835, w40836, w40837, w40838, w40839, w40840, w40841, w40842, w40843, w40844, w40845, w40846, w40847, w40848, w40849, w40850, w40851, w40852, w40853, w40854, w40855, w40856, w40857, w40858, w40859, w40860, w40861, w40862, w40863, w40864, w40865, w40866, w40867, w40868, w40869, w40870, w40871, w40872, w40873, w40874, w40875, w40876, w40877, w40878, w40879, w40880, w40881, w40882, w40883, w40884, w40885, w40886, w40887, w40888, w40889, w40890, w40891, w40892, w40893, w40894, w40895, w40896, w40897, w40898, w40899, w40900, w40901, w40902, w40903, w40904, w40905, w40906, w40907, w40908, w40909, w40910, w40911, w40912, w40913, w40914, w40915, w40916, w40917, w40918, w40919, w40920, w40921, w40922, w40923, w40924, w40925, w40926, w40927, w40928, w40929, w40930, w40931, w40932, w40933, w40934, w40935, w40936, w40937, w40938, w40939, w40940, w40941, w40942, w40943, w40944, w40945, w40946, w40947, w40948, w40949, w40950, w40951, w40952, w40953, w40954, w40955, w40956, w40957, w40958, w40959, w40960, w40961, w40962, w40963, w40964, w40965, w40966, w40967, w40968, w40969, w40970, w40971, w40972, w40973, w40974, w40975, w40976, w40977, w40978, w40979, w40980, w40981, w40982, w40983, w40984, w40985, w40986, w40987, w40988, w40989, w40990, w40991, w40992, w40993, w40994, w40995, w40996, w40997, w40998, w40999, w41000, w41001, w41002, w41003, w41004, w41005, w41006, w41007, w41008, w41009, w41010, w41011, w41012, w41013, w41014, w41015, w41016, w41017, w41018, w41019, w41020, w41021, w41022, w41023, w41024, w41025, w41026, w41027, w41028, w41029, w41030, w41031, w41032, w41033, w41034, w41035, w41036, w41037, w41038, w41039, w41040, w41041, w41042, w41043, w41044, w41045, w41046, w41047, w41048, w41049, w41050, w41051, w41052, w41053, w41054, w41055, w41056, w41057, w41058, w41059, w41060, w41061, w41062, w41063, w41064, w41065, w41066, w41067, w41068, w41069, w41070, w41071, w41072, w41073, w41074, w41075, w41076, w41077, w41078, w41079, w41080, w41081, w41082, w41083, w41084, w41085, w41086, w41087, w41088, w41089, w41090, w41091, w41092, w41093, w41094, w41095, w41096, w41097, w41098, w41099, w41100, w41101, w41102, w41103, w41104, w41105, w41106, w41107, w41108, w41109, w41110, w41111, w41112, w41113, w41114, w41115, w41116, w41117, w41118, w41119, w41120, w41121, w41122, w41123, w41124, w41125, w41126, w41127, w41128, w41129, w41130, w41131, w41132, w41133, w41134, w41135, w41136, w41137, w41138, w41139, w41140, w41141, w41142, w41143, w41144, w41145, w41146, w41147, w41148, w41149, w41150, w41151, w41152, w41153, w41154, w41155, w41156, w41157, w41158, w41159, w41160, w41161, w41162, w41163, w41164, w41165, w41166, w41167, w41168, w41169, w41170, w41171, w41172, w41173, w41174, w41175, w41176, w41177, w41178, w41179, w41180, w41181, w41182, w41183, w41184, w41185, w41186, w41187, w41188, w41189, w41190, w41191, w41192, w41193, w41194, w41195, w41196, w41197, w41198, w41199, w41200, w41201, w41202, w41203, w41204, w41205, w41206, w41207, w41208, w41209, w41210, w41211, w41212, w41213, w41214, w41215, w41216, w41217, w41218, w41219, w41220, w41221, w41222, w41223, w41224, w41225, w41226, w41227, w41228, w41229, w41230, w41231, w41232, w41233, w41234, w41235, w41236, w41237, w41238, w41239, w41240, w41241, w41242, w41243, w41244, w41245, w41246, w41247, w41248, w41249, w41250, w41251, w41252, w41253, w41254, w41255, w41256, w41257, w41258, w41259, w41260, w41261, w41262, w41263, w41264, w41265, w41266, w41267, w41268, w41269, w41270, w41271, w41272, w41273, w41274, w41275, w41276, w41277, w41278, w41279, w41280, w41281, w41282, w41283, w41284, w41285, w41286, w41287, w41288, w41289, w41290, w41291, w41292, w41293, w41294, w41295, w41296, w41297, w41298, w41299, w41300, w41301, w41302, w41303, w41304, w41305, w41306, w41307, w41308, w41309, w41310, w41311, w41312, w41313, w41314, w41315, w41316, w41317, w41318, w41319, w41320, w41321, w41322, w41323, w41324, w41325, w41326, w41327, w41328, w41329, w41330, w41331, w41332, w41333, w41334, w41335, w41336, w41337, w41338, w41339, w41340, w41341, w41342, w41343, w41344, w41345, w41346, w41347, w41348, w41349, w41350, w41351, w41352, w41353, w41354, w41355, w41356, w41357, w41358, w41359, w41360, w41361, w41362, w41363, w41364, w41365, w41366, w41367, w41368, w41369, w41370, w41371, w41372, w41373, w41374, w41375, w41376, w41377, w41378, w41379, w41380, w41381, w41382, w41383, w41384, w41385, w41386, w41387, w41388, w41389, w41390, w41391, w41392, w41393, w41394, w41395, w41396, w41397, w41398, w41399, w41400, w41401, w41402, w41403, w41404, w41405, w41406, w41407, w41408, w41409, w41410, w41411, w41412, w41413, w41414, w41415, w41416, w41417, w41418, w41419, w41420, w41421, w41422, w41423, w41424, w41425, w41426, w41427, w41428, w41429, w41430, w41431, w41432, w41433, w41434, w41435, w41436, w41437, w41438, w41439, w41440, w41441, w41442, w41443, w41444, w41445, w41446, w41447, w41448, w41449, w41450, w41451, w41452, w41453, w41454, w41455, w41456, w41457, w41458, w41459, w41460, w41461, w41462, w41463, w41464, w41465, w41466, w41467, w41468, w41469, w41470, w41471, w41472, w41473, w41474, w41475, w41476, w41477, w41478, w41479, w41480, w41481, w41482, w41483, w41484, w41485, w41486, w41487, w41488, w41489, w41490, w41491, w41492, w41493, w41494, w41495, w41496, w41497, w41498, w41499, w41500, w41501, w41502, w41503, w41504, w41505, w41506, w41507, w41508, w41509, w41510, w41511, w41512, w41513, w41514, w41515, w41516, w41517, w41518, w41519, w41520, w41521, w41522, w41523, w41524, w41525, w41526, w41527, w41528, w41529, w41530, w41531, w41532, w41533, w41534, w41535, w41536, w41537, w41538, w41539, w41540, w41541, w41542, w41543, w41544, w41545, w41546, w41547, w41548, w41549, w41550, w41551, w41552, w41553, w41554, w41555, w41556, w41557, w41558, w41559, w41560, w41561, w41562, w41563, w41564, w41565, w41566, w41567, w41568, w41569, w41570, w41571, w41572, w41573, w41574, w41575, w41576, w41577, w41578, w41579, w41580, w41581, w41582, w41583, w41584, w41585, w41586, w41587, w41588, w41589, w41590, w41591, w41592, w41593, w41594, w41595, w41596, w41597, w41598, w41599, w41600, w41601, w41602, w41603, w41604, w41605, w41606, w41607, w41608, w41609, w41610, w41611, w41612, w41613, w41614, w41615, w41616, w41617, w41618, w41619, w41620, w41621, w41622, w41623, w41624, w41625, w41626, w41627, w41628, w41629, w41630, w41631, w41632, w41633, w41634, w41635, w41636, w41637, w41638, w41639, w41640, w41641, w41642, w41643, w41644, w41645, w41646, w41647, w41648, w41649, w41650, w41651, w41652, w41653, w41654, w41655, w41656, w41657, w41658, w41659, w41660, w41661, w41662, w41663, w41664, w41665, w41666, w41667, w41668, w41669, w41670, w41671, w41672, w41673, w41674, w41675, w41676, w41677, w41678, w41679, w41680, w41681, w41682, w41683, w41684, w41685, w41686, w41687, w41688, w41689, w41690, w41691, w41692, w41693, w41694, w41695, w41696, w41697, w41698, w41699, w41700, w41701, w41702, w41703, w41704, w41705, w41706, w41707, w41708, w41709, w41710, w41711, w41712, w41713, w41714, w41715, w41716, w41717, w41718, w41719, w41720, w41721, w41722, w41723, w41724, w41725, w41726, w41727, w41728, w41729, w41730, w41731, w41732, w41733, w41734, w41735, w41736, w41737, w41738, w41739, w41740, w41741, w41742, w41743, w41744, w41745, w41746, w41747, w41748, w41749, w41750, w41751, w41752, w41753, w41754, w41755, w41756, w41757, w41758, w41759, w41760, w41761, w41762, w41763, w41764, w41765, w41766, w41767, w41768, w41769, w41770, w41771, w41772, w41773, w41774, w41775, w41776, w41777, w41778, w41779, w41780, w41781, w41782, w41783, w41784, w41785, w41786, w41787, w41788, w41789, w41790, w41791, w41792, w41793, w41794, w41795, w41796, w41797, w41798, w41799, w41800, w41801, w41802, w41803, w41804, w41805, w41806, w41807, w41808, w41809, w41810, w41811, w41812, w41813, w41814, w41815, w41816, w41817, w41818, w41819, w41820, w41821, w41822, w41823, w41824, w41825, w41826, w41827, w41828, w41829, w41830, w41831, w41832, w41833, w41834, w41835, w41836, w41837, w41838, w41839, w41840, w41841, w41842, w41843, w41844, w41845, w41846, w41847, w41848, w41849, w41850, w41851, w41852, w41853, w41854, w41855, w41856, w41857, w41858, w41859, w41860, w41861, w41862, w41863, w41864, w41865, w41866, w41867, w41868, w41869, w41870, w41871, w41872, w41873, w41874, w41875, w41876, w41877, w41878, w41879, w41880, w41881, w41882, w41883, w41884, w41885, w41886, w41887, w41888, w41889, w41890, w41891, w41892, w41893, w41894, w41895, w41896, w41897, w41898, w41899, w41900, w41901, w41902, w41903, w41904, w41905, w41906, w41907, w41908, w41909, w41910, w41911, w41912, w41913, w41914, w41915, w41916, w41917, w41918, w41919, w41920, w41921, w41922, w41923, w41924, w41925, w41926, w41927, w41928, w41929, w41930, w41931, w41932, w41933, w41934, w41935, w41936, w41937, w41938, w41939, w41940, w41941, w41942, w41943, w41944, w41945, w41946, w41947, w41948, w41949, w41950, w41951, w41952, w41953, w41954, w41955, w41956, w41957, w41958, w41959, w41960, w41961, w41962, w41963, w41964, w41965, w41966, w41967, w41968, w41969, w41970, w41971, w41972, w41973, w41974, w41975, w41976, w41977, w41978, w41979, w41980, w41981, w41982, w41983, w41984, w41985, w41986, w41987, w41988, w41989, w41990, w41991, w41992, w41993, w41994, w41995, w41996, w41997, w41998, w41999, w42000, w42001, w42002, w42003, w42004, w42005, w42006, w42007, w42008, w42009, w42010, w42011, w42012, w42013, w42014, w42015, w42016, w42017, w42018, w42019, w42020, w42021, w42022, w42023, w42024, w42025, w42026, w42027, w42028, w42029, w42030, w42031, w42032, w42033, w42034, w42035, w42036, w42037, w42038, w42039, w42040, w42041, w42042, w42043, w42044, w42045, w42046, w42047, w42048, w42049, w42050, w42051, w42052, w42053, w42054, w42055, w42056, w42057, w42058, w42059, w42060, w42061, w42062, w42063, w42064, w42065, w42066, w42067, w42068, w42069, w42070, w42071, w42072, w42073, w42074, w42075, w42076, w42077, w42078, w42079, w42080, w42081, w42082, w42083, w42084, w42085, w42086, w42087, w42088, w42089, w42090, w42091, w42092, w42093, w42094, w42095, w42096, w42097, w42098, w42099, w42100, w42101, w42102, w42103, w42104, w42105, w42106, w42107, w42108, w42109, w42110, w42111, w42112, w42113, w42114, w42115, w42116, w42117, w42118, w42119, w42120, w42121, w42122, w42123, w42124, w42125, w42126, w42127, w42128, w42129, w42130, w42131, w42132, w42133, w42134, w42135, w42136, w42137, w42138, w42139, w42140, w42141, w42142, w42143, w42144, w42145, w42146, w42147, w42148, w42149, w42150, w42151, w42152, w42153, w42154, w42155, w42156, w42157, w42158, w42159, w42160, w42161, w42162, w42163, w42164, w42165, w42166, w42167, w42168, w42169, w42170, w42171, w42172, w42173, w42174, w42175, w42176, w42177, w42178, w42179, w42180, w42181, w42182, w42183, w42184, w42185, w42186, w42187, w42188, w42189, w42190, w42191, w42192, w42193, w42194, w42195, w42196, w42197, w42198, w42199, w42200, w42201, w42202, w42203, w42204, w42205, w42206, w42207, w42208, w42209, w42210, w42211, w42212, w42213, w42214, w42215, w42216, w42217, w42218, w42219, w42220, w42221, w42222, w42223, w42224, w42225, w42226, w42227, w42228, w42229, w42230, w42231, w42232, w42233, w42234, w42235, w42236, w42237, w42238, w42239, w42240, w42241, w42242, w42243, w42244, w42245, w42246, w42247, w42248, w42249, w42250, w42251, w42252, w42253, w42254, w42255, w42256, w42257, w42258, w42259, w42260, w42261, w42262, w42263, w42264, w42265, w42266, w42267, w42268, w42269, w42270, w42271, w42272, w42273, w42274, w42275, w42276, w42277, w42278, w42279, w42280, w42281, w42282, w42283, w42284, w42285, w42286, w42287, w42288, w42289, w42290, w42291, w42292, w42293, w42294, w42295, w42296, w42297, w42298, w42299, w42300, w42301, w42302, w42303, w42304, w42305, w42306, w42307, w42308, w42309, w42310, w42311, w42312, w42313, w42314, w42315, w42316, w42317, w42318, w42319, w42320, w42321, w42322, w42323, w42324, w42325, w42326, w42327, w42328, w42329, w42330, w42331, w42332, w42333, w42334, w42335, w42336, w42337, w42338, w42339, w42340, w42341, w42342, w42343, w42344, w42345, w42346, w42347, w42348, w42349, w42350, w42351, w42352, w42353, w42354, w42355, w42356, w42357, w42358, w42359, w42360, w42361, w42362, w42363, w42364, w42365, w42366, w42367, w42368, w42369, w42370, w42371, w42372, w42373, w42374, w42375, w42376, w42377, w42378, w42379, w42380, w42381, w42382, w42383, w42384, w42385, w42386, w42387, w42388, w42389, w42390, w42391, w42392, w42393, w42394, w42395, w42396, w42397, w42398, w42399, w42400, w42401, w42402, w42403, w42404, w42405, w42406, w42407, w42408, w42409, w42410, w42411, w42412, w42413, w42414, w42415, w42416, w42417, w42418, w42419, w42420, w42421, w42422, w42423, w42424, w42425, w42426, w42427, w42428, w42429, w42430, w42431, w42432, w42433, w42434, w42435, w42436, w42437, w42438, w42439, w42440, w42441, w42442, w42443, w42444, w42445, w42446, w42447, w42448, w42449, w42450, w42451, w42452, w42453, w42454, w42455, w42456, w42457, w42458, w42459, w42460, w42461, w42462, w42463, w42464, w42465, w42466, w42467, w42468, w42469, w42470, w42471, w42472, w42473, w42474, w42475, w42476, w42477, w42478, w42479, w42480, w42481, w42482, w42483, w42484, w42485, w42486, w42487, w42488, w42489, w42490, w42491, w42492, w42493, w42494, w42495, w42496, w42497, w42498, w42499, w42500, w42501, w42502, w42503, w42504, w42505, w42506, w42507, w42508, w42509, w42510, w42511, w42512, w42513, w42514, w42515, w42516, w42517, w42518, w42519, w42520, w42521, w42522, w42523, w42524, w42525, w42526, w42527, w42528, w42529, w42530, w42531, w42532, w42533, w42534, w42535, w42536, w42537, w42538, w42539, w42540, w42541, w42542, w42543, w42544, w42545, w42546, w42547, w42548, w42549, w42550, w42551, w42552, w42553, w42554, w42555, w42556, w42557, w42558, w42559, w42560, w42561, w42562, w42563, w42564, w42565, w42566, w42567, w42568, w42569, w42570, w42571, w42572, w42573, w42574, w42575, w42576, w42577, w42578, w42579, w42580, w42581, w42582, w42583, w42584, w42585, w42586, w42587, w42588, w42589, w42590, w42591, w42592, w42593, w42594, w42595, w42596, w42597, w42598, w42599, w42600, w42601, w42602, w42603, w42604, w42605, w42606, w42607, w42608, w42609, w42610, w42611, w42612, w42613, w42614, w42615, w42616, w42617, w42618, w42619, w42620, w42621, w42622, w42623, w42624, w42625, w42626, w42627, w42628, w42629, w42630, w42631, w42632, w42633, w42634, w42635, w42636, w42637, w42638, w42639, w42640, w42641, w42642, w42643, w42644, w42645, w42646, w42647, w42648, w42649, w42650, w42651, w42652, w42653, w42654, w42655, w42656, w42657, w42658, w42659, w42660, w42661, w42662, w42663, w42664, w42665, w42666, w42667, w42668, w42669, w42670, w42671, w42672, w42673, w42674, w42675, w42676, w42677, w42678, w42679, w42680, w42681, w42682, w42683, w42684, w42685, w42686, w42687, w42688, w42689, w42690, w42691, w42692, w42693, w42694, w42695, w42696, w42697, w42698, w42699, w42700, w42701, w42702, w42703, w42704, w42705, w42706, w42707, w42708, w42709, w42710, w42711, w42712, w42713, w42714, w42715, w42716, w42717, w42718, w42719, w42720, w42721, w42722, w42723, w42724, w42725, w42726, w42727, w42728, w42729, w42730, w42731, w42732, w42733, w42734, w42735, w42736, w42737, w42738, w42739, w42740, w42741, w42742, w42743, w42744, w42745, w42746, w42747, w42748, w42749, w42750, w42751, w42752, w42753, w42754, w42755, w42756, w42757, w42758, w42759, w42760, w42761, w42762, w42763, w42764, w42765, w42766, w42767, w42768, w42769, w42770, w42771, w42772, w42773, w42774, w42775, w42776, w42777, w42778, w42779, w42780, w42781, w42782, w42783, w42784, w42785, w42786, w42787, w42788, w42789, w42790, w42791, w42792, w42793, w42794, w42795, w42796, w42797, w42798, w42799, w42800, w42801, w42802, w42803, w42804, w42805, w42806, w42807, w42808, w42809, w42810, w42811, w42812, w42813, w42814, w42815, w42816, w42817, w42818, w42819, w42820, w42821, w42822, w42823, w42824, w42825, w42826, w42827, w42828, w42829, w42830, w42831, w42832, w42833, w42834, w42835, w42836, w42837, w42838, w42839, w42840, w42841, w42842, w42843, w42844, w42845, w42846, w42847, w42848, w42849, w42850, w42851, w42852, w42853, w42854, w42855, w42856, w42857, w42858, w42859, w42860, w42861, w42862, w42863, w42864, w42865, w42866, w42867, w42868, w42869, w42870, w42871, w42872, w42873, w42874, w42875, w42876, w42877, w42878, w42879, w42880, w42881, w42882, w42883, w42884, w42885, w42886, w42887, w42888, w42889, w42890, w42891, w42892, w42893, w42894, w42895, w42896, w42897, w42898, w42899, w42900, w42901, w42902, w42903, w42904, w42905, w42906, w42907, w42908, w42909, w42910, w42911, w42912, w42913, w42914, w42915, w42916, w42917, w42918, w42919, w42920, w42921, w42922, w42923, w42924, w42925, w42926, w42927, w42928, w42929, w42930, w42931, w42932, w42933, w42934, w42935, w42936, w42937, w42938, w42939, w42940, w42941, w42942, w42943, w42944, w42945, w42946, w42947, w42948, w42949, w42950, w42951, w42952, w42953, w42954, w42955, w42956, w42957, w42958, w42959, w42960, w42961, w42962, w42963, w42964, w42965, w42966, w42967, w42968, w42969, w42970, w42971, w42972, w42973, w42974, w42975, w42976, w42977, w42978, w42979, w42980, w42981, w42982, w42983, w42984, w42985, w42986, w42987, w42988, w42989, w42990, w42991, w42992, w42993, w42994, w42995, w42996, w42997, w42998, w42999, w43000, w43001, w43002, w43003, w43004, w43005, w43006, w43007, w43008, w43009, w43010, w43011, w43012, w43013, w43014, w43015, w43016, w43017, w43018, w43019, w43020, w43021, w43022, w43023, w43024, w43025, w43026, w43027, w43028, w43029, w43030, w43031, w43032, w43033, w43034, w43035, w43036, w43037, w43038, w43039, w43040, w43041, w43042, w43043, w43044, w43045, w43046, w43047, w43048, w43049, w43050, w43051, w43052, w43053, w43054, w43055, w43056, w43057, w43058, w43059, w43060, w43061, w43062, w43063, w43064, w43065, w43066, w43067, w43068, w43069, w43070, w43071, w43072, w43073, w43074, w43075, w43076, w43077, w43078, w43079, w43080, w43081, w43082, w43083, w43084, w43085, w43086, w43087, w43088, w43089, w43090, w43091, w43092, w43093, w43094, w43095, w43096, w43097, w43098, w43099, w43100, w43101, w43102, w43103, w43104, w43105, w43106, w43107, w43108, w43109, w43110, w43111, w43112, w43113, w43114, w43115, w43116, w43117, w43118, w43119, w43120, w43121, w43122, w43123, w43124, w43125, w43126, w43127, w43128, w43129, w43130, w43131, w43132, w43133, w43134, w43135, w43136, w43137, w43138, w43139, w43140, w43141, w43142, w43143, w43144, w43145, w43146, w43147, w43148, w43149, w43150, w43151, w43152, w43153, w43154, w43155, w43156, w43157, w43158, w43159, w43160, w43161, w43162, w43163, w43164, w43165, w43166, w43167, w43168, w43169, w43170, w43171, w43172, w43173, w43174, w43175, w43176, w43177, w43178, w43179, w43180, w43181, w43182, w43183, w43184, w43185, w43186, w43187, w43188, w43189, w43190, w43191, w43192, w43193, w43194, w43195, w43196, w43197, w43198, w43199, w43200, w43201, w43202, w43203, w43204, w43205, w43206, w43207, w43208, w43209, w43210, w43211, w43212, w43213, w43214, w43215, w43216, w43217, w43218, w43219, w43220, w43221, w43222, w43223, w43224, w43225, w43226, w43227, w43228, w43229, w43230, w43231, w43232, w43233, w43234, w43235, w43236, w43237, w43238, w43239, w43240, w43241, w43242, w43243, w43244, w43245, w43246, w43247, w43248, w43249, w43250, w43251, w43252, w43253, w43254, w43255, w43256, w43257, w43258, w43259, w43260, w43261, w43262, w43263, w43264, w43265, w43266, w43267, w43268, w43269, w43270, w43271, w43272, w43273, w43274, w43275, w43276, w43277, w43278, w43279, w43280, w43281, w43282, w43283, w43284, w43285, w43286, w43287, w43288, w43289, w43290, w43291, w43292, w43293, w43294, w43295, w43296, w43297, w43298, w43299, w43300, w43301, w43302, w43303, w43304, w43305, w43306, w43307, w43308, w43309, w43310, w43311, w43312, w43313, w43314, w43315, w43316, w43317, w43318, w43319, w43320, w43321, w43322, w43323, w43324, w43325, w43326, w43327, w43328, w43329, w43330, w43331, w43332, w43333, w43334, w43335, w43336, w43337, w43338, w43339, w43340, w43341, w43342, w43343, w43344, w43345, w43346, w43347, w43348, w43349, w43350, w43351, w43352, w43353, w43354, w43355, w43356, w43357, w43358, w43359, w43360, w43361, w43362, w43363, w43364, w43365, w43366, w43367, w43368, w43369, w43370, w43371, w43372, w43373, w43374, w43375, w43376, w43377, w43378, w43379, w43380, w43381, w43382, w43383, w43384, w43385, w43386, w43387, w43388, w43389, w43390, w43391, w43392, w43393, w43394, w43395, w43396, w43397, w43398, w43399, w43400, w43401, w43402, w43403, w43404, w43405, w43406, w43407, w43408, w43409, w43410, w43411, w43412, w43413, w43414, w43415, w43416, w43417, w43418, w43419, w43420, w43421, w43422, w43423, w43424, w43425, w43426, w43427, w43428, w43429, w43430, w43431, w43432, w43433, w43434, w43435, w43436, w43437, w43438, w43439, w43440, w43441, w43442, w43443, w43444, w43445, w43446, w43447, w43448, w43449, w43450, w43451, w43452, w43453, w43454, w43455, w43456, w43457, w43458, w43459, w43460, w43461, w43462, w43463, w43464, w43465, w43466, w43467, w43468, w43469, w43470, w43471, w43472, w43473, w43474, w43475, w43476, w43477, w43478, w43479, w43480, w43481, w43482, w43483, w43484, w43485, w43486, w43487, w43488, w43489, w43490, w43491, w43492, w43493, w43494, w43495, w43496, w43497, w43498, w43499, w43500, w43501, w43502, w43503, w43504, w43505, w43506, w43507, w43508, w43509, w43510, w43511, w43512, w43513, w43514, w43515, w43516, w43517, w43518, w43519, w43520, w43521, w43522, w43523, w43524, w43525, w43526, w43527, w43528, w43529, w43530, w43531, w43532, w43533, w43534, w43535, w43536, w43537, w43538, w43539, w43540, w43541, w43542, w43543, w43544, w43545, w43546, w43547, w43548, w43549, w43550, w43551, w43552, w43553, w43554, w43555, w43556, w43557, w43558, w43559, w43560, w43561, w43562, w43563, w43564, w43565, w43566, w43567, w43568, w43569, w43570, w43571, w43572, w43573, w43574, w43575, w43576, w43577, w43578, w43579, w43580, w43581, w43582, w43583, w43584, w43585, w43586, w43587, w43588, w43589, w43590, w43591, w43592, w43593, w43594, w43595, w43596, w43597, w43598, w43599, w43600, w43601, w43602, w43603, w43604, w43605, w43606, w43607, w43608, w43609, w43610, w43611, w43612, w43613, w43614, w43615, w43616, w43617, w43618, w43619, w43620, w43621, w43622, w43623, w43624, w43625, w43626, w43627, w43628, w43629, w43630, w43631, w43632, w43633, w43634, w43635, w43636, w43637, w43638, w43639, w43640, w43641, w43642, w43643, w43644, w43645, w43646, w43647, w43648, w43649, w43650, w43651, w43652, w43653, w43654, w43655, w43656, w43657, w43658, w43659, w43660, w43661, w43662, w43663, w43664, w43665, w43666, w43667, w43668, w43669, w43670, w43671, w43672, w43673, w43674, w43675, w43676, w43677, w43678, w43679, w43680, w43681, w43682, w43683, w43684, w43685, w43686, w43687, w43688, w43689, w43690, w43691, w43692, w43693, w43694, w43695, w43696, w43697, w43698, w43699, w43700, w43701, w43702, w43703, w43704, w43705, w43706, w43707, w43708, w43709, w43710, w43711, w43712, w43713, w43714, w43715, w43716, w43717, w43718, w43719, w43720, w43721, w43722, w43723, w43724, w43725, w43726, w43727, w43728, w43729, w43730, w43731, w43732, w43733, w43734, w43735, w43736, w43737, w43738, w43739, w43740, w43741, w43742, w43743, w43744, w43745, w43746, w43747, w43748, w43749, w43750, w43751, w43752, w43753, w43754, w43755, w43756, w43757, w43758, w43759, w43760, w43761, w43762, w43763, w43764, w43765, w43766, w43767, w43768, w43769, w43770, w43771, w43772, w43773, w43774, w43775, w43776, w43777, w43778, w43779, w43780, w43781, w43782, w43783, w43784, w43785, w43786, w43787, w43788, w43789, w43790, w43791, w43792, w43793, w43794, w43795, w43796, w43797, w43798, w43799, w43800, w43801, w43802, w43803, w43804, w43805, w43806, w43807, w43808, w43809, w43810, w43811, w43812, w43813, w43814, w43815, w43816, w43817, w43818, w43819, w43820, w43821, w43822, w43823, w43824, w43825, w43826, w43827, w43828, w43829, w43830, w43831, w43832, w43833, w43834, w43835, w43836, w43837, w43838, w43839, w43840, w43841, w43842, w43843, w43844, w43845, w43846, w43847, w43848, w43849, w43850, w43851, w43852, w43853, w43854, w43855, w43856, w43857, w43858, w43859, w43860, w43861, w43862, w43863, w43864, w43865, w43866, w43867, w43868, w43869, w43870, w43871, w43872, w43873, w43874, w43875, w43876, w43877, w43878, w43879, w43880, w43881, w43882, w43883, w43884, w43885, w43886, w43887, w43888, w43889, w43890, w43891, w43892, w43893, w43894, w43895, w43896, w43897, w43898, w43899, w43900, w43901, w43902, w43903, w43904, w43905, w43906, w43907, w43908, w43909, w43910, w43911, w43912, w43913, w43914, w43915, w43916, w43917, w43918, w43919, w43920, w43921, w43922, w43923, w43924, w43925, w43926, w43927, w43928, w43929, w43930, w43931, w43932, w43933, w43934, w43935, w43936, w43937, w43938, w43939, w43940, w43941, w43942, w43943, w43944, w43945, w43946, w43947, w43948, w43949, w43950, w43951, w43952, w43953, w43954, w43955, w43956, w43957, w43958, w43959, w43960, w43961, w43962, w43963, w43964, w43965, w43966, w43967, w43968, w43969, w43970, w43971, w43972, w43973, w43974, w43975, w43976, w43977, w43978, w43979, w43980, w43981, w43982, w43983, w43984, w43985, w43986, w43987, w43988, w43989, w43990, w43991, w43992, w43993, w43994, w43995, w43996, w43997, w43998, w43999, w44000, w44001, w44002, w44003, w44004, w44005, w44006, w44007, w44008, w44009, w44010, w44011, w44012, w44013, w44014, w44015, w44016, w44017, w44018, w44019, w44020, w44021, w44022, w44023, w44024, w44025, w44026, w44027, w44028, w44029, w44030, w44031, w44032, w44033, w44034, w44035, w44036, w44037, w44038, w44039, w44040, w44041, w44042, w44043, w44044, w44045, w44046, w44047, w44048, w44049, w44050, w44051, w44052, w44053, w44054, w44055, w44056, w44057, w44058, w44059, w44060, w44061, w44062, w44063, w44064, w44065, w44066, w44067, w44068, w44069, w44070, w44071, w44072, w44073, w44074, w44075, w44076, w44077, w44078, w44079, w44080, w44081, w44082, w44083, w44084, w44085, w44086, w44087, w44088, w44089, w44090, w44091, w44092, w44093, w44094, w44095, w44096, w44097, w44098, w44099, w44100, w44101, w44102, w44103, w44104, w44105, w44106, w44107, w44108, w44109, w44110, w44111, w44112, w44113, w44114, w44115, w44116, w44117, w44118, w44119, w44120, w44121, w44122, w44123, w44124, w44125, w44126, w44127, w44128, w44129, w44130, w44131, w44132, w44133, w44134, w44135, w44136, w44137, w44138, w44139, w44140, w44141, w44142, w44143, w44144, w44145, w44146, w44147, w44148, w44149, w44150, w44151, w44152, w44153, w44154, w44155, w44156, w44157, w44158, w44159, w44160, w44161, w44162, w44163, w44164, w44165, w44166, w44167, w44168, w44169, w44170, w44171, w44172, w44173, w44174, w44175, w44176, w44177, w44178, w44179, w44180, w44181, w44182, w44183, w44184, w44185, w44186, w44187, w44188, w44189, w44190, w44191, w44192, w44193, w44194, w44195, w44196, w44197, w44198, w44199, w44200, w44201, w44202, w44203, w44204, w44205, w44206, w44207, w44208, w44209, w44210, w44211, w44212, w44213, w44214, w44215, w44216, w44217, w44218, w44219, w44220, w44221, w44222, w44223, w44224, w44225, w44226, w44227, w44228, w44229, w44230, w44231, w44232, w44233, w44234, w44235, w44236, w44237, w44238, w44239, w44240, w44241, w44242, w44243, w44244, w44245, w44246, w44247, w44248, w44249, w44250, w44251, w44252, w44253, w44254, w44255, w44256, w44257, w44258, w44259, w44260, w44261, w44262, w44263, w44264, w44265, w44266, w44267, w44268, w44269, w44270, w44271, w44272, w44273, w44274, w44275, w44276, w44277, w44278, w44279, w44280, w44281, w44282, w44283, w44284, w44285, w44286, w44287, w44288, w44289, w44290, w44291, w44292, w44293, w44294, w44295, w44296, w44297, w44298, w44299, w44300, w44301, w44302, w44303, w44304, w44305, w44306, w44307, w44308, w44309, w44310, w44311, w44312, w44313, w44314, w44315, w44316, w44317, w44318, w44319, w44320, w44321, w44322, w44323, w44324, w44325, w44326, w44327, w44328, w44329, w44330, w44331, w44332, w44333, w44334, w44335, w44336, w44337, w44338, w44339, w44340, w44341, w44342, w44343, w44344, w44345, w44346, w44347, w44348, w44349, w44350, w44351, w44352, w44353, w44354, w44355, w44356, w44357, w44358, w44359, w44360, w44361, w44362, w44363, w44364, w44365, w44366, w44367, w44368, w44369, w44370, w44371, w44372, w44373, w44374, w44375, w44376, w44377, w44378, w44379, w44380, w44381, w44382, w44383, w44384, w44385, w44386, w44387, w44388, w44389, w44390, w44391, w44392, w44393, w44394, w44395, w44396, w44397, w44398, w44399, w44400, w44401, w44402, w44403, w44404, w44405, w44406, w44407, w44408, w44409, w44410, w44411, w44412, w44413, w44414, w44415, w44416, w44417, w44418, w44419, w44420, w44421, w44422, w44423, w44424, w44425, w44426, w44427, w44428, w44429, w44430, w44431, w44432, w44433, w44434, w44435, w44436, w44437, w44438, w44439, w44440, w44441, w44442, w44443, w44444, w44445, w44446, w44447, w44448, w44449, w44450, w44451, w44452, w44453, w44454, w44455, w44456, w44457, w44458, w44459, w44460, w44461, w44462, w44463, w44464, w44465, w44466, w44467, w44468, w44469, w44470, w44471, w44472, w44473, w44474, w44475, w44476, w44477, w44478, w44479, w44480, w44481, w44482, w44483, w44484, w44485, w44486, w44487, w44488, w44489, w44490, w44491, w44492, w44493, w44494, w44495, w44496, w44497, w44498, w44499, w44500, w44501, w44502, w44503, w44504, w44505, w44506, w44507, w44508, w44509, w44510, w44511, w44512, w44513, w44514, w44515, w44516, w44517, w44518, w44519, w44520, w44521, w44522, w44523, w44524, w44525, w44526, w44527, w44528, w44529, w44530, w44531, w44532, w44533, w44534, w44535, w44536, w44537, w44538, w44539, w44540, w44541, w44542, w44543, w44544, w44545, w44546, w44547, w44548, w44549, w44550, w44551, w44552, w44553, w44554, w44555, w44556, w44557, w44558, w44559, w44560, w44561, w44562, w44563, w44564, w44565, w44566, w44567, w44568, w44569, w44570, w44571, w44572, w44573, w44574, w44575, w44576, w44577, w44578, w44579, w44580, w44581, w44582, w44583, w44584, w44585, w44586, w44587, w44588, w44589, w44590, w44591, w44592, w44593, w44594, w44595, w44596, w44597, w44598, w44599, w44600, w44601, w44602, w44603, w44604, w44605, w44606, w44607, w44608, w44609, w44610, w44611, w44612, w44613, w44614, w44615, w44616, w44617, w44618, w44619, w44620, w44621, w44622, w44623, w44624, w44625, w44626, w44627, w44628, w44629, w44630, w44631, w44632, w44633, w44634, w44635, w44636, w44637, w44638, w44639, w44640, w44641, w44642, w44643, w44644, w44645, w44646, w44647, w44648, w44649, w44650, w44651, w44652, w44653, w44654, w44655, w44656, w44657, w44658, w44659, w44660, w44661, w44662, w44663, w44664, w44665, w44666, w44667, w44668, w44669, w44670, w44671, w44672, w44673, w44674, w44675, w44676, w44677, w44678, w44679, w44680, w44681, w44682, w44683, w44684, w44685, w44686, w44687, w44688, w44689, w44690, w44691, w44692, w44693, w44694, w44695, w44696, w44697, w44698, w44699, w44700, w44701, w44702, w44703, w44704, w44705, w44706, w44707, w44708, w44709, w44710, w44711, w44712, w44713, w44714, w44715, w44716, w44717, w44718, w44719, w44720, w44721, w44722, w44723, w44724, w44725, w44726, w44727, w44728, w44729, w44730, w44731, w44732, w44733, w44734, w44735, w44736, w44737, w44738, w44739, w44740, w44741, w44742, w44743, w44744, w44745, w44746, w44747, w44748, w44749, w44750, w44751, w44752, w44753, w44754, w44755, w44756, w44757, w44758, w44759, w44760, w44761, w44762, w44763, w44764, w44765, w44766, w44767, w44768, w44769, w44770, w44771, w44772, w44773, w44774, w44775, w44776, w44777, w44778, w44779, w44780, w44781, w44782, w44783, w44784, w44785, w44786, w44787, w44788, w44789, w44790, w44791, w44792, w44793, w44794, w44795, w44796, w44797, w44798, w44799, w44800, w44801, w44802, w44803, w44804, w44805, w44806, w44807, w44808, w44809, w44810, w44811, w44812, w44813, w44814, w44815, w44816, w44817, w44818, w44819, w44820, w44821, w44822, w44823, w44824, w44825, w44826, w44827, w44828, w44829, w44830, w44831, w44832, w44833, w44834, w44835, w44836, w44837, w44838, w44839, w44840, w44841, w44842, w44843, w44844, w44845, w44846, w44847, w44848, w44849, w44850, w44851, w44852, w44853, w44854, w44855, w44856, w44857, w44858, w44859, w44860, w44861, w44862, w44863, w44864, w44865, w44866, w44867, w44868, w44869, w44870, w44871, w44872, w44873, w44874, w44875, w44876, w44877, w44878, w44879, w44880, w44881, w44882, w44883, w44884, w44885, w44886, w44887, w44888, w44889, w44890, w44891, w44892, w44893, w44894, w44895, w44896, w44897, w44898, w44899, w44900, w44901, w44902, w44903, w44904, w44905, w44906, w44907, w44908, w44909, w44910, w44911, w44912, w44913, w44914, w44915, w44916, w44917, w44918, w44919, w44920, w44921, w44922, w44923, w44924, w44925, w44926, w44927, w44928, w44929, w44930, w44931, w44932, w44933, w44934, w44935, w44936, w44937, w44938, w44939, w44940, w44941, w44942, w44943, w44944, w44945, w44946, w44947, w44948, w44949, w44950, w44951, w44952, w44953, w44954, w44955, w44956, w44957, w44958, w44959, w44960, w44961, w44962, w44963, w44964, w44965, w44966, w44967, w44968, w44969, w44970, w44971, w44972, w44973, w44974, w44975, w44976, w44977, w44978, w44979, w44980, w44981, w44982, w44983, w44984, w44985, w44986, w44987, w44988, w44989, w44990, w44991, w44992, w44993, w44994, w44995, w44996, w44997, w44998, w44999, w45000, w45001, w45002, w45003, w45004, w45005, w45006, w45007, w45008, w45009, w45010, w45011, w45012, w45013, w45014, w45015, w45016, w45017, w45018, w45019, w45020, w45021, w45022, w45023, w45024, w45025, w45026, w45027, w45028, w45029, w45030, w45031, w45032, w45033, w45034, w45035, w45036, w45037, w45038, w45039, w45040, w45041, w45042, w45043, w45044, w45045, w45046, w45047, w45048, w45049, w45050, w45051, w45052, w45053, w45054, w45055, w45056, w45057, w45058, w45059, w45060, w45061, w45062, w45063, w45064, w45065, w45066, w45067, w45068, w45069, w45070, w45071, w45072, w45073, w45074, w45075, w45076, w45077, w45078, w45079, w45080, w45081, w45082, w45083, w45084, w45085, w45086, w45087, w45088, w45089, w45090, w45091, w45092, w45093, w45094, w45095, w45096, w45097, w45098, w45099, w45100, w45101, w45102, w45103, w45104, w45105, w45106, w45107, w45108, w45109, w45110, w45111, w45112, w45113, w45114, w45115, w45116, w45117, w45118, w45119, w45120, w45121, w45122, w45123, w45124, w45125, w45126, w45127, w45128, w45129, w45130, w45131, w45132, w45133, w45134, w45135, w45136, w45137, w45138, w45139, w45140, w45141, w45142, w45143, w45144, w45145, w45146, w45147, w45148, w45149, w45150, w45151, w45152, w45153, w45154, w45155, w45156, w45157, w45158, w45159, w45160, w45161, w45162, w45163, w45164, w45165, w45166, w45167, w45168, w45169, w45170, w45171, w45172, w45173, w45174, w45175, w45176, w45177, w45178, w45179, w45180, w45181, w45182, w45183, w45184, w45185, w45186, w45187, w45188, w45189, w45190, w45191, w45192, w45193, w45194, w45195, w45196, w45197, w45198, w45199, w45200, w45201, w45202, w45203, w45204, w45205, w45206, w45207, w45208, w45209, w45210, w45211, w45212, w45213, w45214, w45215, w45216, w45217, w45218, w45219, w45220, w45221, w45222, w45223, w45224, w45225, w45226, w45227, w45228, w45229, w45230, w45231, w45232, w45233, w45234, w45235, w45236, w45237, w45238, w45239, w45240, w45241, w45242, w45243, w45244, w45245, w45246, w45247, w45248, w45249, w45250, w45251, w45252, w45253, w45254, w45255, w45256, w45257, w45258, w45259, w45260, w45261, w45262, w45263, w45264, w45265, w45266, w45267, w45268, w45269, w45270, w45271, w45272, w45273, w45274, w45275, w45276, w45277, w45278, w45279, w45280, w45281, w45282, w45283, w45284, w45285, w45286, w45287, w45288, w45289, w45290, w45291, w45292, w45293, w45294, w45295, w45296, w45297, w45298, w45299, w45300, w45301, w45302, w45303, w45304, w45305, w45306, w45307, w45308, w45309, w45310, w45311, w45312, w45313, w45314, w45315, w45316, w45317, w45318, w45319, w45320, w45321, w45322, w45323, w45324, w45325, w45326, w45327, w45328, w45329, w45330, w45331, w45332, w45333, w45334, w45335, w45336, w45337, w45338, w45339, w45340, w45341, w45342, w45343, w45344, w45345, w45346, w45347, w45348, w45349, w45350, w45351, w45352, w45353, w45354, w45355, w45356, w45357, w45358, w45359, w45360, w45361, w45362, w45363, w45364, w45365, w45366, w45367, w45368, w45369, w45370, w45371, w45372, w45373, w45374, w45375, w45376, w45377, w45378, w45379, w45380, w45381, w45382, w45383, w45384, w45385, w45386, w45387, w45388, w45389, w45390, w45391, w45392, w45393, w45394, w45395, w45396, w45397, w45398, w45399, w45400, w45401, w45402, w45403, w45404, w45405, w45406, w45407, w45408, w45409, w45410, w45411, w45412, w45413, w45414, w45415, w45416, w45417, w45418, w45419, w45420, w45421, w45422, w45423, w45424, w45425, w45426, w45427, w45428, w45429, w45430, w45431, w45432, w45433, w45434, w45435, w45436, w45437, w45438, w45439, w45440, w45441, w45442, w45443, w45444, w45445, w45446, w45447, w45448, w45449, w45450, w45451, w45452, w45453, w45454, w45455, w45456, w45457, w45458, w45459, w45460, w45461, w45462, w45463, w45464, w45465, w45466, w45467, w45468, w45469, w45470, w45471, w45472, w45473, w45474, w45475, w45476, w45477, w45478, w45479, w45480, w45481, w45482, w45483, w45484, w45485, w45486, w45487, w45488, w45489, w45490, w45491, w45492, w45493, w45494, w45495, w45496, w45497, w45498, w45499, w45500, w45501, w45502, w45503, w45504, w45505, w45506, w45507, w45508, w45509, w45510, w45511, w45512, w45513, w45514, w45515, w45516, w45517, w45518, w45519, w45520, w45521, w45522, w45523, w45524, w45525, w45526, w45527, w45528, w45529, w45530, w45531, w45532, w45533, w45534, w45535, w45536, w45537, w45538, w45539, w45540, w45541, w45542, w45543, w45544, w45545, w45546, w45547, w45548, w45549, w45550, w45551, w45552, w45553, w45554, w45555, w45556, w45557, w45558, w45559, w45560, w45561, w45562, w45563, w45564, w45565, w45566, w45567, w45568, w45569, w45570, w45571, w45572, w45573, w45574, w45575, w45576, w45577, w45578, w45579, w45580, w45581, w45582, w45583, w45584, w45585, w45586, w45587, w45588, w45589, w45590, w45591, w45592, w45593, w45594, w45595, w45596, w45597, w45598, w45599, w45600, w45601, w45602, w45603, w45604, w45605, w45606, w45607, w45608, w45609, w45610, w45611, w45612, w45613, w45614, w45615, w45616, w45617, w45618, w45619, w45620, w45621, w45622, w45623, w45624, w45625, w45626, w45627, w45628, w45629, w45630, w45631, w45632, w45633, w45634, w45635, w45636, w45637, w45638, w45639, w45640, w45641, w45642, w45643, w45644, w45645, w45646, w45647, w45648, w45649, w45650, w45651, w45652, w45653, w45654, w45655, w45656, w45657, w45658, w45659, w45660, w45661, w45662, w45663, w45664, w45665, w45666, w45667, w45668, w45669, w45670, w45671, w45672, w45673, w45674, w45675, w45676, w45677, w45678, w45679, w45680, w45681, w45682, w45683, w45684, w45685, w45686, w45687, w45688, w45689, w45690, w45691, w45692, w45693, w45694, w45695, w45696, w45697, w45698, w45699, w45700, w45701, w45702, w45703, w45704, w45705, w45706, w45707, w45708, w45709, w45710, w45711, w45712, w45713, w45714, w45715, w45716, w45717, w45718, w45719, w45720, w45721, w45722, w45723, w45724, w45725, w45726, w45727, w45728, w45729, w45730, w45731, w45732, w45733, w45734, w45735, w45736, w45737, w45738, w45739, w45740, w45741, w45742, w45743, w45744, w45745, w45746, w45747, w45748, w45749, w45750, w45751, w45752, w45753, w45754, w45755, w45756, w45757, w45758, w45759, w45760, w45761, w45762, w45763, w45764, w45765, w45766, w45767, w45768, w45769, w45770, w45771, w45772, w45773, w45774, w45775, w45776, w45777, w45778, w45779, w45780, w45781, w45782, w45783, w45784, w45785, w45786, w45787, w45788, w45789, w45790, w45791, w45792, w45793, w45794, w45795, w45796, w45797, w45798, w45799, w45800, w45801, w45802, w45803, w45804, w45805, w45806, w45807, w45808, w45809, w45810, w45811, w45812, w45813, w45814, w45815, w45816, w45817, w45818, w45819, w45820, w45821, w45822, w45823, w45824, w45825, w45826, w45827, w45828, w45829, w45830, w45831, w45832, w45833, w45834, w45835, w45836, w45837, w45838, w45839, w45840, w45841, w45842, w45843, w45844, w45845, w45846, w45847, w45848, w45849, w45850, w45851, w45852, w45853, w45854, w45855, w45856, w45857, w45858, w45859, w45860, w45861, w45862, w45863, w45864, w45865, w45866, w45867, w45868, w45869, w45870, w45871, w45872, w45873, w45874, w45875, w45876, w45877, w45878, w45879, w45880, w45881, w45882, w45883, w45884, w45885, w45886, w45887, w45888, w45889, w45890, w45891, w45892, w45893, w45894, w45895, w45896, w45897, w45898, w45899, w45900, w45901, w45902, w45903, w45904, w45905, w45906, w45907, w45908, w45909, w45910, w45911, w45912, w45913, w45914, w45915, w45916, w45917, w45918, w45919, w45920, w45921, w45922, w45923, w45924, w45925, w45926, w45927, w45928, w45929, w45930, w45931, w45932, w45933, w45934, w45935, w45936, w45937, w45938, w45939, w45940, w45941, w45942, w45943, w45944, w45945, w45946, w45947, w45948, w45949, w45950, w45951, w45952, w45953, w45954, w45955, w45956, w45957, w45958, w45959, w45960, w45961, w45962, w45963, w45964, w45965, w45966, w45967, w45968, w45969, w45970, w45971, w45972, w45973, w45974, w45975, w45976, w45977, w45978, w45979, w45980, w45981, w45982, w45983, w45984, w45985, w45986, w45987, w45988, w45989, w45990, w45991, w45992, w45993, w45994, w45995, w45996, w45997, w45998, w45999, w46000, w46001, w46002, w46003, w46004, w46005, w46006, w46007, w46008, w46009, w46010, w46011, w46012, w46013, w46014, w46015, w46016, w46017, w46018, w46019, w46020, w46021, w46022, w46023, w46024, w46025, w46026, w46027, w46028, w46029, w46030, w46031, w46032, w46033, w46034, w46035, w46036, w46037, w46038, w46039, w46040, w46041, w46042, w46043, w46044, w46045, w46046, w46047, w46048, w46049, w46050, w46051, w46052, w46053, w46054, w46055, w46056, w46057, w46058, w46059, w46060, w46061, w46062, w46063, w46064, w46065, w46066, w46067, w46068, w46069, w46070, w46071, w46072, w46073, w46074, w46075, w46076, w46077, w46078, w46079, w46080, w46081, w46082, w46083, w46084, w46085, w46086, w46087, w46088, w46089, w46090, w46091, w46092, w46093, w46094, w46095, w46096, w46097, w46098, w46099, w46100, w46101, w46102, w46103, w46104, w46105, w46106, w46107, w46108, w46109, w46110, w46111, w46112, w46113, w46114, w46115, w46116, w46117, w46118, w46119, w46120, w46121, w46122, w46123, w46124, w46125, w46126, w46127, w46128, w46129, w46130, w46131, w46132, w46133, w46134, w46135, w46136, w46137, w46138, w46139, w46140, w46141, w46142, w46143, w46144, w46145, w46146, w46147, w46148, w46149, w46150, w46151, w46152, w46153, w46154, w46155, w46156, w46157, w46158, w46159, w46160, w46161, w46162, w46163, w46164, w46165, w46166, w46167, w46168, w46169, w46170, w46171, w46172, w46173, w46174, w46175, w46176, w46177, w46178, w46179, w46180, w46181, w46182, w46183, w46184, w46185, w46186, w46187, w46188, w46189, w46190, w46191, w46192, w46193, w46194, w46195, w46196, w46197, w46198, w46199, w46200, w46201, w46202, w46203, w46204, w46205, w46206, w46207, w46208, w46209, w46210, w46211, w46212, w46213, w46214, w46215, w46216, w46217, w46218, w46219, w46220, w46221, w46222, w46223, w46224, w46225, w46226, w46227, w46228, w46229, w46230, w46231, w46232, w46233, w46234, w46235, w46236, w46237, w46238, w46239, w46240, w46241, w46242, w46243, w46244, w46245, w46246, w46247, w46248, w46249, w46250, w46251, w46252, w46253, w46254, w46255, w46256, w46257, w46258, w46259, w46260, w46261, w46262, w46263, w46264, w46265, w46266, w46267, w46268, w46269, w46270, w46271, w46272, w46273, w46274, w46275, w46276, w46277, w46278, w46279, w46280, w46281, w46282, w46283, w46284, w46285, w46286, w46287, w46288, w46289, w46290, w46291, w46292, w46293, w46294, w46295, w46296, w46297, w46298, w46299, w46300, w46301, w46302, w46303, w46304, w46305, w46306, w46307, w46308, w46309, w46310, w46311, w46312, w46313, w46314, w46315, w46316, w46317, w46318, w46319, w46320, w46321, w46322, w46323, w46324, w46325, w46326, w46327, w46328, w46329, w46330, w46331, w46332, w46333, w46334, w46335, w46336, w46337, w46338, w46339, w46340, w46341, w46342, w46343, w46344, w46345, w46346, w46347, w46348, w46349, w46350, w46351, w46352, w46353, w46354, w46355, w46356, w46357, w46358, w46359, w46360, w46361, w46362, w46363, w46364, w46365, w46366, w46367, w46368, w46369, w46370, w46371, w46372, w46373, w46374, w46375, w46376, w46377, w46378, w46379, w46380, w46381, w46382, w46383, w46384, w46385, w46386, w46387, w46388, w46389, w46390, w46391, w46392, w46393, w46394, w46395, w46396, w46397, w46398, w46399, w46400, w46401, w46402, w46403, w46404, w46405, w46406, w46407, w46408, w46409, w46410, w46411, w46412, w46413, w46414, w46415, w46416, w46417, w46418, w46419, w46420, w46421, w46422, w46423, w46424, w46425, w46426, w46427, w46428, w46429, w46430, w46431, w46432, w46433, w46434, w46435, w46436, w46437, w46438, w46439, w46440, w46441, w46442, w46443, w46444, w46445, w46446, w46447, w46448, w46449, w46450, w46451, w46452, w46453, w46454, w46455, w46456, w46457, w46458, w46459, w46460, w46461, w46462, w46463, w46464, w46465, w46466, w46467, w46468, w46469, w46470, w46471, w46472, w46473, w46474, w46475, w46476, w46477, w46478, w46479, w46480, w46481, w46482, w46483, w46484, w46485, w46486, w46487, w46488, w46489, w46490, w46491, w46492, w46493, w46494, w46495, w46496, w46497, w46498, w46499, w46500, w46501, w46502, w46503, w46504, w46505, w46506, w46507, w46508, w46509, w46510, w46511, w46512, w46513, w46514, w46515, w46516, w46517, w46518, w46519, w46520, w46521, w46522, w46523, w46524, w46525, w46526, w46527, w46528, w46529, w46530, w46531, w46532, w46533, w46534, w46535, w46536, w46537, w46538, w46539, w46540, w46541, w46542, w46543, w46544, w46545, w46546, w46547, w46548, w46549, w46550, w46551, w46552, w46553, w46554, w46555, w46556, w46557, w46558, w46559, w46560, w46561, w46562, w46563, w46564, w46565, w46566, w46567, w46568, w46569, w46570, w46571, w46572, w46573, w46574, w46575, w46576, w46577, w46578, w46579, w46580, w46581, w46582, w46583, w46584, w46585, w46586, w46587, w46588, w46589, w46590, w46591, w46592, w46593, w46594, w46595, w46596, w46597, w46598, w46599, w46600, w46601, w46602, w46603, w46604, w46605, w46606, w46607, w46608, w46609, w46610, w46611, w46612, w46613, w46614, w46615, w46616, w46617, w46618, w46619, w46620, w46621, w46622, w46623, w46624, w46625, w46626, w46627, w46628, w46629, w46630, w46631, w46632, w46633, w46634, w46635, w46636, w46637, w46638, w46639, w46640, w46641, w46642, w46643, w46644, w46645, w46646, w46647, w46648, w46649, w46650, w46651, w46652, w46653, w46654, w46655, w46656, w46657, w46658, w46659, w46660, w46661, w46662, w46663, w46664, w46665, w46666, w46667, w46668, w46669, w46670, w46671, w46672, w46673, w46674, w46675, w46676, w46677, w46678, w46679, w46680, w46681, w46682, w46683, w46684, w46685, w46686, w46687, w46688, w46689, w46690, w46691, w46692, w46693, w46694, w46695, w46696, w46697, w46698, w46699, w46700, w46701, w46702, w46703, w46704, w46705, w46706, w46707, w46708, w46709, w46710, w46711, w46712, w46713, w46714, w46715, w46716, w46717, w46718, w46719, w46720, w46721, w46722, w46723, w46724, w46725, w46726, w46727, w46728, w46729, w46730, w46731, w46732, w46733, w46734, w46735, w46736, w46737, w46738, w46739, w46740, w46741, w46742, w46743, w46744, w46745, w46746, w46747, w46748, w46749, w46750, w46751, w46752, w46753, w46754, w46755, w46756, w46757, w46758, w46759, w46760, w46761, w46762, w46763, w46764, w46765, w46766, w46767, w46768, w46769, w46770, w46771, w46772, w46773, w46774, w46775, w46776, w46777, w46778, w46779, w46780, w46781, w46782, w46783, w46784, w46785, w46786, w46787, w46788, w46789, w46790, w46791, w46792, w46793, w46794, w46795, w46796, w46797, w46798, w46799, w46800, w46801, w46802, w46803, w46804, w46805, w46806, w46807, w46808, w46809, w46810, w46811, w46812, w46813, w46814, w46815, w46816, w46817, w46818, w46819, w46820, w46821, w46822, w46823, w46824, w46825, w46826, w46827, w46828, w46829, w46830, w46831, w46832, w46833, w46834, w46835: std_logic;

begin

w0 <= not pi0332 and not pi1144;
w1 <= pi0215 and not w0;
w2 <= pi0265 and not pi0332;
w3 <= pi0216 and not w2;
w4 <= pi0105 and pi0228;
w5 <= pi0095 and not pi0479;
w6 <= pi0234 and w5;
w7 <= not pi0332 and not w6;
w8 <= w4 and w7;
w9 <= pi0153 and not pi0332;
w10 <= not w4 and w9;
w11 <= not pi0216 and not w10;
w12 <= not w8 and w11;
w13 <= not w3 and not w12;
w14 <= not pi0221 and not w13;
w15 <= not pi0216 and pi0833;
w16 <= pi1144 and not w15;
w17 <= pi0929 and w15;
w18 <= not pi0332 and not w16;
w19 <= not w17 and w18;
w20 <= pi0221 and not w19;
w21 <= not w14 and not w20;
w22 <= not pi0215 and not w21;
w23 <= not w1 and not w22;
w24 <= not pi0058 and not pi0090;
w25 <= not pi0088 and not pi0098;
w26 <= not pi0077 and w25;
w27 <= not pi0050 and w26;
w28 <= not pi0102 and w27;
w29 <= not pi0065 and not pi0071;
w30 <= not pi0083 and not pi0103;
w31 <= not pi0067 and not pi0069;
w32 <= not pi0066 and not pi0073;
w33 <= not pi0061 and not pi0076;
w34 <= not pi0085 and not pi0106;
w35 <= w33 and w34;
w36 <= not pi0048 and w35;
w37 <= not pi0089 and w36;
w38 <= not pi0049 and w37;
w39 <= not pi0104 and w38;
w40 <= not pi0045 and w39;
w41 <= not pi0068 and not pi0084;
w42 <= not pi0082 and not pi0111;
w43 <= not pi0036 and w42;
w44 <= w41 and w43;
w45 <= w40 and w44;
w46 <= w32 and w45;
w47 <= w31 and w46;
w48 <= w30 and w47;
w49 <= w29 and w48;
w50 <= not pi0063 and not pi0107;
w51 <= w49 and w50;
w52 <= not pi0064 and w51;
w53 <= not pi0081 and w52;
w54 <= w28 and w53;
w55 <= not pi0047 and not pi0091;
w56 <= not pi0109 and not pi0110;
w57 <= not pi0053 and not pi0060;
w58 <= not pi0086 and w57;
w59 <= not pi0097 and not pi0108;
w60 <= not pi0094 and w59;
w61 <= not pi0046 and w58;
w62 <= w60 and w61;
w63 <= w56 and w62;
w64 <= w55 and w63;
w65 <= w54 and w64;
w66 <= w24 and w65;
w67 <= not pi0035 and not pi0093;
w68 <= w66 and w67;
w69 <= not pi0072 and not pi0096;
w70 <= not pi0051 and not pi0070;
w71 <= w69 and w70;
w72 <= w68 and w71;
w73 <= not pi0032 and not pi0040;
w74 <= w72 and w73;
w75 <= not pi0095 and w74;
w76 <= not w5 and not w75;
w77 <= pi0234 and not w76;
w78 <= not pi0070 and w68;
w79 <= not pi0051 and not pi0096;
w80 <= not pi0040 and not pi0072;
w81 <= not pi0032 and not pi0095;
w82 <= w80 and w81;
w83 <= w79 and w82;
w84 <= w78 and w83;
w85 <= not pi0234 and w84;
w86 <= not w77 and not w85;
w87 <= pi0137 and not w86;
w88 <= w7 and not w87;
w89 <= not pi0215 and not pi0221;
w90 <= w11 and w89;
w91 <= not w88 and w90;
w92 <= not pi0056 and not pi0062;
w93 <= not pi0038 and not pi0039;
w94 <= not pi0100 and w93;
w95 <= not pi0054 and not pi0074;
w96 <= not pi0075 and not pi0087;
w97 <= not pi0092 and w96;
w98 <= w95 and w97;
w99 <= not pi0055 and w98;
w100 <= w94 and w99;
w101 <= w92 and w100;
w102 <= w91 and w101;
w103 <= pi0059 and w23;
w104 <= not w102 and w103;
w105 <= w23 and not w100;
w106 <= not pi0105 and not w9;
w107 <= pi0105 and not w88;
w108 <= not w106 and not w107;
w109 <= pi0228 and not w108;
w110 <= pi0137 and w84;
w111 <= w9 and not w110;
w112 <= not pi0332 and w75;
w113 <= not pi0137 and not pi0153;
w114 <= w112 and w113;
w115 <= not pi0228 and not w111;
w116 <= not w114 and w115;
w117 <= not w109 and not w116;
w118 <= not pi0216 and not w117;
w119 <= not w3 and not w118;
w120 <= not pi0221 and not w119;
w121 <= not w20 and not w120;
w122 <= not pi0215 and not w121;
w123 <= not w1 and not w122;
w124 <= w100 and w123;
w125 <= not w105 and not w124;
w126 <= not pi0056 and not w125;
w127 <= pi0056 and w23;
w128 <= pi0062 and not w127;
w129 <= not w126 and w128;
w130 <= pi0056 and not w125;
w131 <= not pi0087 and not pi0100;
w132 <= not pi0075 and not pi0092;
w133 <= w95 and w132;
w134 <= w131 and w133;
w135 <= w93 and w134;
w136 <= w23 and not w135;
w137 <= pi0228 and not w106;
w138 <= not pi0332 and w86;
w139 <= pi0105 and not w138;
w140 <= w137 and not w139;
w141 <= not pi0228 and w9;
w142 <= not w84 and w141;
w143 <= not pi0216 and not w142;
w144 <= not w140 and w143;
w145 <= not w3 and not w144;
w146 <= not pi0221 and not w145;
w147 <= not w20 and not w146;
w148 <= not pi0215 and not w147;
w149 <= not w1 and w135;
w150 <= not w148 and w149;
w151 <= pi0055 and not w136;
w152 <= not w150 and w151;
w153 <= pi0299 and w23;
w154 <= not pi0224 and pi0833;
w155 <= pi0222 and not w154;
w156 <= not pi0223 and not w155;
w157 <= w0 and not w156;
w158 <= pi0224 and not w2;
w159 <= not pi0222 and not w158;
w160 <= not pi0332 and not pi0929;
w161 <= w154 and w160;
w162 <= not w159 and not w161;
w163 <= not pi0223 and not w162;
w164 <= not w157 and not w163;
w165 <= not pi0299 and not w164;
w166 <= not pi0222 and not pi0224;
w167 <= not pi0223 and w166;
w168 <= not w7 and w167;
w169 <= w165 and not w168;
w170 <= not w153 and not w169;
w171 <= not pi0038 and not pi0100;
w172 <= not pi0039 and not pi0087;
w173 <= w171 and w172;
w174 <= w132 and w173;
w175 <= w170 and not w174;
w176 <= not w88 and w167;
w177 <= not w164 and not w176;
w178 <= not pi0299 and not w177;
w179 <= w23 and not w91;
w180 <= pi0299 and not w179;
w181 <= not w178 and not w180;
w182 <= not pi0039 and not w181;
w183 <= not pi0038 and w131;
w184 <= w132 and w183;
w185 <= w182 and w184;
w186 <= not w175 and not w185;
w187 <= pi0054 and w186;
w188 <= not pi0039 and w171;
w189 <= not w170 and not w188;
w190 <= pi0299 and not w123;
w191 <= not w178 and not w190;
w192 <= w188 and w191;
w193 <= not w189 and not w192;
w194 <= w96 and not w193;
w195 <= not w96 and not w170;
w196 <= pi0092 and not w195;
w197 <= not w194 and w196;
w198 <= pi0087 and not w193;
w199 <= not w93 and not w170;
w200 <= pi0095 and pi0234;
w201 <= not pi0152 and not pi0161;
w202 <= not pi0166 and w201;
w203 <= not pi0146 and not w202;
w204 <= not pi0210 and not w203;
w205 <= not pi0137 and not w200;
w206 <= not w204 and w205;
w207 <= not w86 and not w206;
w208 <= not pi0332 and not w207;
w209 <= pi0105 and not w208;
w210 <= w137 and not w209;
w211 <= w110 and w203;
w212 <= not pi0137 and pi0210;
w213 <= not pi0252 and not w212;
w214 <= not w203 and w213;
w215 <= w112 and w214;
w216 <= w9 and not w211;
w217 <= not w215 and w216;
w218 <= pi0252 and not w203;
w219 <= not w204 and not w218;
w220 <= w114 and w219;
w221 <= not w217 and not w220;
w222 <= not pi0228 and not w221;
w223 <= not pi0216 and not w222;
w224 <= not w210 and w223;
w225 <= not w3 and not w224;
w226 <= not pi0221 and not w225;
w227 <= not w20 and not w226;
w228 <= not pi0215 and not w227;
w229 <= not w1 and not w228;
w230 <= pi0299 and not w229;
w231 <= not pi0144 and not pi0174;
w232 <= not pi0189 and w231;
w233 <= not pi0223 and not w232;
w234 <= pi0142 and not pi0198;
w235 <= not pi0137 and not w234;
w236 <= not w86 and not w235;
w237 <= w7 and not w236;
w238 <= w233 and not w237;
w239 <= not pi0234 and not pi0332;
w240 <= not pi0137 and pi0198;
w241 <= w84 and not w240;
w242 <= w239 and not w241;
w243 <= not pi0223 and w232;
w244 <= pi0234 and not pi0332;
w245 <= not pi0095 and w240;
w246 <= not w76 and not w245;
w247 <= w244 and not w246;
w248 <= not w242 and w243;
w249 <= not w247 and w248;
w250 <= not w238 and not w249;
w251 <= w166 and not w250;
w252 <= not w164 and not w251;
w253 <= not pi0299 and not w252;
w254 <= w93 and not w253;
w255 <= not w230 and w254;
w256 <= pi0100 and not w199;
w257 <= not w255 and w256;
w258 <= pi0039 and w170;
w259 <= pi0038 and not w258;
w260 <= not w182 and w259;
w261 <= pi0039 and not w191;
w262 <= w54 and w62;
w263 <= not pi0058 and not pi0091;
w264 <= not pi0047 and w263;
w265 <= w56 and w264;
w266 <= w262 and w265;
w267 <= not pi0090 and not pi0093;
w268 <= not pi0070 and not pi0096;
w269 <= not pi0035 and not pi0051;
w270 <= w268 and w269;
w271 <= w267 and w270;
w272 <= w266 and w271;
w273 <= w80 and w272;
w274 <= pi0225 and w273;
w275 <= pi0032 and not w274;
w276 <= not pi0095 and not w275;
w277 <= not pi0046 and w56;
w278 <= w55 and w59;
w279 <= w277 and w278;
w280 <= not pi0058 and w279;
w281 <= pi0060 and w54;
w282 <= not pi0053 and not w281;
w283 <= not pi0086 and not pi0094;
w284 <= not pi0060 and w54;
w285 <= pi0053 and not w284;
w286 <= w283 and not w285;
w287 <= not w282 and w286;
w288 <= w267 and w280;
w289 <= w287 and w288;
w290 <= not pi0035 and not w289;
w291 <= not pi0093 and w66;
w292 <= pi0035 and not w291;
w293 <= pi0035 and w291;
w294 <= not pi0225 and w293;
w295 <= not pi0070 and not w294;
w296 <= not pi0051 and w295;
w297 <= not w292 and w296;
w298 <= not w290 and w297;
w299 <= not pi0040 and w69;
w300 <= w298 and w299;
w301 <= not pi0032 and not w300;
w302 <= w276 and not w301;
w303 <= not pi0137 and not w302;
w304 <= pi0095 and not w74;
w305 <= not w5 and not w304;
w306 <= pi0040 and w72;
w307 <= not pi0032 and not w306;
w308 <= pi0072 and not w272;
w309 <= not pi0040 and not w308;
w310 <= pi0051 and not w78;
w311 <= not pi0096 and not w310;
w312 <= not pi0051 and pi0070;
w313 <= w311 and not w312;
w314 <= not w292 and not w294;
w315 <= pi0093 and w66;
w316 <= not pi0035 and not w315;
w317 <= not pi0047 and w63;
w318 <= w54 and w317;
w319 <= pi0091 and w318;
w320 <= w24 and not w319;
w321 <= not pi0109 and w262;
w322 <= pi0110 and not w321;
w323 <= pi0047 and w54;
w324 <= w63 and w323;
w325 <= pi0047 and not w324;
w326 <= not pi0091 and not w325;
w327 <= not w322 and w326;
w328 <= not pi0047 and not pi0110;
w329 <= pi0109 and not w262;
w330 <= not pi0102 and w53;
w331 <= w25 and w330;
w332 <= not pi0050 and w57;
w333 <= not pi0077 and w332;
w334 <= w283 and w333;
w335 <= w331 and w334;
w336 <= not pi0097 and w335;
w337 <= pi0108 and not w336;
w338 <= not pi0046 and not w337;
w339 <= pi0097 and not w335;
w340 <= w26 and w330;
w341 <= w332 and w340;
w342 <= not pi0086 and pi0094;
w343 <= w341 and w342;
w344 <= not pi0097 and not w343;
w345 <= pi0086 and not w341;
w346 <= not pi0094 and not w345;
w347 <= pi0077 and w331;
w348 <= not pi0050 and not w347;
w349 <= pi0081 and not w52;
w350 <= pi0102 and not w53;
w351 <= not w349 and not w350;
w352 <= pi0064 and not w51;
w353 <= pi0071 and not w48;
w354 <= not pi0065 and not w353;
w355 <= not pi0067 and w46;
w356 <= pi0069 and not w355;
w357 <= pi0083 and not w47;
w358 <= not pi0103 and not w357;
w359 <= not w356 and w358;
w360 <= not pi0069 and not pi0083;
w361 <= pi0067 and not w46;
w362 <= w32 and w40;
w363 <= not pi0084 and w362;
w364 <= not pi0068 and w363;
w365 <= w42 and w364;
w366 <= pi0036 and not w365;
w367 <= not pi0036 and not pi0067;
w368 <= not pi0068 and not pi0111;
w369 <= pi0082 and w368;
w370 <= w363 and w369;
w371 <= pi0111 and not w364;
w372 <= not pi0082 and not w371;
w373 <= pi0068 and not w363;
w374 <= pi0084 and not w362;
w375 <= pi0104 and not w38;
w376 <= pi0085 and pi0106;
w377 <= w33 and not w376;
w378 <= pi0061 and pi0076;
w379 <= w34 and not w378;
w380 <= not w377 and not w379;
w381 <= not pi0048 and not w380;
w382 <= not w35 and not w381;
w383 <= pi0089 and not w36;
w384 <= not pi0049 and not w383;
w385 <= not w382 and w384;
w386 <= not w37 and not w385;
w387 <= not pi0045 and not w375;
w388 <= not w386 and w387;
w389 <= not w39 and not w388;
w390 <= not w40 and not w389;
w391 <= w32 and not w390;
w392 <= pi0066 and pi0073;
w393 <= not w32 and not w40;
w394 <= not w392 and not w393;
w395 <= not w391 and w394;
w396 <= not pi0084 and not w395;
w397 <= not w374 and not w396;
w398 <= w368 and not w397;
w399 <= w372 and not w373;
w400 <= not w398 and w399;
w401 <= w367 and not w370;
w402 <= not w400 and w401;
w403 <= not w361 and not w366;
w404 <= not w402 and w403;
w405 <= w360 and not w404;
w406 <= w359 and not w405;
w407 <= pi0103 and w360;
w408 <= w355 and w407;
w409 <= not pi0071 and not w408;
w410 <= not w406 and w409;
w411 <= w354 and not w410;
w412 <= not pi0107 and not w411;
w413 <= pi0065 and not pi0071;
w414 <= w48 and w413;
w415 <= w412 and not w414;
w416 <= pi0107 and not w49;
w417 <= not pi0063 and not w416;
w418 <= not w415 and w417;
w419 <= not pi0064 and not w418;
w420 <= not w352 and not w419;
w421 <= not pi0081 and not pi0102;
w422 <= not w420 and w421;
w423 <= not w412 and w417;
w424 <= pi0063 and not pi0107;
w425 <= w49 and w424;
w426 <= not pi0064 and not w425;
w427 <= not w423 and w426;
w428 <= not w352 and not w427;
w429 <= w422 and not w428;
w430 <= w351 and not w429;
w431 <= w25 and not w430;
w432 <= pi0098 and not w330;
w433 <= not pi0098 and w330;
w434 <= pi0088 and not w433;
w435 <= not pi0077 and not w432;
w436 <= not w434 and w435;
w437 <= not w431 and w436;
w438 <= w348 and not w437;
w439 <= pi0050 and not w340;
w440 <= not pi0060 and not w439;
w441 <= not w438 and w440;
w442 <= w282 and not w441;
w443 <= not w285 and not w442;
w444 <= not pi0086 and not w443;
w445 <= w346 and not w444;
w446 <= w344 and not w445;
w447 <= not w339 and not w446;
w448 <= not pi0108 and not w447;
w449 <= w338 and not w448;
w450 <= pi0046 and w59;
w451 <= w335 and w450;
w452 <= not pi0109 and not w451;
w453 <= not w449 and w452;
w454 <= not w329 and not w453;
w455 <= w328 and not w454;
w456 <= w327 and not w455;
w457 <= w320 and not w456;
w458 <= pi0058 and not w65;
w459 <= pi0090 and not w266;
w460 <= not pi0093 and not w459;
w461 <= not w458 and w460;
w462 <= not w457 and w461;
w463 <= w316 and not w462;
w464 <= w314 and not w463;
w465 <= not pi0051 and not w464;
w466 <= w313 and not w465;
w467 <= not pi0072 and not w466;
w468 <= w309 and not w467;
w469 <= w307 and not w468;
w470 <= not w275 and not w469;
w471 <= not pi0095 and not w470;
w472 <= w305 and not w471;
w473 <= pi0137 and not w472;
w474 <= not w303 and not w473;
w475 <= pi0210 and not w474;
w476 <= not pi0051 and not pi0072;
w477 <= pi0841 and w66;
w478 <= not pi0093 and w477;
w479 <= w476 and w478;
w480 <= not pi0035 and not pi0040;
w481 <= pi0225 and w480;
w482 <= w268 and w481;
w483 <= w479 and w482;
w484 <= pi0032 and not w483;
w485 <= not pi0095 and not w484;
w486 <= not pi0833 and pi0957;
w487 <= pi1091 and not w486;
w488 <= pi0829 and pi0950;
w489 <= pi1092 and pi1093;
w490 <= w488 and w489;
w491 <= w487 and w490;
w492 <= not w290 and not w491;
w493 <= pi1091 and pi1093;
w494 <= not w486 and w493;
w495 <= pi0950 and pi1092;
w496 <= pi0829 and w495;
w497 <= not pi0046 and not pi0109;
w498 <= w55 and w497;
w499 <= not pi0108 and not w339;
w500 <= not pi0110 and w499;
w501 <= not pi0093 and w24;
w502 <= not pi0097 and not w287;
w503 <= w498 and w501;
w504 <= w500 and w503;
w505 <= not w502 and w504;
w506 <= not pi0035 and not w505;
w507 <= w494 and w496;
w508 <= not w506 and w507;
w509 <= not w492 and not w508;
w510 <= w297 and w299;
w511 <= not w509 and w510;
w512 <= not pi0032 and not w511;
w513 <= w485 and not w512;
w514 <= not pi0137 and not w513;
w515 <= not w469 and not w484;
w516 <= not pi0095 and not w515;
w517 <= w305 and not w516;
w518 <= pi0137 and not w517;
w519 <= not w514 and not w518;
w520 <= not pi0210 and not w519;
w521 <= not w475 and not w520;
w522 <= not pi0234 and w521;
w523 <= not pi0096 and not w298;
w524 <= not pi0035 and not pi0070;
w525 <= not pi0051 and w524;
w526 <= not pi0091 and w501;
w527 <= w525 and w526;
w528 <= w318 and w527;
w529 <= pi0096 and not w528;
w530 <= w80 and not w529;
w531 <= not w523 and w530;
w532 <= not pi0032 and not w531;
w533 <= w276 and not w532;
w534 <= not w5 and not w533;
w535 <= not pi0137 and w534;
w536 <= pi0096 and w528;
w537 <= not pi0040 and w476;
w538 <= w68 and w537;
w539 <= w536 and w538;
w540 <= w469 and not w539;
w541 <= not w275 and not w540;
w542 <= not pi0095 and not w541;
w543 <= pi0479 and w304;
w544 <= not w542 and not w543;
w545 <= pi0137 and not w544;
w546 <= not w535 and not w545;
w547 <= pi0210 and not w546;
w548 <= not w484 and not w540;
w549 <= not pi0095 and not w548;
w550 <= not w543 and not w549;
w551 <= pi0137 and not w550;
w552 <= pi0095 and pi0479;
w553 <= not w484 and not w532;
w554 <= not pi0095 and not w553;
w555 <= not w552 and not w554;
w556 <= not pi0137 and not w555;
w557 <= not w551 and not w556;
w558 <= not w487 and w557;
w559 <= w297 and not w506;
w560 <= not pi0096 and not w559;
w561 <= w530 and not w560;
w562 <= not pi0032 and not w561;
w563 <= not w484 and not w562;
w564 <= not pi0095 and not w563;
w565 <= w490 and not w552;
w566 <= not w564 and w565;
w567 <= not w490 and w555;
w568 <= not pi0137 and not w566;
w569 <= not w567 and w568;
w570 <= w487 and not w569;
w571 <= not w551 and w570;
w572 <= not w558 and not w571;
w573 <= not pi0210 and w572;
w574 <= not w547 and not w573;
w575 <= pi0234 and w574;
w576 <= not pi0332 and not w522;
w577 <= not w575 and w576;
w578 <= w202 and not w577;
w579 <= pi0146 and w574;
w580 <= not pi0210 and not w557;
w581 <= not pi0146 and not w547;
w582 <= not w580 and w581;
w583 <= w244 and not w582;
w584 <= not w579 and w583;
w585 <= pi0146 and w521;
w586 <= not w301 and w485;
w587 <= not pi0137 and not w586;
w588 <= not w518 and not w587;
w589 <= not pi0210 and not w588;
w590 <= not pi0146 and not w475;
w591 <= not w589 and w590;
w592 <= w239 and not w585;
w593 <= not w591 and w592;
w594 <= not w202 and not w593;
w595 <= not w584 and w594;
w596 <= not w578 and not w595;
w597 <= pi0105 and not w596;
w598 <= not w106 and not w597;
w599 <= pi0228 and not w598;
w600 <= not pi0109 and not w449;
w601 <= not w329 and not w600;
w602 <= w328 and not w601;
w603 <= w327 and not w602;
w604 <= w320 and not w603;
w605 <= w461 and not w604;
w606 <= w316 and not w605;
w607 <= w314 and not w606;
w608 <= not pi0051 and not w607;
w609 <= w313 and not w608;
w610 <= not pi0072 and not w609;
w611 <= w309 and not w610;
w612 <= w307 and not w611;
w613 <= not w484 and not w612;
w614 <= not pi0095 and not w613;
w615 <= w305 and not w614;
w616 <= pi0137 and not w615;
w617 <= w203 and w587;
w618 <= not w203 and w514;
w619 <= not pi0210 and not pi0234;
w620 <= not w617 and w619;
w621 <= not w618 and w620;
w622 <= not w616 and w621;
w623 <= not w275 and not w612;
w624 <= not pi0095 and not w623;
w625 <= w305 and not w624;
w626 <= pi0137 and not w625;
w627 <= pi0210 and not w303;
w628 <= not w626 and w627;
w629 <= not w539 and w612;
w630 <= not w484 and not w629;
w631 <= not pi0095 and not w630;
w632 <= not w304 and not w631;
w633 <= pi0137 and not w632;
w634 <= not w203 and w487;
w635 <= not w567 and w634;
w636 <= not w304 and w555;
w637 <= not w635 and w636;
w638 <= not w304 and w634;
w639 <= w566 and w638;
w640 <= not pi0137 and not w639;
w641 <= not w637 and w640;
w642 <= not w633 and not w641;
w643 <= not pi0210 and not w642;
w644 <= pi0234 and not w643;
w645 <= not w622 and not w628;
w646 <= not w644 and w645;
w647 <= not pi0137 and not w304;
w648 <= not w534 and w647;
w649 <= not w275 and not w629;
w650 <= not pi0095 and not w649;
w651 <= pi0137 and not w304;
w652 <= not w650 and w651;
w653 <= pi0210 and pi0234;
w654 <= not w648 and w653;
w655 <= not w652 and w654;
w656 <= not w646 and not w655;
w657 <= w9 and not w656;
w658 <= pi0225 and pi0841;
w659 <= w273 and not w658;
w660 <= pi0032 and not w659;
w661 <= not pi0095 and not w660;
w662 <= pi0070 and not w68;
w663 <= w79 and not w662;
w664 <= w80 and w663;
w665 <= not w295 and w664;
w666 <= not pi0032 and not w665;
w667 <= w661 and not w666;
w668 <= pi0137 and not w667;
w669 <= pi0093 and not w66;
w670 <= not pi0035 and not w669;
w671 <= not w458 and not w459;
w672 <= not pi0053 and w441;
w673 <= not pi0086 and not w672;
w674 <= w346 and not w673;
w675 <= w344 and not w674;
w676 <= not w339 and not w675;
w677 <= not pi0108 and not w676;
w678 <= w338 and not w677;
w679 <= not pi0109 and not w678;
w680 <= not w329 and not w679;
w681 <= w328 and not w680;
w682 <= w327 and not w681;
w683 <= w320 and not w682;
w684 <= w671 and not w683;
w685 <= not pi0093 and not w684;
w686 <= w670 and not w685;
w687 <= w296 and not w686;
w688 <= w311 and not w662;
w689 <= not w687 and w688;
w690 <= not pi0072 and not w689;
w691 <= w309 and not w690;
w692 <= w307 and not w691;
w693 <= not w491 and w692;
w694 <= w307 and w491;
w695 <= not pi0097 and not w675;
w696 <= not pi0108 and not w695;
w697 <= w338 and not w696;
w698 <= not pi0109 and not w697;
w699 <= not w329 and not w698;
w700 <= w328 and not w699;
w701 <= w327 and not w700;
w702 <= w320 and not w701;
w703 <= w671 and not w702;
w704 <= not pi0093 and not w703;
w705 <= w670 and not w704;
w706 <= w296 and not w705;
w707 <= w688 and not w706;
w708 <= not pi0072 and not w707;
w709 <= w309 and not w708;
w710 <= w694 and not w709;
w711 <= not w660 and not w710;
w712 <= not w693 and w711;
w713 <= not pi0095 and not w712;
w714 <= w305 and not w713;
w715 <= not pi0137 and not w714;
w716 <= not w668 and not w715;
w717 <= not pi0210 and not w716;
w718 <= not pi0225 and w273;
w719 <= pi0032 and not w718;
w720 <= not pi0095 and not w719;
w721 <= pi0137 and w720;
w722 <= not w666 and w721;
w723 <= not w692 and not w719;
w724 <= not pi0095 and not w723;
w725 <= not pi0137 and w305;
w726 <= not w724 and w725;
w727 <= pi0210 and not w722;
w728 <= not w726 and w727;
w729 <= w244 and not w728;
w730 <= not w717 and w729;
w731 <= not pi0072 and not w536;
w732 <= not w689 and w731;
w733 <= w309 and not w732;
w734 <= w307 and not w733;
w735 <= not w491 and w734;
w736 <= not w707 and w731;
w737 <= w309 and not w736;
w738 <= w694 and not w737;
w739 <= not w660 and not w738;
w740 <= not w735 and w739;
w741 <= not pi0095 and not w740;
w742 <= not w304 and not w741;
w743 <= not pi0137 and not w742;
w744 <= w5 and w74;
w745 <= not pi0072 and w73;
w746 <= w536 and w745;
w747 <= w666 and not w746;
w748 <= w661 and not w747;
w749 <= pi0137 and not w744;
w750 <= not w748 and w749;
w751 <= not w743 and not w750;
w752 <= not pi0210 and not w751;
w753 <= not w719 and not w734;
w754 <= not pi0095 and not w753;
w755 <= w647 and not w754;
w756 <= w720 and not w747;
w757 <= not w744 and not w756;
w758 <= pi0137 and not w757;
w759 <= pi0210 and not w758;
w760 <= not w755 and w759;
w761 <= w239 and not w760;
w762 <= not w752 and w761;
w763 <= w202 and not w730;
w764 <= not w762 and w763;
w765 <= pi0146 and w752;
w766 <= not pi0146 and not pi0210;
w767 <= not w660 and not w734;
w768 <= not pi0095 and not w767;
w769 <= not w304 and not w768;
w770 <= not pi0137 and not w769;
w771 <= not w750 and not w770;
w772 <= w766 and not w771;
w773 <= w761 and not w772;
w774 <= not w765 and w773;
w775 <= not w660 and not w692;
w776 <= not pi0095 and not w775;
w777 <= w305 and not w776;
w778 <= not pi0137 and not w777;
w779 <= not w668 and not w778;
w780 <= w766 and not w779;
w781 <= pi0146 and w717;
w782 <= w729 and not w780;
w783 <= not w781 and w782;
w784 <= not w202 and not w774;
w785 <= not w783 and w784;
w786 <= not pi0153 and not w764;
w787 <= not w785 and w786;
w788 <= not pi0228 and not w657;
w789 <= not w787 and w788;
w790 <= not w599 and not w789;
w791 <= not pi0216 and not w790;
w792 <= not w3 and not w791;
w793 <= not pi0221 and not w792;
w794 <= not w20 and not w793;
w795 <= not pi0215 and not w794;
w796 <= pi0299 and not w1;
w797 <= not w795 and w796;
w798 <= pi0198 and not w546;
w799 <= not pi0198 and w572;
w800 <= not w798 and not w799;
w801 <= pi0142 and w800;
w802 <= not pi0198 and not w557;
w803 <= not pi0142 and not w798;
w804 <= not w802 and w803;
w805 <= w244 and not w804;
w806 <= not w801 and w805;
w807 <= pi0198 and not w474;
w808 <= not pi0198 and not w519;
w809 <= not w807 and not w808;
w810 <= pi0142 and w809;
w811 <= not pi0198 and not w588;
w812 <= not pi0142 and not w807;
w813 <= not w811 and w812;
w814 <= w239 and not w810;
w815 <= not w813 and w814;
w816 <= w233 and not w815;
w817 <= not w806 and w816;
w818 <= not pi0234 and w809;
w819 <= pi0234 and w800;
w820 <= not pi0332 and not w818;
w821 <= not w819 and w820;
w822 <= w243 and not w821;
w823 <= not w817 and not w822;
w824 <= w166 and not w823;
w825 <= w165 and not w824;
w826 <= not pi0039 and not w825;
w827 <= not w797 and w826;
w828 <= not pi0038 and not w261;
w829 <= not w827 and w828;
w830 <= not pi0100 and not w260;
w831 <= not w829 and w830;
w832 <= not pi0087 and not w257;
w833 <= not w831 and w832;
w834 <= not pi0075 and not w198;
w835 <= not w833 and w834;
w836 <= not w170 and not w173;
w837 <= w11 and not w210;
w838 <= not w3 and not w837;
w839 <= not pi0221 and not w838;
w840 <= not w20 and not w839;
w841 <= not pi0215 and not w840;
w842 <= not w1 and not w841;
w843 <= pi0299 and not w842;
w844 <= w173 and not w253;
w845 <= not w843 and w844;
w846 <= pi0075 and not w836;
w847 <= not w845 and w846;
w848 <= not w835 and not w847;
w849 <= not pi0092 and not w848;
w850 <= not pi0054 and not w197;
w851 <= not w849 and w850;
w852 <= not pi0074 and not w187;
w853 <= not w851 and w852;
w854 <= pi0054 and not w170;
w855 <= not pi0054 and w186;
w856 <= pi0074 and not w854;
w857 <= not w855 and w856;
w858 <= not w853 and not w857;
w859 <= not pi0055 and not w858;
w860 <= not pi0056 and not w152;
w861 <= not w859 and w860;
w862 <= not pi0062 and not w130;
w863 <= not w861 and w862;
w864 <= not pi0059 and not w129;
w865 <= not w863 and w864;
w866 <= not pi0057 and not w104;
w867 <= not w865 and w866;
w868 <= not pi0059 and w102;
w869 <= w23 and not w868;
w870 <= pi0057 and not w869;
w871 <= not w867 and not w870;
w872 <= pi0215 and pi1146;
w873 <= pi0216 and not pi0221;
w874 <= pi0276 and w873;
w875 <= not pi1146 and not w15;
w876 <= not pi0939 and w15;
w877 <= pi0221 and not w875;
w878 <= not w876 and w877;
w879 <= not w874 and not w878;
w880 <= not pi0215 and not w879;
w881 <= not w872 and not w880;
w882 <= pi0154 and not w881;
w883 <= not pi0216 and not w4;
w884 <= not w874 and not w883;
w885 <= not pi0221 and not w884;
w886 <= not w878 and not w885;
w887 <= not pi0215 and not w886;
w888 <= not w872 and not w887;
w889 <= not pi0154 and not w888;
w890 <= not w882 and not w889;
w891 <= not pi0057 and not pi0059;
w892 <= w890 and not w891;
w893 <= not pi0056 and w99;
w894 <= w94 and w893;
w895 <= not w890 and not w894;
w896 <= not pi0055 and w135;
w897 <= not w872 and not w878;
w898 <= not pi0228 and w84;
w899 <= not pi0216 and w898;
w900 <= w897 and w899;
w901 <= not w882 and w900;
w902 <= not w890 and w896;
w903 <= not w901 and w902;
w904 <= not w895 and not w903;
w905 <= pi0062 and not w904;
w906 <= not w100 and not w890;
w907 <= pi0056 and not w906;
w908 <= not w903 and w907;
w909 <= w135 and w901;
w910 <= pi0055 and not w890;
w911 <= not w909 and w910;
w912 <= pi0299 and not w890;
w913 <= pi0223 and not pi1146;
w914 <= not pi0222 and pi0224;
w915 <= pi0276 and w914;
w916 <= not pi1146 and not w154;
w917 <= not pi0939 and w154;
w918 <= pi0222 and not w916;
w919 <= not w917 and w918;
w920 <= not pi0223 and not w915;
w921 <= not w919 and w920;
w922 <= not pi0299 and not w913;
w923 <= not w921 and w922;
w924 <= not w912 and not w923;
w925 <= not w95 and w924;
w926 <= pi0299 and not w881;
w927 <= not w923 and not w926;
w928 <= pi0154 and not w927;
w929 <= pi0299 and not w888;
w930 <= not w900 and w929;
w931 <= not w923 and not w930;
w932 <= not pi0154 and not w931;
w933 <= w188 and not w928;
w934 <= not w932 and w933;
w935 <= w96 and w934;
w936 <= w94 and w96;
w937 <= w924 and not w936;
w938 <= pi0092 and not w937;
w939 <= not w935 and w938;
w940 <= pi0075 and w924;
w941 <= not w188 and w924;
w942 <= not w934 and not w941;
w943 <= pi0087 and not w942;
w944 <= not pi0038 and not pi0216;
w945 <= not pi0228 and w944;
w946 <= not pi0154 and pi0299;
w947 <= not pi0146 and not w84;
w948 <= not pi0252 and w84;
w949 <= pi0146 and not w948;
w950 <= not w947 and not w949;
w951 <= pi0152 and not w950;
w952 <= not pi0161 and not pi0166;
w953 <= w948 and w952;
w954 <= w950 and not w952;
w955 <= not pi0152 and not w953;
w956 <= not w954 and w955;
w957 <= not w951 and not w956;
w958 <= not pi0039 and w946;
w959 <= w945 and w958;
w960 <= w897 and w959;
w961 <= w957 and w960;
w962 <= pi0100 and not w924;
w963 <= not w961 and w962;
w964 <= pi0038 and w924;
w965 <= pi0039 and not w84;
w966 <= not pi0070 and w606;
w967 <= not w292 and not w662;
w968 <= not w966 and w967;
w969 <= not pi0051 and not w968;
w970 <= w311 and not w969;
w971 <= w731 and not w970;
w972 <= not w308 and not w971;
w973 <= w73 and not w972;
w974 <= pi0040 and not w72;
w975 <= pi0032 and not w273;
w976 <= not w974 and not w975;
w977 <= not w973 and w976;
w978 <= not pi0095 and not w977;
w979 <= not w304 and not w978;
w980 <= not pi0039 and not w979;
w981 <= not w965 and not w980;
w982 <= not pi0216 and not pi0228;
w983 <= w897 and w982;
w984 <= w981 and w983;
w985 <= w929 and not w984;
w986 <= not w923 and not w985;
w987 <= not pi0154 and not w986;
w988 <= not pi0038 and not w928;
w989 <= not w987 and w988;
w990 <= not pi0100 and not w964;
w991 <= not w989 and w990;
w992 <= not pi0087 and not w963;
w993 <= not w991 and w992;
w994 <= not w943 and not w993;
w995 <= not pi0075 and not w994;
w996 <= not pi0092 and not w940;
w997 <= not w995 and w996;
w998 <= w95 and not w939;
w999 <= not w997 and w998;
w1000 <= not pi0055 and not w925;
w1001 <= not w999 and w1000;
w1002 <= not pi0056 and not w911;
w1003 <= not w1001 and w1002;
w1004 <= not pi0062 and not w908;
w1005 <= not w1003 and w1004;
w1006 <= w891 and not w905;
w1007 <= not w1005 and w1006;
w1008 <= not pi0239 and not w892;
w1009 <= not w1007 and w1008;
w1010 <= w4 and w5;
w1011 <= not pi0216 and not pi0221;
w1012 <= not pi0215 and w1011;
w1013 <= w1010 and w1012;
w1014 <= w881 and not w1013;
w1015 <= not pi0215 and not w1014;
w1016 <= pi0154 and not w1014;
w1017 <= not w889 and not w1015;
w1018 <= not w1016 and w1017;
w1019 <= not w891 and w1018;
w1020 <= not w894 and not w1018;
w1021 <= w900 and not w1016;
w1022 <= not w1018 and not w1021;
w1023 <= w896 and w1022;
w1024 <= not pi0056 and w1023;
w1025 <= not w1020 and not w1024;
w1026 <= pi0062 and not w1025;
w1027 <= not w100 and not w1018;
w1028 <= pi0056 and not w1027;
w1029 <= not w1023 and w1028;
w1030 <= w135 and w1021;
w1031 <= pi0055 and not w1018;
w1032 <= not w1030 and w1031;
w1033 <= not pi0223 and not pi0299;
w1034 <= w166 and w1033;
w1035 <= w5 and w1034;
w1036 <= pi0299 and not w1018;
w1037 <= not w923 and not w1035;
w1038 <= not w1036 and w1037;
w1039 <= not w95 and w1038;
w1040 <= pi0299 and not w1022;
w1041 <= w936 and w1040;
w1042 <= pi0092 and not w1038;
w1043 <= not w1041 and w1042;
w1044 <= pi0075 and w1038;
w1045 <= w188 and w1040;
w1046 <= pi0087 and not w1038;
w1047 <= not w1045 and w1046;
w1048 <= not w1038 and not w1040;
w1049 <= pi0039 and not w1048;
w1050 <= w82 and w536;
w1051 <= not w5 and not w1050;
w1052 <= not pi0224 and w1051;
w1053 <= pi0224 and not pi0276;
w1054 <= not pi0222 and not w1053;
w1055 <= not w1052 and w1054;
w1056 <= not pi0223 and not w919;
w1057 <= not w1055 and w1056;
w1058 <= not w913 and not w1057;
w1059 <= not pi0299 and not w1058;
w1060 <= pi0105 and not w1051;
w1061 <= pi0228 and not w1060;
w1062 <= not w304 and not w1051;
w1063 <= not pi0228 and not w1062;
w1064 <= not w1061 and not w1063;
w1065 <= pi0154 and not w1064;
w1066 <= not pi0072 and not w970;
w1067 <= not w308 and not w1066;
w1068 <= w73 and not w1067;
w1069 <= w976 and not w1068;
w1070 <= not pi0095 and not w1069;
w1071 <= w305 and not w1070;
w1072 <= not pi0228 and w1071;
w1073 <= w4 and w1051;
w1074 <= not w1072 and not w1073;
w1075 <= not pi0154 and not w1074;
w1076 <= w1012 and not w1065;
w1077 <= not w1075 and w1076;
w1078 <= pi0299 and w881;
w1079 <= not w1077 and w1078;
w1080 <= not w1059 and not w1079;
w1081 <= not pi0039 and not w1080;
w1082 <= w171 and not w1049;
w1083 <= not w1081 and w1082;
w1084 <= pi0100 and w961;
w1085 <= not w171 and not w1038;
w1086 <= not w1084 and w1085;
w1087 <= not w1083 and not w1086;
w1088 <= not pi0087 and not w1087;
w1089 <= not pi0075 and not w1047;
w1090 <= not w1088 and w1089;
w1091 <= not pi0092 and not w1044;
w1092 <= not w1090 and w1091;
w1093 <= w95 and not w1043;
w1094 <= not w1092 and w1093;
w1095 <= not pi0055 and not w1039;
w1096 <= not w1094 and w1095;
w1097 <= not pi0056 and not w1032;
w1098 <= not w1096 and w1097;
w1099 <= not pi0062 and not w1029;
w1100 <= not w1098 and w1099;
w1101 <= w891 and not w1026;
w1102 <= not w1100 and w1101;
w1103 <= pi0239 and not w1019;
w1104 <= not w1102 and w1103;
w1105 <= not w1009 and not w1104;
w1106 <= pi0215 and pi1145;
w1107 <= pi0216 and pi0274;
w1108 <= not pi0221 and not w1107;
w1109 <= not pi0151 and not w4;
w1110 <= not pi0216 and not w1109;
w1111 <= w1108 and not w1110;
w1112 <= not pi1145 and not w15;
w1113 <= not pi0927 and w15;
w1114 <= pi0221 and not w1112;
w1115 <= not w1113 and w1114;
w1116 <= not w1111 and not w1115;
w1117 <= not pi0215 and not w1116;
w1118 <= not w1106 and not w1117;
w1119 <= w89 and w1010;
w1120 <= not w1107 and w1119;
w1121 <= w1118 and not w1120;
w1122 <= not w894 and w1121;
w1123 <= not w1010 and not w1109;
w1124 <= not pi0151 and w898;
w1125 <= not w1123 and not w1124;
w1126 <= not pi0216 and not w1125;
w1127 <= w1108 and not w1126;
w1128 <= not w1115 and not w1127;
w1129 <= not pi0215 and not w1128;
w1130 <= not w1106 and not w1129;
w1131 <= w894 and w1130;
w1132 <= pi0062 and not w1122;
w1133 <= not w1131 and w1132;
w1134 <= not w100 and not w1121;
w1135 <= w100 and not w1130;
w1136 <= pi0056 and not w1134;
w1137 <= not w1135 and w1136;
w1138 <= not w135 and w1121;
w1139 <= w135 and w1130;
w1140 <= pi0055 and not w1138;
w1141 <= not w1139 and w1140;
w1142 <= pi0223 and pi1145;
w1143 <= not pi1145 and not w154;
w1144 <= not pi0927 and w154;
w1145 <= pi0222 and not w1143;
w1146 <= not w1144 and w1145;
w1147 <= pi0224 and pi0274;
w1148 <= w914 and not w1147;
w1149 <= not w1146 and not w1148;
w1150 <= not pi0223 and not w1149;
w1151 <= not w1142 and not w1150;
w1152 <= not pi0299 and not w1151;
w1153 <= not w1035 and not w1152;
w1154 <= pi0299 and not w1121;
w1155 <= w1153 and not w1154;
w1156 <= not w95 and w1155;
w1157 <= not w188 and w1155;
w1158 <= pi0299 and not w1130;
w1159 <= w1153 and not w1158;
w1160 <= w188 and w1159;
w1161 <= not w1157 and not w1160;
w1162 <= w96 and not w1161;
w1163 <= not w96 and w1155;
w1164 <= pi0092 and not w1163;
w1165 <= not w1162 and w1164;
w1166 <= pi0075 and w1155;
w1167 <= pi0087 and w1161;
w1168 <= pi0038 and w1155;
w1169 <= pi0039 and not w1159;
w1170 <= not pi0222 and not w1147;
w1171 <= not w1052 and w1170;
w1172 <= not w1146 and not w1171;
w1173 <= not pi0223 and not w1172;
w1174 <= not pi0299 and not w1142;
w1175 <= not w1173 and w1174;
w1176 <= not pi0151 and w1074;
w1177 <= pi0151 and w1064;
w1178 <= not pi0216 and not w1177;
w1179 <= not w1176 and w1178;
w1180 <= w1108 and not w1179;
w1181 <= not w1115 and not w1180;
w1182 <= not pi0215 and not w1181;
w1183 <= pi0299 and not w1106;
w1184 <= not w1182 and w1183;
w1185 <= not pi0039 and not w1175;
w1186 <= not w1184 and w1185;
w1187 <= not pi0038 and not w1169;
w1188 <= not w1186 and w1187;
w1189 <= not pi0100 and not w1168;
w1190 <= not w1188 and w1189;
w1191 <= not w93 and w1155;
w1192 <= not pi0228 and w957;
w1193 <= w4 and not w5;
w1194 <= not w1192 and not w1193;
w1195 <= not pi0151 and w1194;
w1196 <= w1126 and not w1195;
w1197 <= w1108 and not w1196;
w1198 <= not w1115 and not w1197;
w1199 <= not pi0215 and not w1198;
w1200 <= not w1106 and not w1199;
w1201 <= pi0299 and not w1200;
w1202 <= w93 and w1153;
w1203 <= not w1201 and w1202;
w1204 <= pi0100 and not w1191;
w1205 <= not w1203 and w1204;
w1206 <= not w1190 and not w1205;
w1207 <= not pi0087 and not w1206;
w1208 <= not pi0075 and not w1167;
w1209 <= not w1207 and w1208;
w1210 <= not pi0092 and not w1166;
w1211 <= not w1209 and w1210;
w1212 <= w95 and not w1165;
w1213 <= not w1211 and w1212;
w1214 <= not pi0055 and not w1156;
w1215 <= not w1213 and w1214;
w1216 <= not pi0056 and not w1141;
w1217 <= not w1215 and w1216;
w1218 <= not pi0062 and not w1137;
w1219 <= not w1217 and w1218;
w1220 <= pi0235 and w891;
w1221 <= not w1133 and w1220;
w1222 <= not w1219 and w1221;
w1223 <= not w1106 and not w1115;
w1224 <= w899 and w1223;
w1225 <= w100 and w1224;
w1226 <= not pi0056 and w1225;
w1227 <= pi0062 and not w1118;
w1228 <= not w1226 and w1227;
w1229 <= not w1118 and not w1225;
w1230 <= pi0056 and not w1229;
w1231 <= w135 and w1224;
w1232 <= pi0055 and not w1118;
w1233 <= not w1231 and w1232;
w1234 <= pi0299 and not w1118;
w1235 <= not w1152 and not w1234;
w1236 <= not w95 and w1235;
w1237 <= not w1224 and w1234;
w1238 <= w94 and not w1152;
w1239 <= not w1237 and w1238;
w1240 <= w96 and w1239;
w1241 <= not w936 and w1235;
w1242 <= pi0092 and not w1241;
w1243 <= not w1240 and w1242;
w1244 <= pi0075 and w1235;
w1245 <= not w188 and w1235;
w1246 <= not w1239 and not w1245;
w1247 <= pi0087 and not w1246;
w1248 <= not pi0100 and w981;
w1249 <= not pi0039 and pi0100;
w1250 <= w957 and w1249;
w1251 <= not w1248 and not w1250;
w1252 <= w945 and w1223;
w1253 <= not w1251 and w1252;
w1254 <= w1234 and not w1253;
w1255 <= not pi0087 and not w1152;
w1256 <= not w1254 and w1255;
w1257 <= not w1247 and not w1256;
w1258 <= not pi0075 and not w1257;
w1259 <= not pi0092 and not w1244;
w1260 <= not w1258 and w1259;
w1261 <= w95 and not w1243;
w1262 <= not w1260 and w1261;
w1263 <= not pi0055 and not w1236;
w1264 <= not w1262 and w1263;
w1265 <= not pi0056 and not w1233;
w1266 <= not w1264 and w1265;
w1267 <= not pi0062 and not w1230;
w1268 <= not w1266 and w1267;
w1269 <= not pi0235 and w891;
w1270 <= not w1228 and w1269;
w1271 <= not w1268 and w1270;
w1272 <= pi0235 and w1120;
w1273 <= not w891 and not w1272;
w1274 <= w1118 and w1273;
w1275 <= not w1271 and not w1274;
w1276 <= not w1222 and w1275;
w1277 <= pi0215 and pi1143;
w1278 <= pi0216 and pi0264;
w1279 <= not pi0221 and not w1278;
w1280 <= not pi0105 and pi0146;
w1281 <= pi0284 and not w5;
w1282 <= pi0105 and not w1281;
w1283 <= pi0228 and not w1280;
w1284 <= not w1282 and w1283;
w1285 <= not w1010 and not w1284;
w1286 <= not pi0146 and not pi0228;
w1287 <= w1285 and not w1286;
w1288 <= not pi0216 and not w1287;
w1289 <= w1279 and not w1288;
w1290 <= not pi1143 and not w15;
w1291 <= not pi0944 and w15;
w1292 <= pi0221 and not w1290;
w1293 <= not w1291 and w1292;
w1294 <= not w1289 and not w1293;
w1295 <= not pi0215 and not w1294;
w1296 <= not w1277 and not w1295;
w1297 <= not w894 and w1296;
w1298 <= pi0284 and w84;
w1299 <= not w947 and not w1298;
w1300 <= not pi0228 and not w1299;
w1301 <= w1285 and not w1300;
w1302 <= not pi0216 and not w1301;
w1303 <= w1279 and not w1302;
w1304 <= not w1293 and not w1303;
w1305 <= not pi0215 and not w1304;
w1306 <= not w1277 and not w1305;
w1307 <= w894 and w1306;
w1308 <= pi0062 and not w1297;
w1309 <= not w1307 and w1308;
w1310 <= not w100 and not w1296;
w1311 <= w100 and not w1306;
w1312 <= pi0056 and not w1310;
w1313 <= not w1311 and w1312;
w1314 <= not w135 and w1296;
w1315 <= w135 and w1306;
w1316 <= pi0055 and not w1314;
w1317 <= not w1315 and w1316;
w1318 <= w5 and w167;
w1319 <= pi0223 and pi1143;
w1320 <= pi0224 and pi0264;
w1321 <= not pi0222 and not w1320;
w1322 <= not pi0224 and w1281;
w1323 <= w1321 and not w1322;
w1324 <= not pi1143 and not w154;
w1325 <= not pi0944 and w154;
w1326 <= pi0222 and not w1324;
w1327 <= not w1325 and w1326;
w1328 <= not w1323 and not w1327;
w1329 <= not pi0223 and not w1328;
w1330 <= not w1319 and not w1329;
w1331 <= not pi0299 and not w1330;
w1332 <= not w1318 and w1331;
w1333 <= pi0299 and not w1296;
w1334 <= not w1332 and not w1333;
w1335 <= not w95 and w1334;
w1336 <= not w188 and w1334;
w1337 <= pi0299 and not w1306;
w1338 <= not w1332 and not w1337;
w1339 <= w188 and w1338;
w1340 <= not w1336 and not w1339;
w1341 <= w96 and not w1340;
w1342 <= not w96 and w1334;
w1343 <= pi0092 and not w1342;
w1344 <= not w1341 and w1343;
w1345 <= pi0075 and w1334;
w1346 <= pi0087 and w1340;
w1347 <= pi0038 and w1334;
w1348 <= pi0039 and not w1338;
w1349 <= not pi0299 and not w1319;
w1350 <= not pi0284 and w1051;
w1351 <= not pi0224 and not w1350;
w1352 <= w1321 and not w1351;
w1353 <= not w1327 and not w1352;
w1354 <= w1349 and w1353;
w1355 <= pi0299 and not w1277;
w1356 <= w4 and not w1051;
w1357 <= not pi0146 and not w1071;
w1358 <= pi0146 and w1062;
w1359 <= not pi0284 and not w1358;
w1360 <= pi0146 and pi0284;
w1361 <= not w979 and w1360;
w1362 <= not w1359 and not w1361;
w1363 <= not w1357 and not w1362;
w1364 <= not pi0228 and not w1363;
w1365 <= not w1284 and not w1356;
w1366 <= not w1364 and w1365;
w1367 <= not pi0216 and not w1366;
w1368 <= w1279 and not w1367;
w1369 <= not w1293 and not w1368;
w1370 <= not pi0215 and not w1369;
w1371 <= w1355 and not w1370;
w1372 <= not w1051 and w1321;
w1373 <= w1353 and not w1372;
w1374 <= not pi0223 and not w1373;
w1375 <= w1349 and not w1374;
w1376 <= not pi0039 and not w1375;
w1377 <= not w1354 and w1376;
w1378 <= not w1371 and w1377;
w1379 <= not pi0038 and not w1348;
w1380 <= not w1378 and w1379;
w1381 <= not pi0100 and not w1347;
w1382 <= not w1380 and w1381;
w1383 <= not w93 and w1334;
w1384 <= pi0252 and w202;
w1385 <= not pi0284 and not w1384;
w1386 <= w84 and w1385;
w1387 <= not pi0228 and not w1386;
w1388 <= not w949 and w1387;
w1389 <= w1285 and not w1388;
w1390 <= not pi0216 and not w1389;
w1391 <= w1279 and not w1390;
w1392 <= not w1293 and not w1391;
w1393 <= not pi0215 and not w1392;
w1394 <= not w1277 and not w1393;
w1395 <= pi0299 and not w1394;
w1396 <= w93 and not w1332;
w1397 <= not w1395 and w1396;
w1398 <= pi0100 and not w1383;
w1399 <= not w1397 and w1398;
w1400 <= not w1382 and not w1399;
w1401 <= not pi0087 and not w1400;
w1402 <= not pi0075 and not w1346;
w1403 <= not w1401 and w1402;
w1404 <= not pi0092 and not w1345;
w1405 <= not w1403 and w1404;
w1406 <= w95 and not w1344;
w1407 <= not w1405 and w1406;
w1408 <= not pi0055 and not w1335;
w1409 <= not w1407 and w1408;
w1410 <= not pi0056 and not w1317;
w1411 <= not w1409 and w1410;
w1412 <= not pi0062 and not w1313;
w1413 <= not w1411 and w1412;
w1414 <= not pi0238 and w891;
w1415 <= not w1309 and w1414;
w1416 <= not w1413 and w1415;
w1417 <= not w1284 and not w1300;
w1418 <= not pi0216 and not w1417;
w1419 <= w1279 and not w1418;
w1420 <= not w1293 and not w1419;
w1421 <= not pi0215 and not w1420;
w1422 <= not w1277 and not w1421;
w1423 <= w894 and w1422;
w1424 <= w1119 and not w1278;
w1425 <= w1296 and not w1424;
w1426 <= not w894 and w1425;
w1427 <= pi0062 and not w1426;
w1428 <= not w1423 and w1427;
w1429 <= not w100 and not w1425;
w1430 <= w100 and not w1422;
w1431 <= pi0056 and not w1429;
w1432 <= not w1430 and w1431;
w1433 <= w135 and w1422;
w1434 <= not w135 and w1425;
w1435 <= pi0055 and not w1434;
w1436 <= not w1433 and w1435;
w1437 <= pi0299 and not w1425;
w1438 <= not w1331 and not w1437;
w1439 <= not w95 and w1438;
w1440 <= not w188 and w1438;
w1441 <= pi0299 and not w1422;
w1442 <= not w1331 and not w1441;
w1443 <= w188 and w1442;
w1444 <= not w1440 and not w1443;
w1445 <= w96 and not w1444;
w1446 <= not w96 and w1438;
w1447 <= pi0092 and not w1446;
w1448 <= not w1445 and w1447;
w1449 <= pi0075 and w1438;
w1450 <= pi0087 and w1444;
w1451 <= pi0038 and w1438;
w1452 <= pi0039 and not w1442;
w1453 <= not w1060 and w1284;
w1454 <= not pi0146 and w1062;
w1455 <= pi0146 and not w1071;
w1456 <= pi0284 and not w1454;
w1457 <= not w1455 and w1456;
w1458 <= not pi0146 and not pi0284;
w1459 <= not w979 and w1458;
w1460 <= not w1457 and not w1459;
w1461 <= not pi0228 and not w1460;
w1462 <= not w1453 and not w1461;
w1463 <= not pi0216 and not w1462;
w1464 <= w1279 and not w1463;
w1465 <= not w1293 and not w1464;
w1466 <= not pi0215 and not w1465;
w1467 <= w1355 and not w1466;
w1468 <= w1376 and not w1467;
w1469 <= not pi0038 and not w1452;
w1470 <= not w1468 and w1469;
w1471 <= not pi0100 and not w1451;
w1472 <= not w1470 and w1471;
w1473 <= not w93 and w1438;
w1474 <= not w1284 and not w1388;
w1475 <= not pi0216 and not w1474;
w1476 <= w1279 and not w1475;
w1477 <= not w1293 and not w1476;
w1478 <= not pi0215 and not w1477;
w1479 <= not w1277 and not w1478;
w1480 <= pi0299 and not w1479;
w1481 <= w93 and not w1331;
w1482 <= not w1480 and w1481;
w1483 <= pi0100 and not w1473;
w1484 <= not w1482 and w1483;
w1485 <= not w1472 and not w1484;
w1486 <= not pi0087 and not w1485;
w1487 <= not pi0075 and not w1450;
w1488 <= not w1486 and w1487;
w1489 <= not pi0092 and not w1449;
w1490 <= not w1488 and w1489;
w1491 <= w95 and not w1448;
w1492 <= not w1490 and w1491;
w1493 <= not pi0055 and not w1439;
w1494 <= not w1492 and w1493;
w1495 <= not pi0056 and not w1436;
w1496 <= not w1494 and w1495;
w1497 <= not pi0062 and not w1432;
w1498 <= not w1496 and w1497;
w1499 <= pi0238 and w891;
w1500 <= not w1428 and w1499;
w1501 <= not w1498 and w1500;
w1502 <= pi0238 and w1424;
w1503 <= not w891 and not w1502;
w1504 <= w1296 and w1503;
w1505 <= not w1416 and not w1504;
w1506 <= not w1501 and w1505;
w1507 <= pi0215 and pi1142;
w1508 <= pi0216 and pi0277;
w1509 <= not pi0221 and not w1508;
w1510 <= pi0172 and not pi0228;
w1511 <= not pi0105 and pi0172;
w1512 <= pi0262 and not w5;
w1513 <= pi0105 and w1512;
w1514 <= not w1511 and not w1513;
w1515 <= pi0228 and not w1514;
w1516 <= not w1510 and not w1515;
w1517 <= not pi0216 and not w1516;
w1518 <= w1509 and not w1517;
w1519 <= not pi1142 and not w15;
w1520 <= not pi0932 and w15;
w1521 <= pi0221 and not w1519;
w1522 <= not w1520 and w1521;
w1523 <= not w1518 and not w1522;
w1524 <= not pi0215 and not w1523;
w1525 <= not w1507 and not w1524;
w1526 <= not w1013 and not w1525;
w1527 <= not w891 and not w1526;
w1528 <= not w894 and not w1526;
w1529 <= not pi0262 and w84;
w1530 <= not w898 and not w1510;
w1531 <= not w1529 and not w1530;
w1532 <= not w1010 and not w1515;
w1533 <= not w1531 and w1532;
w1534 <= not pi0216 and not w1533;
w1535 <= w1509 and not w1534;
w1536 <= not w1522 and not w1535;
w1537 <= not pi0215 and not w1536;
w1538 <= not w1507 and not w1537;
w1539 <= w894 and w1538;
w1540 <= pi0062 and not w1528;
w1541 <= not w1539 and w1540;
w1542 <= w100 and not w1538;
w1543 <= not w100 and w1526;
w1544 <= pi0056 and not w1543;
w1545 <= not w1542 and w1544;
w1546 <= not w135 and not w1526;
w1547 <= w135 and w1538;
w1548 <= pi0055 and not w1546;
w1549 <= not w1547 and w1548;
w1550 <= pi0223 and pi1142;
w1551 <= pi0224 and pi0277;
w1552 <= not pi0222 and not w1551;
w1553 <= not pi0224 and w1512;
w1554 <= w1552 and not w1553;
w1555 <= not pi1142 and not w154;
w1556 <= not pi0932 and w154;
w1557 <= pi0222 and not w1555;
w1558 <= not w1556 and w1557;
w1559 <= not w1554 and not w1558;
w1560 <= not pi0223 and not w1559;
w1561 <= not w1550 and not w1560;
w1562 <= not pi0299 and not w1561;
w1563 <= not w1318 and w1562;
w1564 <= pi0299 and w1526;
w1565 <= not w1563 and not w1564;
w1566 <= not w95 and w1565;
w1567 <= not w188 and w1565;
w1568 <= pi0299 and not w1538;
w1569 <= not w1563 and not w1568;
w1570 <= w188 and w1569;
w1571 <= not w1567 and not w1570;
w1572 <= w96 and not w1571;
w1573 <= not w96 and w1565;
w1574 <= pi0092 and not w1573;
w1575 <= not w1572 and w1574;
w1576 <= pi0075 and w1565;
w1577 <= pi0087 and w1571;
w1578 <= pi0038 and w1565;
w1579 <= pi0039 and not w1569;
w1580 <= not pi0299 and not w1550;
w1581 <= not pi0262 and w1051;
w1582 <= not pi0224 and not w1581;
w1583 <= w1552 and not w1582;
w1584 <= not w1558 and not w1583;
w1585 <= w1580 and w1584;
w1586 <= pi0299 and not w1507;
w1587 <= pi0262 and w979;
w1588 <= not pi0262 and w1062;
w1589 <= not pi0172 and not w1588;
w1590 <= pi0172 and not pi0262;
w1591 <= w1071 and w1590;
w1592 <= not w1589 and not w1591;
w1593 <= not pi0228 and not w1587;
w1594 <= not w1592 and w1593;
w1595 <= not w1050 and w1513;
w1596 <= pi0228 and not w1511;
w1597 <= not w1595 and w1596;
w1598 <= not w1060 and w1597;
w1599 <= not pi0216 and not w1598;
w1600 <= not w1594 and w1599;
w1601 <= w1509 and not w1600;
w1602 <= not w1522 and not w1601;
w1603 <= not pi0215 and not w1602;
w1604 <= w1586 and not w1603;
w1605 <= not w1051 and w1552;
w1606 <= w1584 and not w1605;
w1607 <= not pi0223 and not w1606;
w1608 <= w1580 and not w1607;
w1609 <= not pi0039 and not w1608;
w1610 <= not w1585 and w1609;
w1611 <= not w1604 and w1610;
w1612 <= not pi0038 and not w1579;
w1613 <= not w1611 and w1612;
w1614 <= not pi0100 and not w1578;
w1615 <= not w1613 and w1614;
w1616 <= not w93 and w1565;
w1617 <= not pi0262 and w957;
w1618 <= not w1192 and not w1510;
w1619 <= not w1617 and not w1618;
w1620 <= w1532 and not w1619;
w1621 <= not pi0216 and not w1620;
w1622 <= w1509 and not w1621;
w1623 <= not w1522 and not w1622;
w1624 <= not pi0215 and not w1623;
w1625 <= not w1507 and not w1624;
w1626 <= pi0299 and not w1625;
w1627 <= w93 and not w1563;
w1628 <= not w1626 and w1627;
w1629 <= pi0100 and not w1616;
w1630 <= not w1628 and w1629;
w1631 <= not w1615 and not w1630;
w1632 <= not pi0087 and not w1631;
w1633 <= not pi0075 and not w1577;
w1634 <= not w1632 and w1633;
w1635 <= not pi0092 and not w1576;
w1636 <= not w1634 and w1635;
w1637 <= w95 and not w1575;
w1638 <= not w1636 and w1637;
w1639 <= not pi0055 and not w1566;
w1640 <= not w1638 and w1639;
w1641 <= not pi0056 and not w1549;
w1642 <= not w1640 and w1641;
w1643 <= not pi0062 and not w1545;
w1644 <= not w1642 and w1643;
w1645 <= w891 and not w1541;
w1646 <= not w1644 and w1645;
w1647 <= not pi0249 and not w1527;
w1648 <= not w1646 and w1647;
w1649 <= not w891 and w1525;
w1650 <= not w894 and w1525;
w1651 <= not w1515 and not w1531;
w1652 <= not pi0216 and not w1651;
w1653 <= w1509 and not w1652;
w1654 <= not w1522 and not w1653;
w1655 <= not pi0215 and not w1654;
w1656 <= not w1507 and not w1655;
w1657 <= w894 and w1656;
w1658 <= pi0062 and not w1650;
w1659 <= not w1657 and w1658;
w1660 <= not w100 and not w1525;
w1661 <= w100 and not w1656;
w1662 <= pi0056 and not w1660;
w1663 <= not w1661 and w1662;
w1664 <= not w135 and w1525;
w1665 <= w135 and w1656;
w1666 <= pi0055 and not w1664;
w1667 <= not w1665 and w1666;
w1668 <= pi0299 and not w1525;
w1669 <= not w1562 and not w1668;
w1670 <= not w95 and w1669;
w1671 <= not w188 and w1669;
w1672 <= pi0299 and not w1656;
w1673 <= not w1562 and not w1672;
w1674 <= w188 and w1673;
w1675 <= not w1671 and not w1674;
w1676 <= w96 and not w1675;
w1677 <= not w96 and w1669;
w1678 <= pi0092 and not w1677;
w1679 <= not w1676 and w1678;
w1680 <= pi0075 and w1669;
w1681 <= pi0087 and w1675;
w1682 <= pi0038 and w1669;
w1683 <= pi0039 and not w1673;
w1684 <= pi0262 and w1071;
w1685 <= not pi0172 and not w1684;
w1686 <= pi0262 and not w1062;
w1687 <= not pi0262 and not w979;
w1688 <= pi0172 and not w1686;
w1689 <= not w1687 and w1688;
w1690 <= not w1685 and not w1689;
w1691 <= not pi0228 and not w1690;
w1692 <= not pi0216 and not w1597;
w1693 <= not w1691 and w1692;
w1694 <= w1509 and not w1693;
w1695 <= not w1522 and not w1694;
w1696 <= not pi0215 and not w1695;
w1697 <= w1586 and not w1696;
w1698 <= w1609 and not w1697;
w1699 <= not pi0038 and not w1683;
w1700 <= not w1698 and w1699;
w1701 <= not pi0100 and not w1682;
w1702 <= not w1700 and w1701;
w1703 <= not w93 and w1669;
w1704 <= not w1515 and not w1619;
w1705 <= not pi0216 and not w1704;
w1706 <= w1509 and not w1705;
w1707 <= not w1522 and not w1706;
w1708 <= not pi0215 and not w1707;
w1709 <= not w1507 and not w1708;
w1710 <= pi0299 and not w1709;
w1711 <= w93 and not w1562;
w1712 <= not w1710 and w1711;
w1713 <= pi0100 and not w1703;
w1714 <= not w1712 and w1713;
w1715 <= not w1702 and not w1714;
w1716 <= not pi0087 and not w1715;
w1717 <= not pi0075 and not w1681;
w1718 <= not w1716 and w1717;
w1719 <= not pi0092 and not w1680;
w1720 <= not w1718 and w1719;
w1721 <= w95 and not w1679;
w1722 <= not w1720 and w1721;
w1723 <= not pi0055 and not w1670;
w1724 <= not w1722 and w1723;
w1725 <= not pi0056 and not w1667;
w1726 <= not w1724 and w1725;
w1727 <= not pi0062 and not w1663;
w1728 <= not w1726 and w1727;
w1729 <= w891 and not w1659;
w1730 <= not w1728 and w1729;
w1731 <= pi0249 and not w1649;
w1732 <= not w1730 and w1731;
w1733 <= not w1648 and not w1732;
w1734 <= pi0215 and pi1141;
w1735 <= pi0216 and pi0270;
w1736 <= not pi0221 and not w1735;
w1737 <= not pi0105 and pi0171;
w1738 <= pi0861 and not w5;
w1739 <= pi0105 and not w1738;
w1740 <= pi0228 and not w1737;
w1741 <= not w1739 and w1740;
w1742 <= not pi0216 and not w1741;
w1743 <= not pi0171 and not pi0228;
w1744 <= w1742 and not w1743;
w1745 <= w1736 and not w1744;
w1746 <= not pi1141 and not w15;
w1747 <= not pi0935 and w15;
w1748 <= pi0221 and not w1746;
w1749 <= not w1747 and w1748;
w1750 <= not w1745 and not w1749;
w1751 <= not pi0215 and not w1750;
w1752 <= not w1734 and not w1751;
w1753 <= not w894 and w1752;
w1754 <= not pi0861 and w84;
w1755 <= pi0171 and not w84;
w1756 <= not pi0228 and not w1754;
w1757 <= not w1755 and w1756;
w1758 <= w1742 and not w1757;
w1759 <= w1736 and not w1758;
w1760 <= not w1749 and not w1759;
w1761 <= not pi0215 and not w1760;
w1762 <= not w1734 and not w1761;
w1763 <= w894 and w1762;
w1764 <= pi0062 and not w1753;
w1765 <= not w1763 and w1764;
w1766 <= not w100 and not w1752;
w1767 <= w100 and not w1762;
w1768 <= pi0056 and not w1766;
w1769 <= not w1767 and w1768;
w1770 <= not w135 and w1752;
w1771 <= w135 and w1762;
w1772 <= pi0055 and not w1770;
w1773 <= not w1771 and w1772;
w1774 <= pi0223 and pi1141;
w1775 <= pi0224 and pi0270;
w1776 <= not pi0222 and not w1775;
w1777 <= not pi0224 and not w1738;
w1778 <= w1776 and not w1777;
w1779 <= not pi1141 and not w154;
w1780 <= not pi0935 and w154;
w1781 <= pi0222 and not w1779;
w1782 <= not w1780 and w1781;
w1783 <= not w1778 and not w1782;
w1784 <= not pi0223 and not w1783;
w1785 <= not w1774 and not w1784;
w1786 <= not pi0299 and not w1785;
w1787 <= pi0299 and not w1752;
w1788 <= not w1786 and not w1787;
w1789 <= not w95 and w1788;
w1790 <= not w188 and w1788;
w1791 <= pi0299 and not w1762;
w1792 <= not w1786 and not w1791;
w1793 <= w188 and w1792;
w1794 <= not w1790 and not w1793;
w1795 <= w96 and not w1794;
w1796 <= not w96 and w1788;
w1797 <= pi0092 and not w1796;
w1798 <= not w1795 and w1797;
w1799 <= pi0075 and w1788;
w1800 <= pi0087 and w1794;
w1801 <= pi0038 and w1788;
w1802 <= pi0039 and not w1792;
w1803 <= not pi0299 and not w1774;
w1804 <= pi0861 and w1051;
w1805 <= not pi0224 and not w1804;
w1806 <= w1776 and not w1805;
w1807 <= not w1782 and not w1806;
w1808 <= w1803 and w1807;
w1809 <= pi0299 and not w1734;
w1810 <= pi0861 and w1062;
w1811 <= not pi0171 and not w1810;
w1812 <= pi0171 and w1071;
w1813 <= not w1811 and not w1812;
w1814 <= pi0861 and not w1813;
w1815 <= not w979 and w1811;
w1816 <= not w1814 and not w1815;
w1817 <= not pi0228 and not w1816;
w1818 <= not w1060 and w1741;
w1819 <= not pi0216 and not w1818;
w1820 <= not w1817 and w1819;
w1821 <= w1736 and not w1820;
w1822 <= not w1749 and not w1821;
w1823 <= not pi0215 and not w1822;
w1824 <= w1809 and not w1823;
w1825 <= not w1051 and w1776;
w1826 <= w1807 and not w1825;
w1827 <= not pi0223 and not w1826;
w1828 <= w1803 and not w1827;
w1829 <= not pi0039 and not w1828;
w1830 <= not w1808 and w1829;
w1831 <= not w1824 and w1830;
w1832 <= not pi0038 and not w1802;
w1833 <= not w1831 and w1832;
w1834 <= not pi0100 and not w1801;
w1835 <= not w1833 and w1834;
w1836 <= not w93 and w1788;
w1837 <= not pi0861 and w957;
w1838 <= pi0171 and not w957;
w1839 <= not pi0228 and not w1837;
w1840 <= not w1838 and w1839;
w1841 <= w1742 and not w1840;
w1842 <= w1736 and not w1841;
w1843 <= not w1749 and not w1842;
w1844 <= not pi0215 and not w1843;
w1845 <= not w1734 and not w1844;
w1846 <= pi0299 and not w1845;
w1847 <= w93 and not w1786;
w1848 <= not w1846 and w1847;
w1849 <= pi0100 and not w1836;
w1850 <= not w1848 and w1849;
w1851 <= not w1835 and not w1850;
w1852 <= not pi0087 and not w1851;
w1853 <= not pi0075 and not w1800;
w1854 <= not w1852 and w1853;
w1855 <= not pi0092 and not w1799;
w1856 <= not w1854 and w1855;
w1857 <= w95 and not w1798;
w1858 <= not w1856 and w1857;
w1859 <= not pi0055 and not w1789;
w1860 <= not w1858 and w1859;
w1861 <= not pi0056 and not w1773;
w1862 <= not w1860 and w1861;
w1863 <= not pi0062 and not w1769;
w1864 <= not w1862 and w1863;
w1865 <= not pi0241 and w891;
w1866 <= not w1765 and w1865;
w1867 <= not w1864 and w1866;
w1868 <= not w1010 and w1742;
w1869 <= not w1757 and w1868;
w1870 <= w1736 and not w1869;
w1871 <= not w1749 and not w1870;
w1872 <= not pi0215 and not w1871;
w1873 <= not w1734 and not w1872;
w1874 <= w894 and w1873;
w1875 <= w1119 and not w1735;
w1876 <= w1752 and not w1875;
w1877 <= not w894 and w1876;
w1878 <= pi0062 and not w1877;
w1879 <= not w1874 and w1878;
w1880 <= not w100 and not w1876;
w1881 <= w100 and not w1873;
w1882 <= pi0056 and not w1880;
w1883 <= not w1881 and w1882;
w1884 <= w135 and w1873;
w1885 <= not w135 and w1876;
w1886 <= pi0055 and not w1885;
w1887 <= not w1884 and w1886;
w1888 <= not w1035 and not w1786;
w1889 <= pi0299 and not w1876;
w1890 <= w1888 and not w1889;
w1891 <= not w95 and w1890;
w1892 <= not w188 and w1890;
w1893 <= pi0299 and not w1873;
w1894 <= w1888 and not w1893;
w1895 <= w188 and w1894;
w1896 <= not w1892 and not w1895;
w1897 <= w96 and not w1896;
w1898 <= not w96 and w1890;
w1899 <= pi0092 and not w1898;
w1900 <= not w1897 and w1899;
w1901 <= pi0075 and w1890;
w1902 <= pi0087 and w1896;
w1903 <= pi0038 and w1890;
w1904 <= pi0039 and not w1894;
w1905 <= not pi0861 and w1071;
w1906 <= not pi0171 and not w1905;
w1907 <= not pi0861 and not w1062;
w1908 <= pi0861 and not w979;
w1909 <= pi0171 and not w1907;
w1910 <= not w1908 and w1909;
w1911 <= not w1906 and not w1910;
w1912 <= not pi0228 and not w1911;
w1913 <= not w1356 and w1742;
w1914 <= not w1912 and w1913;
w1915 <= w1736 and not w1914;
w1916 <= not w1749 and not w1915;
w1917 <= not pi0215 and not w1916;
w1918 <= w1809 and not w1917;
w1919 <= w1829 and not w1918;
w1920 <= not pi0038 and not w1904;
w1921 <= not w1919 and w1920;
w1922 <= not pi0100 and not w1903;
w1923 <= not w1921 and w1922;
w1924 <= not w93 and w1890;
w1925 <= not w1840 and w1868;
w1926 <= w1736 and not w1925;
w1927 <= not w1749 and not w1926;
w1928 <= not pi0215 and not w1927;
w1929 <= not w1734 and not w1928;
w1930 <= pi0299 and not w1929;
w1931 <= w93 and w1888;
w1932 <= not w1930 and w1931;
w1933 <= pi0100 and not w1924;
w1934 <= not w1932 and w1933;
w1935 <= not w1923 and not w1934;
w1936 <= not pi0087 and not w1935;
w1937 <= not pi0075 and not w1902;
w1938 <= not w1936 and w1937;
w1939 <= not pi0092 and not w1901;
w1940 <= not w1938 and w1939;
w1941 <= w95 and not w1900;
w1942 <= not w1940 and w1941;
w1943 <= not pi0055 and not w1891;
w1944 <= not w1942 and w1943;
w1945 <= not pi0056 and not w1887;
w1946 <= not w1944 and w1945;
w1947 <= not pi0062 and not w1883;
w1948 <= not w1946 and w1947;
w1949 <= pi0241 and w891;
w1950 <= not w1879 and w1949;
w1951 <= not w1948 and w1950;
w1952 <= pi0241 and w1875;
w1953 <= not w891 and not w1952;
w1954 <= w1752 and w1953;
w1955 <= not w1951 and not w1954;
w1956 <= not w1867 and w1955;
w1957 <= pi0215 and pi1140;
w1958 <= pi0216 and pi0282;
w1959 <= not pi0221 and not w1958;
w1960 <= not pi0105 and pi0170;
w1961 <= pi0869 and not w5;
w1962 <= pi0105 and not w1961;
w1963 <= pi0228 and not w1960;
w1964 <= not w1962 and w1963;
w1965 <= not pi0216 and not w1964;
w1966 <= not pi0170 and not pi0228;
w1967 <= w1965 and not w1966;
w1968 <= w1959 and not w1967;
w1969 <= not pi1140 and not w15;
w1970 <= not pi0921 and w15;
w1971 <= pi0221 and not w1969;
w1972 <= not w1970 and w1971;
w1973 <= not w1968 and not w1972;
w1974 <= not pi0215 and not w1973;
w1975 <= not w1957 and not w1974;
w1976 <= not w894 and w1975;
w1977 <= not pi0869 and w84;
w1978 <= pi0170 and not w84;
w1979 <= not pi0228 and not w1977;
w1980 <= not w1978 and w1979;
w1981 <= w1965 and not w1980;
w1982 <= w1959 and not w1981;
w1983 <= not w1972 and not w1982;
w1984 <= not pi0215 and not w1983;
w1985 <= not w1957 and not w1984;
w1986 <= w894 and w1985;
w1987 <= pi0062 and not w1976;
w1988 <= not w1986 and w1987;
w1989 <= not w100 and not w1975;
w1990 <= w100 and not w1985;
w1991 <= pi0056 and not w1989;
w1992 <= not w1990 and w1991;
w1993 <= not w135 and w1975;
w1994 <= w135 and w1985;
w1995 <= pi0055 and not w1993;
w1996 <= not w1994 and w1995;
w1997 <= pi0223 and pi1140;
w1998 <= pi0224 and pi0282;
w1999 <= not pi0222 and not w1998;
w2000 <= not pi0224 and not w1961;
w2001 <= w1999 and not w2000;
w2002 <= not pi1140 and not w154;
w2003 <= not pi0921 and w154;
w2004 <= pi0222 and not w2002;
w2005 <= not w2003 and w2004;
w2006 <= not w2001 and not w2005;
w2007 <= not pi0223 and not w2006;
w2008 <= not w1997 and not w2007;
w2009 <= not pi0299 and not w2008;
w2010 <= pi0299 and not w1975;
w2011 <= not w2009 and not w2010;
w2012 <= not w95 and w2011;
w2013 <= not w188 and w2011;
w2014 <= pi0299 and not w1985;
w2015 <= not w2009 and not w2014;
w2016 <= w188 and w2015;
w2017 <= not w2013 and not w2016;
w2018 <= w96 and not w2017;
w2019 <= not w96 and w2011;
w2020 <= pi0092 and not w2019;
w2021 <= not w2018 and w2020;
w2022 <= pi0075 and w2011;
w2023 <= pi0087 and w2017;
w2024 <= pi0038 and w2011;
w2025 <= pi0039 and not w2015;
w2026 <= not pi0299 and not w1997;
w2027 <= pi0869 and w1051;
w2028 <= not pi0224 and not w2027;
w2029 <= w1999 and not w2028;
w2030 <= not w2005 and not w2029;
w2031 <= w2026 and w2030;
w2032 <= pi0299 and not w1957;
w2033 <= pi0869 and w1062;
w2034 <= not pi0170 and not w2033;
w2035 <= pi0170 and w1071;
w2036 <= not w2034 and not w2035;
w2037 <= pi0869 and not w2036;
w2038 <= not w979 and w2034;
w2039 <= not w2037 and not w2038;
w2040 <= not pi0228 and not w2039;
w2041 <= not w1060 and w1964;
w2042 <= not pi0216 and not w2041;
w2043 <= not w2040 and w2042;
w2044 <= w1959 and not w2043;
w2045 <= not w1972 and not w2044;
w2046 <= not pi0215 and not w2045;
w2047 <= w2032 and not w2046;
w2048 <= not w1051 and w1999;
w2049 <= w2030 and not w2048;
w2050 <= not pi0223 and not w2049;
w2051 <= w2026 and not w2050;
w2052 <= not pi0039 and not w2051;
w2053 <= not w2031 and w2052;
w2054 <= not w2047 and w2053;
w2055 <= not pi0038 and not w2025;
w2056 <= not w2054 and w2055;
w2057 <= not pi0100 and not w2024;
w2058 <= not w2056 and w2057;
w2059 <= not w93 and w2011;
w2060 <= not pi0869 and w957;
w2061 <= pi0170 and not w957;
w2062 <= not pi0228 and not w2060;
w2063 <= not w2061 and w2062;
w2064 <= w1965 and not w2063;
w2065 <= w1959 and not w2064;
w2066 <= not w1972 and not w2065;
w2067 <= not pi0215 and not w2066;
w2068 <= not w1957 and not w2067;
w2069 <= pi0299 and not w2068;
w2070 <= w93 and not w2009;
w2071 <= not w2069 and w2070;
w2072 <= pi0100 and not w2059;
w2073 <= not w2071 and w2072;
w2074 <= not w2058 and not w2073;
w2075 <= not pi0087 and not w2074;
w2076 <= not pi0075 and not w2023;
w2077 <= not w2075 and w2076;
w2078 <= not pi0092 and not w2022;
w2079 <= not w2077 and w2078;
w2080 <= w95 and not w2021;
w2081 <= not w2079 and w2080;
w2082 <= not pi0055 and not w2012;
w2083 <= not w2081 and w2082;
w2084 <= not pi0056 and not w1996;
w2085 <= not w2083 and w2084;
w2086 <= not pi0062 and not w1992;
w2087 <= not w2085 and w2086;
w2088 <= not pi0248 and w891;
w2089 <= not w1988 and w2088;
w2090 <= not w2087 and w2089;
w2091 <= not w1010 and w1965;
w2092 <= not w1980 and w2091;
w2093 <= w1959 and not w2092;
w2094 <= not w1972 and not w2093;
w2095 <= not pi0215 and not w2094;
w2096 <= not w1957 and not w2095;
w2097 <= w894 and w2096;
w2098 <= w1119 and not w1958;
w2099 <= w1975 and not w2098;
w2100 <= not w894 and w2099;
w2101 <= pi0062 and not w2100;
w2102 <= not w2097 and w2101;
w2103 <= not w100 and not w2099;
w2104 <= w100 and not w2096;
w2105 <= pi0056 and not w2103;
w2106 <= not w2104 and w2105;
w2107 <= w135 and w2096;
w2108 <= not w135 and w2099;
w2109 <= pi0055 and not w2108;
w2110 <= not w2107 and w2109;
w2111 <= not w1035 and not w2009;
w2112 <= pi0299 and not w2099;
w2113 <= w2111 and not w2112;
w2114 <= not w95 and w2113;
w2115 <= not w188 and w2113;
w2116 <= pi0299 and not w2096;
w2117 <= w2111 and not w2116;
w2118 <= w188 and w2117;
w2119 <= not w2115 and not w2118;
w2120 <= w96 and not w2119;
w2121 <= not w96 and w2113;
w2122 <= pi0092 and not w2121;
w2123 <= not w2120 and w2122;
w2124 <= pi0075 and w2113;
w2125 <= pi0087 and w2119;
w2126 <= pi0038 and w2113;
w2127 <= pi0039 and not w2117;
w2128 <= not pi0869 and w1071;
w2129 <= not pi0170 and not w2128;
w2130 <= not pi0869 and not w1062;
w2131 <= pi0869 and not w979;
w2132 <= pi0170 and not w2130;
w2133 <= not w2131 and w2132;
w2134 <= not w2129 and not w2133;
w2135 <= not pi0228 and not w2134;
w2136 <= not w1356 and w1965;
w2137 <= not w2135 and w2136;
w2138 <= w1959 and not w2137;
w2139 <= not w1972 and not w2138;
w2140 <= not pi0215 and not w2139;
w2141 <= w2032 and not w2140;
w2142 <= w2052 and not w2141;
w2143 <= not pi0038 and not w2127;
w2144 <= not w2142 and w2143;
w2145 <= not pi0100 and not w2126;
w2146 <= not w2144 and w2145;
w2147 <= not w93 and w2113;
w2148 <= not w2063 and w2091;
w2149 <= w1959 and not w2148;
w2150 <= not w1972 and not w2149;
w2151 <= not pi0215 and not w2150;
w2152 <= not w1957 and not w2151;
w2153 <= pi0299 and not w2152;
w2154 <= w93 and w2111;
w2155 <= not w2153 and w2154;
w2156 <= pi0100 and not w2147;
w2157 <= not w2155 and w2156;
w2158 <= not w2146 and not w2157;
w2159 <= not pi0087 and not w2158;
w2160 <= not pi0075 and not w2125;
w2161 <= not w2159 and w2160;
w2162 <= not pi0092 and not w2124;
w2163 <= not w2161 and w2162;
w2164 <= w95 and not w2123;
w2165 <= not w2163 and w2164;
w2166 <= not pi0055 and not w2114;
w2167 <= not w2165 and w2166;
w2168 <= not pi0056 and not w2110;
w2169 <= not w2167 and w2168;
w2170 <= not pi0062 and not w2106;
w2171 <= not w2169 and w2170;
w2172 <= pi0248 and w891;
w2173 <= not w2102 and w2172;
w2174 <= not w2171 and w2173;
w2175 <= pi0248 and w2098;
w2176 <= not w891 and not w2175;
w2177 <= w1975 and w2176;
w2178 <= not w2174 and not w2177;
w2179 <= not w2090 and w2178;
w2180 <= pi0215 and pi1139;
w2181 <= pi0216 and not pi1139;
w2182 <= pi0833 and pi0920;
w2183 <= not pi0833 and pi1139;
w2184 <= not pi0216 and not w2182;
w2185 <= not w2183 and w2184;
w2186 <= pi0221 and not w2185;
w2187 <= not w2181 and w2186;
w2188 <= pi0216 and pi0281;
w2189 <= not pi0221 and not w2188;
w2190 <= not pi0216 and not pi0862;
w2191 <= w1193 and w2190;
w2192 <= w2189 and not w2191;
w2193 <= not w2187 and not w2192;
w2194 <= not pi0216 and not w2186;
w2195 <= pi0148 and not w4;
w2196 <= w2194 and w2195;
w2197 <= not pi0215 and not w2196;
w2198 <= not w2193 and w2197;
w2199 <= not w2180 and not w2198;
w2200 <= not w1013 and not w2199;
w2201 <= not w891 and not w2200;
w2202 <= not w894 and not w2200;
w2203 <= not pi0148 and not pi0215;
w2204 <= pi0862 and not w1010;
w2205 <= not w4 and not w898;
w2206 <= not pi0216 and not w2204;
w2207 <= not w2205 and w2206;
w2208 <= w2189 and not w2207;
w2209 <= not w2187 and not w2208;
w2210 <= w2203 and not w2209;
w2211 <= pi0148 and not pi0215;
w2212 <= not w898 and not w1193;
w2213 <= w2190 and not w2212;
w2214 <= w2189 and not w2213;
w2215 <= not w2187 and not w2214;
w2216 <= w2194 and w2212;
w2217 <= w2211 and not w2216;
w2218 <= not w2215 and w2217;
w2219 <= not w2180 and not w2218;
w2220 <= not w2210 and w2219;
w2221 <= w894 and w2220;
w2222 <= pi0062 and not w2202;
w2223 <= not w2221 and w2222;
w2224 <= w100 and not w2220;
w2225 <= not w100 and w2200;
w2226 <= pi0056 and not w2225;
w2227 <= not w2224 and w2226;
w2228 <= not w135 and not w2200;
w2229 <= w135 and w2220;
w2230 <= pi0055 and not w2228;
w2231 <= not w2229 and w2230;
w2232 <= pi0223 and pi1139;
w2233 <= not pi1139 and not w154;
w2234 <= not pi0920 and w154;
w2235 <= pi0222 and not w2233;
w2236 <= not w2234 and w2235;
w2237 <= not pi0224 and not w2232;
w2238 <= not w2236 and w2237;
w2239 <= w5 and w2238;
w2240 <= not pi0862 and w2238;
w2241 <= pi0224 and pi0281;
w2242 <= not pi0222 and not w2241;
w2243 <= not w2236 and not w2242;
w2244 <= not pi0223 and not w2243;
w2245 <= not w2232 and not w2244;
w2246 <= not pi0299 and not w2245;
w2247 <= not w2240 and w2246;
w2248 <= not w2239 and w2247;
w2249 <= pi0299 and w2200;
w2250 <= not w2248 and not w2249;
w2251 <= not w95 and w2250;
w2252 <= not w188 and w2250;
w2253 <= pi0299 and not w2220;
w2254 <= not w2248 and not w2253;
w2255 <= w188 and w2254;
w2256 <= not w2252 and not w2255;
w2257 <= w96 and not w2256;
w2258 <= not w96 and w2250;
w2259 <= pi0092 and not w2258;
w2260 <= not w2257 and w2259;
w2261 <= pi0075 and w2250;
w2262 <= pi0087 and w2256;
w2263 <= not w93 and w2250;
w2264 <= not w4 and not w1192;
w2265 <= w2189 and w2264;
w2266 <= w2209 and not w2265;
w2267 <= w2203 and not w2266;
w2268 <= w1194 and w2189;
w2269 <= w2215 and not w2268;
w2270 <= w1194 and w2194;
w2271 <= w2211 and not w2270;
w2272 <= not w2269 and w2271;
w2273 <= not w2180 and not w2267;
w2274 <= not w2272 and w2273;
w2275 <= pi0299 and not w2274;
w2276 <= w93 and not w2248;
w2277 <= not w2275 and w2276;
w2278 <= pi0100 and not w2263;
w2279 <= not w2277 and w2278;
w2280 <= pi0038 and w2250;
w2281 <= pi0039 and not w2254;
w2282 <= not w1051 and w2238;
w2283 <= not w2240 and not w2245;
w2284 <= not w2282 and w2283;
w2285 <= not pi0299 and not w2284;
w2286 <= not w1074 and w2190;
w2287 <= w2189 and not w2286;
w2288 <= not w2187 and not w2287;
w2289 <= w1074 and w2194;
w2290 <= w2211 and not w2289;
w2291 <= not w2288 and w2290;
w2292 <= pi0862 and not w1064;
w2293 <= not pi0228 and w979;
w2294 <= not w4 and not w2293;
w2295 <= not pi0862 and w2294;
w2296 <= not pi0216 and not w2292;
w2297 <= not w2295 and w2296;
w2298 <= w2189 and not w2297;
w2299 <= not w2187 and not w2298;
w2300 <= w2203 and not w2299;
w2301 <= pi0299 and not w2180;
w2302 <= not w2291 and w2301;
w2303 <= not w2300 and w2302;
w2304 <= not pi0039 and not w2285;
w2305 <= not w2303 and w2304;
w2306 <= not pi0038 and not w2281;
w2307 <= not w2305 and w2306;
w2308 <= not pi0100 and not w2280;
w2309 <= not w2307 and w2308;
w2310 <= not w2279 and not w2309;
w2311 <= not pi0087 and not w2310;
w2312 <= not pi0075 and not w2262;
w2313 <= not w2311 and w2312;
w2314 <= not pi0092 and not w2261;
w2315 <= not w2313 and w2314;
w2316 <= w95 and not w2260;
w2317 <= not w2315 and w2316;
w2318 <= not pi0055 and not w2251;
w2319 <= not w2317 and w2318;
w2320 <= not pi0056 and not w2231;
w2321 <= not w2319 and w2320;
w2322 <= not pi0062 and not w2227;
w2323 <= not w2321 and w2322;
w2324 <= w891 and not w2223;
w2325 <= not w2323 and w2324;
w2326 <= not pi0247 and not w2201;
w2327 <= not w2325 and w2326;
w2328 <= not w891 and w2199;
w2329 <= not w894 and w2199;
w2330 <= w2197 and not w2215;
w2331 <= w2219 and not w2330;
w2332 <= w894 and w2331;
w2333 <= pi0062 and not w2329;
w2334 <= not w2332 and w2333;
w2335 <= not w100 and not w2199;
w2336 <= w100 and not w2331;
w2337 <= pi0056 and not w2335;
w2338 <= not w2336 and w2337;
w2339 <= not w135 and w2199;
w2340 <= w135 and w2331;
w2341 <= pi0055 and not w2339;
w2342 <= not w2340 and w2341;
w2343 <= not w1035 and not w2247;
w2344 <= pi0299 and not w2199;
w2345 <= w2343 and not w2344;
w2346 <= not w95 and w2345;
w2347 <= not w188 and w2345;
w2348 <= pi0299 and not w2331;
w2349 <= w2343 and not w2348;
w2350 <= w188 and w2349;
w2351 <= not w2347 and not w2350;
w2352 <= w96 and not w2351;
w2353 <= not w96 and w2345;
w2354 <= pi0092 and not w2353;
w2355 <= not w2352 and w2354;
w2356 <= pi0075 and w2345;
w2357 <= pi0087 and w2351;
w2358 <= not w93 and w2345;
w2359 <= w2203 and not w2269;
w2360 <= not pi0216 and not w2187;
w2361 <= w2264 and w2360;
w2362 <= w2211 and not w2215;
w2363 <= not w2361 and w2362;
w2364 <= not w2180 and not w2363;
w2365 <= not w2359 and w2364;
w2366 <= pi0299 and not w2365;
w2367 <= w93 and w2343;
w2368 <= not w2366 and w2367;
w2369 <= pi0100 and not w2358;
w2370 <= not w2368 and w2369;
w2371 <= pi0038 and w2345;
w2372 <= pi0039 and not w2349;
w2373 <= w1051 and w2240;
w2374 <= w2246 and not w2373;
w2375 <= pi0862 and not w2294;
w2376 <= not pi0862 and w1064;
w2377 <= not pi0216 and not w2376;
w2378 <= not w2375 and w2377;
w2379 <= w2189 and not w2378;
w2380 <= not w2187 and not w2379;
w2381 <= w2211 and not w2380;
w2382 <= w2203 and not w2288;
w2383 <= not w2180 and not w2382;
w2384 <= not w2381 and w2383;
w2385 <= pi0299 and not w2384;
w2386 <= not w2374 and not w2385;
w2387 <= not pi0039 and not w2386;
w2388 <= not pi0038 and not w2372;
w2389 <= not w2387 and w2388;
w2390 <= not pi0100 and not w2371;
w2391 <= not w2389 and w2390;
w2392 <= not w2370 and not w2391;
w2393 <= not pi0087 and not w2392;
w2394 <= not pi0075 and not w2357;
w2395 <= not w2393 and w2394;
w2396 <= not pi0092 and not w2356;
w2397 <= not w2395 and w2396;
w2398 <= w95 and not w2355;
w2399 <= not w2397 and w2398;
w2400 <= not pi0055 and not w2346;
w2401 <= not w2399 and w2400;
w2402 <= not pi0056 and not w2342;
w2403 <= not w2401 and w2402;
w2404 <= not pi0062 and not w2338;
w2405 <= not w2403 and w2404;
w2406 <= w891 and not w2334;
w2407 <= not w2405 and w2406;
w2408 <= pi0247 and not w2328;
w2409 <= not w2407 and w2408;
w2410 <= not w2327 and not w2409;
w2411 <= pi0215 and pi1138;
w2412 <= pi0216 and pi0269;
w2413 <= not pi0221 and not w2412;
w2414 <= not pi0105 and pi0169;
w2415 <= pi0877 and not w5;
w2416 <= pi0105 and not w2415;
w2417 <= pi0228 and not w2414;
w2418 <= not w2416 and w2417;
w2419 <= not pi0216 and not w2418;
w2420 <= not pi0169 and not pi0228;
w2421 <= w2419 and not w2420;
w2422 <= w2413 and not w2421;
w2423 <= not pi1138 and not w15;
w2424 <= not pi0940 and w15;
w2425 <= pi0221 and not w2423;
w2426 <= not w2424 and w2425;
w2427 <= not w2422 and not w2426;
w2428 <= not pi0215 and not w2427;
w2429 <= not w2411 and not w2428;
w2430 <= not w894 and w2429;
w2431 <= not pi0877 and w84;
w2432 <= pi0169 and not w84;
w2433 <= not pi0228 and not w2431;
w2434 <= not w2432 and w2433;
w2435 <= w2419 and not w2434;
w2436 <= w2413 and not w2435;
w2437 <= not w2426 and not w2436;
w2438 <= not pi0215 and not w2437;
w2439 <= not w2411 and not w2438;
w2440 <= w894 and w2439;
w2441 <= pi0062 and not w2430;
w2442 <= not w2440 and w2441;
w2443 <= not w100 and not w2429;
w2444 <= w100 and not w2439;
w2445 <= pi0056 and not w2443;
w2446 <= not w2444 and w2445;
w2447 <= not w135 and w2429;
w2448 <= w135 and w2439;
w2449 <= pi0055 and not w2447;
w2450 <= not w2448 and w2449;
w2451 <= pi0223 and pi1138;
w2452 <= pi0224 and pi0269;
w2453 <= not pi0222 and not w2452;
w2454 <= not pi0224 and not w2415;
w2455 <= w2453 and not w2454;
w2456 <= not pi1138 and not w154;
w2457 <= not pi0940 and w154;
w2458 <= pi0222 and not w2456;
w2459 <= not w2457 and w2458;
w2460 <= not w2455 and not w2459;
w2461 <= not pi0223 and not w2460;
w2462 <= not w2451 and not w2461;
w2463 <= not pi0299 and not w2462;
w2464 <= pi0299 and not w2429;
w2465 <= not w2463 and not w2464;
w2466 <= not w95 and w2465;
w2467 <= not w188 and w2465;
w2468 <= pi0299 and not w2439;
w2469 <= not w2463 and not w2468;
w2470 <= w188 and w2469;
w2471 <= not w2467 and not w2470;
w2472 <= w96 and not w2471;
w2473 <= not w96 and w2465;
w2474 <= pi0092 and not w2473;
w2475 <= not w2472 and w2474;
w2476 <= pi0075 and w2465;
w2477 <= pi0087 and w2471;
w2478 <= pi0038 and w2465;
w2479 <= pi0039 and not w2469;
w2480 <= not pi0299 and not w2451;
w2481 <= pi0877 and w1051;
w2482 <= not pi0224 and not w2481;
w2483 <= w2453 and not w2482;
w2484 <= not w2459 and not w2483;
w2485 <= w2480 and w2484;
w2486 <= pi0299 and not w2411;
w2487 <= pi0877 and w1062;
w2488 <= not pi0169 and not w2487;
w2489 <= pi0169 and w1071;
w2490 <= not w2488 and not w2489;
w2491 <= pi0877 and not w2490;
w2492 <= not w979 and w2488;
w2493 <= not w2491 and not w2492;
w2494 <= not pi0228 and not w2493;
w2495 <= not w1060 and w2418;
w2496 <= not pi0216 and not w2495;
w2497 <= not w2494 and w2496;
w2498 <= w2413 and not w2497;
w2499 <= not w2426 and not w2498;
w2500 <= not pi0215 and not w2499;
w2501 <= w2486 and not w2500;
w2502 <= not w1051 and w2453;
w2503 <= w2484 and not w2502;
w2504 <= not pi0223 and not w2503;
w2505 <= w2480 and not w2504;
w2506 <= not pi0039 and not w2505;
w2507 <= not w2485 and w2506;
w2508 <= not w2501 and w2507;
w2509 <= not pi0038 and not w2479;
w2510 <= not w2508 and w2509;
w2511 <= not pi0100 and not w2478;
w2512 <= not w2510 and w2511;
w2513 <= not w93 and w2465;
w2514 <= not pi0877 and w957;
w2515 <= pi0169 and not w957;
w2516 <= not pi0228 and not w2514;
w2517 <= not w2515 and w2516;
w2518 <= w2419 and not w2517;
w2519 <= w2413 and not w2518;
w2520 <= not w2426 and not w2519;
w2521 <= not pi0215 and not w2520;
w2522 <= not w2411 and not w2521;
w2523 <= pi0299 and not w2522;
w2524 <= w93 and not w2463;
w2525 <= not w2523 and w2524;
w2526 <= pi0100 and not w2513;
w2527 <= not w2525 and w2526;
w2528 <= not w2512 and not w2527;
w2529 <= not pi0087 and not w2528;
w2530 <= not pi0075 and not w2477;
w2531 <= not w2529 and w2530;
w2532 <= not pi0092 and not w2476;
w2533 <= not w2531 and w2532;
w2534 <= w95 and not w2475;
w2535 <= not w2533 and w2534;
w2536 <= not pi0055 and not w2466;
w2537 <= not w2535 and w2536;
w2538 <= not pi0056 and not w2450;
w2539 <= not w2537 and w2538;
w2540 <= not pi0062 and not w2446;
w2541 <= not w2539 and w2540;
w2542 <= not pi0246 and w891;
w2543 <= not w2442 and w2542;
w2544 <= not w2541 and w2543;
w2545 <= not w1010 and w2419;
w2546 <= not w2434 and w2545;
w2547 <= w2413 and not w2546;
w2548 <= not w2426 and not w2547;
w2549 <= not pi0215 and not w2548;
w2550 <= not w2411 and not w2549;
w2551 <= w894 and w2550;
w2552 <= w1119 and not w2412;
w2553 <= w2429 and not w2552;
w2554 <= not w894 and w2553;
w2555 <= pi0062 and not w2554;
w2556 <= not w2551 and w2555;
w2557 <= not w100 and not w2553;
w2558 <= w100 and not w2550;
w2559 <= pi0056 and not w2557;
w2560 <= not w2558 and w2559;
w2561 <= w135 and w2550;
w2562 <= not w135 and w2553;
w2563 <= pi0055 and not w2562;
w2564 <= not w2561 and w2563;
w2565 <= not w1035 and not w2463;
w2566 <= pi0299 and not w2553;
w2567 <= w2565 and not w2566;
w2568 <= not w95 and w2567;
w2569 <= not w188 and w2567;
w2570 <= pi0299 and not w2550;
w2571 <= w2565 and not w2570;
w2572 <= w188 and w2571;
w2573 <= not w2569 and not w2572;
w2574 <= w96 and not w2573;
w2575 <= not w96 and w2567;
w2576 <= pi0092 and not w2575;
w2577 <= not w2574 and w2576;
w2578 <= pi0075 and w2567;
w2579 <= pi0087 and w2573;
w2580 <= pi0038 and w2567;
w2581 <= pi0039 and not w2571;
w2582 <= not pi0877 and w1071;
w2583 <= not pi0169 and not w2582;
w2584 <= not pi0877 and not w1062;
w2585 <= pi0877 and not w979;
w2586 <= pi0169 and not w2584;
w2587 <= not w2585 and w2586;
w2588 <= not w2583 and not w2587;
w2589 <= not pi0228 and not w2588;
w2590 <= not w1356 and w2419;
w2591 <= not w2589 and w2590;
w2592 <= w2413 and not w2591;
w2593 <= not w2426 and not w2592;
w2594 <= not pi0215 and not w2593;
w2595 <= w2486 and not w2594;
w2596 <= w2506 and not w2595;
w2597 <= not pi0038 and not w2581;
w2598 <= not w2596 and w2597;
w2599 <= not pi0100 and not w2580;
w2600 <= not w2598 and w2599;
w2601 <= not w93 and w2567;
w2602 <= not w2517 and w2545;
w2603 <= w2413 and not w2602;
w2604 <= not w2426 and not w2603;
w2605 <= not pi0215 and not w2604;
w2606 <= not w2411 and not w2605;
w2607 <= pi0299 and not w2606;
w2608 <= w93 and w2565;
w2609 <= not w2607 and w2608;
w2610 <= pi0100 and not w2601;
w2611 <= not w2609 and w2610;
w2612 <= not w2600 and not w2611;
w2613 <= not pi0087 and not w2612;
w2614 <= not pi0075 and not w2579;
w2615 <= not w2613 and w2614;
w2616 <= not pi0092 and not w2578;
w2617 <= not w2615 and w2616;
w2618 <= w95 and not w2577;
w2619 <= not w2617 and w2618;
w2620 <= not pi0055 and not w2568;
w2621 <= not w2619 and w2620;
w2622 <= not pi0056 and not w2564;
w2623 <= not w2621 and w2622;
w2624 <= not pi0062 and not w2560;
w2625 <= not w2623 and w2624;
w2626 <= pi0246 and w891;
w2627 <= not w2556 and w2626;
w2628 <= not w2625 and w2627;
w2629 <= pi0246 and w2552;
w2630 <= not w891 and not w2629;
w2631 <= w2429 and w2630;
w2632 <= not w2628 and not w2631;
w2633 <= not w2544 and w2632;
w2634 <= pi0215 and pi1137;
w2635 <= pi0216 and pi0280;
w2636 <= not pi0221 and not w2635;
w2637 <= not pi0105 and pi0168;
w2638 <= pi0878 and not w5;
w2639 <= pi0105 and not w2638;
w2640 <= pi0228 and not w2637;
w2641 <= not w2639 and w2640;
w2642 <= not pi0216 and not w2641;
w2643 <= not pi0168 and not pi0228;
w2644 <= w2642 and not w2643;
w2645 <= w2636 and not w2644;
w2646 <= not pi1137 and not w15;
w2647 <= not pi0933 and w15;
w2648 <= pi0221 and not w2646;
w2649 <= not w2647 and w2648;
w2650 <= not w2645 and not w2649;
w2651 <= not pi0215 and not w2650;
w2652 <= not w2634 and not w2651;
w2653 <= not w894 and w2652;
w2654 <= not pi0878 and w84;
w2655 <= pi0168 and not w84;
w2656 <= not pi0228 and not w2654;
w2657 <= not w2655 and w2656;
w2658 <= w2642 and not w2657;
w2659 <= w2636 and not w2658;
w2660 <= not w2649 and not w2659;
w2661 <= not pi0215 and not w2660;
w2662 <= not w2634 and not w2661;
w2663 <= w894 and w2662;
w2664 <= pi0062 and not w2653;
w2665 <= not w2663 and w2664;
w2666 <= not w100 and not w2652;
w2667 <= w100 and not w2662;
w2668 <= pi0056 and not w2666;
w2669 <= not w2667 and w2668;
w2670 <= not w135 and w2652;
w2671 <= w135 and w2662;
w2672 <= pi0055 and not w2670;
w2673 <= not w2671 and w2672;
w2674 <= pi0223 and pi1137;
w2675 <= pi0224 and pi0280;
w2676 <= not pi0222 and not w2675;
w2677 <= not pi0224 and not w2638;
w2678 <= w2676 and not w2677;
w2679 <= not pi1137 and not w154;
w2680 <= not pi0933 and w154;
w2681 <= pi0222 and not w2679;
w2682 <= not w2680 and w2681;
w2683 <= not w2678 and not w2682;
w2684 <= not pi0223 and not w2683;
w2685 <= not w2674 and not w2684;
w2686 <= not pi0299 and not w2685;
w2687 <= pi0299 and not w2652;
w2688 <= not w2686 and not w2687;
w2689 <= not w95 and w2688;
w2690 <= not w188 and w2688;
w2691 <= pi0299 and not w2662;
w2692 <= not w2686 and not w2691;
w2693 <= w188 and w2692;
w2694 <= not w2690 and not w2693;
w2695 <= w96 and not w2694;
w2696 <= not w96 and w2688;
w2697 <= pi0092 and not w2696;
w2698 <= not w2695 and w2697;
w2699 <= pi0075 and w2688;
w2700 <= pi0087 and w2694;
w2701 <= pi0038 and w2688;
w2702 <= pi0039 and not w2692;
w2703 <= not pi0299 and not w2674;
w2704 <= pi0878 and w1051;
w2705 <= not pi0224 and not w2704;
w2706 <= w2676 and not w2705;
w2707 <= not w2682 and not w2706;
w2708 <= w2703 and w2707;
w2709 <= pi0299 and not w2634;
w2710 <= pi0878 and w1062;
w2711 <= not pi0168 and not w2710;
w2712 <= pi0168 and w1071;
w2713 <= not w2711 and not w2712;
w2714 <= pi0878 and not w2713;
w2715 <= not w979 and w2711;
w2716 <= not w2714 and not w2715;
w2717 <= not pi0228 and not w2716;
w2718 <= not w1060 and w2641;
w2719 <= not pi0216 and not w2718;
w2720 <= not w2717 and w2719;
w2721 <= w2636 and not w2720;
w2722 <= not w2649 and not w2721;
w2723 <= not pi0215 and not w2722;
w2724 <= w2709 and not w2723;
w2725 <= not w1051 and w2676;
w2726 <= w2707 and not w2725;
w2727 <= not pi0223 and not w2726;
w2728 <= w2703 and not w2727;
w2729 <= not pi0039 and not w2728;
w2730 <= not w2708 and w2729;
w2731 <= not w2724 and w2730;
w2732 <= not pi0038 and not w2702;
w2733 <= not w2731 and w2732;
w2734 <= not pi0100 and not w2701;
w2735 <= not w2733 and w2734;
w2736 <= not w93 and w2688;
w2737 <= not pi0878 and w957;
w2738 <= pi0168 and not w957;
w2739 <= not pi0228 and not w2737;
w2740 <= not w2738 and w2739;
w2741 <= w2642 and not w2740;
w2742 <= w2636 and not w2741;
w2743 <= not w2649 and not w2742;
w2744 <= not pi0215 and not w2743;
w2745 <= not w2634 and not w2744;
w2746 <= pi0299 and not w2745;
w2747 <= w93 and not w2686;
w2748 <= not w2746 and w2747;
w2749 <= pi0100 and not w2736;
w2750 <= not w2748 and w2749;
w2751 <= not w2735 and not w2750;
w2752 <= not pi0087 and not w2751;
w2753 <= not pi0075 and not w2700;
w2754 <= not w2752 and w2753;
w2755 <= not pi0092 and not w2699;
w2756 <= not w2754 and w2755;
w2757 <= w95 and not w2698;
w2758 <= not w2756 and w2757;
w2759 <= not pi0055 and not w2689;
w2760 <= not w2758 and w2759;
w2761 <= not pi0056 and not w2673;
w2762 <= not w2760 and w2761;
w2763 <= not pi0062 and not w2669;
w2764 <= not w2762 and w2763;
w2765 <= not pi0240 and w891;
w2766 <= not w2665 and w2765;
w2767 <= not w2764 and w2766;
w2768 <= not w1010 and w2642;
w2769 <= not w2657 and w2768;
w2770 <= w2636 and not w2769;
w2771 <= not w2649 and not w2770;
w2772 <= not pi0215 and not w2771;
w2773 <= not w2634 and not w2772;
w2774 <= w894 and w2773;
w2775 <= w1119 and not w2635;
w2776 <= w2652 and not w2775;
w2777 <= not w894 and w2776;
w2778 <= pi0062 and not w2777;
w2779 <= not w2774 and w2778;
w2780 <= not w100 and not w2776;
w2781 <= w100 and not w2773;
w2782 <= pi0056 and not w2780;
w2783 <= not w2781 and w2782;
w2784 <= w135 and w2773;
w2785 <= not w135 and w2776;
w2786 <= pi0055 and not w2785;
w2787 <= not w2784 and w2786;
w2788 <= not w1035 and not w2686;
w2789 <= pi0299 and not w2776;
w2790 <= w2788 and not w2789;
w2791 <= not w95 and w2790;
w2792 <= not w188 and w2790;
w2793 <= pi0299 and not w2773;
w2794 <= w2788 and not w2793;
w2795 <= w188 and w2794;
w2796 <= not w2792 and not w2795;
w2797 <= w96 and not w2796;
w2798 <= not w96 and w2790;
w2799 <= pi0092 and not w2798;
w2800 <= not w2797 and w2799;
w2801 <= pi0075 and w2790;
w2802 <= pi0087 and w2796;
w2803 <= pi0038 and w2790;
w2804 <= pi0039 and not w2794;
w2805 <= not pi0878 and w1071;
w2806 <= not pi0168 and not w2805;
w2807 <= not pi0878 and not w1062;
w2808 <= pi0878 and not w979;
w2809 <= pi0168 and not w2807;
w2810 <= not w2808 and w2809;
w2811 <= not w2806 and not w2810;
w2812 <= not pi0228 and not w2811;
w2813 <= not w1356 and w2642;
w2814 <= not w2812 and w2813;
w2815 <= w2636 and not w2814;
w2816 <= not w2649 and not w2815;
w2817 <= not pi0215 and not w2816;
w2818 <= w2709 and not w2817;
w2819 <= w2729 and not w2818;
w2820 <= not pi0038 and not w2804;
w2821 <= not w2819 and w2820;
w2822 <= not pi0100 and not w2803;
w2823 <= not w2821 and w2822;
w2824 <= not w93 and w2790;
w2825 <= not w2740 and w2768;
w2826 <= w2636 and not w2825;
w2827 <= not w2649 and not w2826;
w2828 <= not pi0215 and not w2827;
w2829 <= not w2634 and not w2828;
w2830 <= pi0299 and not w2829;
w2831 <= w93 and w2788;
w2832 <= not w2830 and w2831;
w2833 <= pi0100 and not w2824;
w2834 <= not w2832 and w2833;
w2835 <= not w2823 and not w2834;
w2836 <= not pi0087 and not w2835;
w2837 <= not pi0075 and not w2802;
w2838 <= not w2836 and w2837;
w2839 <= not pi0092 and not w2801;
w2840 <= not w2838 and w2839;
w2841 <= w95 and not w2800;
w2842 <= not w2840 and w2841;
w2843 <= not pi0055 and not w2791;
w2844 <= not w2842 and w2843;
w2845 <= not pi0056 and not w2787;
w2846 <= not w2844 and w2845;
w2847 <= not pi0062 and not w2783;
w2848 <= not w2846 and w2847;
w2849 <= pi0240 and w891;
w2850 <= not w2779 and w2849;
w2851 <= not w2848 and w2850;
w2852 <= pi0240 and w2775;
w2853 <= not w891 and not w2852;
w2854 <= w2652 and w2853;
w2855 <= not w2851 and not w2854;
w2856 <= not w2767 and w2855;
w2857 <= pi0215 and pi1136;
w2858 <= pi0216 and pi0266;
w2859 <= pi0875 and not w5;
w2860 <= pi0105 and not w2859;
w2861 <= not pi0105 and not pi0166;
w2862 <= not w2860 and not w2861;
w2863 <= pi0228 and w2862;
w2864 <= pi0166 and not pi0228;
w2865 <= not w2863 and not w2864;
w2866 <= not pi0216 and not w2865;
w2867 <= not w2858 and not w2866;
w2868 <= not pi0221 and not w2867;
w2869 <= not pi1136 and not w15;
w2870 <= not pi0928 and w15;
w2871 <= pi0221 and not w2869;
w2872 <= not w2870 and w2871;
w2873 <= not w2868 and not w2872;
w2874 <= not pi0215 and not w2873;
w2875 <= not w2857 and not w2874;
w2876 <= not w891 and w2875;
w2877 <= not w894 and w2875;
w2878 <= not pi0166 and not w84;
w2879 <= not pi0875 and w84;
w2880 <= not pi0228 and not w2878;
w2881 <= not w2879 and w2880;
w2882 <= not w2863 and not w2881;
w2883 <= not pi0216 and not w2882;
w2884 <= not w2858 and not w2883;
w2885 <= not pi0221 and not w2884;
w2886 <= not w2872 and not w2885;
w2887 <= not pi0215 and not w2886;
w2888 <= not w2857 and not w2887;
w2889 <= w894 and w2888;
w2890 <= pi0062 and not w2877;
w2891 <= not w2889 and w2890;
w2892 <= not w100 and not w2875;
w2893 <= w100 and not w2888;
w2894 <= pi0056 and not w2892;
w2895 <= not w2893 and w2894;
w2896 <= not w135 and w2875;
w2897 <= w135 and w2888;
w2898 <= pi0055 and not w2896;
w2899 <= not w2897 and w2898;
w2900 <= pi0223 and pi1136;
w2901 <= pi0224 and not pi0266;
w2902 <= not pi0224 and not pi0875;
w2903 <= not w5 and w2902;
w2904 <= not pi0222 and not w2901;
w2905 <= not w2903 and w2904;
w2906 <= not pi1136 and not w154;
w2907 <= not pi0928 and w154;
w2908 <= pi0222 and not w2906;
w2909 <= not w2907 and w2908;
w2910 <= not w2905 and not w2909;
w2911 <= not pi0223 and not w2910;
w2912 <= not w2900 and not w2911;
w2913 <= not pi0299 and not w2912;
w2914 <= w167 and not w2859;
w2915 <= w2913 and not w2914;
w2916 <= pi0299 and not w2875;
w2917 <= not w2915 and not w2916;
w2918 <= not w95 and w2917;
w2919 <= not w188 and w2917;
w2920 <= pi0299 and not w2888;
w2921 <= not w2915 and not w2920;
w2922 <= w188 and w2921;
w2923 <= not w2919 and not w2922;
w2924 <= w96 and not w2923;
w2925 <= not w96 and w2917;
w2926 <= pi0092 and not w2925;
w2927 <= not w2924 and w2926;
w2928 <= pi0075 and w2917;
w2929 <= pi0087 and w2923;
w2930 <= pi0038 and w2917;
w2931 <= pi0039 and not w2921;
w2932 <= w166 and not w1051;
w2933 <= w2905 and not w2932;
w2934 <= not pi0299 and not w2900;
w2935 <= not w2909 and w2934;
w2936 <= not w2933 and w2935;
w2937 <= w1061 and not w2862;
w2938 <= not pi0216 and not w2937;
w2939 <= pi0166 and w1062;
w2940 <= not pi0166 and not w1071;
w2941 <= pi0875 and not w2939;
w2942 <= not w2940 and w2941;
w2943 <= pi0166 and not pi0875;
w2944 <= not w979 and w2943;
w2945 <= not w2942 and not w2944;
w2946 <= not pi0228 and not w2945;
w2947 <= not w1061 and not w2946;
w2948 <= w2938 and not w2947;
w2949 <= not w2858 and not w2948;
w2950 <= not pi0221 and not w2949;
w2951 <= not w2872 and not w2950;
w2952 <= not pi0215 and not w2951;
w2953 <= pi0299 and not w2857;
w2954 <= not w2952 and w2953;
w2955 <= w2910 and not w2932;
w2956 <= not pi0223 and not w2955;
w2957 <= w2934 and not w2956;
w2958 <= not pi0039 and not w2957;
w2959 <= not w2936 and w2958;
w2960 <= not w2954 and w2959;
w2961 <= not pi0038 and not w2931;
w2962 <= not w2960 and w2961;
w2963 <= not pi0100 and not w2930;
w2964 <= not w2962 and w2963;
w2965 <= not w93 and w2917;
w2966 <= not pi0875 and w950;
w2967 <= pi0166 and not w2966;
w2968 <= not w201 and not w950;
w2969 <= w201 and not w948;
w2970 <= pi0875 and not w2969;
w2971 <= not w2968 and w2970;
w2972 <= not w2967 and not w2971;
w2973 <= not pi0228 and not w2972;
w2974 <= not w2863 and not w2973;
w2975 <= not pi0216 and not w2974;
w2976 <= not w2858 and not w2975;
w2977 <= not pi0221 and not w2976;
w2978 <= not w2872 and not w2977;
w2979 <= not pi0215 and not w2978;
w2980 <= not w2857 and not w2979;
w2981 <= pi0299 and not w2980;
w2982 <= w93 and not w2915;
w2983 <= not w2981 and w2982;
w2984 <= pi0100 and not w2965;
w2985 <= not w2983 and w2984;
w2986 <= not w2964 and not w2985;
w2987 <= not pi0087 and not w2986;
w2988 <= not pi0075 and not w2929;
w2989 <= not w2987 and w2988;
w2990 <= not pi0092 and not w2928;
w2991 <= not w2989 and w2990;
w2992 <= w95 and not w2927;
w2993 <= not w2991 and w2992;
w2994 <= not pi0055 and not w2918;
w2995 <= not w2993 and w2994;
w2996 <= not pi0056 and not w2899;
w2997 <= not w2995 and w2996;
w2998 <= not pi0062 and not w2895;
w2999 <= not w2997 and w2998;
w3000 <= w891 and not w2891;
w3001 <= not w2999 and w3000;
w3002 <= not pi0245 and not w2876;
w3003 <= not w3001 and w3002;
w3004 <= not w1013 and w2875;
w3005 <= not w891 and w3004;
w3006 <= not w1010 and not w2863;
w3007 <= not w2881 and w3006;
w3008 <= not pi0216 and not w3007;
w3009 <= not w2858 and not w3008;
w3010 <= not pi0221 and not w3009;
w3011 <= not w2872 and not w3010;
w3012 <= not pi0215 and not w3011;
w3013 <= not w2857 and not w3012;
w3014 <= w894 and w3013;
w3015 <= not w894 and w3004;
w3016 <= pi0062 and not w3015;
w3017 <= not w3014 and w3016;
w3018 <= not w100 and not w3004;
w3019 <= w100 and not w3013;
w3020 <= pi0056 and not w3018;
w3021 <= not w3019 and w3020;
w3022 <= w135 and w3013;
w3023 <= not w135 and w3004;
w3024 <= pi0055 and not w3023;
w3025 <= not w3022 and w3024;
w3026 <= pi0299 and not w3004;
w3027 <= not w2913 and not w3026;
w3028 <= not w95 and w3027;
w3029 <= not w188 and w3027;
w3030 <= pi0299 and not w3013;
w3031 <= not w2913 and not w3030;
w3032 <= w188 and w3031;
w3033 <= not w3029 and not w3032;
w3034 <= w96 and not w3033;
w3035 <= not w96 and w3027;
w3036 <= pi0092 and not w3035;
w3037 <= not w3034 and w3036;
w3038 <= pi0075 and w3027;
w3039 <= pi0087 and w3033;
w3040 <= pi0038 and w3027;
w3041 <= pi0039 and not w3031;
w3042 <= not pi0166 and not w1062;
w3043 <= pi0166 and w1071;
w3044 <= not pi0875 and not w3042;
w3045 <= not w3043 and w3044;
w3046 <= not pi0166 and not w979;
w3047 <= pi0875 and not w3046;
w3048 <= not pi0228 and not w3045;
w3049 <= not w3047 and w3048;
w3050 <= w2938 and not w3049;
w3051 <= not w2858 and not w3050;
w3052 <= not pi0221 and not w3051;
w3053 <= not w2872 and not w3052;
w3054 <= not pi0215 and not w3053;
w3055 <= w2953 and not w3054;
w3056 <= w2958 and not w3055;
w3057 <= not pi0038 and not w3041;
w3058 <= not w3056 and w3057;
w3059 <= not pi0100 and not w3040;
w3060 <= not w3058 and w3059;
w3061 <= not w93 and w3027;
w3062 <= not w2973 and w3006;
w3063 <= not pi0216 and not w3062;
w3064 <= not w2858 and not w3063;
w3065 <= not pi0221 and not w3064;
w3066 <= not w2872 and not w3065;
w3067 <= not pi0215 and not w3066;
w3068 <= not w2857 and not w3067;
w3069 <= pi0299 and not w3068;
w3070 <= w93 and not w2913;
w3071 <= not w3069 and w3070;
w3072 <= pi0100 and not w3061;
w3073 <= not w3071 and w3072;
w3074 <= not w3060 and not w3073;
w3075 <= not pi0087 and not w3074;
w3076 <= not pi0075 and not w3039;
w3077 <= not w3075 and w3076;
w3078 <= not pi0092 and not w3038;
w3079 <= not w3077 and w3078;
w3080 <= w95 and not w3037;
w3081 <= not w3079 and w3080;
w3082 <= not pi0055 and not w3028;
w3083 <= not w3081 and w3082;
w3084 <= not pi0056 and not w3025;
w3085 <= not w3083 and w3084;
w3086 <= not pi0062 and not w3021;
w3087 <= not w3085 and w3086;
w3088 <= w891 and not w3017;
w3089 <= not w3087 and w3088;
w3090 <= pi0245 and not w3005;
w3091 <= not w3089 and w3090;
w3092 <= not w3003 and not w3091;
w3093 <= pi0215 and pi1135;
w3094 <= pi0216 and pi0279;
w3095 <= pi0879 and not w5;
w3096 <= pi0105 and not w3095;
w3097 <= not pi0105 and not pi0161;
w3098 <= not w3096 and not w3097;
w3099 <= pi0228 and w3098;
w3100 <= pi0161 and not pi0228;
w3101 <= not w3099 and not w3100;
w3102 <= not pi0216 and not w3101;
w3103 <= not w3094 and not w3102;
w3104 <= not pi0221 and not w3103;
w3105 <= not pi1135 and not w15;
w3106 <= not pi0938 and w15;
w3107 <= pi0221 and not w3105;
w3108 <= not w3106 and w3107;
w3109 <= not w3104 and not w3108;
w3110 <= not pi0215 and not w3109;
w3111 <= not w3093 and not w3110;
w3112 <= not w891 and w3111;
w3113 <= not w894 and w3111;
w3114 <= not pi0879 and w84;
w3115 <= not w898 and not w3100;
w3116 <= not w3114 and not w3115;
w3117 <= not w3099 and not w3116;
w3118 <= not pi0216 and not w3117;
w3119 <= not w3094 and not w3118;
w3120 <= not pi0221 and not w3119;
w3121 <= not w3108 and not w3120;
w3122 <= not pi0215 and not w3121;
w3123 <= not w3093 and not w3122;
w3124 <= w894 and w3123;
w3125 <= pi0062 and not w3113;
w3126 <= not w3124 and w3125;
w3127 <= not w100 and not w3111;
w3128 <= w100 and not w3123;
w3129 <= pi0056 and not w3127;
w3130 <= not w3128 and w3129;
w3131 <= not w135 and w3111;
w3132 <= w135 and w3123;
w3133 <= pi0055 and not w3131;
w3134 <= not w3132 and w3133;
w3135 <= pi0223 and pi1135;
w3136 <= not pi1135 and not w154;
w3137 <= not pi0938 and w154;
w3138 <= pi0222 and not w3136;
w3139 <= not w3137 and w3138;
w3140 <= pi0224 and not pi0279;
w3141 <= not pi0224 and not pi0879;
w3142 <= not w5 and w3141;
w3143 <= not pi0222 and not w3140;
w3144 <= not w3142 and w3143;
w3145 <= not w3139 and not w3144;
w3146 <= not pi0223 and not w3145;
w3147 <= not w3135 and not w3146;
w3148 <= not pi0299 and not w3147;
w3149 <= w167 and not w3095;
w3150 <= w3148 and not w3149;
w3151 <= pi0299 and not w3111;
w3152 <= not w3150 and not w3151;
w3153 <= not w95 and w3152;
w3154 <= not w188 and w3152;
w3155 <= pi0299 and not w3123;
w3156 <= not w3150 and not w3155;
w3157 <= w188 and w3156;
w3158 <= not w3154 and not w3157;
w3159 <= w96 and not w3158;
w3160 <= not w96 and w3152;
w3161 <= pi0092 and not w3160;
w3162 <= not w3159 and w3161;
w3163 <= pi0075 and w3152;
w3164 <= pi0087 and w3158;
w3165 <= pi0038 and w3152;
w3166 <= pi0039 and not w3156;
w3167 <= not pi0299 and not w3135;
w3168 <= w2932 and not w3139;
w3169 <= w3146 and not w3168;
w3170 <= w3167 and not w3169;
w3171 <= w1061 and not w3098;
w3172 <= not pi0216 and not w3171;
w3173 <= pi0161 and w1062;
w3174 <= not pi0161 and not w1071;
w3175 <= pi0879 and not w3173;
w3176 <= not w3174 and w3175;
w3177 <= pi0161 and not pi0879;
w3178 <= not w979 and w3177;
w3179 <= not w3176 and not w3178;
w3180 <= not pi0228 and not w3179;
w3181 <= not w1061 and not w3180;
w3182 <= w3172 and not w3181;
w3183 <= not w3094 and not w3182;
w3184 <= not pi0221 and not w3183;
w3185 <= not w3108 and not w3184;
w3186 <= not pi0215 and not w3185;
w3187 <= pi0299 and not w3093;
w3188 <= not w3186 and w3187;
w3189 <= not pi0039 and not w3170;
w3190 <= not w3188 and w3189;
w3191 <= not pi0038 and not w3166;
w3192 <= not w3190 and w3191;
w3193 <= not pi0100 and not w3165;
w3194 <= not w3192 and w3193;
w3195 <= not w93 and w3152;
w3196 <= not pi0879 and w950;
w3197 <= pi0161 and not w3196;
w3198 <= not pi0152 and not pi0166;
w3199 <= not w948 and w3198;
w3200 <= not w950 and not w3198;
w3201 <= pi0879 and not w3199;
w3202 <= not w3200 and w3201;
w3203 <= not w3197 and not w3202;
w3204 <= not pi0228 and not w3203;
w3205 <= not w3099 and not w3204;
w3206 <= not pi0216 and not w3205;
w3207 <= not w3094 and not w3206;
w3208 <= not pi0221 and not w3207;
w3209 <= not w3108 and not w3208;
w3210 <= not pi0215 and not w3209;
w3211 <= not w3093 and not w3210;
w3212 <= pi0299 and not w3211;
w3213 <= w93 and not w3150;
w3214 <= not w3212 and w3213;
w3215 <= pi0100 and not w3195;
w3216 <= not w3214 and w3215;
w3217 <= not w3194 and not w3216;
w3218 <= not pi0087 and not w3217;
w3219 <= not pi0075 and not w3164;
w3220 <= not w3218 and w3219;
w3221 <= not pi0092 and not w3163;
w3222 <= not w3220 and w3221;
w3223 <= w95 and not w3162;
w3224 <= not w3222 and w3223;
w3225 <= not pi0055 and not w3153;
w3226 <= not w3224 and w3225;
w3227 <= not pi0056 and not w3134;
w3228 <= not w3226 and w3227;
w3229 <= not pi0062 and not w3130;
w3230 <= not w3228 and w3229;
w3231 <= w891 and not w3126;
w3232 <= not w3230 and w3231;
w3233 <= not pi0244 and not w3112;
w3234 <= not w3232 and w3233;
w3235 <= not w1013 and w3111;
w3236 <= not w891 and w3235;
w3237 <= not w1010 and not w3099;
w3238 <= not w3116 and w3237;
w3239 <= not pi0216 and not w3238;
w3240 <= not w3094 and not w3239;
w3241 <= not pi0221 and not w3240;
w3242 <= not w3108 and not w3241;
w3243 <= not pi0215 and not w3242;
w3244 <= not w3093 and not w3243;
w3245 <= w894 and w3244;
w3246 <= not w894 and w3235;
w3247 <= pi0062 and not w3246;
w3248 <= not w3245 and w3247;
w3249 <= not w100 and not w3235;
w3250 <= w100 and not w3244;
w3251 <= pi0056 and not w3249;
w3252 <= not w3250 and w3251;
w3253 <= w135 and w3244;
w3254 <= not w135 and w3235;
w3255 <= pi0055 and not w3254;
w3256 <= not w3253 and w3255;
w3257 <= pi0299 and not w3235;
w3258 <= not w3148 and not w3257;
w3259 <= not w95 and w3258;
w3260 <= not w188 and w3258;
w3261 <= pi0299 and not w3244;
w3262 <= not w3148 and not w3261;
w3263 <= w188 and w3262;
w3264 <= not w3260 and not w3263;
w3265 <= w96 and not w3264;
w3266 <= not w96 and w3258;
w3267 <= pi0092 and not w3266;
w3268 <= not w3265 and w3267;
w3269 <= pi0075 and w3258;
w3270 <= pi0087 and w3264;
w3271 <= pi0038 and w3258;
w3272 <= pi0039 and not w3262;
w3273 <= not w2932 and w3145;
w3274 <= not pi0223 and not w3273;
w3275 <= w3167 and not w3274;
w3276 <= not pi0161 and not w1062;
w3277 <= pi0161 and w1071;
w3278 <= not pi0879 and not w3276;
w3279 <= not w3277 and w3278;
w3280 <= not pi0161 and not w979;
w3281 <= pi0879 and not w3280;
w3282 <= not pi0228 and not w3279;
w3283 <= not w3281 and w3282;
w3284 <= w3172 and not w3283;
w3285 <= not w3094 and not w3284;
w3286 <= not pi0221 and not w3285;
w3287 <= not w3108 and not w3286;
w3288 <= not pi0215 and not w3287;
w3289 <= w3187 and not w3288;
w3290 <= not pi0039 and not w3275;
w3291 <= not w3289 and w3290;
w3292 <= not pi0038 and not w3272;
w3293 <= not w3291 and w3292;
w3294 <= not pi0100 and not w3271;
w3295 <= not w3293 and w3294;
w3296 <= not w93 and w3258;
w3297 <= not w3204 and w3237;
w3298 <= not pi0216 and not w3297;
w3299 <= not w3094 and not w3298;
w3300 <= not pi0221 and not w3299;
w3301 <= not w3108 and not w3300;
w3302 <= not pi0215 and not w3301;
w3303 <= not w3093 and not w3302;
w3304 <= pi0299 and not w3303;
w3305 <= w93 and not w3148;
w3306 <= not w3304 and w3305;
w3307 <= pi0100 and not w3296;
w3308 <= not w3306 and w3307;
w3309 <= not w3295 and not w3308;
w3310 <= not pi0087 and not w3309;
w3311 <= not pi0075 and not w3270;
w3312 <= not w3310 and w3311;
w3313 <= not pi0092 and not w3269;
w3314 <= not w3312 and w3313;
w3315 <= w95 and not w3268;
w3316 <= not w3314 and w3315;
w3317 <= not pi0055 and not w3259;
w3318 <= not w3316 and w3317;
w3319 <= not pi0056 and not w3256;
w3320 <= not w3318 and w3319;
w3321 <= not pi0062 and not w3252;
w3322 <= not w3320 and w3321;
w3323 <= w891 and not w3248;
w3324 <= not w3322 and w3323;
w3325 <= pi0244 and not w3236;
w3326 <= not w3324 and w3325;
w3327 <= not w3234 and not w3326;
w3328 <= pi0216 and pi0278;
w3329 <= not pi0221 and not w3328;
w3330 <= not pi0105 and pi0152;
w3331 <= pi0846 and not w5;
w3332 <= pi0105 and w3331;
w3333 <= not w3330 and not w3332;
w3334 <= pi0228 and not w3333;
w3335 <= pi0152 and not pi0228;
w3336 <= not w3334 and not w3335;
w3337 <= not pi0216 and not w3336;
w3338 <= w3329 and not w3337;
w3339 <= pi0833 and not pi0930;
w3340 <= not pi0216 and pi0221;
w3341 <= w3339 and w3340;
w3342 <= pi0221 and not w15;
w3343 <= not pi0215 and not w3342;
w3344 <= not w3341 and w3343;
w3345 <= not w3338 and w3344;
w3346 <= not w1013 and not w3345;
w3347 <= not w891 and not w3346;
w3348 <= not w894 and not w3346;
w3349 <= not w1010 and not w3334;
w3350 <= not pi0152 and not w84;
w3351 <= not pi0846 and w84;
w3352 <= not pi0228 and not w3350;
w3353 <= not w3351 and w3352;
w3354 <= w3349 and not w3353;
w3355 <= not pi0216 and not w3354;
w3356 <= w3329 and not w3355;
w3357 <= w3344 and not w3356;
w3358 <= w894 and w3357;
w3359 <= pi0062 and not w3348;
w3360 <= not w3358 and w3359;
w3361 <= w100 and not w3357;
w3362 <= not w100 and w3346;
w3363 <= pi0056 and not w3362;
w3364 <= not w3361 and w3363;
w3365 <= not w135 and not w3346;
w3366 <= w135 and w3357;
w3367 <= pi0055 and not w3365;
w3368 <= not w3366 and w3367;
w3369 <= pi0224 and pi0278;
w3370 <= not pi0222 and not w3369;
w3371 <= not pi0224 and w3331;
w3372 <= w3370 and not w3371;
w3373 <= pi0222 and not pi0224;
w3374 <= w3339 and w3373;
w3375 <= w156 and not w3374;
w3376 <= not w3372 and w3375;
w3377 <= not pi0299 and not w3376;
w3378 <= not w1318 and w3377;
w3379 <= pi0299 and w3346;
w3380 <= not w3378 and not w3379;
w3381 <= not w95 and w3380;
w3382 <= not w188 and w3380;
w3383 <= pi0299 and not w3357;
w3384 <= not w3378 and not w3383;
w3385 <= w188 and w3384;
w3386 <= not w3382 and not w3385;
w3387 <= w96 and not w3386;
w3388 <= not w96 and w3380;
w3389 <= pi0092 and not w3388;
w3390 <= not w3387 and w3389;
w3391 <= pi0075 and w3380;
w3392 <= pi0087 and w3386;
w3393 <= pi0038 and w3380;
w3394 <= pi0039 and not w3384;
w3395 <= not pi0846 and w1051;
w3396 <= not pi0224 and not w3395;
w3397 <= w3370 and not w3396;
w3398 <= not w3374 and not w3397;
w3399 <= not w155 and w1033;
w3400 <= w3398 and w3399;
w3401 <= pi0228 and not w3330;
w3402 <= pi0105 and not w3395;
w3403 <= w3401 and not w3402;
w3404 <= not pi0216 and not w3403;
w3405 <= not pi0152 and w1062;
w3406 <= pi0152 and not w1071;
w3407 <= not pi0846 and not w3405;
w3408 <= not w3406 and w3407;
w3409 <= not pi0152 and pi0846;
w3410 <= not w979 and w3409;
w3411 <= not w3408 and not w3410;
w3412 <= not pi0228 and not w3411;
w3413 <= w3404 and not w3412;
w3414 <= w3329 and not w3413;
w3415 <= not w3341 and not w3414;
w3416 <= not pi0215 and pi0299;
w3417 <= not w3342 and w3416;
w3418 <= w3415 and w3417;
w3419 <= not pi0039 and not w3400;
w3420 <= not w3418 and w3419;
w3421 <= not pi0038 and not w3394;
w3422 <= not w3420 and w3421;
w3423 <= not pi0100 and not w3393;
w3424 <= not w3422 and w3423;
w3425 <= not w93 and w3380;
w3426 <= pi0846 and not w956;
w3427 <= not w951 and not w3426;
w3428 <= not pi0228 and not w3427;
w3429 <= w3349 and not w3428;
w3430 <= not pi0216 and not w3429;
w3431 <= w3329 and not w3430;
w3432 <= w3344 and not w3431;
w3433 <= pi0299 and not w3432;
w3434 <= w93 and not w3378;
w3435 <= not w3433 and w3434;
w3436 <= pi0100 and not w3425;
w3437 <= not w3435 and w3436;
w3438 <= not w3424 and not w3437;
w3439 <= not pi0087 and not w3438;
w3440 <= not pi0075 and not w3392;
w3441 <= not w3439 and w3440;
w3442 <= not pi0092 and not w3391;
w3443 <= not w3441 and w3442;
w3444 <= w95 and not w3390;
w3445 <= not w3443 and w3444;
w3446 <= not pi0055 and not w3381;
w3447 <= not w3445 and w3446;
w3448 <= not pi0056 and not w3368;
w3449 <= not w3447 and w3448;
w3450 <= not pi0062 and not w3364;
w3451 <= not w3449 and w3450;
w3452 <= w891 and not w3360;
w3453 <= not w3451 and w3452;
w3454 <= pi0242 and not w3347;
w3455 <= not w3453 and w3454;
w3456 <= not w891 and w3345;
w3457 <= not w894 and w3345;
w3458 <= not w3334 and not w3353;
w3459 <= not pi0216 and not w3458;
w3460 <= w3329 and not w3459;
w3461 <= w3344 and not w3460;
w3462 <= w894 and w3461;
w3463 <= pi0062 and not w3457;
w3464 <= not w3462 and w3463;
w3465 <= not w100 and not w3345;
w3466 <= w100 and not w3461;
w3467 <= pi0056 and not w3465;
w3468 <= not w3466 and w3467;
w3469 <= not w135 and w3345;
w3470 <= w135 and w3461;
w3471 <= pi0055 and not w3469;
w3472 <= not w3470 and w3471;
w3473 <= pi0299 and not w3345;
w3474 <= not w3377 and not w3473;
w3475 <= not w95 and w3474;
w3476 <= not w188 and w3474;
w3477 <= pi0299 and not w3461;
w3478 <= not w3377 and not w3477;
w3479 <= w188 and w3478;
w3480 <= not w3476 and not w3479;
w3481 <= w96 and not w3480;
w3482 <= not w96 and w3474;
w3483 <= pi0092 and not w3482;
w3484 <= not w3481 and w3483;
w3485 <= pi0075 and w3474;
w3486 <= pi0087 and w3480;
w3487 <= pi0038 and w3474;
w3488 <= pi0039 and not w3478;
w3489 <= not w1050 and w3371;
w3490 <= w3370 and not w3489;
w3491 <= not w3374 and w3399;
w3492 <= not w3490 and w3491;
w3493 <= not w1051 and w3401;
w3494 <= pi0152 and not pi0846;
w3495 <= not w979 and w3494;
w3496 <= pi0152 and w1062;
w3497 <= not pi0152 and not w1071;
w3498 <= pi0846 and not w3496;
w3499 <= not w3497 and w3498;
w3500 <= not pi0228 and not w3495;
w3501 <= not w3499 and w3500;
w3502 <= w3404 and not w3493;
w3503 <= not w3501 and w3502;
w3504 <= w3329 and not w3503;
w3505 <= not w3341 and not w3504;
w3506 <= w3417 and w3505;
w3507 <= not pi0039 and not w3492;
w3508 <= not w3506 and w3507;
w3509 <= not pi0038 and not w3488;
w3510 <= not w3508 and w3509;
w3511 <= not pi0100 and not w3487;
w3512 <= not w3510 and w3511;
w3513 <= not w93 and w3474;
w3514 <= not w3334 and not w3428;
w3515 <= not pi0216 and not w3514;
w3516 <= w3329 and not w3515;
w3517 <= w3344 and not w3516;
w3518 <= pi0299 and not w3517;
w3519 <= w93 and not w3377;
w3520 <= not w3518 and w3519;
w3521 <= pi0100 and not w3513;
w3522 <= not w3520 and w3521;
w3523 <= not w3512 and not w3522;
w3524 <= not pi0087 and not w3523;
w3525 <= not pi0075 and not w3486;
w3526 <= not w3524 and w3525;
w3527 <= not pi0092 and not w3485;
w3528 <= not w3526 and w3527;
w3529 <= w95 and not w3484;
w3530 <= not w3528 and w3529;
w3531 <= not pi0055 and not w3475;
w3532 <= not w3530 and w3531;
w3533 <= not pi0056 and not w3472;
w3534 <= not w3532 and w3533;
w3535 <= not pi0062 and not w3468;
w3536 <= not w3534 and w3535;
w3537 <= w891 and not w3464;
w3538 <= not w3536 and w3537;
w3539 <= not pi0242 and not w3456;
w3540 <= not w3538 and w3539;
w3541 <= not w3455 and not w3540;
w3542 <= not pi1134 and not w3541;
w3543 <= not w3338 and not w3341;
w3544 <= not pi0215 and not w3543;
w3545 <= not w891 and w3544;
w3546 <= not w894 and w3544;
w3547 <= not w3341 and not w3460;
w3548 <= not pi0215 and not w3547;
w3549 <= w894 and w3548;
w3550 <= pi0062 and not w3546;
w3551 <= not w3549 and w3550;
w3552 <= not w100 and not w3544;
w3553 <= w100 and not w3548;
w3554 <= pi0056 and not w3552;
w3555 <= not w3553 and w3554;
w3556 <= not w135 and w3544;
w3557 <= w135 and w3548;
w3558 <= pi0055 and not w3556;
w3559 <= not w3557 and w3558;
w3560 <= w156 and w3378;
w3561 <= not pi0299 and not w3560;
w3562 <= not pi0223 and w3372;
w3563 <= w3561 and not w3562;
w3564 <= pi0299 and not w3544;
w3565 <= not w3563 and not w3564;
w3566 <= not w95 and w3565;
w3567 <= not w188 and w3565;
w3568 <= pi0299 and not w3548;
w3569 <= not w3563 and not w3568;
w3570 <= w188 and w3569;
w3571 <= not w3567 and not w3570;
w3572 <= w96 and not w3571;
w3573 <= not w96 and w3565;
w3574 <= pi0092 and not w3573;
w3575 <= not w3572 and w3574;
w3576 <= pi0075 and w3565;
w3577 <= pi0087 and w3571;
w3578 <= pi0038 and w3565;
w3579 <= pi0039 and not w3569;
w3580 <= w1033 and w3490;
w3581 <= w3416 and not w3505;
w3582 <= w1033 and not w3398;
w3583 <= not pi0039 and not w3582;
w3584 <= not w3580 and w3583;
w3585 <= not w3581 and w3584;
w3586 <= not pi0038 and not w3579;
w3587 <= not w3585 and w3586;
w3588 <= not pi0100 and not w3578;
w3589 <= not w3587 and w3588;
w3590 <= not w93 and w3565;
w3591 <= not w3341 and not w3516;
w3592 <= not pi0215 and not w3591;
w3593 <= pi0299 and not w3592;
w3594 <= w93 and not w3563;
w3595 <= not w3593 and w3594;
w3596 <= pi0100 and not w3590;
w3597 <= not w3595 and w3596;
w3598 <= not w3589 and not w3597;
w3599 <= not pi0087 and not w3598;
w3600 <= not pi0075 and not w3577;
w3601 <= not w3599 and w3600;
w3602 <= not pi0092 and not w3576;
w3603 <= not w3601 and w3602;
w3604 <= w95 and not w3575;
w3605 <= not w3603 and w3604;
w3606 <= not pi0055 and not w3566;
w3607 <= not w3605 and w3606;
w3608 <= not pi0056 and not w3559;
w3609 <= not w3607 and w3608;
w3610 <= not pi0062 and not w3555;
w3611 <= not w3609 and w3610;
w3612 <= w891 and not w3551;
w3613 <= not w3611 and w3612;
w3614 <= not pi0242 and not w3545;
w3615 <= not w3613 and w3614;
w3616 <= not w1013 and w3544;
w3617 <= not w891 and w3616;
w3618 <= not w3341 and not w3356;
w3619 <= not pi0215 and not w3618;
w3620 <= w894 and w3619;
w3621 <= not w894 and w3616;
w3622 <= pi0062 and not w3621;
w3623 <= not w3620 and w3622;
w3624 <= not w100 and not w3616;
w3625 <= w100 and not w3619;
w3626 <= pi0056 and not w3624;
w3627 <= not w3625 and w3626;
w3628 <= w135 and w3619;
w3629 <= not w135 and w3616;
w3630 <= pi0055 and not w3629;
w3631 <= not w3628 and w3630;
w3632 <= pi0299 and not w3616;
w3633 <= not w3561 and not w3632;
w3634 <= not w95 and w3633;
w3635 <= not w188 and w3633;
w3636 <= pi0299 and not w3619;
w3637 <= not w3561 and not w3636;
w3638 <= w188 and w3637;
w3639 <= not w3635 and not w3638;
w3640 <= w96 and not w3639;
w3641 <= not w96 and w3633;
w3642 <= pi0092 and not w3641;
w3643 <= not w3640 and w3642;
w3644 <= pi0075 and w3633;
w3645 <= pi0087 and w3639;
w3646 <= pi0038 and w3633;
w3647 <= pi0039 and not w3637;
w3648 <= not w3415 and w3416;
w3649 <= w3583 and not w3648;
w3650 <= not pi0038 and not w3647;
w3651 <= not w3649 and w3650;
w3652 <= not pi0100 and not w3646;
w3653 <= not w3651 and w3652;
w3654 <= not w93 and w3633;
w3655 <= not w3341 and not w3431;
w3656 <= not pi0215 and not w3655;
w3657 <= pi0299 and not w3656;
w3658 <= w93 and not w3561;
w3659 <= not w3657 and w3658;
w3660 <= pi0100 and not w3654;
w3661 <= not w3659 and w3660;
w3662 <= not w3653 and not w3661;
w3663 <= not pi0087 and not w3662;
w3664 <= not pi0075 and not w3645;
w3665 <= not w3663 and w3664;
w3666 <= not pi0092 and not w3644;
w3667 <= not w3665 and w3666;
w3668 <= w95 and not w3643;
w3669 <= not w3667 and w3668;
w3670 <= not pi0055 and not w3634;
w3671 <= not w3669 and w3670;
w3672 <= not pi0056 and not w3631;
w3673 <= not w3671 and w3672;
w3674 <= not pi0062 and not w3627;
w3675 <= not w3673 and w3674;
w3676 <= w891 and not w3623;
w3677 <= not w3675 and w3676;
w3678 <= pi0242 and not w3617;
w3679 <= not w3677 and w3678;
w3680 <= pi1134 and not w3615;
w3681 <= not w3679 and w3680;
w3682 <= not w3542 and not w3681;
w3683 <= pi0057 and pi0059;
w3684 <= w84 and w101;
w3685 <= not w891 and not w3684;
w3686 <= not w3683 and not w3685;
w3687 <= pi0057 and not w3686;
w3688 <= w75 and w188;
w3689 <= w99 and w3688;
w3690 <= pi0056 and not w3689;
w3691 <= not pi0054 and w97;
w3692 <= w3688 and w3691;
w3693 <= pi0074 and not w3692;
w3694 <= not pi0055 and not w3693;
w3695 <= pi0087 and not w3688;
w3696 <= not pi0075 and not w3695;
w3697 <= not pi0054 and not pi0092;
w3698 <= not pi0039 and w75;
w3699 <= pi0038 and not w3698;
w3700 <= not pi0100 and not w3699;
w3701 <= pi0058 and w65;
w3702 <= not pi0090 and not w3701;
w3703 <= w283 and w332;
w3704 <= w437 and w3703;
w3705 <= w344 and not w3704;
w3706 <= not w339 and not w3705;
w3707 <= not pi0108 and not w3706;
w3708 <= w338 and not w3707;
w3709 <= not pi0110 and w452;
w3710 <= not w3708 and w3709;
w3711 <= not w322 and not w329;
w3712 <= not w3710 and w3711;
w3713 <= not pi0047 and not w3712;
w3714 <= w263 and not w325;
w3715 <= not w3713 and w3714;
w3716 <= w3702 and not w3715;
w3717 <= not w459 and not w3716;
w3718 <= not pi0093 and not w3717;
w3719 <= not pi0841 and w66;
w3720 <= pi0093 and not w3719;
w3721 <= not w3718 and not w3720;
w3722 <= not pi0035 and not w3721;
w3723 <= not pi0070 and not w292;
w3724 <= not w3722 and w3723;
w3725 <= not pi0051 and not w3724;
w3726 <= w311 and not w3725;
w3727 <= w731 and not w3726;
w3728 <= w309 and not w3727;
w3729 <= w307 and not w3728;
w3730 <= not pi0198 and not pi0299;
w3731 <= not pi0210 and pi0299;
w3732 <= not w3730 and not w3731;
w3733 <= not pi0035 and w71;
w3734 <= not pi0040 and w3733;
w3735 <= w478 and w3734;
w3736 <= pi0032 and not w3735;
w3737 <= not w3732 and not w3736;
w3738 <= not w975 and w3732;
w3739 <= not w3737 and not w3738;
w3740 <= not w3729 and not w3739;
w3741 <= not pi0095 and not w3740;
w3742 <= not w304 and not w3741;
w3743 <= not pi0039 and not w3742;
w3744 <= pi0835 and pi0984;
w3745 <= not pi0252 and not pi1001;
w3746 <= not pi0979 and not w3745;
w3747 <= not w3744 and w3746;
w3748 <= not pi0287 and w3747;
w3749 <= pi0835 and pi0950;
w3750 <= w3748 and w3749;
w3751 <= w491 and w3750;
w3752 <= pi0222 and pi0224;
w3753 <= pi0603 and not pi0642;
w3754 <= not pi0614 and not pi0616;
w3755 <= w3753 and w3754;
w3756 <= not pi0662 and pi0680;
w3757 <= not pi0661 and w3756;
w3758 <= not pi0681 and w3757;
w3759 <= not w3755 and not w3758;
w3760 <= not pi0332 and not pi0468;
w3761 <= not w3759 and not w3760;
w3762 <= not pi0587 and not pi0602;
w3763 <= not pi0961 and not pi0967;
w3764 <= not pi0969 and not pi0971;
w3765 <= not pi0974 and not pi0977;
w3766 <= w3764 and w3765;
w3767 <= w3762 and w3763;
w3768 <= w3766 and w3767;
w3769 <= w3760 and not w3768;
w3770 <= not w3761 and not w3769;
w3771 <= w3751 and w3752;
w3772 <= not w3770 and w3771;
w3773 <= w84 and not w3772;
w3774 <= not pi0223 and not w3773;
w3775 <= pi1092 and w3750;
w3776 <= not pi0824 and not pi0829;
w3777 <= pi0824 and not pi1091;
w3778 <= pi1093 and not w487;
w3779 <= not w3777 and w3778;
w3780 <= not w3776 and not w3779;
w3781 <= w3775 and w3780;
w3782 <= not w3760 and not w3781;
w3783 <= not w3759 and not w3782;
w3784 <= w84 and not w3783;
w3785 <= w75 and w3760;
w3786 <= not w3759 and w3785;
w3787 <= not w3784 and not w3786;
w3788 <= w3768 and not w3787;
w3789 <= not w3755 and not w3760;
w3790 <= not w3758 and w3789;
w3791 <= w3781 and not w3790;
w3792 <= w84 and not w3791;
w3793 <= not w3768 and w3792;
w3794 <= pi0223 and not w3793;
w3795 <= not w3788 and w3794;
w3796 <= not pi0299 and not w3774;
w3797 <= not w3795 and w3796;
w3798 <= pi0216 and pi0221;
w3799 <= not pi0907 and not pi0947;
w3800 <= not pi0960 and not pi0963;
w3801 <= not pi0970 and not pi0972;
w3802 <= not pi0975 and not pi0978;
w3803 <= w3801 and w3802;
w3804 <= w3800 and w3803;
w3805 <= w3799 and w3804;
w3806 <= w3760 and not w3805;
w3807 <= not w3761 and not w3806;
w3808 <= w3751 and w3798;
w3809 <= not w3807 and w3808;
w3810 <= w84 and not w3809;
w3811 <= not pi0215 and not w3810;
w3812 <= w3792 and not w3805;
w3813 <= not w3787 and w3805;
w3814 <= pi0215 and not w3812;
w3815 <= not w3813 and w3814;
w3816 <= pi0299 and not w3811;
w3817 <= not w3815 and w3816;
w3818 <= pi0039 and not w3797;
w3819 <= not w3817 and w3818;
w3820 <= not w3743 and not w3819;
w3821 <= not pi0038 and not w3820;
w3822 <= w3700 and not w3821;
w3823 <= not pi0142 and not w232;
w3824 <= not pi0299 and w3823;
w3825 <= pi0299 and w203;
w3826 <= not w3824 and not w3825;
w3827 <= not w948 and w3826;
w3828 <= not pi0041 and not pi0099;
w3829 <= not pi0101 and w3828;
w3830 <= not pi0042 and not pi0043;
w3831 <= not pi0052 and w3830;
w3832 <= not pi0113 and not pi0116;
w3833 <= not pi0114 and not pi0115;
w3834 <= w3832 and w3833;
w3835 <= w3831 and w3834;
w3836 <= w3829 and w3835;
w3837 <= not pi0044 and w3836;
w3838 <= not pi0683 and not w3837;
w3839 <= pi0129 and pi0250;
w3840 <= w495 and not w3776;
w3841 <= not pi1093 and w3840;
w3842 <= not pi0250 and not w3841;
w3843 <= not w3839 and not w3842;
w3844 <= not w3838 and not w3843;
w3845 <= not w3826 and not w3837;
w3846 <= w3844 and w3845;
w3847 <= not pi0039 and w84;
w3848 <= not pi0038 and pi0100;
w3849 <= w3847 and w3848;
w3850 <= not w3827 and not w3846;
w3851 <= w3849 and w3850;
w3852 <= not pi0087 and not w3851;
w3853 <= not w3822 and w3852;
w3854 <= w3696 and w3697;
w3855 <= not w3853 and w3854;
w3856 <= not pi0074 and not w3855;
w3857 <= w3694 and not w3856;
w3858 <= not pi0056 and not w3857;
w3859 <= not w3690 and not w3858;
w3860 <= not pi0062 and not w3859;
w3861 <= w893 and w3688;
w3862 <= pi0062 and not w3861;
w3863 <= not pi0059 and not w3862;
w3864 <= not w3860 and w3863;
w3865 <= not pi0057 and not w3864;
w3866 <= not w3687 and not w3865;
w3867 <= not pi0055 and w92;
w3868 <= not pi0059 and w3867;
w3869 <= not pi0228 and not w3868;
w3870 <= pi0057 and not w3869;
w3871 <= not w3758 and not w3760;
w3872 <= not pi0907 and w3760;
w3873 <= not w3871 and not w3872;
w3874 <= not pi0228 and not w135;
w3875 <= pi0030 and pi0228;
w3876 <= not w898 and not w3875;
w3877 <= not w3874 and not w3876;
w3878 <= w3873 and w3877;
w3879 <= w3870 and w3878;
w3880 <= not pi0228 and not w3867;
w3881 <= w3878 and not w3880;
w3882 <= pi0059 and not w3881;
w3883 <= w3873 and w3875;
w3884 <= not w92 and w3883;
w3885 <= pi0055 and not w3878;
w3886 <= not pi0054 and w132;
w3887 <= pi0299 and w3873;
w3888 <= not pi0602 and w3760;
w3889 <= not w3871 and not w3888;
w3890 <= not pi0299 and w3889;
w3891 <= not w3887 and not w3890;
w3892 <= w3875 and not w3891;
w3893 <= not w3886 and not w3892;
w3894 <= not w173 and w3892;
w3895 <= not pi0039 and not w3876;
w3896 <= not w3891 and w3895;
w3897 <= w183 and w3896;
w3898 <= not w3894 and not w3897;
w3899 <= w132 and w3898;
w3900 <= not pi0054 and w3899;
w3901 <= pi0074 and not w3893;
w3902 <= not w3900 and w3901;
w3903 <= not w132 and not w3892;
w3904 <= not w3899 and not w3903;
w3905 <= pi0054 and not w3904;
w3906 <= not pi0075 and w3898;
w3907 <= pi0075 and not w3892;
w3908 <= pi0092 and not w3907;
w3909 <= not w3906 and w3908;
w3910 <= pi0075 and w3898;
w3911 <= pi0087 and w3892;
w3912 <= not w93 and w3892;
w3913 <= w3875 and w3889;
w3914 <= w84 and not w3843;
w3915 <= pi0683 and not w3837;
w3916 <= w3914 and w3915;
w3917 <= not w3871 and w3916;
w3918 <= w3823 and w3917;
w3919 <= pi0252 and not w3823;
w3920 <= pi0252 and w3785;
w3921 <= not w3758 and w3920;
w3922 <= pi0252 and w84;
w3923 <= w3758 and w3922;
w3924 <= not w3921 and not w3923;
w3925 <= w3919 and not w3924;
w3926 <= not w3918 and not w3925;
w3927 <= not pi0228 and not w3888;
w3928 <= not w3926 and w3927;
w3929 <= not pi0299 and not w3913;
w3930 <= not w3928 and w3929;
w3931 <= pi0299 and not w3883;
w3932 <= w203 and not w3917;
w3933 <= not w203 and w3924;
w3934 <= not pi0228 and not w3872;
w3935 <= not w3932 and w3934;
w3936 <= not w3933 and w3935;
w3937 <= w3931 and not w3936;
w3938 <= w93 and not w3937;
w3939 <= not w3930 and w3938;
w3940 <= pi0100 and not w3912;
w3941 <= not w3939 and w3940;
w3942 <= not pi0215 and pi0221;
w3943 <= not pi0287 and w84;
w3944 <= pi0835 and w3747;
w3945 <= w3943 and w3944;
w3946 <= pi0824 and pi1093;
w3947 <= w495 and w3946;
w3948 <= w3945 and w3947;
w3949 <= not pi1091 and w3948;
w3950 <= pi1091 and w486;
w3951 <= w3947 and not w3950;
w3952 <= not w491 and not w3951;
w3953 <= pi1091 and not w3952;
w3954 <= w3945 and w3953;
w3955 <= not w3949 and not w3954;
w3956 <= pi0216 and not w3955;
w3957 <= not pi0829 and not w486;
w3958 <= pi1091 and not w3957;
w3959 <= w3948 and not w3958;
w3960 <= not pi0216 and w3959;
w3961 <= not w3956 and not w3960;
w3962 <= not pi0228 and not w3961;
w3963 <= not w3875 and not w3962;
w3964 <= w3942 and not w3963;
w3965 <= not w3875 and not w3964;
w3966 <= w3873 and not w3965;
w3967 <= pi0299 and not w3966;
w3968 <= pi0222 and not pi0223;
w3969 <= not pi0224 and not w3959;
w3970 <= pi0224 and w3955;
w3971 <= w3968 and not w3969;
w3972 <= not w3970 and w3971;
w3973 <= not pi0228 and w3972;
w3974 <= not w3875 and not w3973;
w3975 <= w3889 and not w3974;
w3976 <= not pi0299 and not w3975;
w3977 <= pi0039 and not w3976;
w3978 <= not w3967 and w3977;
w3979 <= pi0158 and pi0159;
w3980 <= pi0160 and pi0197;
w3981 <= w3979 and w3980;
w3982 <= pi0091 and not w318;
w3983 <= not pi0058 and not w3982;
w3984 <= not pi0091 and not pi0314;
w3985 <= w328 and not w329;
w3986 <= pi0067 and w46;
w3987 <= pi0085 and w390;
w3988 <= w32 and not w3987;
w3989 <= w394 and not w3988;
w3990 <= w41 and not w3989;
w3991 <= not w373 and not w374;
w3992 <= not w3990 and w3991;
w3993 <= w42 and w3992;
w3994 <= not w370 and not w3993;
w3995 <= w367 and not w3994;
w3996 <= w360 and not w3986;
w3997 <= not w3995 and w3996;
w3998 <= w359 and not w3997;
w3999 <= not pi0071 and not w3998;
w4000 <= not pi0064 and w50;
w4001 <= w354 and w4000;
w4002 <= not w3999 and w4001;
w4003 <= not pi0081 and not w4002;
w4004 <= w408 and w4001;
w4005 <= w4003 and not w4004;
w4006 <= not pi0102 and not w349;
w4007 <= w26 and w4006;
w4008 <= not w4005 and w4007;
w4009 <= w348 and not w4008;
w4010 <= w440 and not w4009;
w4011 <= w282 and not w4010;
w4012 <= not w285 and not w4011;
w4013 <= not pi0086 and not w4012;
w4014 <= not pi0046 and w59;
w4015 <= w346 and w4014;
w4016 <= not w4013 and w4015;
w4017 <= w452 and not w4016;
w4018 <= w3985 and not w4017;
w4019 <= w3984 and not w4018;
w4020 <= not pi0091 and pi0314;
w4021 <= not w4003 and w4007;
w4022 <= w348 and not w4021;
w4023 <= w440 and not w4022;
w4024 <= w282 and not w4023;
w4025 <= not w285 and not w4024;
w4026 <= not pi0086 and not w4025;
w4027 <= w4015 and not w4026;
w4028 <= w452 and not w4027;
w4029 <= w3985 and not w4028;
w4030 <= w4020 and not w4029;
w4031 <= w3983 and not w4030;
w4032 <= not w4019 and w4031;
w4033 <= not pi0090 and not w4032;
w4034 <= not w459 and not w4033;
w4035 <= not pi0093 and not w4034;
w4036 <= pi0093 and not w477;
w4037 <= not pi0035 and not w4036;
w4038 <= not w4035 and w4037;
w4039 <= not pi0070 and not w4038;
w4040 <= w663 and not w4039;
w4041 <= not pi0072 and not w4040;
w4042 <= not pi0095 and w73;
w4043 <= not w308 and w4042;
w4044 <= not w4041 and w4043;
w4045 <= not w744 and not w4044;
w4046 <= not pi0841 and w291;
w4047 <= w525 and w4046;
w4048 <= w299 and w4047;
w4049 <= pi0032 and w4048;
w4050 <= not pi0095 and w4049;
w4051 <= not pi0210 and w4050;
w4052 <= w4045 and not w4051;
w4053 <= not w3760 and not w4052;
w4054 <= not pi0047 and w56;
w4055 <= not w451 and not w4016;
w4056 <= w4054 and not w4055;
w4057 <= w3984 and not w4056;
w4058 <= not w451 and not w4027;
w4059 <= w4054 and not w4058;
w4060 <= w4020 and not w4059;
w4061 <= w3983 and not w4060;
w4062 <= not w4057 and w4061;
w4063 <= not pi0090 and not w4062;
w4064 <= not w459 and not w4063;
w4065 <= not pi0093 and not w4064;
w4066 <= w4037 and not w4065;
w4067 <= not pi0070 and not w4066;
w4068 <= w663 and not w4067;
w4069 <= not pi0072 and not w4068;
w4070 <= w4043 and not w4069;
w4071 <= not w744 and not w4070;
w4072 <= not w4051 and w4071;
w4073 <= w3760 and not w4072;
w4074 <= not w4053 and not w4073;
w4075 <= w3873 and not w4074;
w4076 <= w3981 and not w4075;
w4077 <= w3873 and not w4052;
w4078 <= not w3981 and not w4077;
w4079 <= not pi0228 and not w4078;
w4080 <= not w4076 and w4079;
w4081 <= w3931 and not w4080;
w4082 <= not pi0198 and w4050;
w4083 <= w4045 and not w4082;
w4084 <= not pi0228 and not w4083;
w4085 <= not w3875 and not w4084;
w4086 <= w3889 and not w4085;
w4087 <= not pi0299 and not w4086;
w4088 <= pi0145 and pi0180;
w4089 <= pi0181 and pi0182;
w4090 <= w4088 and w4089;
w4091 <= not pi0299 and w4090;
w4092 <= not w4087 and not w4091;
w4093 <= not w3760 and not w4083;
w4094 <= w4071 and not w4082;
w4095 <= w3760 and not w4094;
w4096 <= not w4093 and not w4095;
w4097 <= not pi0228 and w3889;
w4098 <= not w4096 and w4097;
w4099 <= not w3913 and not w4098;
w4100 <= w4090 and not w4099;
w4101 <= not w4092 and not w4100;
w4102 <= pi0232 and not w4081;
w4103 <= not w4101 and w4102;
w4104 <= not pi0228 and w4077;
w4105 <= w3931 and not w4104;
w4106 <= not pi0232 and not w4105;
w4107 <= not w4087 and w4106;
w4108 <= not w4103 and not w4107;
w4109 <= not pi0039 and not w4108;
w4110 <= not pi0038 and not w3978;
w4111 <= not w4109 and w4110;
w4112 <= pi0038 and not w3892;
w4113 <= not w3896 and w4112;
w4114 <= not w4111 and not w4113;
w4115 <= not pi0100 and not w4114;
w4116 <= not pi0087 and not w3941;
w4117 <= not w4115 and w4116;
w4118 <= not pi0075 and not w3911;
w4119 <= not w4117 and w4118;
w4120 <= not pi0092 and not w3910;
w4121 <= not w4119 and w4120;
w4122 <= not pi0054 and not w3909;
w4123 <= not w4121 and w4122;
w4124 <= not pi0074 and not w3905;
w4125 <= not w4123 and w4124;
w4126 <= not pi0055 and not w3902;
w4127 <= not w4125 and w4126;
w4128 <= w92 and not w3885;
w4129 <= not w4127 and w4128;
w4130 <= not pi0059 and not w3884;
w4131 <= not w4129 and w4130;
w4132 <= not pi0057 and not w3882;
w4133 <= not w4131 and w4132;
w4134 <= not w3879 and not w4133;
w4135 <= not pi0947 and w3760;
w4136 <= not w3789 and not w4135;
w4137 <= w3877 and w4136;
w4138 <= w3870 and w4137;
w4139 <= not w3880 and w4137;
w4140 <= pi0059 and not w4139;
w4141 <= w3875 and w4136;
w4142 <= not w92 and w4141;
w4143 <= pi0055 and not w4137;
w4144 <= pi0299 and not w4136;
w4145 <= not pi0587 and w3760;
w4146 <= not w3789 and not w4145;
w4147 <= not pi0299 and not w4146;
w4148 <= not w4144 and not w4147;
w4149 <= w3875 and w4148;
w4150 <= not w3886 and not w4149;
w4151 <= not w173 and w4149;
w4152 <= w3895 and w4148;
w4153 <= w183 and w4152;
w4154 <= not w4151 and not w4153;
w4155 <= w132 and w4154;
w4156 <= not pi0054 and w4155;
w4157 <= pi0074 and not w4150;
w4158 <= not w4156 and w4157;
w4159 <= not w132 and not w4149;
w4160 <= not w4155 and not w4159;
w4161 <= pi0054 and not w4160;
w4162 <= not pi0075 and w4154;
w4163 <= pi0075 and not w4149;
w4164 <= pi0092 and not w4163;
w4165 <= not w4162 and w4164;
w4166 <= pi0075 and w4154;
w4167 <= pi0087 and w4149;
w4168 <= not w93 and w4149;
w4169 <= pi0299 and not w4141;
w4170 <= not w3789 and w3916;
w4171 <= w203 and not w4135;
w4172 <= w4170 and w4171;
w4173 <= not w3755 and not w3920;
w4174 <= w3755 and not w3922;
w4175 <= not w4173 and not w4174;
w4176 <= w3755 and not w3760;
w4177 <= not pi0947 and not w4176;
w4178 <= not w203 and not w4177;
w4179 <= w4175 and w4178;
w4180 <= not w4172 and not w4179;
w4181 <= not pi0228 and not w4180;
w4182 <= w4169 and not w4181;
w4183 <= not pi0228 and w232;
w4184 <= not w4145 and w4175;
w4185 <= w4183 and not w4184;
w4186 <= not pi0587 and not w4176;
w4187 <= pi0142 and not w4175;
w4188 <= not pi0142 and not w4170;
w4189 <= not pi0228 and not w4186;
w4190 <= not w4188 and w4189;
w4191 <= not w4187 and w4190;
w4192 <= w3875 and w4146;
w4193 <= not w4183 and not w4192;
w4194 <= not w4191 and w4193;
w4195 <= not w4185 and not w4194;
w4196 <= not pi0299 and not w4195;
w4197 <= w93 and not w4182;
w4198 <= not w4196 and w4197;
w4199 <= pi0100 and not w4168;
w4200 <= not w4198 and w4199;
w4201 <= not w3974 and w4146;
w4202 <= not pi0299 and not w4201;
w4203 <= pi0299 and w3942;
w4204 <= not w4169 and not w4203;
w4205 <= w3964 and w4136;
w4206 <= not w4204 and not w4205;
w4207 <= pi0039 and not w4202;
w4208 <= not w4206 and w4207;
w4209 <= not w4074 and w4136;
w4210 <= w3981 and not w4209;
w4211 <= not w4052 and w4136;
w4212 <= not w3981 and not w4211;
w4213 <= not pi0228 and not w4212;
w4214 <= not w4210 and w4213;
w4215 <= w4169 and not w4214;
w4216 <= not w4085 and w4146;
w4217 <= not w4090 and w4216;
w4218 <= not pi0228 and w4146;
w4219 <= not w4096 and w4218;
w4220 <= not w4192 and not w4219;
w4221 <= w4090 and not w4220;
w4222 <= not pi0299 and not w4217;
w4223 <= not w4221 and w4222;
w4224 <= pi0232 and not w4215;
w4225 <= not w4223 and w4224;
w4226 <= not pi0228 and w4211;
w4227 <= w4169 and not w4226;
w4228 <= not pi0299 and not w4216;
w4229 <= not pi0232 and not w4227;
w4230 <= not w4228 and w4229;
w4231 <= not w4225 and not w4230;
w4232 <= not pi0039 and not w4231;
w4233 <= not pi0038 and not w4208;
w4234 <= not w4232 and w4233;
w4235 <= pi0038 and not w4149;
w4236 <= not w4152 and w4235;
w4237 <= not w4234 and not w4236;
w4238 <= not pi0100 and not w4237;
w4239 <= not pi0087 and not w4200;
w4240 <= not w4238 and w4239;
w4241 <= not pi0075 and not w4167;
w4242 <= not w4240 and w4241;
w4243 <= not pi0092 and not w4166;
w4244 <= not w4242 and w4243;
w4245 <= not pi0054 and not w4165;
w4246 <= not w4244 and w4245;
w4247 <= not pi0074 and not w4161;
w4248 <= not w4246 and w4247;
w4249 <= not pi0055 and not w4158;
w4250 <= not w4248 and w4249;
w4251 <= w92 and not w4143;
w4252 <= not w4250 and w4251;
w4253 <= not pi0059 and not w4142;
w4254 <= not w4252 and w4253;
w4255 <= not pi0057 and not w4140;
w4256 <= not w4254 and w4255;
w4257 <= not w4138 and not w4256;
w4258 <= pi0030 and w3760;
w4259 <= pi0228 and w4258;
w4260 <= pi0970 and w4259;
w4261 <= not pi0228 and pi0970;
w4262 <= w3785 and w4261;
w4263 <= w135 and w4262;
w4264 <= w3868 and w4263;
w4265 <= not w4260 and not w4264;
w4266 <= pi0057 and not w4265;
w4267 <= w3867 and w4263;
w4268 <= pi0059 and not w4260;
w4269 <= not w4267 and w4268;
w4270 <= not w92 and w4260;
w4271 <= pi0055 and not w4260;
w4272 <= not w4263 and w4271;
w4273 <= pi0299 and pi0970;
w4274 <= not pi0299 and pi0967;
w4275 <= not w4273 and not w4274;
w4276 <= w4259 and not w4275;
w4277 <= not w3886 and not w4276;
w4278 <= not w173 and w4276;
w4279 <= pi0299 and not w4260;
w4280 <= not w4262 and w4279;
w4281 <= pi0228 and not w4258;
w4282 <= not pi0228 and not w3785;
w4283 <= not w4281 and not w4282;
w4284 <= pi0967 and w4283;
w4285 <= not pi0299 and not w4284;
w4286 <= not pi0039 and not w4280;
w4287 <= not w4285 and w4286;
w4288 <= w183 and w4287;
w4289 <= not w4278 and not w4288;
w4290 <= w132 and w4289;
w4291 <= not pi0054 and w4290;
w4292 <= pi0074 and not w4277;
w4293 <= not w4291 and w4292;
w4294 <= not w132 and not w4276;
w4295 <= not w4290 and not w4294;
w4296 <= pi0054 and not w4295;
w4297 <= not pi0075 and w4289;
w4298 <= pi0075 and not w4276;
w4299 <= pi0092 and not w4298;
w4300 <= not w4297 and w4299;
w4301 <= pi0075 and w4289;
w4302 <= pi0087 and w4276;
w4303 <= not w93 and w4276;
w4304 <= not w203 and not w3920;
w4305 <= w3760 and w3916;
w4306 <= w203 and not w4305;
w4307 <= not pi0228 and not w4304;
w4308 <= not w4306 and w4307;
w4309 <= pi0970 and w4308;
w4310 <= w4279 and not w4309;
w4311 <= not w3823 and w3920;
w4312 <= w3823 and w4305;
w4313 <= not pi0228 and not w4311;
w4314 <= not w4312 and w4313;
w4315 <= not w4281 and not w4314;
w4316 <= pi0967 and w4315;
w4317 <= not pi0299 and not w4316;
w4318 <= w93 and not w4310;
w4319 <= not w4317 and w4318;
w4320 <= pi0100 and not w4303;
w4321 <= not w4319 and w4320;
w4322 <= w3942 and not w3961;
w4323 <= w3760 and w4322;
w4324 <= not pi0228 and not w4323;
w4325 <= w4273 and not w4324;
w4326 <= w3760 and w3972;
w4327 <= not pi0228 and not w4326;
w4328 <= w4274 and not w4327;
w4329 <= not w4325 and not w4328;
w4330 <= pi0039 and not w4281;
w4331 <= not w4329 and w4330;
w4332 <= w3760 and not w4085;
w4333 <= not w4090 and not w4332;
w4334 <= not w4083 and not w4090;
w4335 <= not pi0228 and w4095;
w4336 <= not w4259 and not w4334;
w4337 <= not w4335 and w4336;
w4338 <= not w4333 and not w4337;
w4339 <= pi0967 and w4338;
w4340 <= not pi0299 and not w4339;
w4341 <= w3760 and not w4052;
w4342 <= w4261 and w4341;
w4343 <= w4279 and not w4342;
w4344 <= pi0299 and w3979;
w4345 <= not w4343 and not w4344;
w4346 <= w3980 and not w4073;
w4347 <= not w3980 and w4052;
w4348 <= not w4346 and not w4347;
w4349 <= w3760 and w4348;
w4350 <= w4261 and w4349;
w4351 <= not w4260 and not w4350;
w4352 <= w3979 and not w4351;
w4353 <= not w4345 and not w4352;
w4354 <= pi0232 and not w4340;
w4355 <= not w4353 and w4354;
w4356 <= pi0967 and w4332;
w4357 <= not pi0299 and not w4356;
w4358 <= not pi0232 and not w4343;
w4359 <= not w4357 and w4358;
w4360 <= not w4355 and not w4359;
w4361 <= not pi0039 and not w4360;
w4362 <= not pi0038 and not w4331;
w4363 <= not w4361 and w4362;
w4364 <= pi0039 and w4276;
w4365 <= pi0038 and not w4364;
w4366 <= not w4287 and w4365;
w4367 <= not w4363 and not w4366;
w4368 <= not pi0100 and not w4367;
w4369 <= not pi0087 and not w4321;
w4370 <= not w4368 and w4369;
w4371 <= not pi0075 and not w4302;
w4372 <= not w4370 and w4371;
w4373 <= not pi0092 and not w4301;
w4374 <= not w4372 and w4373;
w4375 <= not pi0054 and not w4300;
w4376 <= not w4374 and w4375;
w4377 <= not pi0074 and not w4296;
w4378 <= not w4376 and w4377;
w4379 <= not pi0055 and not w4293;
w4380 <= not w4378 and w4379;
w4381 <= w92 and not w4272;
w4382 <= not w4380 and w4381;
w4383 <= not pi0059 and not w4270;
w4384 <= not w4382 and w4383;
w4385 <= not pi0057 and not w4269;
w4386 <= not w4384 and w4385;
w4387 <= not w4266 and not w4386;
w4388 <= pi0972 and w4259;
w4389 <= not pi0228 and pi0972;
w4390 <= w3785 and w4389;
w4391 <= w135 and w4390;
w4392 <= w3868 and w4391;
w4393 <= not w4388 and not w4392;
w4394 <= pi0057 and not w4393;
w4395 <= w3867 and w4391;
w4396 <= pi0059 and not w4388;
w4397 <= not w4395 and w4396;
w4398 <= not w92 and w4388;
w4399 <= pi0055 and not w4388;
w4400 <= not w4391 and w4399;
w4401 <= not pi0299 and pi0961;
w4402 <= pi0299 and pi0972;
w4403 <= not w4401 and not w4402;
w4404 <= w4259 and not w4403;
w4405 <= not w3886 and not w4404;
w4406 <= not w173 and w4404;
w4407 <= pi0299 and not w4388;
w4408 <= not w4390 and w4407;
w4409 <= pi0961 and w4283;
w4410 <= not pi0299 and not w4409;
w4411 <= not pi0039 and not w4408;
w4412 <= not w4410 and w4411;
w4413 <= w183 and w4412;
w4414 <= not w4406 and not w4413;
w4415 <= w132 and w4414;
w4416 <= not pi0054 and w4415;
w4417 <= pi0074 and not w4405;
w4418 <= not w4416 and w4417;
w4419 <= not w132 and not w4404;
w4420 <= not w4415 and not w4419;
w4421 <= pi0054 and not w4420;
w4422 <= not pi0075 and w4414;
w4423 <= pi0075 and not w4404;
w4424 <= pi0092 and not w4423;
w4425 <= not w4422 and w4424;
w4426 <= pi0075 and w4414;
w4427 <= pi0087 and w4404;
w4428 <= not w93 and w4404;
w4429 <= pi0972 and w4308;
w4430 <= w4407 and not w4429;
w4431 <= pi0961 and w4315;
w4432 <= not pi0299 and not w4431;
w4433 <= w93 and not w4430;
w4434 <= not w4432 and w4433;
w4435 <= pi0100 and not w4428;
w4436 <= not w4434 and w4435;
w4437 <= not w4327 and w4401;
w4438 <= not w4324 and w4402;
w4439 <= not w4437 and not w4438;
w4440 <= w4330 and not w4439;
w4441 <= pi0961 and w4338;
w4442 <= not pi0299 and not w4441;
w4443 <= w4341 and w4389;
w4444 <= w4407 and not w4443;
w4445 <= not w4344 and not w4444;
w4446 <= w4349 and w4389;
w4447 <= not w4388 and not w4446;
w4448 <= w3979 and not w4447;
w4449 <= not w4445 and not w4448;
w4450 <= pi0232 and not w4442;
w4451 <= not w4449 and w4450;
w4452 <= pi0961 and w4332;
w4453 <= not pi0299 and not w4452;
w4454 <= not pi0232 and not w4444;
w4455 <= not w4453 and w4454;
w4456 <= not w4451 and not w4455;
w4457 <= not pi0039 and not w4456;
w4458 <= not pi0038 and not w4440;
w4459 <= not w4457 and w4458;
w4460 <= pi0039 and w4404;
w4461 <= pi0038 and not w4460;
w4462 <= not w4412 and w4461;
w4463 <= not w4459 and not w4462;
w4464 <= not pi0100 and not w4463;
w4465 <= not pi0087 and not w4436;
w4466 <= not w4464 and w4465;
w4467 <= not pi0075 and not w4427;
w4468 <= not w4466 and w4467;
w4469 <= not pi0092 and not w4426;
w4470 <= not w4468 and w4469;
w4471 <= not pi0054 and not w4425;
w4472 <= not w4470 and w4471;
w4473 <= not pi0074 and not w4421;
w4474 <= not w4472 and w4473;
w4475 <= not pi0055 and not w4418;
w4476 <= not w4474 and w4475;
w4477 <= w92 and not w4400;
w4478 <= not w4476 and w4477;
w4479 <= not pi0059 and not w4398;
w4480 <= not w4478 and w4479;
w4481 <= not pi0057 and not w4397;
w4482 <= not w4480 and w4481;
w4483 <= not w4394 and not w4482;
w4484 <= pi0960 and w4259;
w4485 <= not pi0228 and pi0960;
w4486 <= w3785 and w4485;
w4487 <= w135 and w4486;
w4488 <= w3868 and w4487;
w4489 <= not w4484 and not w4488;
w4490 <= pi0057 and not w4489;
w4491 <= w3867 and w4487;
w4492 <= pi0059 and not w4484;
w4493 <= not w4491 and w4492;
w4494 <= not w92 and w4484;
w4495 <= pi0055 and not w4484;
w4496 <= not w4487 and w4495;
w4497 <= not pi0299 and pi0977;
w4498 <= pi0299 and pi0960;
w4499 <= not w4497 and not w4498;
w4500 <= w4259 and not w4499;
w4501 <= not w3886 and not w4500;
w4502 <= not w173 and w4500;
w4503 <= pi0299 and not w4484;
w4504 <= not w4486 and w4503;
w4505 <= pi0977 and w4283;
w4506 <= not pi0299 and not w4505;
w4507 <= not pi0039 and not w4504;
w4508 <= not w4506 and w4507;
w4509 <= w183 and w4508;
w4510 <= not w4502 and not w4509;
w4511 <= w132 and w4510;
w4512 <= not pi0054 and w4511;
w4513 <= pi0074 and not w4501;
w4514 <= not w4512 and w4513;
w4515 <= not w132 and not w4500;
w4516 <= not w4511 and not w4515;
w4517 <= pi0054 and not w4516;
w4518 <= not pi0075 and w4510;
w4519 <= pi0075 and not w4500;
w4520 <= pi0092 and not w4519;
w4521 <= not w4518 and w4520;
w4522 <= pi0075 and w4510;
w4523 <= pi0087 and w4500;
w4524 <= not w93 and w4500;
w4525 <= pi0960 and w4308;
w4526 <= w4503 and not w4525;
w4527 <= pi0977 and w4315;
w4528 <= not pi0299 and not w4527;
w4529 <= w93 and not w4526;
w4530 <= not w4528 and w4529;
w4531 <= pi0100 and not w4524;
w4532 <= not w4530 and w4531;
w4533 <= not w4327 and w4497;
w4534 <= not w4324 and w4498;
w4535 <= not w4533 and not w4534;
w4536 <= w4330 and not w4535;
w4537 <= pi0977 and w4338;
w4538 <= not pi0299 and not w4537;
w4539 <= w4341 and w4485;
w4540 <= w4503 and not w4539;
w4541 <= not w4344 and not w4540;
w4542 <= w4349 and w4485;
w4543 <= not w4484 and not w4542;
w4544 <= w3979 and not w4543;
w4545 <= not w4541 and not w4544;
w4546 <= pi0232 and not w4538;
w4547 <= not w4545 and w4546;
w4548 <= pi0977 and w4332;
w4549 <= not pi0299 and not w4548;
w4550 <= not pi0232 and not w4540;
w4551 <= not w4549 and w4550;
w4552 <= not w4547 and not w4551;
w4553 <= not pi0039 and not w4552;
w4554 <= not pi0038 and not w4536;
w4555 <= not w4553 and w4554;
w4556 <= pi0039 and w4500;
w4557 <= pi0038 and not w4556;
w4558 <= not w4508 and w4557;
w4559 <= not w4555 and not w4558;
w4560 <= not pi0100 and not w4559;
w4561 <= not pi0087 and not w4532;
w4562 <= not w4560 and w4561;
w4563 <= not pi0075 and not w4523;
w4564 <= not w4562 and w4563;
w4565 <= not pi0092 and not w4522;
w4566 <= not w4564 and w4565;
w4567 <= not pi0054 and not w4521;
w4568 <= not w4566 and w4567;
w4569 <= not pi0074 and not w4517;
w4570 <= not w4568 and w4569;
w4571 <= not pi0055 and not w4514;
w4572 <= not w4570 and w4571;
w4573 <= w92 and not w4496;
w4574 <= not w4572 and w4573;
w4575 <= not pi0059 and not w4494;
w4576 <= not w4574 and w4575;
w4577 <= not pi0057 and not w4493;
w4578 <= not w4576 and w4577;
w4579 <= not w4490 and not w4578;
w4580 <= pi0963 and w4259;
w4581 <= not pi0228 and pi0963;
w4582 <= w3785 and w4581;
w4583 <= w135 and w4582;
w4584 <= w3868 and w4583;
w4585 <= not w4580 and not w4584;
w4586 <= pi0057 and not w4585;
w4587 <= w3867 and w4583;
w4588 <= pi0059 and not w4580;
w4589 <= not w4587 and w4588;
w4590 <= not w92 and w4580;
w4591 <= pi0055 and not w4580;
w4592 <= not w4583 and w4591;
w4593 <= not pi0299 and pi0969;
w4594 <= pi0299 and pi0963;
w4595 <= not w4593 and not w4594;
w4596 <= w4259 and not w4595;
w4597 <= not w3886 and not w4596;
w4598 <= not w173 and w4596;
w4599 <= pi0299 and not w4580;
w4600 <= not w4582 and w4599;
w4601 <= pi0969 and w4283;
w4602 <= not pi0299 and not w4601;
w4603 <= not pi0039 and not w4600;
w4604 <= not w4602 and w4603;
w4605 <= w183 and w4604;
w4606 <= not w4598 and not w4605;
w4607 <= w132 and w4606;
w4608 <= not pi0054 and w4607;
w4609 <= pi0074 and not w4597;
w4610 <= not w4608 and w4609;
w4611 <= not w132 and not w4596;
w4612 <= not w4607 and not w4611;
w4613 <= pi0054 and not w4612;
w4614 <= not pi0075 and w4606;
w4615 <= pi0075 and not w4596;
w4616 <= pi0092 and not w4615;
w4617 <= not w4614 and w4616;
w4618 <= pi0075 and w4606;
w4619 <= pi0087 and w4596;
w4620 <= not w93 and w4596;
w4621 <= pi0963 and w4308;
w4622 <= w4599 and not w4621;
w4623 <= pi0969 and w4315;
w4624 <= not pi0299 and not w4623;
w4625 <= w93 and not w4622;
w4626 <= not w4624 and w4625;
w4627 <= pi0100 and not w4620;
w4628 <= not w4626 and w4627;
w4629 <= not w4327 and w4593;
w4630 <= not w4324 and w4594;
w4631 <= not w4629 and not w4630;
w4632 <= w4330 and not w4631;
w4633 <= pi0969 and w4338;
w4634 <= not pi0299 and not w4633;
w4635 <= w4341 and w4581;
w4636 <= w4599 and not w4635;
w4637 <= not w4344 and not w4636;
w4638 <= w4349 and w4581;
w4639 <= not w4580 and not w4638;
w4640 <= w3979 and not w4639;
w4641 <= not w4637 and not w4640;
w4642 <= pi0232 and not w4634;
w4643 <= not w4641 and w4642;
w4644 <= pi0969 and w4332;
w4645 <= not pi0299 and not w4644;
w4646 <= not pi0232 and not w4636;
w4647 <= not w4645 and w4646;
w4648 <= not w4643 and not w4647;
w4649 <= not pi0039 and not w4648;
w4650 <= not pi0038 and not w4632;
w4651 <= not w4649 and w4650;
w4652 <= pi0039 and w4596;
w4653 <= pi0038 and not w4652;
w4654 <= not w4604 and w4653;
w4655 <= not w4651 and not w4654;
w4656 <= not pi0100 and not w4655;
w4657 <= not pi0087 and not w4628;
w4658 <= not w4656 and w4657;
w4659 <= not pi0075 and not w4619;
w4660 <= not w4658 and w4659;
w4661 <= not pi0092 and not w4618;
w4662 <= not w4660 and w4661;
w4663 <= not pi0054 and not w4617;
w4664 <= not w4662 and w4663;
w4665 <= not pi0074 and not w4613;
w4666 <= not w4664 and w4665;
w4667 <= not pi0055 and not w4610;
w4668 <= not w4666 and w4667;
w4669 <= w92 and not w4592;
w4670 <= not w4668 and w4669;
w4671 <= not pi0059 and not w4590;
w4672 <= not w4670 and w4671;
w4673 <= not pi0057 and not w4589;
w4674 <= not w4672 and w4673;
w4675 <= not w4586 and not w4674;
w4676 <= pi0975 and w4259;
w4677 <= not pi0228 and pi0975;
w4678 <= w3785 and w4677;
w4679 <= w135 and w4678;
w4680 <= w3868 and w4679;
w4681 <= not w4676 and not w4680;
w4682 <= pi0057 and not w4681;
w4683 <= w3867 and w4679;
w4684 <= pi0059 and not w4676;
w4685 <= not w4683 and w4684;
w4686 <= not w92 and w4676;
w4687 <= pi0055 and not w4676;
w4688 <= not w4679 and w4687;
w4689 <= not pi0299 and pi0971;
w4690 <= pi0299 and pi0975;
w4691 <= not w4689 and not w4690;
w4692 <= w4259 and not w4691;
w4693 <= not w3886 and not w4692;
w4694 <= not w173 and w4692;
w4695 <= pi0299 and not w4676;
w4696 <= not w4678 and w4695;
w4697 <= pi0971 and w4283;
w4698 <= not pi0299 and not w4697;
w4699 <= not pi0039 and not w4696;
w4700 <= not w4698 and w4699;
w4701 <= w183 and w4700;
w4702 <= not w4694 and not w4701;
w4703 <= w132 and w4702;
w4704 <= not pi0054 and w4703;
w4705 <= pi0074 and not w4693;
w4706 <= not w4704 and w4705;
w4707 <= not w132 and not w4692;
w4708 <= not w4703 and not w4707;
w4709 <= pi0054 and not w4708;
w4710 <= not pi0075 and w4702;
w4711 <= pi0075 and not w4692;
w4712 <= pi0092 and not w4711;
w4713 <= not w4710 and w4712;
w4714 <= pi0075 and w4702;
w4715 <= pi0087 and w4692;
w4716 <= not w93 and w4692;
w4717 <= pi0975 and w4308;
w4718 <= w4695 and not w4717;
w4719 <= pi0971 and w4315;
w4720 <= not pi0299 and not w4719;
w4721 <= w93 and not w4718;
w4722 <= not w4720 and w4721;
w4723 <= pi0100 and not w4716;
w4724 <= not w4722 and w4723;
w4725 <= not w4327 and w4689;
w4726 <= not w4324 and w4690;
w4727 <= not w4725 and not w4726;
w4728 <= w4330 and not w4727;
w4729 <= pi0971 and w4338;
w4730 <= not pi0299 and not w4729;
w4731 <= w4341 and w4677;
w4732 <= w4695 and not w4731;
w4733 <= not w4344 and not w4732;
w4734 <= w4349 and w4677;
w4735 <= not w4676 and not w4734;
w4736 <= w3979 and not w4735;
w4737 <= not w4733 and not w4736;
w4738 <= pi0232 and not w4730;
w4739 <= not w4737 and w4738;
w4740 <= pi0971 and w4332;
w4741 <= not pi0299 and not w4740;
w4742 <= not pi0232 and not w4732;
w4743 <= not w4741 and w4742;
w4744 <= not w4739 and not w4743;
w4745 <= not pi0039 and not w4744;
w4746 <= not pi0038 and not w4728;
w4747 <= not w4745 and w4746;
w4748 <= pi0039 and w4692;
w4749 <= pi0038 and not w4748;
w4750 <= not w4700 and w4749;
w4751 <= not w4747 and not w4750;
w4752 <= not pi0100 and not w4751;
w4753 <= not pi0087 and not w4724;
w4754 <= not w4752 and w4753;
w4755 <= not pi0075 and not w4715;
w4756 <= not w4754 and w4755;
w4757 <= not pi0092 and not w4714;
w4758 <= not w4756 and w4757;
w4759 <= not pi0054 and not w4713;
w4760 <= not w4758 and w4759;
w4761 <= not pi0074 and not w4709;
w4762 <= not w4760 and w4761;
w4763 <= not pi0055 and not w4706;
w4764 <= not w4762 and w4763;
w4765 <= w92 and not w4688;
w4766 <= not w4764 and w4765;
w4767 <= not pi0059 and not w4686;
w4768 <= not w4766 and w4767;
w4769 <= not pi0057 and not w4685;
w4770 <= not w4768 and w4769;
w4771 <= not w4682 and not w4770;
w4772 <= pi0978 and w4259;
w4773 <= not pi0228 and pi0978;
w4774 <= w135 and w4773;
w4775 <= w3785 and w4774;
w4776 <= w3868 and w4775;
w4777 <= not w4772 and not w4776;
w4778 <= pi0057 and not w4777;
w4779 <= w3867 and w4775;
w4780 <= pi0059 and not w4772;
w4781 <= not w4779 and w4780;
w4782 <= not w92 and w4772;
w4783 <= pi0055 and not w4772;
w4784 <= not w4775 and w4783;
w4785 <= not pi0299 and pi0974;
w4786 <= pi0299 and pi0978;
w4787 <= not w4785 and not w4786;
w4788 <= w4259 and not w4787;
w4789 <= not w3886 and not w4788;
w4790 <= w4283 and not w4787;
w4791 <= not pi0228 and not w173;
w4792 <= w4790 and not w4791;
w4793 <= w132 and not w4792;
w4794 <= not pi0054 and w4793;
w4795 <= pi0074 and not w4789;
w4796 <= not w4794 and w4795;
w4797 <= not w132 and not w4788;
w4798 <= not w4793 and not w4797;
w4799 <= pi0054 and not w4798;
w4800 <= not pi0075 and not w4792;
w4801 <= pi0075 and not w4788;
w4802 <= pi0092 and not w4801;
w4803 <= not w4800 and w4802;
w4804 <= pi0075 and not w4792;
w4805 <= pi0087 and w4788;
w4806 <= not w93 and w4788;
w4807 <= pi0299 and not w4772;
w4808 <= pi0978 and w4308;
w4809 <= w4807 and not w4808;
w4810 <= pi0974 and w4315;
w4811 <= not pi0299 and not w4810;
w4812 <= w93 and not w4809;
w4813 <= not w4811 and w4812;
w4814 <= pi0100 and not w4806;
w4815 <= not w4813 and w4814;
w4816 <= pi0039 and w4788;
w4817 <= not pi0039 and w4790;
w4818 <= pi0038 and not w4816;
w4819 <= not w4817 and w4818;
w4820 <= not w4327 and w4785;
w4821 <= not w4324 and w4786;
w4822 <= not w4820 and not w4821;
w4823 <= w4330 and not w4822;
w4824 <= pi0974 and w4338;
w4825 <= not pi0299 and not w4824;
w4826 <= w4341 and w4773;
w4827 <= w4807 and not w4826;
w4828 <= not w4344 and not w4827;
w4829 <= w4349 and w4773;
w4830 <= not w4772 and not w4829;
w4831 <= w3979 and not w4830;
w4832 <= not w4828 and not w4831;
w4833 <= pi0232 and not w4825;
w4834 <= not w4832 and w4833;
w4835 <= pi0974 and w4332;
w4836 <= not pi0299 and not w4835;
w4837 <= not pi0232 and not w4827;
w4838 <= not w4836 and w4837;
w4839 <= not w4834 and not w4838;
w4840 <= not pi0039 and not w4839;
w4841 <= not pi0038 and not w4823;
w4842 <= not w4840 and w4841;
w4843 <= not w4819 and not w4842;
w4844 <= not pi0100 and not w4843;
w4845 <= not pi0087 and not w4815;
w4846 <= not w4844 and w4845;
w4847 <= not pi0075 and not w4805;
w4848 <= not w4846 and w4847;
w4849 <= not pi0092 and not w4804;
w4850 <= not w4848 and w4849;
w4851 <= not pi0054 and not w4803;
w4852 <= not w4850 and w4851;
w4853 <= not pi0074 and not w4799;
w4854 <= not w4852 and w4853;
w4855 <= not pi0055 and not w4796;
w4856 <= not w4854 and w4855;
w4857 <= w92 and not w4784;
w4858 <= not w4856 and w4857;
w4859 <= not pi0059 and not w4782;
w4860 <= not w4858 and w4859;
w4861 <= not pi0057 and not w4781;
w4862 <= not w4860 and w4861;
w4863 <= not w4778 and not w4862;
w4864 <= w183 and w3847;
w4865 <= pi0075 and not w4864;
w4866 <= w96 and w171;
w4867 <= w3847 and w4866;
w4868 <= pi0092 and not w4867;
w4869 <= not w4865 and not w4868;
w4870 <= pi0299 and not w3807;
w4871 <= w4322 and w4870;
w4872 <= not pi0299 and not w3770;
w4873 <= w3972 and w4872;
w4874 <= pi0039 and not w4873;
w4875 <= not w4871 and w4874;
w4876 <= pi0299 and w4052;
w4877 <= not pi0299 and w4083;
w4878 <= not pi0232 and not w4876;
w4879 <= not w4877 and w4878;
w4880 <= w4090 and w4095;
w4881 <= not pi0299 and not w4093;
w4882 <= not w4334 and w4881;
w4883 <= not w4880 and w4882;
w4884 <= not w3979 and w4876;
w4885 <= not w4053 and w4344;
w4886 <= not w4348 and w4885;
w4887 <= pi0232 and not w4884;
w4888 <= not w4883 and w4887;
w4889 <= not w4886 and w4888;
w4890 <= not pi0039 and not w4879;
w4891 <= not w4889 and w4890;
w4892 <= not w4875 and not w4891;
w4893 <= not pi0038 and not w4892;
w4894 <= not w3699 and not w4893;
w4895 <= not pi0100 and not w4894;
w4896 <= not pi0038 and w3847;
w4897 <= pi0100 and not w4896;
w4898 <= w3852 and not w4897;
w4899 <= not w4895 and w4898;
w4900 <= w132 and not w4899;
w4901 <= w4869 and not w4900;
w4902 <= not pi0054 and not w4901;
w4903 <= not pi0092 and w4867;
w4904 <= pi0054 and not w4903;
w4905 <= not w4902 and not w4904;
w4906 <= not pi0074 and not w4905;
w4907 <= not w3693 and not w4906;
w4908 <= not pi0055 and not w4907;
w4909 <= w98 and w3688;
w4910 <= pi0055 and not w4909;
w4911 <= not pi0056 and not w4910;
w4912 <= not pi0062 and w4911;
w4913 <= not w4908 and w4912;
w4914 <= w891 and not w4913;
w4915 <= w3686 and not w4914;
w4916 <= not pi0954 and not w4915;
w4917 <= pi0024 and pi0954;
w4918 <= not w4916 and not w4917;
w4919 <= w94 and w898;
w4920 <= w893 and w4919;
w4921 <= not w4 and not w4920;
w4922 <= pi0062 and not w4921;
w4923 <= w100 and w898;
w4924 <= pi0056 and not w4;
w4925 <= not w4923 and w4924;
w4926 <= w94 and w3691;
w4927 <= w898 and w4926;
w4928 <= not pi0074 and w4927;
w4929 <= not w4 and not w4928;
w4930 <= pi0055 and not w4929;
w4931 <= not w4 and not w95;
w4932 <= w898 and w936;
w4933 <= not w4 and not w4932;
w4934 <= pi0092 and not w4933;
w4935 <= pi0075 and not w4;
w4936 <= not w4 and not w4919;
w4937 <= pi0087 and not w4936;
w4938 <= not pi0100 and w2293;
w4939 <= w84 and not w3919;
w4940 <= not pi0299 and not w4939;
w4941 <= pi0299 and not w957;
w4942 <= not w4940 and not w4941;
w4943 <= pi0100 and w898;
w4944 <= w4942 and w4943;
w4945 <= not pi0039 and not w4944;
w4946 <= not w4938 and w4945;
w4947 <= not pi0100 and w898;
w4948 <= pi0039 and not w4947;
w4949 <= not pi0038 and not w4948;
w4950 <= not w4946 and w4949;
w4951 <= not w4 and not w4950;
w4952 <= not pi0087 and not w4951;
w4953 <= not pi0075 and not w4937;
w4954 <= not w4952 and w4953;
w4955 <= not pi0092 and not w4935;
w4956 <= not w4954 and w4955;
w4957 <= w95 and not w4934;
w4958 <= not w4956 and w4957;
w4959 <= not pi0055 and not w4931;
w4960 <= not w4958 and w4959;
w4961 <= not pi0056 and not w4930;
w4962 <= not w4960 and w4961;
w4963 <= not pi0062 and not w4925;
w4964 <= not w4962 and w4963;
w4965 <= not w4922 and not w4964;
w4966 <= w891 and not w4965;
w4967 <= w4 and not w891;
w4968 <= not w4966 and not w4967;
w4969 <= pi0119 and pi1056;
w4970 <= not pi0228 and pi0252;
w4971 <= not pi0119 and not w4970;
w4972 <= not pi0468 and not w4971;
w4973 <= not w4969 and w4972;
w4974 <= pi0119 and pi1077;
w4975 <= w4972 and not w4974;
w4976 <= pi0119 and pi1073;
w4977 <= w4972 and not w4976;
w4978 <= pi0119 and pi1041;
w4979 <= w4972 and not w4978;
w4980 <= pi0824 and w495;
w4981 <= not pi0122 and pi1093;
w4982 <= w4980 and w4981;
w4983 <= not pi1091 and w4982;
w4984 <= not pi0098 and w4983;
w4985 <= pi0567 and w4984;
w4986 <= not pi0285 and not pi0286;
w4987 <= not pi0289 and w4986;
w4988 <= not pi0288 and w4987;
w4989 <= not pi0057 and w3868;
w4990 <= not w4988 and not w4989;
w4991 <= w4985 and w4990;
w4992 <= not pi0074 and w3697;
w4993 <= not pi0122 and pi0829;
w4994 <= w524 and not w3720;
w4995 <= not pi0841 and w266;
w4996 <= pi0090 and w4995;
w4997 <= not pi0093 and not w4996;
w4998 <= w4994 and not w4997;
w4999 <= not pi0051 and not w4998;
w5000 <= not pi0088 and pi0098;
w5001 <= not pi0050 and not pi0077;
w5002 <= not pi0094 and w5001;
w5003 <= w330 and w5002;
w5004 <= w58 and w5000;
w5005 <= w5003 and w5004;
w5006 <= not pi0097 and not w5005;
w5007 <= w280 and not w5006;
w5008 <= not pi0035 and w267;
w5009 <= not pi0070 and w5008;
w5010 <= w5007 and w5009;
w5011 <= w4999 and not w5010;
w5012 <= not w310 and not w5011;
w5013 <= not pi0096 and w82;
w5014 <= w5012 and w5013;
w5015 <= w3840 and w5014;
w5016 <= not w4993 and w5015;
w5017 <= not pi0096 and not w5012;
w5018 <= pi0096 and not w4047;
w5019 <= w82 and not w5018;
w5020 <= w495 and w4993;
w5021 <= w5019 and w5020;
w5022 <= not w5017 and w5021;
w5023 <= not w5016 and not w5022;
w5024 <= not pi1093 and not w5023;
w5025 <= not pi0087 and not w5024;
w5026 <= w84 and w3841;
w5027 <= pi0087 and not w5026;
w5028 <= not pi0075 and w94;
w5029 <= not w5027 and w5028;
w5030 <= not w5025 and w5029;
w5031 <= not pi0567 and not w5030;
w5032 <= w4992 and not w5031;
w5033 <= not pi0299 and not w232;
w5034 <= pi0299 and not w202;
w5035 <= not w5033 and not w5034;
w5036 <= pi0232 and w3760;
w5037 <= w5035 and w5036;
w5038 <= w173 and not w5037;
w5039 <= w4984 and not w5038;
w5040 <= not pi0024 and w3922;
w5041 <= not w486 and not w3837;
w5042 <= pi1093 and w5020;
w5043 <= w5041 and w5042;
w5044 <= w5040 and w5043;
w5045 <= pi1091 and not w5044;
w5046 <= w5038 and not w5045;
w5047 <= not pi0098 and w4980;
w5048 <= w4981 and w5047;
w5049 <= not pi1091 and not w5048;
w5050 <= w5046 and not w5049;
w5051 <= pi0075 and not w5039;
w5052 <= not w5050 and w5051;
w5053 <= pi1093 and w486;
w5054 <= w3840 and not w5053;
w5055 <= w84 and w5054;
w5056 <= pi1091 and not w5055;
w5057 <= not pi1091 and not w5026;
w5058 <= w84 and w4980;
w5059 <= pi0122 and w5058;
w5060 <= not pi0122 and w5047;
w5061 <= not w5059 and not w5060;
w5062 <= pi1093 and not w5061;
w5063 <= w5057 and not w5062;
w5064 <= w188 and not w5056;
w5065 <= not w5063 and w5064;
w5066 <= not w4984 and not w5065;
w5067 <= pi0087 and not w5066;
w5068 <= not w93 and w4984;
w5069 <= pi0228 and not w5037;
w5070 <= not w4984 and not w5069;
w5071 <= w84 and w5043;
w5072 <= pi1091 and not w5071;
w5073 <= not w5049 and not w5072;
w5074 <= w5069 and not w5073;
w5075 <= w93 and not w5070;
w5076 <= not w5074 and w5075;
w5077 <= pi0100 and not w5068;
w5078 <= not w5076 and w5077;
w5079 <= pi0038 and w4984;
w5080 <= pi1093 and not w486;
w5081 <= not w310 and w5013;
w5082 <= not w4999 and w5081;
w5083 <= w4980 and w5082;
w5084 <= not pi0829 and w5083;
w5085 <= not pi0024 and w319;
w5086 <= not pi0046 and pi0097;
w5087 <= not pi0108 and w5086;
w5088 <= w4054 and w5087;
w5089 <= w335 and w5088;
w5090 <= not pi0091 and w5089;
w5091 <= not w5085 and not w5090;
w5092 <= w24 and w4994;
w5093 <= not w5091 and w5092;
w5094 <= w4999 and not w5093;
w5095 <= not w310 and not w5094;
w5096 <= not pi0096 and not w5095;
w5097 <= w496 and w5019;
w5098 <= not w5096 and w5097;
w5099 <= not w5084 and not w5098;
w5100 <= not pi0122 and not w5099;
w5101 <= pi0122 and w3840;
w5102 <= w5082 and w5101;
w5103 <= not w5100 and not w5102;
w5104 <= w5080 and not w5103;
w5105 <= pi1091 and not w5104;
w5106 <= not w5024 and w5105;
w5107 <= not pi0039 and not w5106;
w5108 <= not pi1091 and not w5024;
w5109 <= pi0122 and w5083;
w5110 <= not w5060 and not w5109;
w5111 <= pi1093 and not w5110;
w5112 <= w5108 and not w5111;
w5113 <= w5107 and not w5112;
w5114 <= not pi0223 and w3373;
w5115 <= w4984 and not w5114;
w5116 <= not w486 and w488;
w5117 <= w3945 and w5116;
w5118 <= w489 and w5117;
w5119 <= pi1091 and not w5118;
w5120 <= not w5049 and not w5119;
w5121 <= w3761 and w5120;
w5122 <= not w3761 and w4984;
w5123 <= not w5121 and not w5122;
w5124 <= w3768 and w5123;
w5125 <= not w3790 and w5120;
w5126 <= w3790 and w4984;
w5127 <= not w5125 and not w5126;
w5128 <= not w3768 and w5127;
w5129 <= w5114 and not w5124;
w5130 <= not w5128 and w5129;
w5131 <= not pi0299 and not w5115;
w5132 <= not w5130 and w5131;
w5133 <= not pi0216 and w3942;
w5134 <= w4984 and not w5133;
w5135 <= w3805 and w5123;
w5136 <= not w3805 and w5127;
w5137 <= w5133 and not w5135;
w5138 <= not w5136 and w5137;
w5139 <= pi0299 and not w5134;
w5140 <= not w5138 and w5139;
w5141 <= pi0039 and not w5132;
w5142 <= not w5140 and w5141;
w5143 <= not w5113 and not w5142;
w5144 <= not pi0038 and not w5143;
w5145 <= not pi0100 and not w5079;
w5146 <= not w5144 and w5145;
w5147 <= not pi0087 and not w5078;
w5148 <= not w5146 and w5147;
w5149 <= not pi0075 and not w5067;
w5150 <= not w5148 and w5149;
w5151 <= not w5052 and not w5150;
w5152 <= pi0567 and not w5151;
w5153 <= w5032 and not w5152;
w5154 <= w4985 and not w4992;
w5155 <= not w5153 and not w5154;
w5156 <= not w4988 and w5155;
w5157 <= pi1091 and w5041;
w5158 <= w5020 and w5157;
w5159 <= w5040 and w5158;
w5160 <= pi1093 and w5159;
w5161 <= w5038 and w5160;
w5162 <= pi0075 and not w5161;
w5163 <= not w5106 and not w5108;
w5164 <= not pi0039 and not w5163;
w5165 <= pi1091 and w5118;
w5166 <= not w3807 and w5165;
w5167 <= not pi0216 and w4203;
w5168 <= w5166 and w5167;
w5169 <= not w3770 and w5165;
w5170 <= not pi0299 and w3968;
w5171 <= not pi0224 and w5170;
w5172 <= w5169 and w5171;
w5173 <= pi0039 and not w5168;
w5174 <= not w5172 and w5173;
w5175 <= not pi0038 and not w5174;
w5176 <= not w5164 and w5175;
w5177 <= not pi0100 and not w5176;
w5178 <= w3947 and w5082;
w5179 <= w5175 and w5178;
w5180 <= not w5105 and w5179;
w5181 <= w5177 and not w5180;
w5182 <= pi1091 and w5071;
w5183 <= pi0228 and w5182;
w5184 <= w93 and not w5037;
w5185 <= w5183 and w5184;
w5186 <= pi0100 and not w5185;
w5187 <= not w5181 and not w5186;
w5188 <= not pi0087 and not w5187;
w5189 <= not pi1091 and pi1093;
w5190 <= not w5058 and w5189;
w5191 <= not w5055 and not w5189;
w5192 <= w188 and not w5191;
w5193 <= not w5190 and w5192;
w5194 <= pi0087 and not w5193;
w5195 <= not w5188 and not w5194;
w5196 <= not pi0075 and not w5195;
w5197 <= not w5162 and not w5196;
w5198 <= pi0567 and not w5197;
w5199 <= w5032 and not w5198;
w5200 <= w4988 and not w5199;
w5201 <= w4989 and not w5156;
w5202 <= not w5200 and w5201;
w5203 <= pi0217 and not w4991;
w5204 <= not w5202 and w5203;
w5205 <= not pi1161 and not pi1162;
w5206 <= not pi1163 and w5205;
w5207 <= not pi0592 and w4985;
w5208 <= pi0592 and w4985;
w5209 <= not pi0363 and not pi0372;
w5210 <= pi0363 and pi0372;
w5211 <= not w5209 and not w5210;
w5212 <= pi0386 and not w5211;
w5213 <= not pi0386 and w5211;
w5214 <= not w5212 and not w5213;
w5215 <= pi0338 and not pi0388;
w5216 <= not pi0338 and pi0388;
w5217 <= not w5215 and not w5216;
w5218 <= pi0337 and not pi0339;
w5219 <= not pi0337 and pi0339;
w5220 <= not w5218 and not w5219;
w5221 <= pi0387 and w5220;
w5222 <= not pi0387 and not w5220;
w5223 <= not w5221 and not w5222;
w5224 <= pi0380 and not w5223;
w5225 <= not pi0380 and w5223;
w5226 <= not w5224 and not w5225;
w5227 <= w5217 and not w5226;
w5228 <= not w5217 and w5226;
w5229 <= not w5227 and not w5228;
w5230 <= w5214 and w5229;
w5231 <= not w5214 and not w5229;
w5232 <= not w5230 and not w5231;
w5233 <= pi1196 and not w5232;
w5234 <= not pi0368 and not pi0389;
w5235 <= pi0368 and pi0389;
w5236 <= not w5234 and not w5235;
w5237 <= pi0365 and not pi0447;
w5238 <= not pi0365 and pi0447;
w5239 <= not w5237 and not w5238;
w5240 <= pi0336 and not pi0383;
w5241 <= not pi0336 and pi0383;
w5242 <= not w5240 and not w5241;
w5243 <= pi0364 and not pi0366;
w5244 <= not pi0364 and pi0366;
w5245 <= not w5243 and not w5244;
w5246 <= w5242 and w5245;
w5247 <= not w5242 and not w5245;
w5248 <= not w5246 and not w5247;
w5249 <= w5239 and w5248;
w5250 <= not w5239 and not w5248;
w5251 <= not w5249 and not w5250;
w5252 <= pi0367 and not w5251;
w5253 <= not pi0367 and w5251;
w5254 <= not w5252 and not w5253;
w5255 <= w5236 and w5254;
w5256 <= not w5236 and not w5254;
w5257 <= pi1197 and not w5255;
w5258 <= not w5256 and w5257;
w5259 <= not w5233 and not w5258;
w5260 <= pi0592 and not w5259;
w5261 <= pi0379 and not pi0382;
w5262 <= not pi0379 and pi0382;
w5263 <= not w5261 and not w5262;
w5264 <= pi0376 and not pi0439;
w5265 <= not pi0376 and pi0439;
w5266 <= not w5264 and not w5265;
w5267 <= pi0381 and w5266;
w5268 <= not pi0381 and not w5266;
w5269 <= not w5267 and not w5268;
w5270 <= pi0317 and not pi0385;
w5271 <= not pi0317 and pi0385;
w5272 <= not w5270 and not w5271;
w5273 <= pi0378 and w5272;
w5274 <= not pi0378 and not w5272;
w5275 <= not w5273 and not w5274;
w5276 <= w5269 and not w5275;
w5277 <= not w5269 and w5275;
w5278 <= not w5276 and not w5277;
w5279 <= w5263 and w5278;
w5280 <= not w5263 and not w5278;
w5281 <= not w5279 and not w5280;
w5282 <= not pi0377 and not w5281;
w5283 <= pi0377 and w5281;
w5284 <= not w5282 and not w5283;
w5285 <= w5259 and not w5284;
w5286 <= pi0592 and not w5285;
w5287 <= w4985 and not w5286;
w5288 <= pi1199 and not w5287;
w5289 <= not w5260 and not w5288;
w5290 <= w5208 and w5289;
w5291 <= not pi1198 and w5290;
w5292 <= pi0384 and not pi0442;
w5293 <= not pi0384 and pi0442;
w5294 <= not w5292 and not w5293;
w5295 <= pi0440 and not w5294;
w5296 <= not pi0440 and w5294;
w5297 <= not w5295 and not w5296;
w5298 <= not pi0369 and not pi0374;
w5299 <= pi0369 and pi0374;
w5300 <= not w5298 and not w5299;
w5301 <= not pi0370 and not w5300;
w5302 <= pi0370 and w5300;
w5303 <= not w5301 and not w5302;
w5304 <= not pi0371 and not w5303;
w5305 <= pi0371 and w5303;
w5306 <= not w5304 and not w5305;
w5307 <= not pi0373 and not w5306;
w5308 <= pi0373 and w5306;
w5309 <= not w5307 and not w5308;
w5310 <= pi0375 and not w5309;
w5311 <= not pi0375 and w5309;
w5312 <= not w5310 and not w5311;
w5313 <= not w5297 and not w5312;
w5314 <= w5297 and w5312;
w5315 <= not w5313 and not w5314;
w5316 <= w5290 and w5315;
w5317 <= not w5207 and not w5291;
w5318 <= not w5316 and w5317;
w5319 <= not pi0590 and not w5318;
w5320 <= pi0351 and pi1199;
w5321 <= pi0345 and not pi0346;
w5322 <= not pi0345 and pi0346;
w5323 <= not w5321 and not w5322;
w5324 <= pi0323 and not w5323;
w5325 <= not pi0323 and w5323;
w5326 <= not w5324 and not w5325;
w5327 <= pi0358 and not pi0450;
w5328 <= not pi0358 and pi0450;
w5329 <= not w5327 and not w5328;
w5330 <= w5326 and not w5329;
w5331 <= not w5326 and w5329;
w5332 <= not w5330 and not w5331;
w5333 <= not pi0327 and not pi0362;
w5334 <= pi0327 and pi0362;
w5335 <= not w5333 and not w5334;
w5336 <= pi0343 and not pi0344;
w5337 <= not pi0343 and pi0344;
w5338 <= not w5336 and not w5337;
w5339 <= w5335 and not w5338;
w5340 <= not w5335 and w5338;
w5341 <= not w5339 and not w5340;
w5342 <= w5332 and w5341;
w5343 <= not w5332 and not w5341;
w5344 <= pi1197 and not w5342;
w5345 <= not w5343 and w5344;
w5346 <= pi0320 and not pi0460;
w5347 <= not pi0320 and pi0460;
w5348 <= not w5346 and not w5347;
w5349 <= pi0342 and not w5348;
w5350 <= not pi0342 and w5348;
w5351 <= not w5349 and not w5350;
w5352 <= pi0452 and not pi0455;
w5353 <= not pi0452 and pi0455;
w5354 <= not w5352 and not w5353;
w5355 <= pi0355 and w5354;
w5356 <= not pi0355 and not w5354;
w5357 <= not w5355 and not w5356;
w5358 <= pi0361 and not pi0458;
w5359 <= not pi0361 and pi0458;
w5360 <= not w5358 and not w5359;
w5361 <= w5357 and w5360;
w5362 <= not w5357 and not w5360;
w5363 <= not w5361 and not w5362;
w5364 <= not pi0441 and w5363;
w5365 <= pi0441 and not w5363;
w5366 <= not pi0592 and not w5364;
w5367 <= not w5365 and w5366;
w5368 <= w4985 and w5351;
w5369 <= not w5367 and w5368;
w5370 <= pi0361 and not pi0441;
w5371 <= not pi0361 and pi0441;
w5372 <= not w5370 and not w5371;
w5373 <= w5351 and w5372;
w5374 <= not w5351 and not w5372;
w5375 <= not w5373 and not w5374;
w5376 <= pi0458 and w5375;
w5377 <= not pi0458 and not w5375;
w5378 <= not w5376 and not w5377;
w5379 <= w5357 and w5378;
w5380 <= not w5357 and not w5378;
w5381 <= not w5379 and not w5380;
w5382 <= not pi0592 and w5381;
w5383 <= w4985 and not w5351;
w5384 <= not w5382 and w5383;
w5385 <= pi1196 and not w5369;
w5386 <= not w5384 and w5385;
w5387 <= not pi1198 and not w5386;
w5388 <= pi1196 and w5381;
w5389 <= pi0321 and not pi0347;
w5390 <= not pi0321 and pi0347;
w5391 <= not w5389 and not w5390;
w5392 <= pi0316 and not pi0349;
w5393 <= not pi0316 and pi0349;
w5394 <= not w5392 and not w5393;
w5395 <= pi0348 and w5394;
w5396 <= not pi0348 and not w5394;
w5397 <= not w5395 and not w5396;
w5398 <= pi0315 and not pi0359;
w5399 <= not pi0315 and pi0359;
w5400 <= not w5398 and not w5399;
w5401 <= pi0322 and w5400;
w5402 <= not pi0322 and not w5400;
w5403 <= not w5401 and not w5402;
w5404 <= w5397 and not w5403;
w5405 <= not w5397 and w5403;
w5406 <= not w5404 and not w5405;
w5407 <= w5391 and w5406;
w5408 <= not w5391 and not w5406;
w5409 <= not w5407 and not w5408;
w5410 <= pi0350 and not w5409;
w5411 <= not pi0350 and w5409;
w5412 <= not w5410 and not w5411;
w5413 <= not w5388 and w5412;
w5414 <= pi1198 and w5207;
w5415 <= w5413 and w5414;
w5416 <= not w5387 and not w5415;
w5417 <= not w5345 and not w5416;
w5418 <= not pi0592 and not w5417;
w5419 <= w4985 and not w5418;
w5420 <= not w5320 and not w5419;
w5421 <= pi1199 and not w5208;
w5422 <= pi0351 and w5421;
w5423 <= not w5420 and not w5422;
w5424 <= not pi0461 and not w5423;
w5425 <= not pi0351 and pi1199;
w5426 <= not w5419 and not w5425;
w5427 <= not pi0351 and w5421;
w5428 <= not w5426 and not w5427;
w5429 <= pi0461 and not w5428;
w5430 <= not w5424 and not w5429;
w5431 <= not pi0357 and not w5430;
w5432 <= not pi0461 and not w5428;
w5433 <= pi0461 and not w5423;
w5434 <= not w5432 and not w5433;
w5435 <= pi0357 and not w5434;
w5436 <= not w5431 and not w5435;
w5437 <= not pi0356 and not w5436;
w5438 <= not pi0357 and not w5434;
w5439 <= pi0357 and not w5430;
w5440 <= not w5438 and not w5439;
w5441 <= pi0356 and not w5440;
w5442 <= pi0360 and not pi0462;
w5443 <= not pi0360 and pi0462;
w5444 <= not w5442 and not w5443;
w5445 <= pi0352 and not pi0353;
w5446 <= not pi0352 and pi0353;
w5447 <= not w5445 and not w5446;
w5448 <= w5444 and w5447;
w5449 <= not w5444 and not w5447;
w5450 <= not w5448 and not w5449;
w5451 <= pi0354 and not w5450;
w5452 <= not pi0354 and w5450;
w5453 <= not w5451 and not w5452;
w5454 <= not w5437 and w5453;
w5455 <= not w5441 and w5454;
w5456 <= not pi0356 and not w5440;
w5457 <= pi0356 and not w5436;
w5458 <= not w5453 and not w5456;
w5459 <= not w5457 and w5458;
w5460 <= not w5455 and not w5459;
w5461 <= pi0590 and not w5460;
w5462 <= not pi0591 and not w5319;
w5463 <= not w5461 and w5462;
w5464 <= pi0590 and w4985;
w5465 <= pi1197 and not w5208;
w5466 <= pi0318 and not pi0409;
w5467 <= not pi0318 and pi0409;
w5468 <= not w5466 and not w5467;
w5469 <= pi0401 and not pi0402;
w5470 <= not pi0401 and pi0402;
w5471 <= not w5469 and not w5470;
w5472 <= pi0406 and w5471;
w5473 <= not pi0406 and not w5471;
w5474 <= not w5472 and not w5473;
w5475 <= not pi0403 and not pi0405;
w5476 <= pi0403 and pi0405;
w5477 <= not w5475 and not w5476;
w5478 <= pi0325 and not pi0326;
w5479 <= not pi0325 and pi0326;
w5480 <= not w5478 and not w5479;
w5481 <= w5477 and w5480;
w5482 <= not w5477 and not w5480;
w5483 <= not w5481 and not w5482;
w5484 <= w5474 and not w5483;
w5485 <= not w5474 and w5483;
w5486 <= not w5484 and not w5485;
w5487 <= w5468 and w5486;
w5488 <= not w5468 and not w5486;
w5489 <= not w5487 and not w5488;
w5490 <= w5048 and not w5489;
w5491 <= not pi1091 and w5490;
w5492 <= pi0567 and w5491;
w5493 <= pi0390 and not pi0410;
w5494 <= not pi0390 and pi0410;
w5495 <= not w5493 and not w5494;
w5496 <= pi0397 and not pi0412;
w5497 <= not pi0397 and pi0412;
w5498 <= not w5496 and not w5497;
w5499 <= pi0404 and w5498;
w5500 <= not pi0404 and not w5498;
w5501 <= not w5499 and not w5500;
w5502 <= pi0319 and not pi0324;
w5503 <= not pi0319 and pi0324;
w5504 <= not w5502 and not w5503;
w5505 <= pi0456 and not w5504;
w5506 <= not pi0456 and w5504;
w5507 <= not w5505 and not w5506;
w5508 <= w5501 and not w5507;
w5509 <= not w5501 and w5507;
w5510 <= not w5508 and not w5509;
w5511 <= w5495 and w5510;
w5512 <= not w5495 and not w5510;
w5513 <= not w5511 and not w5512;
w5514 <= pi0411 and w5513;
w5515 <= not pi0411 and not w5513;
w5516 <= not w5514 and not w5515;
w5517 <= pi1196 and not w5516;
w5518 <= not pi0592 and w5492;
w5519 <= not w5517 and w5518;
w5520 <= w5421 and not w5519;
w5521 <= not pi0592 and pi1196;
w5522 <= w4985 and not w5521;
w5523 <= w5048 and w5516;
w5524 <= not pi1091 and w5523;
w5525 <= pi0567 and w5524;
w5526 <= w5521 and w5525;
w5527 <= not pi1199 and not w5522;
w5528 <= not w5526 and w5527;
w5529 <= not w5520 and not w5528;
w5530 <= not pi1197 and not w5529;
w5531 <= not w5465 and not w5530;
w5532 <= pi0333 and not w5531;
w5533 <= pi1198 and not w5208;
w5534 <= w5529 and not w5533;
w5535 <= pi0328 and not pi0408;
w5536 <= not pi0328 and pi0408;
w5537 <= not w5535 and not w5536;
w5538 <= not pi0394 and not pi0396;
w5539 <= pi0394 and pi0396;
w5540 <= not w5538 and not w5539;
w5541 <= w5537 and not w5540;
w5542 <= not w5537 and w5540;
w5543 <= not w5541 and not w5542;
w5544 <= pi0398 and not pi0399;
w5545 <= not pi0398 and pi0399;
w5546 <= not w5544 and not w5545;
w5547 <= pi0395 and w5546;
w5548 <= not pi0395 and not w5546;
w5549 <= not w5547 and not w5548;
w5550 <= pi0329 and not w5549;
w5551 <= not pi0329 and w5549;
w5552 <= not w5550 and not w5551;
w5553 <= pi0400 and not w5552;
w5554 <= not pi0400 and w5552;
w5555 <= not w5553 and not w5554;
w5556 <= w5543 and w5555;
w5557 <= not w5543 and not w5555;
w5558 <= not w5556 and not w5557;
w5559 <= not w5534 and not w5558;
w5560 <= not pi0333 and not w5529;
w5561 <= not w5559 and not w5560;
w5562 <= not w5532 and w5561;
w5563 <= not pi0391 and not w5562;
w5564 <= not pi0333 and not w5531;
w5565 <= w5529 and not w5559;
w5566 <= not w5564 and w5565;
w5567 <= pi0391 and not w5566;
w5568 <= not w5563 and not w5567;
w5569 <= not pi0392 and not w5568;
w5570 <= not pi0391 and not w5566;
w5571 <= pi0391 and not w5562;
w5572 <= not w5570 and not w5571;
w5573 <= pi0392 and not w5572;
w5574 <= not w5569 and not w5573;
w5575 <= not pi0393 and not w5574;
w5576 <= not pi0392 and not w5572;
w5577 <= pi0392 and not w5568;
w5578 <= not w5576 and not w5577;
w5579 <= pi0393 and not w5578;
w5580 <= pi0407 and not pi0463;
w5581 <= not pi0407 and pi0463;
w5582 <= not w5580 and not w5581;
w5583 <= pi0335 and not pi0413;
w5584 <= not pi0335 and pi0413;
w5585 <= not w5583 and not w5584;
w5586 <= w5582 and w5585;
w5587 <= not w5582 and not w5585;
w5588 <= not w5586 and not w5587;
w5589 <= pi0334 and not w5588;
w5590 <= not pi0334 and w5588;
w5591 <= not w5589 and not w5590;
w5592 <= not w5575 and w5591;
w5593 <= not w5579 and w5592;
w5594 <= not pi0393 and not w5578;
w5595 <= pi0393 and not w5574;
w5596 <= not w5591 and not w5594;
w5597 <= not w5595 and w5596;
w5598 <= not w5593 and not w5597;
w5599 <= not pi0590 and not w5598;
w5600 <= pi0591 and not w5464;
w5601 <= not w5599 and w5600;
w5602 <= not w5463 and not w5601;
w5603 <= not pi0588 and not w5602;
w5604 <= not pi0590 and not pi0591;
w5605 <= w4985 and not w5604;
w5606 <= not pi0417 and not pi0418;
w5607 <= pi0417 and pi0418;
w5608 <= not w5606 and not w5607;
w5609 <= pi0437 and w5608;
w5610 <= not pi0437 and not w5608;
w5611 <= not w5609 and not w5610;
w5612 <= pi0453 and not pi0464;
w5613 <= not pi0453 and pi0464;
w5614 <= not w5612 and not w5613;
w5615 <= w5611 and w5614;
w5616 <= not w5611 and not w5614;
w5617 <= not w5615 and not w5616;
w5618 <= pi0415 and not pi0431;
w5619 <= not pi0415 and pi0431;
w5620 <= not w5618 and not w5619;
w5621 <= pi0416 and not pi0438;
w5622 <= not pi0416 and pi0438;
w5623 <= not w5621 and not w5622;
w5624 <= w5620 and w5623;
w5625 <= not w5620 and not w5623;
w5626 <= not w5624 and not w5625;
w5627 <= w5617 and not w5626;
w5628 <= not w5617 and w5626;
w5629 <= pi1197 and not w5627;
w5630 <= not w5628 and w5629;
w5631 <= pi0421 and not pi0454;
w5632 <= not pi0421 and pi0454;
w5633 <= not w5631 and not w5632;
w5634 <= pi0432 and not pi0459;
w5635 <= not pi0432 and pi0459;
w5636 <= not w5634 and not w5635;
w5637 <= w5633 and not w5636;
w5638 <= not w5633 and w5636;
w5639 <= not w5637 and not w5638;
w5640 <= not pi0419 and not pi0420;
w5641 <= pi0419 and pi0420;
w5642 <= not w5640 and not w5641;
w5643 <= pi0423 and not pi0424;
w5644 <= not pi0423 and pi0424;
w5645 <= not w5643 and not w5644;
w5646 <= w5642 and not w5645;
w5647 <= not w5642 and w5645;
w5648 <= not w5646 and not w5647;
w5649 <= w5639 and w5648;
w5650 <= not w5639 and not w5648;
w5651 <= not w5649 and not w5650;
w5652 <= pi0425 and not w5651;
w5653 <= not pi0425 and w5651;
w5654 <= pi1198 and not w5652;
w5655 <= not w5653 and w5654;
w5656 <= not w5630 and not w5655;
w5657 <= not pi0429 and not pi0435;
w5658 <= pi0429 and pi0435;
w5659 <= not w5657 and not w5658;
w5660 <= pi0434 and not pi0446;
w5661 <= not pi0434 and pi0446;
w5662 <= not w5660 and not w5661;
w5663 <= pi0414 and not pi0422;
w5664 <= not pi0414 and pi0422;
w5665 <= not w5663 and not w5664;
w5666 <= w5662 and w5665;
w5667 <= not w5662 and not w5665;
w5668 <= not w5666 and not w5667;
w5669 <= w5659 and w5668;
w5670 <= not w5659 and not w5668;
w5671 <= not w5669 and not w5670;
w5672 <= pi0436 and not pi0443;
w5673 <= not pi0436 and pi0443;
w5674 <= not w5672 and not w5673;
w5675 <= not pi0444 and w5674;
w5676 <= pi0444 and not w5674;
w5677 <= not w5675 and not w5676;
w5678 <= not w5671 and not w5677;
w5679 <= w5671 and w5677;
w5680 <= w5521 and not w5678;
w5681 <= not w5679 and w5680;
w5682 <= w5656 and not w5681;
w5683 <= w5207 and w5682;
w5684 <= not pi1199 and not w5208;
w5685 <= not w5683 and w5684;
w5686 <= pi0433 and not pi0451;
w5687 <= not pi0433 and pi0451;
w5688 <= not w5686 and not w5687;
w5689 <= pi0449 and w5688;
w5690 <= not pi0449 and not w5688;
w5691 <= not w5689 and not w5690;
w5692 <= not pi0427 and pi0428;
w5693 <= pi0427 and not pi0428;
w5694 <= not w5692 and not w5693;
w5695 <= pi0430 and not w5694;
w5696 <= not pi0430 and w5694;
w5697 <= not w5695 and not w5696;
w5698 <= not pi0426 and not w5697;
w5699 <= pi0426 and w5697;
w5700 <= not w5698 and not w5699;
w5701 <= not pi0445 and not w5700;
w5702 <= pi0445 and w5700;
w5703 <= not w5701 and not w5702;
w5704 <= not pi0448 and not w5703;
w5705 <= pi0448 and w5703;
w5706 <= not w5704 and not w5705;
w5707 <= w5683 and not w5706;
w5708 <= not w5208 and not w5707;
w5709 <= w5691 and not w5708;
w5710 <= w5683 and w5706;
w5711 <= not w5208 and not w5710;
w5712 <= not w5691 and not w5711;
w5713 <= pi1199 and not w5709;
w5714 <= not w5712 and w5713;
w5715 <= w5604 and not w5685;
w5716 <= not w5714 and w5715;
w5717 <= pi0588 and not w5605;
w5718 <= not w5716 and w5717;
w5719 <= w4990 and not w5718;
w5720 <= not w5603 and w5719;
w5721 <= w5199 and not w5604;
w5722 <= not pi0087 and not w5186;
w5723 <= not w5177 and w5722;
w5724 <= pi0087 and not pi0100;
w5725 <= w93 and w5724;
w5726 <= not w5056 and w5725;
w5727 <= not w5057 and w5726;
w5728 <= not pi0075 and not w5727;
w5729 <= not w5723 and w5728;
w5730 <= not w5162 and not w5729;
w5731 <= pi0567 and not w5730;
w5732 <= w5032 and not w5731;
w5733 <= not pi0592 and not w5732;
w5734 <= pi0592 and not w5199;
w5735 <= not w5733 and not w5734;
w5736 <= not w5656 and w5735;
w5737 <= not pi1196 and not w5199;
w5738 <= not pi0443 and not pi0592;
w5739 <= not w5199 and not w5738;
w5740 <= not w5732 and w5738;
w5741 <= not w5739 and not w5740;
w5742 <= not pi0444 and not w5741;
w5743 <= pi0443 and not pi0592;
w5744 <= not w5199 and not w5743;
w5745 <= not w5732 and w5743;
w5746 <= not w5744 and not w5745;
w5747 <= pi0444 and not w5746;
w5748 <= not w5742 and not w5747;
w5749 <= not pi0436 and not w5748;
w5750 <= not pi0444 and not w5746;
w5751 <= pi0444 and not w5741;
w5752 <= not w5750 and not w5751;
w5753 <= pi0436 and not w5752;
w5754 <= w5671 and not w5749;
w5755 <= not w5753 and w5754;
w5756 <= not pi0436 and not w5752;
w5757 <= pi0436 and not w5748;
w5758 <= not w5671 and not w5756;
w5759 <= not w5757 and w5758;
w5760 <= pi1196 and not w5755;
w5761 <= not w5759 and w5760;
w5762 <= w5656 and not w5737;
w5763 <= not w5761 and w5762;
w5764 <= not w5736 and not w5763;
w5765 <= not pi1199 and w5764;
w5766 <= pi0428 and not w5764;
w5767 <= not pi0428 and w5735;
w5768 <= not w5766 and not w5767;
w5769 <= not pi0427 and not w5768;
w5770 <= not pi0428 and not w5764;
w5771 <= pi0428 and w5735;
w5772 <= not w5770 and not w5771;
w5773 <= pi0427 and not w5772;
w5774 <= not w5769 and not w5773;
w5775 <= pi0430 and not w5774;
w5776 <= not pi0427 and not w5772;
w5777 <= pi0427 and not w5768;
w5778 <= not w5776 and not w5777;
w5779 <= not pi0430 and not w5778;
w5780 <= not w5775 and not w5779;
w5781 <= pi0426 and not w5780;
w5782 <= pi0430 and not w5778;
w5783 <= not pi0430 and not w5774;
w5784 <= not w5782 and not w5783;
w5785 <= not pi0426 and not w5784;
w5786 <= not w5781 and not w5785;
w5787 <= pi0445 and not w5786;
w5788 <= pi0426 and not w5784;
w5789 <= not pi0426 and not w5780;
w5790 <= not w5788 and not w5789;
w5791 <= not pi0445 and not w5790;
w5792 <= not w5787 and not w5791;
w5793 <= pi0448 and not w5691;
w5794 <= not pi0448 and w5691;
w5795 <= not w5793 and not w5794;
w5796 <= not w5792 and not w5795;
w5797 <= pi0445 and not w5790;
w5798 <= not pi0445 and not w5786;
w5799 <= not w5797 and not w5798;
w5800 <= w5795 and not w5799;
w5801 <= pi1199 and not w5796;
w5802 <= not w5800 and w5801;
w5803 <= w5604 and not w5765;
w5804 <= not w5802 and w5803;
w5805 <= w4988 and not w5721;
w5806 <= not w5804 and w5805;
w5807 <= not w5155 and not w5604;
w5808 <= not pi1196 and w5155;
w5809 <= w5155 and not w5738;
w5810 <= not pi0436 and pi0444;
w5811 <= pi0436 and not pi0444;
w5812 <= not w5810 and not w5811;
w5813 <= w5671 and not w5812;
w5814 <= not w5671 and w5812;
w5815 <= not w5813 and not w5814;
w5816 <= not w5740 and w5815;
w5817 <= not w5809 and w5816;
w5818 <= w5155 and not w5743;
w5819 <= not w5745 and not w5815;
w5820 <= not w5818 and w5819;
w5821 <= pi1196 and not w5817;
w5822 <= not w5820 and w5821;
w5823 <= not w5808 and not w5822;
w5824 <= w5656 and not w5823;
w5825 <= pi0592 and w5155;
w5826 <= not w5733 and not w5825;
w5827 <= not w5656 and not w5826;
w5828 <= not w5824 and not w5827;
w5829 <= not pi1199 and not w5828;
w5830 <= not pi0428 and w5826;
w5831 <= pi0428 and w5828;
w5832 <= pi0427 and not w5830;
w5833 <= not w5831 and w5832;
w5834 <= not pi0428 and w5828;
w5835 <= pi0428 and w5826;
w5836 <= not pi0427 and not w5835;
w5837 <= not w5834 and w5836;
w5838 <= not w5833 and not w5837;
w5839 <= not pi0430 and not w5838;
w5840 <= w5694 and w5826;
w5841 <= not w5694 and w5828;
w5842 <= not w5840 and not w5841;
w5843 <= pi0430 and w5842;
w5844 <= not w5839 and not w5843;
w5845 <= not pi0426 and not w5844;
w5846 <= pi0430 and not w5838;
w5847 <= not pi0430 and w5842;
w5848 <= not w5846 and not w5847;
w5849 <= pi0426 and not w5848;
w5850 <= not w5845 and not w5849;
w5851 <= not pi0445 and not w5850;
w5852 <= not pi0426 and not w5848;
w5853 <= pi0426 and not w5844;
w5854 <= not w5852 and not w5853;
w5855 <= pi0445 and not w5854;
w5856 <= not w5851 and not w5855;
w5857 <= pi0448 and w5856;
w5858 <= not pi0445 and not w5854;
w5859 <= pi0445 and not w5850;
w5860 <= not w5858 and not w5859;
w5861 <= not pi0448 and w5860;
w5862 <= not w5691 and not w5857;
w5863 <= not w5861 and w5862;
w5864 <= not pi0448 and w5856;
w5865 <= pi0448 and w5860;
w5866 <= w5691 and not w5864;
w5867 <= not w5865 and w5866;
w5868 <= not w5863 and not w5867;
w5869 <= pi1199 and not w5868;
w5870 <= w5604 and not w5829;
w5871 <= not w5869 and w5870;
w5872 <= not w4988 and not w5807;
w5873 <= not w5871 and w5872;
w5874 <= not w5806 and not w5873;
w5875 <= pi0588 and not w5874;
w5876 <= pi0591 and w5199;
w5877 <= w5388 and not w5735;
w5878 <= not pi0350 and not pi0592;
w5879 <= not w5199 and not w5878;
w5880 <= not w5732 and w5878;
w5881 <= w5409 and not w5880;
w5882 <= not w5879 and w5881;
w5883 <= pi0350 and not pi0592;
w5884 <= not w5199 and not w5883;
w5885 <= not w5732 and w5883;
w5886 <= not w5409 and not w5885;
w5887 <= not w5884 and w5886;
w5888 <= not w5388 and not w5882;
w5889 <= not w5887 and w5888;
w5890 <= pi1198 and not w5877;
w5891 <= not w5889 and w5890;
w5892 <= not pi0455 and not w5735;
w5893 <= pi0455 and not w5199;
w5894 <= not w5892 and not w5893;
w5895 <= not pi0452 and not w5894;
w5896 <= pi0455 and not w5735;
w5897 <= not pi0455 and not w5199;
w5898 <= not w5896 and not w5897;
w5899 <= pi0452 and not w5898;
w5900 <= not w5895 and not w5899;
w5901 <= not pi0355 and not w5900;
w5902 <= not pi0452 and not w5898;
w5903 <= pi0452 and not w5894;
w5904 <= not w5902 and not w5903;
w5905 <= pi0355 and not w5904;
w5906 <= not w5901 and not w5905;
w5907 <= pi0458 and not w5906;
w5908 <= not pi0355 and not w5904;
w5909 <= pi0355 and not w5900;
w5910 <= not w5908 and not w5909;
w5911 <= not pi0458 and not w5910;
w5912 <= w5375 and not w5907;
w5913 <= not w5911 and w5912;
w5914 <= pi0458 and not w5910;
w5915 <= not pi0458 and not w5906;
w5916 <= not w5375 and not w5914;
w5917 <= not w5915 and w5916;
w5918 <= pi1196 and not w5913;
w5919 <= not w5917 and w5918;
w5920 <= not pi1198 and not w5737;
w5921 <= not w5919 and w5920;
w5922 <= not w5891 and not w5921;
w5923 <= not w5345 and not w5922;
w5924 <= w5345 and w5735;
w5925 <= not w5923 and not w5924;
w5926 <= not w5425 and w5925;
w5927 <= pi1199 and not w5735;
w5928 <= not pi0351 and w5927;
w5929 <= not w5926 and not w5928;
w5930 <= not pi0461 and not w5929;
w5931 <= not w5320 and w5925;
w5932 <= pi0351 and w5927;
w5933 <= not w5931 and not w5932;
w5934 <= pi0461 and not w5933;
w5935 <= not w5930 and not w5934;
w5936 <= not pi0357 and not w5935;
w5937 <= not pi0461 and not w5933;
w5938 <= pi0461 and not w5929;
w5939 <= not w5937 and not w5938;
w5940 <= pi0357 and not w5939;
w5941 <= not w5936 and not w5940;
w5942 <= not pi0356 and not w5941;
w5943 <= not pi0357 and not w5939;
w5944 <= pi0357 and not w5935;
w5945 <= not w5943 and not w5944;
w5946 <= pi0356 and not w5945;
w5947 <= not w5942 and not w5946;
w5948 <= not w5453 and not w5947;
w5949 <= not pi0356 and not w5945;
w5950 <= pi0356 and not w5941;
w5951 <= not w5949 and not w5950;
w5952 <= w5453 and not w5951;
w5953 <= not pi0591 and not w5948;
w5954 <= not w5952 and w5953;
w5955 <= pi0590 and not w5876;
w5956 <= not w5954 and w5955;
w5957 <= pi1197 and not w5735;
w5958 <= pi1198 and not w5558;
w5959 <= w5735 and w5958;
w5960 <= not pi0075 and w5517;
w5961 <= not w5489 and not w5960;
w5962 <= w5180 and w5961;
w5963 <= w5177 and not w5962;
w5964 <= w5722 and not w5963;
w5965 <= not w5191 and w5725;
w5966 <= w5058 and not w5489;
w5967 <= w5189 and not w5966;
w5968 <= w5965 and not w5967;
w5969 <= not pi1196 and w5968;
w5970 <= w5058 and w5516;
w5971 <= w5189 and not w5970;
w5972 <= w5968 and not w5971;
w5973 <= not pi0075 and not pi0592;
w5974 <= pi1199 and w5973;
w5975 <= not w5969 and w5974;
w5976 <= not w5972 and w5975;
w5977 <= not w5964 and w5976;
w5978 <= not w5197 and not w5973;
w5979 <= w5965 and not w5971;
w5980 <= w5180 and w5516;
w5981 <= w5177 and not w5980;
w5982 <= w5722 and not w5981;
w5983 <= pi1196 and w5973;
w5984 <= not w5979 and w5983;
w5985 <= not w5982 and w5984;
w5986 <= not pi1196 and w5196;
w5987 <= not w5985 and not w5986;
w5988 <= not pi1199 and not w5987;
w5989 <= not w5977 and not w5978;
w5990 <= not w5988 and w5989;
w5991 <= pi0567 and not w5990;
w5992 <= w5032 and not w5958;
w5993 <= not w5991 and w5992;
w5994 <= not w5959 and not w5993;
w5995 <= not pi1197 and w5994;
w5996 <= not w5957 and not w5995;
w5997 <= pi0333 and not w5996;
w5998 <= not pi0333 and w5994;
w5999 <= not w5997 and not w5998;
w6000 <= pi0391 and not w5999;
w6001 <= pi0333 and not w5994;
w6002 <= not pi0333 and w5996;
w6003 <= not w6001 and not w6002;
w6004 <= not pi0391 and w6003;
w6005 <= not w6000 and not w6004;
w6006 <= not pi0392 and not w6005;
w6007 <= not pi0391 and not w5999;
w6008 <= pi0391 and w6003;
w6009 <= not w6007 and not w6008;
w6010 <= pi0392 and not w6009;
w6011 <= not w6006 and not w6010;
w6012 <= not pi0393 and not w6011;
w6013 <= not pi0392 and not w6009;
w6014 <= pi0392 and not w6005;
w6015 <= not w6013 and not w6014;
w6016 <= pi0393 and not w6015;
w6017 <= not w6012 and not w6016;
w6018 <= not pi0334 and w6017;
w6019 <= not pi0393 and not w6015;
w6020 <= pi0393 and not w6011;
w6021 <= not w6019 and not w6020;
w6022 <= pi0334 and w6021;
w6023 <= w5588 and not w6018;
w6024 <= not w6022 and w6023;
w6025 <= not pi0334 and w6021;
w6026 <= pi0334 and w6017;
w6027 <= not w5588 and not w6025;
w6028 <= not w6026 and w6027;
w6029 <= pi0591 and not w6024;
w6030 <= not w6028 and w6029;
w6031 <= pi0377 and pi0592;
w6032 <= not w5199 and not w6031;
w6033 <= not w5732 and w6031;
w6034 <= not w5281 and not w6033;
w6035 <= not w6032 and w6034;
w6036 <= not pi0377 and pi0592;
w6037 <= not w5199 and not w6036;
w6038 <= not w5732 and w6036;
w6039 <= w5281 and not w6038;
w6040 <= not w6037 and w6039;
w6041 <= not w6035 and not w6040;
w6042 <= w5259 and not w6041;
w6043 <= pi0592 and not w5732;
w6044 <= not pi0592 and not w5199;
w6045 <= not w6043 and not w6044;
w6046 <= not w5259 and w6045;
w6047 <= not w6042 and not w6046;
w6048 <= pi1199 and w6047;
w6049 <= w5199 and not w5258;
w6050 <= w5258 and w6045;
w6051 <= not w6049 and not w6050;
w6052 <= w5232 and not w6051;
w6053 <= not pi1196 and not w5258;
w6054 <= w6045 and not w6053;
w6055 <= not pi1196 and w6049;
w6056 <= not w6054 and not w6055;
w6057 <= not w5232 and not w6056;
w6058 <= not pi1199 and not w6052;
w6059 <= not w6057 and w6058;
w6060 <= not w6048 and not w6059;
w6061 <= not pi0374 and not w6060;
w6062 <= not pi1198 and pi1199;
w6063 <= w6047 and w6062;
w6064 <= not pi1198 and w6059;
w6065 <= pi1198 and not w6045;
w6066 <= not w6063 and not w6065;
w6067 <= not w6064 and w6066;
w6068 <= pi0374 and not w6067;
w6069 <= not w6061 and not w6068;
w6070 <= pi0369 and not w6069;
w6071 <= not pi0374 and not w6067;
w6072 <= pi0374 and not w6060;
w6073 <= not w6071 and not w6072;
w6074 <= not pi0369 and not w6073;
w6075 <= not w6070 and not w6074;
w6076 <= not pi0370 and not w6075;
w6077 <= not pi0369 and not w6069;
w6078 <= pi0369 and not w6073;
w6079 <= not w6077 and not w6078;
w6080 <= pi0370 and not w6079;
w6081 <= not w6076 and not w6080;
w6082 <= not pi0371 and not w6081;
w6083 <= not pi0370 and not w6079;
w6084 <= pi0370 and not w6075;
w6085 <= not w6083 and not w6084;
w6086 <= pi0371 and not w6085;
w6087 <= not w6082 and not w6086;
w6088 <= not pi0373 and not w6087;
w6089 <= not pi0371 and not w6085;
w6090 <= pi0371 and not w6081;
w6091 <= not w6089 and not w6090;
w6092 <= pi0373 and not w6091;
w6093 <= not w6088 and not w6092;
w6094 <= not pi0375 and w6093;
w6095 <= not pi0373 and not w6091;
w6096 <= pi0373 and not w6087;
w6097 <= not w6095 and not w6096;
w6098 <= pi0375 and w6097;
w6099 <= w5297 and not w6094;
w6100 <= not w6098 and w6099;
w6101 <= pi0375 and w6093;
w6102 <= not pi0375 and w6097;
w6103 <= not w5297 and not w6101;
w6104 <= not w6102 and w6103;
w6105 <= not pi0591 and not w6100;
w6106 <= not w6104 and w6105;
w6107 <= not pi0590 and not w6030;
w6108 <= not w6106 and w6107;
w6109 <= w4988 and not w6108;
w6110 <= not w5956 and w6109;
w6111 <= pi0591 and not w5155;
w6112 <= w5345 and not w5826;
w6113 <= w5388 and not w5826;
w6114 <= w5155 and not w5883;
w6115 <= w5886 and not w6114;
w6116 <= w5155 and not w5878;
w6117 <= w5881 and not w6116;
w6118 <= not w5388 and not w6115;
w6119 <= not w6117 and w6118;
w6120 <= pi1198 and not w6113;
w6121 <= not w6119 and w6120;
w6122 <= pi0455 and not w5826;
w6123 <= not pi0455 and w5155;
w6124 <= not w6122 and not w6123;
w6125 <= not pi0452 and not w6124;
w6126 <= not pi0455 and not w5826;
w6127 <= pi0455 and w5155;
w6128 <= not w6126 and not w6127;
w6129 <= pi0452 and not w6128;
w6130 <= pi0355 and not w5378;
w6131 <= not pi0355 and w5378;
w6132 <= not w6130 and not w6131;
w6133 <= not w6125 and not w6132;
w6134 <= not w6129 and w6133;
w6135 <= not pi0452 and not w6128;
w6136 <= pi0452 and not w6124;
w6137 <= w6132 and not w6135;
w6138 <= not w6136 and w6137;
w6139 <= pi1196 and not w6134;
w6140 <= not w6138 and w6139;
w6141 <= not pi1198 and not w5808;
w6142 <= not w6140 and w6141;
w6143 <= not w5345 and not w6121;
w6144 <= not w6142 and w6143;
w6145 <= not w6112 and not w6144;
w6146 <= not w5425 and not w6145;
w6147 <= pi1199 and not w5826;
w6148 <= not pi0351 and w6147;
w6149 <= not w6146 and not w6148;
w6150 <= not pi0461 and not w6149;
w6151 <= not w5320 and not w6145;
w6152 <= pi0351 and w6147;
w6153 <= not w6151 and not w6152;
w6154 <= pi0461 and not w6153;
w6155 <= not w6150 and not w6154;
w6156 <= not pi0357 and not w6155;
w6157 <= not pi0461 and not w6153;
w6158 <= pi0461 and not w6149;
w6159 <= not w6157 and not w6158;
w6160 <= pi0357 and not w6159;
w6161 <= not w6156 and not w6160;
w6162 <= not pi0356 and not w6161;
w6163 <= not pi0357 and not w6159;
w6164 <= pi0357 and not w6155;
w6165 <= not w6163 and not w6164;
w6166 <= pi0356 and not w6165;
w6167 <= not w6162 and not w6166;
w6168 <= not w5453 and not w6167;
w6169 <= not pi0356 and not w6165;
w6170 <= pi0356 and not w6161;
w6171 <= not w6169 and not w6170;
w6172 <= w5453 and not w6171;
w6173 <= not pi0591 and not w6168;
w6174 <= not w6172 and w6173;
w6175 <= pi0590 and not w6111;
w6176 <= not w6174 and w6175;
w6177 <= not w4992 and w5525;
w6178 <= pi0038 and w5524;
w6179 <= not pi0100 and not w6178;
w6180 <= w5108 and not w5516;
w6181 <= w5113 and not w6180;
w6182 <= not w5133 and w5524;
w6183 <= pi0299 and not w6182;
w6184 <= not w3790 and w5165;
w6185 <= not w5524 and not w6184;
w6186 <= not w3805 and w6185;
w6187 <= w3761 and w5165;
w6188 <= not w5524 and not w6187;
w6189 <= w3805 and w6188;
w6190 <= w5133 and not w6186;
w6191 <= not w6189 and w6190;
w6192 <= w6183 and not w6191;
w6193 <= not w5114 and w5524;
w6194 <= not pi0299 and not w6193;
w6195 <= not w3768 and w6185;
w6196 <= w3768 and w6188;
w6197 <= w5114 and not w6195;
w6198 <= not w6196 and w6197;
w6199 <= w6194 and not w6198;
w6200 <= pi0039 and not w6192;
w6201 <= not w6199 and w6200;
w6202 <= not w6181 and not w6201;
w6203 <= not pi0038 and not w6202;
w6204 <= w6179 and not w6203;
w6205 <= w5186 and not w5524;
w6206 <= not w6204 and not w6205;
w6207 <= not pi0087 and not w6206;
w6208 <= not w188 and w5524;
w6209 <= pi0087 and not w6208;
w6210 <= w5057 and not w5516;
w6211 <= w5065 and not w6210;
w6212 <= w6209 and not w6211;
w6213 <= not w6207 and not w6212;
w6214 <= not pi0075 and not w6213;
w6215 <= not w5038 and w5524;
w6216 <= pi0075 and not w6215;
w6217 <= not pi1091 and not w5523;
w6218 <= w5046 and not w6217;
w6219 <= w6216 and not w6218;
w6220 <= not w6214 and not w6219;
w6221 <= pi0567 and not w6220;
w6222 <= w5032 and not w6221;
w6223 <= w5521 and not w6177;
w6224 <= not w6222 and w6223;
w6225 <= not pi1199 and not w5808;
w6226 <= not w6224 and w6225;
w6227 <= w5047 and not w5489;
w6228 <= w6177 and w6227;
w6229 <= w5521 and not w6228;
w6230 <= not w4992 and w5492;
w6231 <= not pi0592 and not pi1196;
w6232 <= not w6230 and w6231;
w6233 <= not w6229 and not w6232;
w6234 <= not w5032 and not w6233;
w6235 <= not w5133 and w5491;
w6236 <= pi0299 and not w6235;
w6237 <= not w6183 and not w6236;
w6238 <= not w5489 and w5524;
w6239 <= not w6187 and not w6238;
w6240 <= w3805 and w6239;
w6241 <= not w6184 and not w6238;
w6242 <= not w3805 and w6241;
w6243 <= w5133 and not w6240;
w6244 <= not w6242 and w6243;
w6245 <= not w6237 and not w6244;
w6246 <= not w5114 and w5491;
w6247 <= not pi0299 and not w6246;
w6248 <= not w6194 and not w6247;
w6249 <= w3768 and w6239;
w6250 <= not w3768 and w6241;
w6251 <= w5114 and not w6249;
w6252 <= not w6250 and w6251;
w6253 <= not w6248 and not w6252;
w6254 <= pi0039 and not w6245;
w6255 <= not w6253 and w6254;
w6256 <= w5083 and not w5489;
w6257 <= pi0122 and not w6256;
w6258 <= not pi0122 and not w6227;
w6259 <= pi1093 and not w6258;
w6260 <= not w6257 and w6259;
w6261 <= w5108 and not w6260;
w6262 <= w6181 and not w6261;
w6263 <= not w6255 and not w6262;
w6264 <= not pi0038 and not w6263;
w6265 <= pi0038 and w5491;
w6266 <= not pi0100 and not w6265;
w6267 <= not w6179 and not w6266;
w6268 <= not w6264 and not w6267;
w6269 <= not w93 and w6238;
w6270 <= not pi0232 and not w6238;
w6271 <= not w5183 and w6270;
w6272 <= w3760 and not w5034;
w6273 <= not w5033 and not w6272;
w6274 <= pi0228 and w6273;
w6275 <= w6238 and not w6274;
w6276 <= w5033 and w5182;
w6277 <= not pi1091 and not w6238;
w6278 <= w6273 and not w6277;
w6279 <= not w5072 and w6278;
w6280 <= not w6276 and not w6279;
w6281 <= pi0228 and not w6280;
w6282 <= pi0232 and not w6275;
w6283 <= not w6281 and w6282;
w6284 <= w93 and not w6271;
w6285 <= not w6283 and w6284;
w6286 <= pi0100 and not w6269;
w6287 <= not w6285 and w6286;
w6288 <= not w6268 and not w6287;
w6289 <= not pi0087 and not w6288;
w6290 <= not w188 and w5491;
w6291 <= pi0087 and not w6290;
w6292 <= not w6209 and not w6291;
w6293 <= w5057 and w5489;
w6294 <= w5065 and not w6293;
w6295 <= not w6210 and w6294;
w6296 <= not w6292 and not w6295;
w6297 <= not w6289 and not w6296;
w6298 <= not pi0075 and not w6297;
w6299 <= not w5038 and w5491;
w6300 <= pi0075 and not w6299;
w6301 <= not w6216 and not w6300;
w6302 <= w5046 and not w6277;
w6303 <= not w6301 and not w6302;
w6304 <= not w6298 and not w6303;
w6305 <= w6229 and not w6304;
w6306 <= w6291 and not w6294;
w6307 <= w5186 and not w5491;
w6308 <= w5107 and not w6261;
w6309 <= not w5491 and not w6184;
w6310 <= not w3805 and w6309;
w6311 <= not w5491 and not w6187;
w6312 <= w3805 and w6311;
w6313 <= w5133 and not w6310;
w6314 <= not w6312 and w6313;
w6315 <= w6236 and not w6314;
w6316 <= not w3768 and w6309;
w6317 <= w3768 and w6311;
w6318 <= w5114 and not w6316;
w6319 <= not w6317 and w6318;
w6320 <= w6247 and not w6319;
w6321 <= pi0039 and not w6315;
w6322 <= not w6320 and w6321;
w6323 <= not w6308 and not w6322;
w6324 <= not pi0038 and not w6323;
w6325 <= w6266 and not w6324;
w6326 <= not w6307 and not w6325;
w6327 <= not pi0087 and not w6326;
w6328 <= not w6306 and not w6327;
w6329 <= not pi0075 and not w6328;
w6330 <= not pi1091 and not w5490;
w6331 <= w5046 and not w6330;
w6332 <= w6300 and not w6331;
w6333 <= not w6329 and not w6332;
w6334 <= w6232 and not w6333;
w6335 <= not w6305 and not w6334;
w6336 <= pi0567 and not w6335;
w6337 <= pi1199 and not w6234;
w6338 <= not w6336 and w6337;
w6339 <= not w5958 and not w6226;
w6340 <= not w6338 and w6339;
w6341 <= w5733 and w5958;
w6342 <= not w5825 and not w6341;
w6343 <= not w6340 and w6342;
w6344 <= not pi1197 and not w6343;
w6345 <= pi1197 and not w5826;
w6346 <= not w6344 and not w6345;
w6347 <= not pi0333 and not w6346;
w6348 <= pi0333 and not w6343;
w6349 <= not w6347 and not w6348;
w6350 <= not pi0391 and not w6349;
w6351 <= not pi0333 and not w6343;
w6352 <= pi0333 and not w6346;
w6353 <= not w6351 and not w6352;
w6354 <= pi0391 and not w6353;
w6355 <= not w6350 and not w6354;
w6356 <= not pi0392 and not w6355;
w6357 <= not pi0391 and not w6353;
w6358 <= pi0391 and not w6349;
w6359 <= not w6357 and not w6358;
w6360 <= pi0392 and not w6359;
w6361 <= not w6356 and not w6360;
w6362 <= pi0393 and w5591;
w6363 <= not pi0393 and not w5591;
w6364 <= not w6362 and not w6363;
w6365 <= not w6361 and not w6364;
w6366 <= not pi0392 and not w6359;
w6367 <= pi0392 and not w6355;
w6368 <= not w6366 and not w6367;
w6369 <= w6364 and not w6368;
w6370 <= pi0591 and not w6365;
w6371 <= not w6369 and w6370;
w6372 <= not pi0592 and w5155;
w6373 <= not w6043 and not w6372;
w6374 <= not w5259 and w6373;
w6375 <= not w5155 and w5259;
w6376 <= not pi1199 and not w6375;
w6377 <= not w6374 and w6376;
w6378 <= w5155 and not w6036;
w6379 <= w6039 and not w6378;
w6380 <= w5155 and not w6031;
w6381 <= w6034 and not w6380;
w6382 <= not w6379 and not w6381;
w6383 <= w5259 and not w6382;
w6384 <= pi1199 and not w6374;
w6385 <= not w6383 and w6384;
w6386 <= not w6377 and not w6385;
w6387 <= not pi0374 and not w6386;
w6388 <= not pi1198 and not w6386;
w6389 <= pi1198 and not w6373;
w6390 <= not w6388 and not w6389;
w6391 <= pi0374 and not w6390;
w6392 <= not w6387 and not w6391;
w6393 <= pi0369 and not w6392;
w6394 <= not pi0374 and not w6390;
w6395 <= pi0374 and not w6386;
w6396 <= not w6394 and not w6395;
w6397 <= not pi0369 and not w6396;
w6398 <= not w6393 and not w6397;
w6399 <= not pi0370 and not w6398;
w6400 <= not pi0369 and not w6392;
w6401 <= pi0369 and not w6396;
w6402 <= not w6400 and not w6401;
w6403 <= pi0370 and not w6402;
w6404 <= not w6399 and not w6403;
w6405 <= not pi0371 and not w6404;
w6406 <= not pi0370 and not w6402;
w6407 <= pi0370 and not w6398;
w6408 <= not w6406 and not w6407;
w6409 <= pi0371 and not w6408;
w6410 <= not w6405 and not w6409;
w6411 <= pi0375 and w5297;
w6412 <= not pi0375 and not w5297;
w6413 <= not w6411 and not w6412;
w6414 <= pi0373 and not w6413;
w6415 <= not pi0373 and w6413;
w6416 <= not w6414 and not w6415;
w6417 <= not w6410 and not w6416;
w6418 <= not pi0371 and not w6408;
w6419 <= pi0371 and not w6404;
w6420 <= not w6418 and not w6419;
w6421 <= w6416 and not w6420;
w6422 <= not pi0591 and not w6417;
w6423 <= not w6421 and w6422;
w6424 <= not pi0590 and not w6371;
w6425 <= not w6423 and w6424;
w6426 <= not w4988 and not w6425;
w6427 <= not w6176 and w6426;
w6428 <= not pi0588 and not w6427;
w6429 <= not w6110 and w6428;
w6430 <= w4989 and not w5875;
w6431 <= not w6429 and w6430;
w6432 <= not pi0217 and not w5720;
w6433 <= not w6431 and w6432;
w6434 <= not w5204 and w5206;
w6435 <= not w6433 and w6434;
w6436 <= pi1161 and not pi1163;
w6437 <= w489 and w6436;
w6438 <= not pi0031 and pi1162;
w6439 <= w6437 and w6438;
w6440 <= not w6435 and not w6439;
w6441 <= w92 and w891;
w6442 <= not pi0055 and not pi0074;
w6443 <= w6441 and w6442;
w6444 <= w3697 and w6443;
w6445 <= pi0100 and w93;
w6446 <= not w3826 and w3837;
w6447 <= w3914 and w6446;
w6448 <= not pi0137 and w6447;
w6449 <= not pi0137 and pi0252;
w6450 <= pi0129 and w84;
w6451 <= not w3837 and not w5037;
w6452 <= w3826 and not w6451;
w6453 <= w6449 and w6452;
w6454 <= w6450 and w6453;
w6455 <= not w6448 and not w6454;
w6456 <= w6445 and not w6455;
w6457 <= not pi0024 and not pi0090;
w6458 <= w3734 and w6457;
w6459 <= w60 and w277;
w6460 <= w264 and w6459;
w6461 <= pi0050 and w340;
w6462 <= w58 and w6461;
w6463 <= not pi0093 and w6460;
w6464 <= w6462 and w6463;
w6465 <= w6458 and w6464;
w6466 <= pi0829 and not pi1093;
w6467 <= w495 and w6466;
w6468 <= not w491 and not w6467;
w6469 <= not w4988 and w6468;
w6470 <= not pi0137 and not w6469;
w6471 <= w6465 and not w6470;
w6472 <= not pi0068 and not pi0073;
w6473 <= w25 and w367;
w6474 <= not pi0103 and w34;
w6475 <= w6473 and w6474;
w6476 <= not pi0089 and not pi0102;
w6477 <= w5001 and w6476;
w6478 <= not pi0045 and not pi0048;
w6479 <= w29 and w360;
w6480 <= not pi0061 and not pi0104;
w6481 <= w6478 and w6480;
w6482 <= w6479 and w6481;
w6483 <= not pi0049 and not pi0066;
w6484 <= not pi0064 and not pi0081;
w6485 <= w50 and w6484;
w6486 <= pi0076 and not pi0084;
w6487 <= w42 and w6486;
w6488 <= w6472 and w6483;
w6489 <= w6487 and w6488;
w6490 <= w6477 and w6485;
w6491 <= w6489 and w6490;
w6492 <= w6475 and w6482;
w6493 <= w6491 and w6492;
w6494 <= w58 and w6493;
w6495 <= w6460 and w6494;
w6496 <= pi0024 and not w6495;
w6497 <= not w6461 and not w6493;
w6498 <= w62 and w265;
w6499 <= not w6497 and w6498;
w6500 <= not pi0024 and not w6499;
w6501 <= w70 and w299;
w6502 <= not pi0137 and w5008;
w6503 <= w6501 and w6502;
w6504 <= not w6469 and w6503;
w6505 <= not w6496 and w6504;
w6506 <= not w6500 and w6505;
w6507 <= not w6471 and not w6506;
w6508 <= not pi0032 and not w6507;
w6509 <= not pi0024 and not pi0841;
w6510 <= pi0032 and not w6509;
w6511 <= w273 and w6510;
w6512 <= not w6508 and not w6511;
w6513 <= not w3732 and not w6512;
w6514 <= not pi0032 and not w6465;
w6515 <= w3732 and not w3736;
w6516 <= not w6514 and w6515;
w6517 <= not w6513 and not w6516;
w6518 <= not pi0095 and w94;
w6519 <= not w6517 and w6518;
w6520 <= not w6456 and not w6519;
w6521 <= w96 and not w6520;
w6522 <= not pi0024 and w68;
w6523 <= w82 and w268;
w6524 <= not pi0051 and w6523;
w6525 <= w6522 and w6524;
w6526 <= w6468 and w6525;
w6527 <= pi0252 and not w6451;
w6528 <= not pi0087 and w93;
w6529 <= pi0075 and not pi0100;
w6530 <= w6528 and w6529;
w6531 <= not pi0137 and w6530;
w6532 <= not w3845 and w6531;
w6533 <= not w6527 and w6532;
w6534 <= w6526 and w6533;
w6535 <= not w6521 and not w6534;
w6536 <= w6444 and not w6535;
w6537 <= not pi0195 and not pi0196;
w6538 <= not pi0138 and w6537;
w6539 <= not pi0139 and w6538;
w6540 <= not pi0118 and w6539;
w6541 <= not pi0079 and w6540;
w6542 <= not pi0034 and w6541;
w6543 <= not pi0033 and not w6542;
w6544 <= pi0149 and pi0157;
w6545 <= not pi0149 and not pi0157;
w6546 <= w3760 and not w6545;
w6547 <= not w6544 and w6546;
w6548 <= pi0232 and w6547;
w6549 <= pi0075 and not w6548;
w6550 <= pi0100 and not w6548;
w6551 <= not w6549 and not w6550;
w6552 <= not pi0075 and not pi0100;
w6553 <= w5036 and w6552;
w6554 <= pi0164 and w6553;
w6555 <= w6551 and not w6554;
w6556 <= not pi0074 and not w6555;
w6557 <= pi0169 and w6553;
w6558 <= w6551 and not w6557;
w6559 <= pi0074 and not w6558;
w6560 <= not w891 and not w6556;
w6561 <= not w6559 and w6560;
w6562 <= pi0054 and not w6555;
w6563 <= pi0164 and w5036;
w6564 <= pi0038 and w6563;
w6565 <= w6552 and w6564;
w6566 <= w6551 and not w6565;
w6567 <= not w6562 and w6566;
w6568 <= not pi0074 and not w6567;
w6569 <= not w6559 and not w6568;
w6570 <= not w92 and not w6569;
w6571 <= w891 and not w6570;
w6572 <= pi0299 and not w6547;
w6573 <= pi0178 and pi0183;
w6574 <= not pi0178 and not pi0183;
w6575 <= w3760 and not w6574;
w6576 <= not w6573 and w6575;
w6577 <= not pi0299 and not w6576;
w6578 <= pi0232 and not w6572;
w6579 <= not w6577 and w6578;
w6580 <= pi0100 and not w6579;
w6581 <= pi0075 and not w6579;
w6582 <= not w6580 and not w6581;
w6583 <= pi0191 and not pi0299;
w6584 <= pi0169 and pi0299;
w6585 <= not w6583 and not w6584;
w6586 <= w6553 and not w6585;
w6587 <= w6582 and not w6586;
w6588 <= pi0074 and not w6587;
w6589 <= not pi0055 and not w6588;
w6590 <= not pi0186 and not pi0299;
w6591 <= not pi0164 and pi0299;
w6592 <= not w6590 and not w6591;
w6593 <= w5036 and w6592;
w6594 <= w6552 and w6593;
w6595 <= w6582 and not w6594;
w6596 <= pi0054 and not w6595;
w6597 <= pi0038 and w6593;
w6598 <= pi0087 and not w6597;
w6599 <= pi0216 and w3942;
w6600 <= w3806 and not w3955;
w6601 <= pi0154 and not w6600;
w6602 <= w3806 and w3959;
w6603 <= not pi0154 and not w6602;
w6604 <= not pi0152 and not w6603;
w6605 <= not w6601 and w6604;
w6606 <= w3760 and w5165;
w6607 <= not w3805 and w6606;
w6608 <= pi0152 and pi0154;
w6609 <= w6607 and w6608;
w6610 <= not w6605 and not w6609;
w6611 <= w6599 and not w6610;
w6612 <= pi0299 and not w6611;
w6613 <= not pi0176 and pi0232;
w6614 <= pi0224 and w3968;
w6615 <= w3769 and w3959;
w6616 <= w6614 and w6615;
w6617 <= not pi0174 and w6616;
w6618 <= not pi0299 and not w6617;
w6619 <= w6613 and not w6618;
w6620 <= pi0176 and pi0232;
w6621 <= w3769 and w6614;
w6622 <= w5165 and w6621;
w6623 <= pi0174 and w6622;
w6624 <= not w3955 and w6614;
w6625 <= w3769 and w6624;
w6626 <= not pi0174 and w6625;
w6627 <= not pi0299 and not w6623;
w6628 <= not w6626 and w6627;
w6629 <= w6620 and not w6628;
w6630 <= not w6619 and not w6629;
w6631 <= pi0039 and not w6612;
w6632 <= not w6630 and w6631;
w6633 <= w744 and w3760;
w6634 <= pi0180 and w6633;
w6635 <= pi0090 and not w4995;
w6636 <= not pi0072 and not pi0093;
w6637 <= w270 and w6636;
w6638 <= not w6635 and w6637;
w6639 <= not pi0066 and not pi0084;
w6640 <= not pi0068 and w31;
w6641 <= not pi0111 and w30;
w6642 <= not pi0036 and w6640;
w6643 <= w6641 and w6642;
w6644 <= not pi0102 and w6484;
w6645 <= w29 and w6644;
w6646 <= w27 and w6645;
w6647 <= pi0073 and not pi0082;
w6648 <= w6639 and w6647;
w6649 <= w6643 and w6648;
w6650 <= w6646 and w6649;
w6651 <= w40 and w6650;
w6652 <= w6498 and w6651;
w6653 <= w50 and w6652;
w6654 <= w3702 and not w6653;
w6655 <= w6638 and not w6654;
w6656 <= w81 and w3760;
w6657 <= not pi0040 and w6656;
w6658 <= w6655 and w6657;
w6659 <= not pi0183 and w6658;
w6660 <= pi0183 and w3760;
w6661 <= w67 and not w3702;
w6662 <= not w6635 and w6661;
w6663 <= w48 and w6646;
w6664 <= not pi0060 and w6663;
w6665 <= pi0053 and not w6664;
w6666 <= not pi0060 and w6461;
w6667 <= w282 and not w6666;
w6668 <= not w6665 and not w6667;
w6669 <= w57 and w6651;
w6670 <= w50 and not w6669;
w6671 <= not w6668 and w6670;
w6672 <= w283 and not w6671;
w6673 <= not pi0090 and w280;
w6674 <= w67 and w6673;
w6675 <= w286 and w6674;
w6676 <= w50 and w6675;
w6677 <= w6672 and w6676;
w6678 <= not pi0070 and not w6677;
w6679 <= not w6662 and w6678;
w6680 <= w82 and w663;
w6681 <= not w6679 and w6680;
w6682 <= not w6678 and w6680;
w6683 <= not w4050 and not w6682;
w6684 <= not pi0198 and not w6683;
w6685 <= not w6681 and not w6684;
w6686 <= w6660 and not w6685;
w6687 <= not pi0174 and not w6659;
w6688 <= not w6686 and w6687;
w6689 <= not w6667 and w6675;
w6690 <= not pi0070 and not w6689;
w6691 <= not w6662 and w6690;
w6692 <= w6680 and not w6691;
w6693 <= not w4082 and not w6692;
w6694 <= w3760 and not w6693;
w6695 <= pi0183 and w6694;
w6696 <= not w3702 and w6638;
w6697 <= w6657 and w6696;
w6698 <= not pi0183 and w6697;
w6699 <= pi0174 and not w6698;
w6700 <= not w6695 and w6699;
w6701 <= not w6688 and not w6700;
w6702 <= pi0193 and not w6701;
w6703 <= not pi0040 and w3760;
w6704 <= not pi0090 and w6637;
w6705 <= w6653 and w6704;
w6706 <= w81 and w6705;
w6707 <= w6703 and w6706;
w6708 <= not pi0174 and not pi0183;
w6709 <= w6707 and w6708;
w6710 <= not w4082 and not w6682;
w6711 <= not pi0174 and w6710;
w6712 <= w6680 and not w6690;
w6713 <= not w4082 and not w6712;
w6714 <= pi0174 and w6713;
w6715 <= w6660 and not w6714;
w6716 <= not w6711 and w6715;
w6717 <= not pi0193 and not w6709;
w6718 <= not w6716 and w6717;
w6719 <= not w6702 and not w6718;
w6720 <= not pi0299 and not w6634;
w6721 <= not w6719 and w6720;
w6722 <= not pi0039 and pi0232;
w6723 <= pi0158 and w6633;
w6724 <= pi0172 and w6681;
w6725 <= not w4051 and not w6682;
w6726 <= not pi0152 and w6725;
w6727 <= not w6724 and w6726;
w6728 <= pi0172 and w6692;
w6729 <= not w4051 and not w6712;
w6730 <= pi0152 and not w6728;
w6731 <= w6729 and w6730;
w6732 <= pi0149 and w3760;
w6733 <= not w6731 and w6732;
w6734 <= not w6727 and w6733;
w6735 <= not pi0152 and w6658;
w6736 <= not w6697 and not w6735;
w6737 <= pi0172 and not w6736;
w6738 <= not pi0152 and not pi0172;
w6739 <= w6707 and w6738;
w6740 <= not w6737 and not w6739;
w6741 <= not pi0149 and not w6740;
w6742 <= pi0299 and not w6723;
w6743 <= not w6741 and w6742;
w6744 <= not w6734 and w6743;
w6745 <= w6722 and not w6744;
w6746 <= not w6721 and w6745;
w6747 <= not w6632 and not w6746;
w6748 <= not pi0038 and not w6747;
w6749 <= pi0299 and w5036;
w6750 <= not w3698 and w6749;
w6751 <= not pi0186 and not w6750;
w6752 <= not w3847 and w5036;
w6753 <= pi0186 and not w6752;
w6754 <= pi0164 and not w6753;
w6755 <= not w6751 and w6754;
w6756 <= not pi0299 and w5036;
w6757 <= not w3698 and w6756;
w6758 <= not pi0164 and pi0186;
w6759 <= w6757 and w6758;
w6760 <= not w6755 and not w6759;
w6761 <= pi0038 and not w6760;
w6762 <= not pi0087 and not w6761;
w6763 <= not w6748 and w6762;
w6764 <= not pi0100 and not w6598;
w6765 <= not w6763 and w6764;
w6766 <= not w6580 and not w6765;
w6767 <= w132 and not w6766;
w6768 <= not pi0075 and pi0092;
w6769 <= not pi0100 and w6597;
w6770 <= not w6580 and not w6769;
w6771 <= not pi0038 and not pi0087;
w6772 <= pi0232 and not w946;
w6773 <= not pi0176 and not pi0299;
w6774 <= w3760 and not w6773;
w6775 <= w6772 and w6774;
w6776 <= not pi0100 and w6771;
w6777 <= w6775 and w6776;
w6778 <= w3698 and w6777;
w6779 <= w6770 and not w6778;
w6780 <= w6768 and not w6779;
w6781 <= not w6581 and not w6780;
w6782 <= not w6767 and w6781;
w6783 <= not pi0054 and not w6782;
w6784 <= not w6596 and not w6783;
w6785 <= not pi0074 and not w6784;
w6786 <= w6589 and not w6785;
w6787 <= pi0055 and not w6559;
w6788 <= not pi0092 and not w6549;
w6789 <= pi0038 and not w6563;
w6790 <= w131 and not w6789;
w6791 <= pi0149 and w5036;
w6792 <= w3698 and w6791;
w6793 <= not pi0038 and not w6792;
w6794 <= w6790 and not w6793;
w6795 <= w5724 and w6564;
w6796 <= not w6550 and not w6795;
w6797 <= not w6794 and w6796;
w6798 <= not pi0075 and not w6797;
w6799 <= w6788 and not w6798;
w6800 <= pi0092 and w6566;
w6801 <= not pi0054 and not w6800;
w6802 <= not w6799 and w6801;
w6803 <= not w6562 and not w6802;
w6804 <= not pi0074 and not w6803;
w6805 <= w6787 and not w6804;
w6806 <= w92 and not w6805;
w6807 <= not w6786 and w6806;
w6808 <= w6571 and not w6807;
w6809 <= not w6561 and not w6808;
w6810 <= w6543 and not w6809;
w6811 <= not pi0040 and w50;
w6812 <= not pi0038 and w6811;
w6813 <= w6552 and w6812;
w6814 <= w95 and w6813;
w6815 <= not w92 and w6814;
w6816 <= w279 and w283;
w6817 <= not pi0053 and w6816;
w6818 <= w6664 and w6817;
w6819 <= not pi0058 and w6818;
w6820 <= w5008 and w6819;
w6821 <= not pi0032 and w71;
w6822 <= w6820 and w6821;
w6823 <= not pi0095 and w6822;
w6824 <= not pi0039 and not w6791;
w6825 <= w6823 and w6824;
w6826 <= w6811 and not w6825;
w6827 <= not pi0038 and not w6826;
w6828 <= w6790 and not w6827;
w6829 <= not pi0038 and not w6811;
w6830 <= not pi0100 and not w6829;
w6831 <= not w6789 and w6830;
w6832 <= pi0087 and w6831;
w6833 <= not w6550 and not w6832;
w6834 <= not w6828 and w6833;
w6835 <= not pi0075 and not w6834;
w6836 <= w6788 and not w6835;
w6837 <= not pi0075 and w6831;
w6838 <= pi0092 and w6551;
w6839 <= not w6837 and w6838;
w6840 <= not pi0054 and not w6839;
w6841 <= not w6836 and w6840;
w6842 <= not w6562 and not w6841;
w6843 <= not pi0074 and not w6842;
w6844 <= w6787 and not w6843;
w6845 <= w172 and w6823;
w6846 <= not w6775 and w6845;
w6847 <= w171 and w6811;
w6848 <= not w6846 and w6847;
w6849 <= w6770 and not w6848;
w6850 <= w6768 and not w6849;
w6851 <= pi0087 and not w6847;
w6852 <= w6770 and w6851;
w6853 <= not w6599 and w6811;
w6854 <= pi0299 and not w6853;
w6855 <= w3946 and not w3958;
w6856 <= w3775 and w6855;
w6857 <= not w3751 and not w6856;
w6858 <= w6823 and not w6857;
w6859 <= w3761 and w6858;
w6860 <= w6811 and not w6859;
w6861 <= w3760 and w6858;
w6862 <= w6811 and not w6861;
w6863 <= not w3805 and not w6862;
w6864 <= w6860 and not w6863;
w6865 <= w6854 and not w6864;
w6866 <= not w6614 and w6811;
w6867 <= not w6860 and not w6866;
w6868 <= not w3768 and not w6862;
w6869 <= not w6866 and w6868;
w6870 <= not w6867 and not w6869;
w6871 <= not pi0299 and not w6870;
w6872 <= not w6865 and not w6871;
w6873 <= not pi0232 and not w6872;
w6874 <= w6823 and w6856;
w6875 <= w3760 and w6874;
w6876 <= w6811 and not w6875;
w6877 <= not w3768 and not w6876;
w6878 <= not w6866 and w6877;
w6879 <= pi0174 and w6878;
w6880 <= not w6867 and not w6879;
w6881 <= not pi0299 and not w6880;
w6882 <= w6811 and not w6874;
w6883 <= w3806 and not w6882;
w6884 <= pi0152 and w6883;
w6885 <= w6860 and not w6884;
w6886 <= pi0154 and not w6885;
w6887 <= w3751 and w6823;
w6888 <= not w3790 and w6887;
w6889 <= w6811 and not w6888;
w6890 <= w3760 and w6889;
w6891 <= not pi0152 and w6890;
w6892 <= not pi0154 and not w6864;
w6893 <= not w6891 and w6892;
w6894 <= w6599 and not w6886;
w6895 <= not w6893 and w6894;
w6896 <= w6854 and not w6895;
w6897 <= not w6881 and not w6896;
w6898 <= w3769 and w6887;
w6899 <= w6614 and w6811;
w6900 <= not w6898 and w6899;
w6901 <= not w6866 and not w6900;
w6902 <= not pi0299 and w6901;
w6903 <= w6897 and not w6902;
w6904 <= w6613 and not w6903;
w6905 <= w6620 and not w6897;
w6906 <= pi0039 and not w6873;
w6907 <= not w6905 and w6906;
w6908 <= not w6904 and w6907;
w6909 <= pi0095 and not w6811;
w6910 <= not w5 and not w6909;
w6911 <= not pi0040 and not pi0479;
w6912 <= w50 and not w6822;
w6913 <= w6911 and w6912;
w6914 <= not w6910 and not w6913;
w6915 <= pi0032 and not w6811;
w6916 <= w50 and not w69;
w6917 <= w50 and not w6820;
w6918 <= pi0070 and not w6917;
w6919 <= w50 and not w6818;
w6920 <= pi0058 and not w6919;
w6921 <= w50 and not w279;
w6922 <= not w50 and not w283;
w6923 <= w279 and not w6922;
w6924 <= not w6672 and w6923;
w6925 <= not pi0058 and not w6921;
w6926 <= not w6924 and w6925;
w6927 <= not w6920 and not w6926;
w6928 <= not pi0090 and not w6927;
w6929 <= not pi0841 and w6819;
w6930 <= w50 and not w6929;
w6931 <= pi0090 and not w6930;
w6932 <= w67 and not w6931;
w6933 <= not w6928 and w6932;
w6934 <= w50 and not w67;
w6935 <= not pi0070 and not w6934;
w6936 <= not w6933 and w6935;
w6937 <= not w6918 and not w6936;
w6938 <= not pi0051 and not w6937;
w6939 <= pi0051 and not w50;
w6940 <= w69 and not w6939;
w6941 <= not w6938 and w6940;
w6942 <= not w6916 and not w6941;
w6943 <= not pi0040 and not w6942;
w6944 <= not pi0032 and not w6943;
w6945 <= not w6915 and not w6944;
w6946 <= not pi0095 and not w6945;
w6947 <= not w6914 and not w6946;
w6948 <= w6704 and w6929;
w6949 <= w6811 and not w6948;
w6950 <= pi0032 and not w6949;
w6951 <= not w6944 and not w6950;
w6952 <= not pi0095 and not w6951;
w6953 <= not pi0198 and w6952;
w6954 <= w6947 and not w6953;
w6955 <= not w3760 and w6954;
w6956 <= w6668 and w6816;
w6957 <= w50 and not w6956;
w6958 <= not pi0058 and not w6957;
w6959 <= not w6920 and not w6958;
w6960 <= not pi0090 and not w6959;
w6961 <= w6932 and not w6960;
w6962 <= w6935 and not w6961;
w6963 <= not w6918 and not w6962;
w6964 <= not pi0051 and not w6963;
w6965 <= w6940 and not w6964;
w6966 <= not w6916 and not w6965;
w6967 <= not pi0040 and not w6966;
w6968 <= not pi0032 and not w6967;
w6969 <= not w6950 and not w6968;
w6970 <= not pi0095 and not w6969;
w6971 <= not pi0198 and w6970;
w6972 <= w3760 and not w6909;
w6973 <= not w6915 and not w6968;
w6974 <= not pi0095 and not w6973;
w6975 <= w6972 and not w6974;
w6976 <= not w6971 and w6975;
w6977 <= not w6955 and not w6976;
w6978 <= not pi0183 and not w6977;
w6979 <= not pi0040 and not w6915;
w6980 <= w50 and not w3733;
w6981 <= not pi0032 and not w6980;
w6982 <= pi0093 and not w50;
w6983 <= w3733 and not w6982;
w6984 <= w50 and not w6920;
w6985 <= not pi0090 and not w6984;
w6986 <= not w6931 and not w6985;
w6987 <= not pi0093 and not w6986;
w6988 <= w6983 and not w6987;
w6989 <= w6981 and not w6988;
w6990 <= w6979 and not w6989;
w6991 <= not pi0095 and not w6990;
w6992 <= w6972 and not w6991;
w6993 <= not w6955 and not w6992;
w6994 <= pi0183 and not w6993;
w6995 <= not w6978 and not w6994;
w6996 <= not pi0095 and w6995;
w6997 <= not pi0174 and not w6914;
w6998 <= not w6996 and w6997;
w6999 <= not w6660 and not w6954;
w7000 <= not pi0090 and w6652;
w7001 <= w6986 and not w7000;
w7002 <= not pi0093 and not w7001;
w7003 <= w6983 and not w7002;
w7004 <= w6981 and not w7003;
w7005 <= w6979 and not w7004;
w7006 <= not pi0095 and not w7005;
w7007 <= not w6914 and not w7006;
w7008 <= w3760 and not w7007;
w7009 <= pi0183 and w7008;
w7010 <= pi0174 and not w7009;
w7011 <= not w6999 and w7010;
w7012 <= not pi0180 and not w7011;
w7013 <= not w6998 and w7012;
w7014 <= not pi0174 and not w6995;
w7015 <= w6972 and not w7006;
w7016 <= not w6955 and not w7015;
w7017 <= pi0183 and not w7016;
w7018 <= not w6909 and not w6946;
w7019 <= not w6953 and w7018;
w7020 <= w6703 and w7019;
w7021 <= not w6955 and not w7020;
w7022 <= not pi0183 and not w7021;
w7023 <= not w7017 and not w7022;
w7024 <= pi0174 and not w7023;
w7025 <= pi0180 and not w7014;
w7026 <= not w7024 and w7025;
w7027 <= not w7013 and not w7026;
w7028 <= not pi0193 and not w7027;
w7029 <= not pi0040 and not w50;
w7030 <= pi0032 and not w7029;
w7031 <= w24 and w67;
w7032 <= not w50 and not w7031;
w7033 <= w5008 and w6926;
w7034 <= not w7032 and not w7033;
w7035 <= not pi0070 and not w7034;
w7036 <= not w6918 and not w7035;
w7037 <= not pi0051 and not w7036;
w7038 <= w6940 and not w7037;
w7039 <= not pi0040 and not w6916;
w7040 <= not w7038 and w7039;
w7041 <= not pi0032 and not w7040;
w7042 <= not w7030 and not w7041;
w7043 <= not w299 and not w6811;
w7044 <= not w7042 and not w7043;
w7045 <= not pi0095 and not w7044;
w7046 <= not w6914 and not w7045;
w7047 <= not w6909 and not w7045;
w7048 <= pi0095 and not w7029;
w7049 <= not pi0040 and not w6949;
w7050 <= pi0032 and not w7049;
w7051 <= not w7041 and not w7050;
w7052 <= not pi0095 and not w7051;
w7053 <= not w7048 and not w7052;
w7054 <= w7047 and not w7053;
w7055 <= not pi0198 and not w7054;
w7056 <= w3760 and not w7055;
w7057 <= w3760 and not w6811;
w7058 <= not w7056 and not w7057;
w7059 <= w7046 and not w7058;
w7060 <= not w6955 and not w7059;
w7061 <= not pi0183 and not w7060;
w7062 <= w267 and w3733;
w7063 <= w6498 and w7062;
w7064 <= not pi0032 and w7063;
w7065 <= w6651 and w7064;
w7066 <= w6811 and not w7065;
w7067 <= not pi0095 and not w7066;
w7068 <= w3760 and not w7067;
w7069 <= not w6914 and w7068;
w7070 <= not w6955 and not w7069;
w7071 <= pi0183 and not w7070;
w7072 <= pi0174 and not w7071;
w7073 <= not w7061 and w7072;
w7074 <= not w3760 and not w6954;
w7075 <= w5008 and w6958;
w7076 <= not w7032 and not w7075;
w7077 <= not pi0070 and not w7076;
w7078 <= not w6918 and not w7077;
w7079 <= not pi0051 and not w7078;
w7080 <= w6940 and not w7079;
w7081 <= not w6916 and not w7080;
w7082 <= not pi0040 and not w7081;
w7083 <= not pi0032 and not w7082;
w7084 <= not w6915 and not w7083;
w7085 <= not pi0095 and not w7084;
w7086 <= not w6914 and not w7085;
w7087 <= not w6950 and not w7083;
w7088 <= not pi0095 and not w7087;
w7089 <= not pi0198 and w7088;
w7090 <= w7086 and not w7089;
w7091 <= w3760 and not w7090;
w7092 <= not w7074 and not w7091;
w7093 <= not pi0183 and w7092;
w7094 <= not pi0095 and not w6811;
w7095 <= not w6914 and not w7094;
w7096 <= w3760 and w7095;
w7097 <= not w6955 and not w7096;
w7098 <= pi0183 and not w7097;
w7099 <= not pi0174 and not w7093;
w7100 <= not w7098 and w7099;
w7101 <= not pi0180 and not w7100;
w7102 <= not w7073 and w7101;
w7103 <= w6972 and not w7067;
w7104 <= not w6955 and not w7103;
w7105 <= pi0183 and not w7104;
w7106 <= w7047 and w7056;
w7107 <= not w6955 and not w7106;
w7108 <= not pi0183 and not w7107;
w7109 <= pi0174 and not w7105;
w7110 <= not w7108 and w7109;
w7111 <= not w7057 and not w7074;
w7112 <= pi0183 and w7111;
w7113 <= not pi0040 and w7081;
w7114 <= not pi0032 and not w7113;
w7115 <= not w7030 and not w7114;
w7116 <= not pi0095 and not w7115;
w7117 <= not w7048 and not w7116;
w7118 <= pi0198 and not w7117;
w7119 <= not w7050 and not w7114;
w7120 <= not pi0095 and not w7119;
w7121 <= not w7048 and not w7120;
w7122 <= not pi0198 and not w7121;
w7123 <= not w7118 and not w7122;
w7124 <= w6703 and not w7123;
w7125 <= not w6955 and not w7124;
w7126 <= not pi0183 and not w7125;
w7127 <= not pi0174 and not w7112;
w7128 <= not w7126 and w7127;
w7129 <= pi0180 and not w7110;
w7130 <= not w7128 and w7129;
w7131 <= pi0193 and not w7102;
w7132 <= not w7130 and w7131;
w7133 <= not w7028 and not w7132;
w7134 <= not pi0299 and not w7133;
w7135 <= pi0158 and pi0299;
w7136 <= not pi0210 and w6952;
w7137 <= w6947 and not w7136;
w7138 <= not w3760 and w7137;
w7139 <= not pi0210 and w6970;
w7140 <= w6975 and not w7139;
w7141 <= not w7138 and not w7140;
w7142 <= not pi0152 and not w7141;
w7143 <= not w3760 and not w7137;
w7144 <= w7018 and not w7136;
w7145 <= w3760 and not w7144;
w7146 <= not w7143 and not w7145;
w7147 <= pi0152 and w7146;
w7148 <= not pi0172 and not w7142;
w7149 <= not w7147 and w7148;
w7150 <= not w6909 and not w7088;
w7151 <= not pi0210 and not w7150;
w7152 <= w3760 and not w7151;
w7153 <= not w6909 and not w7085;
w7154 <= w7152 and w7153;
w7155 <= not w7138 and not w7154;
w7156 <= not pi0152 and not w7155;
w7157 <= not pi0210 and not w7054;
w7158 <= w3760 and not w7157;
w7159 <= w7047 and w7158;
w7160 <= not w7138 and not w7159;
w7161 <= pi0152 and not w7160;
w7162 <= pi0172 and not w7156;
w7163 <= not w7161 and w7162;
w7164 <= not w7149 and not w7163;
w7165 <= w7135 and not w7164;
w7166 <= not pi0158 and pi0299;
w7167 <= not w6914 and not w6974;
w7168 <= not w7139 and w7167;
w7169 <= w3760 and w7168;
w7170 <= not pi0152 and not w7169;
w7171 <= pi0152 and not w7137;
w7172 <= not pi0172 and not w7170;
w7173 <= not w7171 and w7172;
w7174 <= not w7057 and not w7158;
w7175 <= w7046 and not w7174;
w7176 <= pi0152 and not w7175;
w7177 <= not w7057 and not w7152;
w7178 <= w7086 and not w7177;
w7179 <= not pi0152 and not w7178;
w7180 <= pi0172 and not w7179;
w7181 <= not w7176 and w7180;
w7182 <= not w7138 and w7166;
w7183 <= not w7173 and w7182;
w7184 <= not w7181 and w7183;
w7185 <= not pi0149 and not w7184;
w7186 <= not w7165 and w7185;
w7187 <= not w7015 and not w7138;
w7188 <= pi0152 and not w7187;
w7189 <= not w6992 and not w7138;
w7190 <= not pi0152 and not w7189;
w7191 <= not pi0172 and not w7188;
w7192 <= not w7190 and w7191;
w7193 <= not w7103 and not w7138;
w7194 <= pi0152 and not w7193;
w7195 <= not w7057 and not w7143;
w7196 <= not pi0152 and w7195;
w7197 <= pi0172 and not w7194;
w7198 <= not w7196 and w7197;
w7199 <= not w7192 and not w7198;
w7200 <= w7135 and not w7199;
w7201 <= not w7069 and not w7138;
w7202 <= pi0152 and not w7201;
w7203 <= not w7096 and not w7138;
w7204 <= not pi0152 and not w7203;
w7205 <= pi0172 and not w7202;
w7206 <= not w7204 and w7205;
w7207 <= not w6914 and not w6991;
w7208 <= w3760 and not w7207;
w7209 <= not w7143 and not w7208;
w7210 <= not pi0152 and w7209;
w7211 <= not w7008 and not w7143;
w7212 <= pi0152 and w7211;
w7213 <= not pi0172 and not w7210;
w7214 <= not w7212 and w7213;
w7215 <= not w7206 and not w7214;
w7216 <= w7166 and not w7215;
w7217 <= pi0149 and not w7200;
w7218 <= not w7216 and w7217;
w7219 <= not w7186 and not w7218;
w7220 <= not w7134 and not w7219;
w7221 <= pi0232 and not w7220;
w7222 <= not w3732 and w6952;
w7223 <= w6947 and not w7222;
w7224 <= not pi0232 and not w7223;
w7225 <= not pi0039 and not w7224;
w7226 <= not w7221 and w7225;
w7227 <= not w6908 and not w7226;
w7228 <= not pi0038 and not w7227;
w7229 <= not w6761 and not w7228;
w7230 <= not pi0100 and not w7229;
w7231 <= not pi0087 and not w6580;
w7232 <= not w7230 and w7231;
w7233 <= w132 and not w6852;
w7234 <= not w7232 and w7233;
w7235 <= not w6581 and not w6850;
w7236 <= not w7234 and w7235;
w7237 <= not pi0054 and not w7236;
w7238 <= not w6596 and not w7237;
w7239 <= not pi0074 and not w7238;
w7240 <= w6589 and not w7239;
w7241 <= w92 and not w6844;
w7242 <= not w7240 and w7241;
w7243 <= w6571 and not w6815;
w7244 <= not w7242 and w7243;
w7245 <= not w6561 and not w7244;
w7246 <= not w6543 and not w7245;
w7247 <= not pi0954 and not w6810;
w7248 <= not w7246 and w7247;
w7249 <= pi0033 and not w6809;
w7250 <= not pi0033 and not w7245;
w7251 <= pi0954 and not w7249;
w7252 <= not w7250 and w7251;
w7253 <= not w7248 and not w7252;
w7254 <= pi0197 and w6545;
w7255 <= not pi0197 and not w6545;
w7256 <= not w7254 and not w7255;
w7257 <= pi0162 and w3760;
w7258 <= w7256 and not w7257;
w7259 <= w7254 and w7257;
w7260 <= not pi0162 and not pi0197;
w7261 <= w6546 and not w7260;
w7262 <= w3760 and not w7261;
w7263 <= not w7259 and w7262;
w7264 <= not w7256 and not w7263;
w7265 <= not w7258 and not w7264;
w7266 <= pi0232 and w7265;
w7267 <= not w6552 and w7266;
w7268 <= pi0167 and w5036;
w7269 <= w6552 and w7268;
w7270 <= not w7267 and not w7269;
w7271 <= not pi0074 and w7270;
w7272 <= pi0148 and w6553;
w7273 <= pi0074 and not w7272;
w7274 <= not w7267 and w7273;
w7275 <= not w7271 and not w7274;
w7276 <= not w891 and w7275;
w7277 <= not pi0054 and not w7267;
w7278 <= pi0038 and w7269;
w7279 <= w7277 and not w7278;
w7280 <= not pi0074 and w7279;
w7281 <= w7275 and not w7280;
w7282 <= not w92 and not w7281;
w7283 <= w891 and not w7282;
w7284 <= pi0140 and pi0145;
w7285 <= w6574 and not w7284;
w7286 <= not pi0140 and not pi0145;
w7287 <= w3760 and not w7286;
w7288 <= w7285 and w7287;
w7289 <= not w7284 and not w7286;
w7290 <= w6575 and not w7289;
w7291 <= not pi0299 and not w7288;
w7292 <= not w7290 and w7291;
w7293 <= pi0299 and not w7265;
w7294 <= pi0232 and not w7292;
w7295 <= not w7293 and w7294;
w7296 <= pi0100 and not w7295;
w7297 <= pi0075 and not w7295;
w7298 <= not w7296 and not w7297;
w7299 <= pi0141 and not pi0299;
w7300 <= pi0148 and pi0299;
w7301 <= not w7299 and not w7300;
w7302 <= w5036 and not w7301;
w7303 <= w6552 and not w7302;
w7304 <= w7298 and not w7303;
w7305 <= pi0074 and not w7304;
w7306 <= not pi0055 and not w7305;
w7307 <= pi0188 and not pi0299;
w7308 <= pi0167 and pi0299;
w7309 <= not w7307 and not w7308;
w7310 <= w5036 and not w7309;
w7311 <= not pi0100 and not w7310;
w7312 <= not pi0075 and w7311;
w7313 <= w7298 and not w7312;
w7314 <= pi0054 and not w7313;
w7315 <= not pi0188 and not w6750;
w7316 <= pi0188 and w6757;
w7317 <= not pi0167 and not w7316;
w7318 <= pi0167 and pi0188;
w7319 <= not w6752 and w7318;
w7320 <= not w7315 and not w7319;
w7321 <= not w7317 and w7320;
w7322 <= pi0038 and not w7321;
w7323 <= not pi0038 and pi0155;
w7324 <= pi0161 and not w6607;
w7325 <= not pi0161 and not w6600;
w7326 <= w6599 and not w7325;
w7327 <= not w7324 and w7326;
w7328 <= w7323 and not w7327;
w7329 <= not pi0038 and not pi0155;
w7330 <= not pi0161 and w6599;
w7331 <= w6602 and w7330;
w7332 <= w7329 and not w7331;
w7333 <= not w7328 and not w7332;
w7334 <= pi0299 and not w7333;
w7335 <= not pi0177 and not pi0299;
w7336 <= not pi0144 and w6616;
w7337 <= w7335 and not w7336;
w7338 <= not pi0144 and w6625;
w7339 <= pi0177 and not pi0299;
w7340 <= pi0144 and w6622;
w7341 <= w7339 and not w7340;
w7342 <= not w7338 and w7341;
w7343 <= pi0232 and not w7337;
w7344 <= not w7342 and w7343;
w7345 <= not pi0038 and not w7344;
w7346 <= not w7334 and not w7345;
w7347 <= pi0039 and not w7346;
w7348 <= not pi0146 and not w6658;
w7349 <= pi0146 and not w6707;
w7350 <= not pi0161 and not w7349;
w7351 <= not w7348 and w7350;
w7352 <= not pi0146 and pi0161;
w7353 <= w6697 and w7352;
w7354 <= not w7351 and not w7353;
w7355 <= not pi0162 and not w7354;
w7356 <= not pi0159 and pi0299;
w7357 <= pi0159 and pi0299;
w7358 <= not pi0162 and w6633;
w7359 <= w7357 and not w7358;
w7360 <= not w7356 and not w7359;
w7361 <= not w7257 and not w7360;
w7362 <= pi0159 and w744;
w7363 <= not pi0146 and w6692;
w7364 <= w6729 and not w7363;
w7365 <= pi0161 and not w7364;
w7366 <= not pi0146 and w6681;
w7367 <= w6725 and not w7366;
w7368 <= not pi0161 and not w7367;
w7369 <= pi0299 and not w7362;
w7370 <= not w7365 and w7369;
w7371 <= not w7368 and w7370;
w7372 <= not w7361 and not w7371;
w7373 <= not w7355 and not w7372;
w7374 <= pi0181 and w6633;
w7375 <= pi0140 and not w3760;
w7376 <= not pi0142 and w6697;
w7377 <= not pi0140 and not w7376;
w7378 <= not pi0142 and w6692;
w7379 <= pi0140 and not w7378;
w7380 <= w6713 and w7379;
w7381 <= not w7377 and not w7380;
w7382 <= pi0144 and not w7381;
w7383 <= not pi0142 and w6658;
w7384 <= pi0142 and w6707;
w7385 <= not pi0140 and not w7384;
w7386 <= not w7383 and w7385;
w7387 <= not pi0142 and w6681;
w7388 <= pi0140 and w6710;
w7389 <= not w7387 and w7388;
w7390 <= not w7386 and not w7389;
w7391 <= not pi0144 and not w7390;
w7392 <= not w7375 and not w7382;
w7393 <= not w7391 and w7392;
w7394 <= not pi0299 and not w7374;
w7395 <= not w7393 and w7394;
w7396 <= pi0232 and not w7373;
w7397 <= not w7395 and w7396;
w7398 <= w93 and not w7397;
w7399 <= not w7322 and not w7347;
w7400 <= not w7398 and w7399;
w7401 <= not pi0100 and not w7400;
w7402 <= not w7296 and not w7401;
w7403 <= not pi0087 and not w7402;
w7404 <= not w171 and not w7311;
w7405 <= not w7296 and w7404;
w7406 <= pi0087 and not w7405;
w7407 <= not w7403 and not w7406;
w7408 <= w132 and not w7407;
w7409 <= pi0038 and not w7309;
w7410 <= pi0155 and pi0299;
w7411 <= not w7339 and not w7410;
w7412 <= w93 and not w7411;
w7413 <= w75 and w7412;
w7414 <= not w7409 and not w7413;
w7415 <= w5036 and not w7414;
w7416 <= not pi0100 and not w7415;
w7417 <= not w7296 and not w7416;
w7418 <= not pi0087 and not w7417;
w7419 <= not w7406 and not w7418;
w7420 <= w6768 and not w7419;
w7421 <= not w7297 and not w7420;
w7422 <= not w7408 and w7421;
w7423 <= not pi0054 and not w7422;
w7424 <= not w7314 and not w7423;
w7425 <= not pi0074 and not w7424;
w7426 <= w7306 and not w7425;
w7427 <= pi0055 and not w7274;
w7428 <= pi0054 and w7270;
w7429 <= pi0038 and w7268;
w7430 <= not pi0092 and pi0162;
w7431 <= w6722 and w7430;
w7432 <= w6771 and w7431;
w7433 <= w3785 and w7432;
w7434 <= not w7429 and not w7433;
w7435 <= w6552 and not w7434;
w7436 <= w7277 and not w7435;
w7437 <= not w7428 and not w7436;
w7438 <= not pi0074 and not w7437;
w7439 <= w7427 and not w7438;
w7440 <= w92 and not w7439;
w7441 <= not w7426 and w7440;
w7442 <= w7283 and not w7441;
w7443 <= not w7276 and not w7442;
w7444 <= pi0034 and w7443;
w7445 <= not w92 and not w6814;
w7446 <= w891 and not w7445;
w7447 <= not w7283 and not w7446;
w7448 <= not w6813 and w7279;
w7449 <= not w3697 and not w7448;
w7450 <= pi0075 and not w7266;
w7451 <= pi0100 and not w7266;
w7452 <= w6845 and not w7257;
w7453 <= w6812 and not w7452;
w7454 <= not pi0100 and not w7453;
w7455 <= not pi0232 and w6845;
w7456 <= not w7454 and not w7455;
w7457 <= not w7429 and not w7456;
w7458 <= not w7451 and not w7457;
w7459 <= not pi0075 and not w7458;
w7460 <= not pi0092 and not w7450;
w7461 <= not w7459 and w7460;
w7462 <= not w7449 and not w7461;
w7463 <= not w7428 and not w7462;
w7464 <= not pi0074 and not w7463;
w7465 <= w7427 and not w7464;
w7466 <= pi0146 and w7209;
w7467 <= not pi0146 and not w7203;
w7468 <= not pi0161 and not w7466;
w7469 <= not w7467 and w7468;
w7470 <= pi0146 and w7211;
w7471 <= not pi0146 and not w7201;
w7472 <= pi0161 and not w7470;
w7473 <= not w7471 and w7472;
w7474 <= not w7469 and not w7473;
w7475 <= pi0162 and not w7474;
w7476 <= not pi0161 and not w7169;
w7477 <= pi0161 and not w7137;
w7478 <= pi0146 and not w7476;
w7479 <= not w7477 and w7478;
w7480 <= not pi0161 and not w7178;
w7481 <= pi0161 and not w7175;
w7482 <= not pi0146 and not w7480;
w7483 <= not w7481 and w7482;
w7484 <= not pi0162 and not w7138;
w7485 <= not w7479 and w7484;
w7486 <= not w7483 and w7485;
w7487 <= not w7475 and not w7486;
w7488 <= w7356 and not w7487;
w7489 <= pi0142 and w6954;
w7490 <= not pi0142 and not w7060;
w7491 <= not pi0140 and not w7489;
w7492 <= not w7490 and w7491;
w7493 <= pi0142 and not w7008;
w7494 <= not w7074 and w7493;
w7495 <= not pi0142 and not w7070;
w7496 <= pi0140 and not w7494;
w7497 <= not w7495 and w7496;
w7498 <= not w7492 and not w7497;
w7499 <= not pi0181 and not w7498;
w7500 <= not pi0142 and not w7107;
w7501 <= pi0142 and not w7021;
w7502 <= not pi0140 and not w7501;
w7503 <= not w7500 and w7502;
w7504 <= pi0142 and not w7016;
w7505 <= not pi0142 and not w7104;
w7506 <= pi0140 and not w7504;
w7507 <= not w7505 and w7506;
w7508 <= not w7503 and not w7507;
w7509 <= pi0181 and not w7508;
w7510 <= pi0144 and not w7509;
w7511 <= not w7499 and w7510;
w7512 <= not w6971 and w7167;
w7513 <= w3760 and not w7512;
w7514 <= pi0142 and not w7513;
w7515 <= not w7074 and w7514;
w7516 <= not pi0142 and w7092;
w7517 <= not pi0140 and not w7515;
w7518 <= not w7516 and w7517;
w7519 <= pi0142 and not w7208;
w7520 <= not w7074 and w7519;
w7521 <= not pi0142 and not w7097;
w7522 <= pi0140 and not w7520;
w7523 <= not w7521 and w7522;
w7524 <= not w7518 and not w7523;
w7525 <= not pi0181 and not w7524;
w7526 <= pi0142 and not w6977;
w7527 <= not pi0142 and not w7125;
w7528 <= not pi0140 and not w7526;
w7529 <= not w7527 and w7528;
w7530 <= not pi0142 and w7111;
w7531 <= pi0142 and not w6993;
w7532 <= pi0140 and not w7530;
w7533 <= not w7531 and w7532;
w7534 <= not w7529 and not w7533;
w7535 <= pi0181 and not w7534;
w7536 <= not pi0144 and not w7525;
w7537 <= not w7535 and w7536;
w7538 <= not pi0299 and not w7537;
w7539 <= not w7511 and w7538;
w7540 <= pi0146 and w7146;
w7541 <= not pi0146 and not w7160;
w7542 <= pi0161 and not w7540;
w7543 <= not w7541 and w7542;
w7544 <= pi0146 and not w7141;
w7545 <= not pi0146 and not w7155;
w7546 <= not pi0161 and not w7544;
w7547 <= not w7545 and w7546;
w7548 <= not pi0162 and not w7543;
w7549 <= not w7547 and w7548;
w7550 <= not pi0146 and w7195;
w7551 <= pi0146 and not w7189;
w7552 <= not pi0161 and not w7550;
w7553 <= not w7551 and w7552;
w7554 <= pi0146 and not w7187;
w7555 <= not pi0146 and not w7193;
w7556 <= pi0161 and not w7554;
w7557 <= not w7555 and w7556;
w7558 <= pi0162 and not w7553;
w7559 <= not w7557 and w7558;
w7560 <= w7357 and not w7549;
w7561 <= not w7559 and w7560;
w7562 <= not w7488 and not w7561;
w7563 <= not w7539 and w7562;
w7564 <= pi0232 and not w7563;
w7565 <= not w7224 and not w7564;
w7566 <= w93 and not w7565;
w7567 <= pi0144 and w6870;
w7568 <= not pi0144 and not w6867;
w7569 <= not w6901 and w7568;
w7570 <= w7335 and not w7569;
w7571 <= not w7567 and w7570;
w7572 <= not w6867 and not w6878;
w7573 <= w7339 and not w7568;
w7574 <= not w7572 and w7573;
w7575 <= not w7571 and not w7574;
w7576 <= pi0232 and not w7575;
w7577 <= not w6873 and not w7576;
w7578 <= not pi0038 and not w7577;
w7579 <= not pi0161 and w6890;
w7580 <= not w6864 and not w7579;
w7581 <= w6599 and not w7580;
w7582 <= w6854 and w7329;
w7583 <= not w7581 and w7582;
w7584 <= pi0161 and w6883;
w7585 <= w6599 and w6860;
w7586 <= not w7584 and w7585;
w7587 <= w6854 and w7323;
w7588 <= not w7586 and w7587;
w7589 <= not w7583 and not w7588;
w7590 <= pi0232 and not w7589;
w7591 <= not w7578 and not w7590;
w7592 <= pi0039 and not w7591;
w7593 <= not pi0087 and not w7322;
w7594 <= not w7592 and w7593;
w7595 <= not w7566 and w7594;
w7596 <= pi0038 and not w7310;
w7597 <= not w6829 and not w7596;
w7598 <= pi0087 and w7597;
w7599 <= not pi0100 and not w7598;
w7600 <= not w7595 and w7599;
w7601 <= not w7296 and not w7600;
w7602 <= w132 and not w7601;
w7603 <= not pi0038 and w7411;
w7604 <= w5036 and not w7603;
w7605 <= w6845 and not w7604;
w7606 <= w7597 and not w7605;
w7607 <= not pi0100 and not w7606;
w7608 <= not w7296 and not w7607;
w7609 <= w6768 and not w7608;
w7610 <= not w7297 and not w7609;
w7611 <= not w7602 and w7610;
w7612 <= not pi0054 and not w7611;
w7613 <= not w7314 and not w7612;
w7614 <= not pi0074 and not w7613;
w7615 <= w7306 and not w7614;
w7616 <= w92 and not w7465;
w7617 <= not w7615 and w7616;
w7618 <= not w7447 and not w7617;
w7619 <= not w7276 and not w7618;
w7620 <= not pi0034 and w7619;
w7621 <= not pi0033 and not pi0954;
w7622 <= not w7444 and not w7621;
w7623 <= not w7620 and w7622;
w7624 <= not pi0034 and not w6541;
w7625 <= w7443 and w7624;
w7626 <= w7619 and not w7624;
w7627 <= w7621 and not w7625;
w7628 <= not w7626 and w7627;
w7629 <= not w7623 and not w7628;
w7630 <= w92 and w135;
w7631 <= w6525 and w7630;
w7632 <= not pi0055 and w7631;
w7633 <= pi0059 and not w7632;
w7634 <= not pi0024 and w4903;
w7635 <= pi0054 and not w7634;
w7636 <= pi0137 and w6447;
w7637 <= w486 and w493;
w7638 <= w4980 and not w7637;
w7639 <= pi0683 and w7638;
w7640 <= pi0252 and not w3837;
w7641 <= not w7639 and w7640;
w7642 <= pi0146 and w5034;
w7643 <= pi0142 and w5033;
w7644 <= not w7642 and not w7643;
w7645 <= not w5035 and w7644;
w7646 <= not w7641 and not w7645;
w7647 <= not w5037 and not w7646;
w7648 <= not w6449 and not w7647;
w7649 <= w3826 and not w6452;
w7650 <= not w7641 and w7649;
w7651 <= not w7648 and not w7650;
w7652 <= w6450 and not w7651;
w7653 <= not w7636 and not w7652;
w7654 <= w6445 and not w7653;
w7655 <= not pi0090 and w3701;
w7656 <= not pi0093 and not w7655;
w7657 <= not w3720 and not w7656;
w7658 <= not pi0035 and not w7657;
w7659 <= pi0035 and not w478;
w7660 <= w6501 and not w7659;
w7661 <= not w7658 and w7660;
w7662 <= not pi0032 and w7661;
w7663 <= pi0032 and not pi0093;
w7664 <= w6458 and w7663;
w7665 <= w4995 and w7664;
w7666 <= not w7662 and not w7665;
w7667 <= not pi0095 and not w3732;
w7668 <= not w7666 and w7667;
w7669 <= w3732 and not w7658;
w7670 <= not pi0137 and not w3732;
w7671 <= w487 and w5042;
w7672 <= not w4988 and not w7670;
w7673 <= w7671 and w7672;
w7674 <= not pi0122 and not w3841;
w7675 <= w4988 and not w7670;
w7676 <= w7674 and w7675;
w7677 <= not w7673 and not w7676;
w7678 <= not w7669 and w7677;
w7679 <= w267 and w6495;
w7680 <= w7658 and not w7679;
w7681 <= w81 and w7660;
w7682 <= not w7680 and w7681;
w7683 <= not w7678 and w7682;
w7684 <= not w306 and not w7661;
w7685 <= pi1082 and w81;
w7686 <= not w7684 and w7685;
w7687 <= not pi0038 and not w7683;
w7688 <= not w7686 and w7687;
w7689 <= not w7668 and w7688;
w7690 <= pi0038 and not w6525;
w7691 <= not pi0039 and not pi0100;
w7692 <= not w7690 and w7691;
w7693 <= not w7689 and w7692;
w7694 <= not w7654 and not w7693;
w7695 <= w96 and not w7694;
w7696 <= pi0137 and w6468;
w7697 <= not w3845 and w7696;
w7698 <= not w6527 and not w7697;
w7699 <= w6530 and not w7698;
w7700 <= w6525 and w7699;
w7701 <= not w7695 and not w7700;
w7702 <= not pi0092 and not w7701;
w7703 <= not pi0054 and not w7702;
w7704 <= w92 and w6442;
w7705 <= not w7635 and w7704;
w7706 <= not w7703 and w7705;
w7707 <= not pi0059 and not w7706;
w7708 <= not pi0057 and not w7633;
w7709 <= not w7707 and w7708;
w7710 <= w280 and w334;
w7711 <= not pi0065 and w25;
w7712 <= w50 and w7711;
w7713 <= w6644 and w7712;
w7714 <= not pi0069 and w7713;
w7715 <= not pi0067 and not pi0071;
w7716 <= not pi0083 and w365;
w7717 <= pi0036 and not pi0103;
w7718 <= w7715 and w7717;
w7719 <= w7714 and w7718;
w7720 <= w7716 and w7719;
w7721 <= w7710 and w7720;
w7722 <= not pi0058 and w5085;
w7723 <= not w7721 and not w7722;
w7724 <= w267 and w4042;
w7725 <= w3733 and w7724;
w7726 <= w95 and w4989;
w7727 <= w936 and w7726;
w7728 <= not pi0092 and w7727;
w7729 <= w7725 and w7728;
w7730 <= w3841 and w7729;
w7731 <= not w7723 and w7730;
w7732 <= not pi0081 and not w352;
w7733 <= not pi0045 and not pi0073;
w7734 <= w6483 and w7733;
w7735 <= not pi0071 and w50;
w7736 <= not pi0104 and w35;
w7737 <= w7735 and w7736;
w7738 <= not pi0048 and not pi0065;
w7739 <= not pi0082 and not pi0084;
w7740 <= pi0089 and w7739;
w7741 <= w7738 and w7740;
w7742 <= w7734 and w7741;
w7743 <= w6643 and w7742;
w7744 <= w7737 and w7743;
w7745 <= pi0332 and w7744;
w7746 <= not pi0064 and not w7745;
w7747 <= w4042 and w7031;
w7748 <= w64 and w7747;
w7749 <= w71 and w7748;
w7750 <= not pi0039 and not pi0841;
w7751 <= w28 and w7750;
w7752 <= not w7746 and w7751;
w7753 <= w7749 and w7752;
w7754 <= w7732 and w7753;
w7755 <= not pi0038 and not w7754;
w7756 <= not pi0039 and w82;
w7757 <= pi0024 and w7756;
w7758 <= w272 and w7757;
w7759 <= pi0038 and not w7758;
w7760 <= w134 and w4989;
w7761 <= not w7755 and w7760;
w7762 <= not w7759 and w7761;
w7763 <= not pi0038 and w7760;
w7764 <= pi0786 and not pi1082;
w7765 <= not pi0984 and not w495;
w7766 <= pi0835 and not w7765;
w7767 <= w3746 and not w7766;
w7768 <= w3780 and not w7767;
w7769 <= pi1093 and w7768;
w7770 <= w3747 and w3943;
w7771 <= not w7769 and w7770;
w7772 <= not pi0223 and w7771;
w7773 <= w3761 and w7768;
w7774 <= w7770 and not w7773;
w7775 <= w3768 and w7774;
w7776 <= not w3790 and w7768;
w7777 <= w7770 and not w7776;
w7778 <= not w3768 and w7777;
w7779 <= not pi0299 and not w7775;
w7780 <= not w7778 and w7779;
w7781 <= not w7772 and w7780;
w7782 <= not pi0215 and w7771;
w7783 <= w3805 and w7774;
w7784 <= not w3805 and w7777;
w7785 <= pi0299 and not w7783;
w7786 <= not w7784 and w7785;
w7787 <= not w7782 and w7786;
w7788 <= not w7764 and not w7781;
w7789 <= not w7787 and w7788;
w7790 <= w3416 and not w3807;
w7791 <= w1033 and not w3770;
w7792 <= not w7790 and not w7791;
w7793 <= w3841 and w7764;
w7794 <= not w7792 and w7793;
w7795 <= w3945 and w7794;
w7796 <= not w7789 and not w7795;
w7797 <= pi0039 and not w7796;
w7798 <= not pi0039 and not pi0095;
w7799 <= w3732 and w4049;
w7800 <= not pi0986 and not w3841;
w7801 <= pi0252 and not w7800;
w7802 <= pi0314 and not w7801;
w7803 <= pi0108 and w277;
w7804 <= w336 and w7803;
w7805 <= not pi0841 and w57;
w7806 <= w283 and w7805;
w7807 <= w277 and not w337;
w7808 <= w6484 and w6639;
w7809 <= not pi0065 and not pi0069;
w7810 <= w7808 and w7809;
w7811 <= pi0048 and not pi0049;
w7812 <= not pi0068 and not pi0082;
w7813 <= w7811 and w7812;
w7814 <= w7733 and w7813;
w7815 <= w6473 and w6477;
w7816 <= w6641 and w7815;
w7817 <= w7810 and w7814;
w7818 <= w7816 and w7817;
w7819 <= w7737 and w7818;
w7820 <= not pi0097 and w7806;
w7821 <= w7819 and w7820;
w7822 <= w7807 and w7821;
w7823 <= not pi0047 and not w7804;
w7824 <= not w7822 and w7823;
w7825 <= w3714 and w7802;
w7826 <= not w7824 and w7825;
w7827 <= not pi0047 and not pi0841;
w7828 <= w7819 and w7827;
w7829 <= not w323 and not w7828;
w7830 <= w63 and w263;
w7831 <= not w7802 and w7830;
w7832 <= not w7829 and w7831;
w7833 <= not w7826 and not w7832;
w7834 <= w267 and not w7833;
w7835 <= not pi0035 and not w7834;
w7836 <= pi0035 and not w4046;
w7837 <= w71 and not w7836;
w7838 <= w73 and w7837;
w7839 <= not w7835 and w7838;
w7840 <= not w7799 and not w7839;
w7841 <= w7798 and not w7840;
w7842 <= not w7797 and not w7841;
w7843 <= w7763 and not w7842;
w7844 <= not pi0093 and pi0102;
w7845 <= w24 and w7844;
w7846 <= w27 and w7845;
w7847 <= w3733 and w7846;
w7848 <= w64 and w7847;
w7849 <= w53 and w7848;
w7850 <= w4042 and w7849;
w7851 <= pi1082 and not w7850;
w7852 <= w81 and not w974;
w7853 <= not pi0040 and not w7849;
w7854 <= w7852 and not w7853;
w7855 <= not pi1082 and not w7854;
w7856 <= w7728 and not w7851;
w7857 <= not w7855 and w7856;
w7858 <= not pi0189 and w3760;
w7859 <= pi0144 and w7858;
w7860 <= not pi0174 and w7859;
w7861 <= not pi0299 and not w7860;
w7862 <= not pi0166 and w3760;
w7863 <= pi0161 and w7862;
w7864 <= not pi0152 and w7863;
w7865 <= not w5033 and not w7864;
w7866 <= pi0232 and not w7861;
w7867 <= not w7865 and w7866;
w7868 <= not pi0072 and not w7867;
w7869 <= pi0039 and not w7868;
w7870 <= not pi0041 and not pi0072;
w7871 <= not pi0039 and not w7870;
w7872 <= not w7869 and not w7871;
w7873 <= not w183 and w7872;
w7874 <= not w5069 and not w7870;
w7875 <= not w487 and w7870;
w7876 <= w5069 and not w7875;
w7877 <= not pi0041 and pi0072;
w7878 <= w487 and not w7877;
w7879 <= not pi0044 and w84;
w7880 <= not pi0101 and w7879;
w7881 <= w5042 and w7880;
w7882 <= w5040 and w7881;
w7883 <= pi0041 and not w7882;
w7884 <= not pi0099 and w3835;
w7885 <= not pi0072 and pi0101;
w7886 <= not pi0041 and not w7885;
w7887 <= pi0252 and w4042;
w7888 <= not pi0024 and w272;
w7889 <= w5042 and w7887;
w7890 <= w7888 and w7889;
w7891 <= not pi0044 and w7890;
w7892 <= w7886 and w7891;
w7893 <= not w7884 and w7892;
w7894 <= w7878 and not w7893;
w7895 <= not w7883 and w7894;
w7896 <= w7876 and not w7895;
w7897 <= not w7874 and not w7896;
w7898 <= not pi0039 and not w7897;
w7899 <= w183 and not w7869;
w7900 <= not w7898 and w7899;
w7901 <= pi0075 and not w7873;
w7902 <= not w7900 and w7901;
w7903 <= not w171 and w7871;
w7904 <= not pi0228 and w7870;
w7905 <= w272 and w4042;
w7906 <= not pi0044 and w7905;
w7907 <= w7886 and w7906;
w7908 <= not w7877 and not w7907;
w7909 <= pi0041 and not w7880;
w7910 <= pi0228 and w7908;
w7911 <= not w7909 and w7910;
w7912 <= w188 and not w7904;
w7913 <= not w7911 and w7912;
w7914 <= pi0087 and not w7903;
w7915 <= not w7869 and w7914;
w7916 <= not w7913 and w7915;
w7917 <= pi0038 and not w7872;
w7918 <= pi0041 and not w7881;
w7919 <= w487 and not w7884;
w7920 <= not w7878 and not w7919;
w7921 <= not pi0072 and not w5042;
w7922 <= not w7908 and not w7921;
w7923 <= not w7884 and w7922;
w7924 <= not w7918 and not w7920;
w7925 <= not w7923 and w7924;
w7926 <= w7876 and not w7925;
w7927 <= not w7874 and not w7926;
w7928 <= not pi0039 and not w7927;
w7929 <= not w7869 and not w7928;
w7930 <= w3848 and not w7929;
w7931 <= pi0287 and w84;
w7932 <= w7867 and w7931;
w7933 <= not w7868 and not w7932;
w7934 <= pi0039 and not w7933;
w7935 <= pi0901 and not pi0959;
w7936 <= not pi0480 and pi0949;
w7937 <= w280 and w343;
w7938 <= w271 and w7937;
w7939 <= not w7936 and w7938;
w7940 <= w271 and w7936;
w7941 <= w263 and not w322;
w7942 <= not pi0109 and w4014;
w7943 <= w343 and w7942;
w7944 <= not pi0110 and not w7943;
w7945 <= not pi0047 and w7940;
w7946 <= w7941 and w7945;
w7947 <= not w7944 and w7946;
w7948 <= w7935 and not w7939;
w7949 <= not w7947 and w7948;
w7950 <= w264 and w321;
w7951 <= pi0110 and w7950;
w7952 <= w7940 and w7951;
w7953 <= not w7935 and not w7952;
w7954 <= not pi0250 and pi0252;
w7955 <= w4042 and w7954;
w7956 <= not w7953 and w7955;
w7957 <= not w7949 and w7956;
w7958 <= not pi0072 and w7957;
w7959 <= w7725 and w7951;
w7960 <= w7936 and not w7954;
w7961 <= w7959 and w7960;
w7962 <= not w7958 and not w7961;
w7963 <= not pi0044 and not w7962;
w7964 <= not pi0101 and w7963;
w7965 <= pi0041 and not w7964;
w7966 <= pi0044 and pi0072;
w7967 <= w4042 and not w7954;
w7968 <= w7952 and w7967;
w7969 <= not pi0072 and not w7968;
w7970 <= not w7957 and w7969;
w7971 <= not pi0044 and not w7970;
w7972 <= not w7966 and not w7971;
w7973 <= not pi0101 and w7972;
w7974 <= w7886 and not w7973;
w7975 <= not w7965 and not w7974;
w7976 <= not pi0228 and not w7975;
w7977 <= not pi0072 and not w5014;
w7978 <= not w5020 and w7977;
w7979 <= w4042 and not w5018;
w7980 <= not w5017 and w7979;
w7981 <= not pi0072 and w5020;
w7982 <= not w7980 and w7981;
w7983 <= not pi1093 and not w7978;
w7984 <= not w7982 and w7983;
w7985 <= w7977 and not w7984;
w7986 <= not pi0044 and not w7985;
w7987 <= not w7966 and not w7986;
w7988 <= not pi0101 and w7987;
w7989 <= w7886 and not w7988;
w7990 <= w5014 and not w5020;
w7991 <= not pi1093 and not w5022;
w7992 <= not w7990 and w7991;
w7993 <= not pi0044 and not w7992;
w7994 <= pi1093 and not w5014;
w7995 <= w7993 and not w7994;
w7996 <= not pi0101 and w7995;
w7997 <= pi0041 and not w7996;
w7998 <= not w487 and not w7997;
w7999 <= not w7989 and w7998;
w8000 <= w498 and not w5006;
w8001 <= w500 and w8000;
w8002 <= not w5085 and not w8001;
w8003 <= w24 and not w8002;
w8004 <= w4997 and not w8003;
w8005 <= w4994 and not w8004;
w8006 <= not pi0051 and not w8005;
w8007 <= not w310 and not w8006;
w8008 <= not pi0096 and not w8007;
w8009 <= w7979 and w7981;
w8010 <= not w8008 and w8009;
w8011 <= not w7990 and not w8010;
w8012 <= pi1093 and w8011;
w8013 <= w7993 and not w8012;
w8014 <= not pi0101 and w8013;
w8015 <= pi0041 and not w8014;
w8016 <= not pi0072 and w8011;
w8017 <= pi1093 and not w8016;
w8018 <= not w7984 and not w8017;
w8019 <= not pi0044 and not w8018;
w8020 <= not w7966 and not w8019;
w8021 <= not pi0101 and w8020;
w8022 <= w7886 and not w8021;
w8023 <= w487 and not w8022;
w8024 <= not w8015 and w8023;
w8025 <= pi0228 and not w7999;
w8026 <= not w8024 and w8025;
w8027 <= not pi0039 and not w7976;
w8028 <= not w8026 and w8027;
w8029 <= w171 and not w7934;
w8030 <= not w8028 and w8029;
w8031 <= not pi0087 and not w7917;
w8032 <= not w7930 and w8031;
w8033 <= not w8030 and w8032;
w8034 <= not pi0075 and not w7916;
w8035 <= not w8033 and w8034;
w8036 <= not w7902 and not w8035;
w8037 <= w4992 and not w8036;
w8038 <= not w4992 and not w7872;
w8039 <= w4989 and not w8038;
w8040 <= not w8037 and w8039;
w8041 <= pi0039 and pi0232;
w8042 <= w7864 and w8041;
w8043 <= not pi0072 and not w7871;
w8044 <= not w4989 and w8043;
w8045 <= not w8042 and w8044;
w8046 <= not w8040 and not w8045;
w8047 <= pi0211 and pi0214;
w8048 <= pi0212 and w8047;
w8049 <= not pi0219 and not w8048;
w8050 <= pi0207 and pi0208;
w8051 <= pi0042 and not pi0072;
w8052 <= not w183 and w8051;
w8053 <= not w5069 and not w8051;
w8054 <= not pi0115 and w487;
w8055 <= w8051 and not w8054;
w8056 <= w5069 and not w8055;
w8057 <= pi0114 and not w8051;
w8058 <= w8054 and not w8057;
w8059 <= w3829 and w7891;
w8060 <= not pi0113 and w8059;
w8061 <= not pi0116 and w8060;
w8062 <= w8051 and not w8061;
w8063 <= w3828 and w7880;
w8064 <= w3832 and w8063;
w8065 <= w5042 and w8064;
w8066 <= not pi0114 and not w3831;
w8067 <= w8065 and w8066;
w8068 <= w5040 and w8067;
w8069 <= not pi0042 and w8068;
w8070 <= not pi0114 and not w8062;
w8071 <= not w8069 and w8070;
w8072 <= w8058 and not w8071;
w8073 <= w8056 and not w8072;
w8074 <= w183 and not w8053;
w8075 <= not w8073 and w8074;
w8076 <= not pi0039 and not w8052;
w8077 <= not w8075 and w8076;
w8078 <= not pi0072 and pi0199;
w8079 <= not pi0232 and not w8078;
w8080 <= not pi0299 and not w8079;
w8081 <= not pi0072 and not w7858;
w8082 <= pi0199 and w8081;
w8083 <= pi0232 and not w8082;
w8084 <= w8080 and not w8083;
w8085 <= not pi0166 and w5036;
w8086 <= not pi0072 and not w8085;
w8087 <= pi0299 and w8086;
w8088 <= pi0039 and not w8087;
w8089 <= not w8084 and w8088;
w8090 <= not w8077 and not w8089;
w8091 <= pi0075 and not w8090;
w8092 <= not pi0039 and not w8051;
w8093 <= not w171 and w8092;
w8094 <= w3829 and w7906;
w8095 <= pi0228 and w8094;
w8096 <= w3834 and w8095;
w8097 <= w8051 and not w8096;
w8098 <= pi0228 and w8064;
w8099 <= not pi0115 and w8098;
w8100 <= not pi0114 and w8099;
w8101 <= not pi0042 and w8100;
w8102 <= w188 and not w8097;
w8103 <= not w8101 and w8102;
w8104 <= pi0087 and not w8093;
w8105 <= not w8103 and w8104;
w8106 <= not w8089 and w8105;
w8107 <= pi0115 and not w8051;
w8108 <= pi0042 and not pi0114;
w8109 <= pi0072 and pi0116;
w8110 <= pi0072 and pi0113;
w8111 <= pi0072 and not w3828;
w8112 <= not pi0099 and w7974;
w8113 <= not w8111 and not w8112;
w8114 <= not pi0113 and not w8113;
w8115 <= not w8110 and not w8114;
w8116 <= not pi0116 and not w8115;
w8117 <= not w8109 and not w8116;
w8118 <= w8108 and not w8117;
w8119 <= w3828 and w7964;
w8120 <= not pi0113 and w8119;
w8121 <= not pi0116 and w8120;
w8122 <= not pi0042 and not w8121;
w8123 <= not w8057 and not w8122;
w8124 <= not w8118 and w8123;
w8125 <= not pi0115 and not w8124;
w8126 <= not pi0228 and not w8107;
w8127 <= not w8125 and w8126;
w8128 <= not pi0099 and w8022;
w8129 <= not w8111 and not w8128;
w8130 <= not pi0113 and not w8129;
w8131 <= not w8110 and not w8130;
w8132 <= not pi0116 and not w8131;
w8133 <= not w8109 and not w8132;
w8134 <= w8108 and not w8133;
w8135 <= w3828 and w8014;
w8136 <= w3832 and w8135;
w8137 <= not pi0042 and not w8136;
w8138 <= not w8057 and not w8137;
w8139 <= not w8134 and w8138;
w8140 <= w8054 and not w8139;
w8141 <= not pi0115 and not w487;
w8142 <= w3828 and w7996;
w8143 <= w3832 and w8142;
w8144 <= not pi0042 and w8143;
w8145 <= not pi0099 and w7989;
w8146 <= not w8111 and not w8145;
w8147 <= not pi0113 and not w8146;
w8148 <= not w8110 and not w8147;
w8149 <= not pi0116 and not w8148;
w8150 <= not w8109 and not w8149;
w8151 <= pi0042 and w8150;
w8152 <= not pi0114 and not w8144;
w8153 <= not w8151 and w8152;
w8154 <= not w8057 and not w8153;
w8155 <= w8141 and not w8154;
w8156 <= pi0228 and not w8107;
w8157 <= not w8155 and w8156;
w8158 <= not w8140 and w8157;
w8159 <= not pi0039 and not w8127;
w8160 <= not w8158 and w8159;
w8161 <= pi0232 and pi0299;
w8162 <= w7862 and w7931;
w8163 <= not w8086 and w8161;
w8164 <= not w8162 and w8163;
w8165 <= pi0232 and not pi0299;
w8166 <= w3760 and w7931;
w8167 <= not pi0189 and w8166;
w8168 <= not w8081 and not w8167;
w8169 <= pi0199 and not w8168;
w8170 <= w8165 and not w8169;
w8171 <= pi0072 and not pi0232;
w8172 <= pi0299 and not w8171;
w8173 <= w8079 and not w8172;
w8174 <= not w8164 and not w8173;
w8175 <= not w8170 and w8174;
w8176 <= pi0039 and not w8175;
w8177 <= not w8160 and not w8176;
w8178 <= w171 and not w8177;
w8179 <= w3832 and w8094;
w8180 <= not pi0072 and not w8179;
w8181 <= not w7921 and not w8180;
w8182 <= pi0042 and not w8181;
w8183 <= not pi0042 and w8067;
w8184 <= not pi0114 and not w8182;
w8185 <= not w8183 and w8184;
w8186 <= w8058 and not w8185;
w8187 <= w8056 and not w8186;
w8188 <= not w8053 and not w8187;
w8189 <= not pi0039 and not w8188;
w8190 <= not w8089 and not w8189;
w8191 <= w3848 and not w8190;
w8192 <= not w8089 and not w8092;
w8193 <= pi0038 and not w8192;
w8194 <= not pi0087 and not w8193;
w8195 <= not w8191 and w8194;
w8196 <= not w8178 and w8195;
w8197 <= not pi0075 and not w8106;
w8198 <= not w8196 and w8197;
w8199 <= w4992 and not w8091;
w8200 <= not w8198 and w8199;
w8201 <= not w8050 and not w8200;
w8202 <= not pi0072 and pi0200;
w8203 <= not pi0232 and not w8202;
w8204 <= not pi0299 and not w8203;
w8205 <= pi0200 and w8081;
w8206 <= pi0232 and not w8205;
w8207 <= w8204 and not w8206;
w8208 <= pi0039 and not w8207;
w8209 <= not w8084 and w8208;
w8210 <= not w8092 and not w8209;
w8211 <= not w4992 and w8210;
w8212 <= w8050 and not w8211;
w8213 <= w8089 and w8208;
w8214 <= not w8077 and not w8213;
w8215 <= pi0075 and not w8214;
w8216 <= not w8189 and not w8213;
w8217 <= w3848 and not w8216;
w8218 <= pi0038 and not w8210;
w8219 <= not pi0087 and not w8218;
w8220 <= not w8194 and not w8219;
w8221 <= pi0232 and not w8169;
w8222 <= pi0200 and not w8168;
w8223 <= w8221 and not w8222;
w8224 <= not pi0299 and w8223;
w8225 <= w8173 and not w8202;
w8226 <= not w8164 and not w8225;
w8227 <= not w8224 and w8226;
w8228 <= pi0039 and not w8227;
w8229 <= not w8160 and not w8228;
w8230 <= w171 and not w8229;
w8231 <= not w8217 and not w8220;
w8232 <= not w8230 and w8231;
w8233 <= w8104 and not w8213;
w8234 <= not w8103 and w8233;
w8235 <= not pi0075 and not w8234;
w8236 <= not w8232 and w8235;
w8237 <= w4992 and not w8215;
w8238 <= not w8236 and w8237;
w8239 <= w8212 and not w8238;
w8240 <= not w8201 and not w8239;
w8241 <= not w4992 and w8192;
w8242 <= not w8049 and not w8241;
w8243 <= not w8240 and w8242;
w8244 <= pi0039 and not w8084;
w8245 <= not w8077 and not w8244;
w8246 <= pi0075 and not w8245;
w8247 <= w8105 and not w8244;
w8248 <= not w8189 and not w8244;
w8249 <= w3848 and not w8248;
w8250 <= not w8092 and not w8244;
w8251 <= pi0038 and not w8250;
w8252 <= w8080 and not w8221;
w8253 <= pi0039 and not w8252;
w8254 <= not w8160 and not w8253;
w8255 <= w171 and not w8254;
w8256 <= not pi0087 and not w8251;
w8257 <= not w8249 and w8256;
w8258 <= not w8255 and w8257;
w8259 <= not pi0075 and not w8247;
w8260 <= not w8258 and w8259;
w8261 <= w4992 and not w8246;
w8262 <= not w8260 and w8261;
w8263 <= not w4992 and w8250;
w8264 <= not w8050 and not w8263;
w8265 <= not w8262 and w8264;
w8266 <= not w8077 and not w8209;
w8267 <= pi0075 and not w8266;
w8268 <= w8105 and not w8209;
w8269 <= not w8080 and not w8204;
w8270 <= not w8223 and not w8269;
w8271 <= pi0039 and not w8270;
w8272 <= not w8160 and not w8271;
w8273 <= w171 and not w8272;
w8274 <= not w8189 and not w8209;
w8275 <= w3848 and not w8274;
w8276 <= w8219 and not w8275;
w8277 <= not w8273 and w8276;
w8278 <= not pi0075 and not w8268;
w8279 <= not w8277 and w8278;
w8280 <= w4992 and not w8267;
w8281 <= not w8279 and w8280;
w8282 <= w8212 and not w8281;
w8283 <= not w8265 and not w8282;
w8284 <= w8049 and not w8283;
w8285 <= w4989 and not w8243;
w8286 <= not w8284 and w8285;
w8287 <= not w8049 and w8086;
w8288 <= pi0039 and not w8287;
w8289 <= not w4989 and not w8092;
w8290 <= not w8288 and w8289;
w8291 <= not w8286 and not w8290;
w8292 <= pi0043 and not pi0072;
w8293 <= not w5069 and not w8292;
w8294 <= not pi0042 and w3833;
w8295 <= w487 and w8294;
w8296 <= w8292 and not w8295;
w8297 <= w5069 and not w8296;
w8298 <= not pi0072 and not w8061;
w8299 <= pi0043 and w8298;
w8300 <= not pi0043 and pi0052;
w8301 <= w5040 and w8065;
w8302 <= w8300 and w8301;
w8303 <= not w8299 and not w8302;
w8304 <= w8295 and not w8303;
w8305 <= w8297 and not w8304;
w8306 <= not w8293 and not w8305;
w8307 <= not pi0039 and not w8306;
w8308 <= w183 and not w8307;
w8309 <= not pi0039 and not w8292;
w8310 <= not w183 and not w8309;
w8311 <= not w8308 and not w8310;
w8312 <= not w8208 and not w8311;
w8313 <= pi0075 and not w8312;
w8314 <= not w171 and w8309;
w8315 <= not pi0043 and not w8064;
w8316 <= pi0043 and not w8180;
w8317 <= pi0228 and w8294;
w8318 <= not w8316 and w8317;
w8319 <= not w8315 and w8318;
w8320 <= w8292 and not w8317;
w8321 <= w188 and not w8320;
w8322 <= not w8319 and w8321;
w8323 <= pi0087 and not w8314;
w8324 <= not w8322 and w8323;
w8325 <= not w8208 and w8324;
w8326 <= w8065 and w8300;
w8327 <= pi0043 and not w8181;
w8328 <= not w8326 and not w8327;
w8329 <= w8295 and not w8328;
w8330 <= w8297 and not w8329;
w8331 <= not w8293 and not w8330;
w8332 <= not pi0039 and not w8331;
w8333 <= not w8208 and not w8332;
w8334 <= w3848 and not w8333;
w8335 <= not w8208 and not w8309;
w8336 <= pi0038 and not w8335;
w8337 <= pi0232 and not w8222;
w8338 <= w8204 and not w8337;
w8339 <= pi0039 and not w8338;
w8340 <= not pi0228 and not w8121;
w8341 <= not w487 and not w8142;
w8342 <= w487 and not w8135;
w8343 <= not w8341 and not w8342;
w8344 <= w3832 and w8343;
w8345 <= pi0228 and not w8344;
w8346 <= not w8340 and not w8345;
w8347 <= not pi0043 and not w8346;
w8348 <= not w8292 and not w8294;
w8349 <= not w487 and not w8150;
w8350 <= w487 and not w8133;
w8351 <= not w8349 and not w8350;
w8352 <= pi0228 and not w8351;
w8353 <= not pi0228 and not w8117;
w8354 <= not w8352 and not w8353;
w8355 <= pi0043 and w8294;
w8356 <= not w8354 and w8355;
w8357 <= not w8347 and not w8348;
w8358 <= not w8356 and w8357;
w8359 <= not pi0039 and not w8358;
w8360 <= not w8339 and not w8359;
w8361 <= w171 and not w8360;
w8362 <= not pi0087 and not w8336;
w8363 <= not w8334 and w8362;
w8364 <= not w8361 and w8363;
w8365 <= not pi0075 and not w8325;
w8366 <= not w8364 and w8365;
w8367 <= w4992 and not w8313;
w8368 <= not w8366 and w8367;
w8369 <= not w4992 and w8335;
w8370 <= not w8050 and not w8369;
w8371 <= not w8368 and w8370;
w8372 <= not pi0199 and not pi0200;
w8373 <= not pi0299 and not w8372;
w8374 <= not pi0072 and not w8373;
w8375 <= not pi0232 and not w8374;
w8376 <= not pi0299 and not w8375;
w8377 <= w8081 and w8372;
w8378 <= pi0232 and not w8377;
w8379 <= w8376 and not w8378;
w8380 <= pi0039 and not w8379;
w8381 <= not w8309 and not w8380;
w8382 <= not w4992 and w8381;
w8383 <= not w8311 and not w8380;
w8384 <= pi0075 and not w8383;
w8385 <= not w8332 and not w8380;
w8386 <= w3848 and not w8385;
w8387 <= pi0038 and not w8381;
w8388 <= not w8168 and w8372;
w8389 <= pi0232 and not w8388;
w8390 <= w8376 and not w8389;
w8391 <= pi0039 and not w8390;
w8392 <= not w8359 and not w8391;
w8393 <= w171 and not w8392;
w8394 <= not pi0087 and not w8387;
w8395 <= not w8386 and w8394;
w8396 <= not w8393 and w8395;
w8397 <= not w94 and not w8381;
w8398 <= w8324 and not w8397;
w8399 <= not pi0075 and not w8398;
w8400 <= not w8396 and w8399;
w8401 <= w4992 and not w8384;
w8402 <= not w8400 and w8401;
w8403 <= w8050 and not w8382;
w8404 <= not w8402 and w8403;
w8405 <= not w8371 and not w8404;
w8406 <= pi0212 and pi0214;
w8407 <= not pi0211 and not pi0219;
w8408 <= w8406 and not w8407;
w8409 <= not pi0211 and not w8406;
w8410 <= not w8408 and not w8409;
w8411 <= not w8405 and not w8410;
w8412 <= w8088 and not w8207;
w8413 <= not w8311 and not w8412;
w8414 <= pi0075 and not w8413;
w8415 <= w8324 and not w8412;
w8416 <= not w8332 and not w8412;
w8417 <= w3848 and not w8416;
w8418 <= not w8309 and not w8412;
w8419 <= pi0038 and not w8418;
w8420 <= w8165 and not w8222;
w8421 <= not w8172 and w8203;
w8422 <= not w8164 and not w8421;
w8423 <= not w8420 and w8422;
w8424 <= pi0039 and not w8423;
w8425 <= not w8359 and not w8424;
w8426 <= w171 and not w8425;
w8427 <= not pi0087 and not w8419;
w8428 <= not w8417 and w8427;
w8429 <= not w8426 and w8428;
w8430 <= not pi0075 and not w8415;
w8431 <= not w8429 and w8430;
w8432 <= w4992 and not w8414;
w8433 <= not w8431 and w8432;
w8434 <= not w4992 and w8418;
w8435 <= not w8050 and not w8434;
w8436 <= not w8433 and w8435;
w8437 <= not w8087 and w8380;
w8438 <= not w8309 and not w8437;
w8439 <= not w4992 and w8438;
w8440 <= not w8311 and not w8437;
w8441 <= pi0075 and not w8440;
w8442 <= w8324 and not w8437;
w8443 <= not w8332 and not w8437;
w8444 <= w3848 and not w8443;
w8445 <= pi0038 and not w8438;
w8446 <= w8165 and not w8388;
w8447 <= not w8164 and not w8375;
w8448 <= not w8446 and w8447;
w8449 <= pi0039 and not w8448;
w8450 <= not w8359 and not w8449;
w8451 <= w171 and not w8450;
w8452 <= not pi0087 and not w8445;
w8453 <= not w8444 and w8452;
w8454 <= not w8451 and w8453;
w8455 <= not pi0075 and not w8442;
w8456 <= not w8454 and w8455;
w8457 <= w4992 and not w8441;
w8458 <= not w8456 and w8457;
w8459 <= w8050 and not w8439;
w8460 <= not w8458 and w8459;
w8461 <= not w8436 and not w8460;
w8462 <= w8410 and not w8461;
w8463 <= w4989 and not w8411;
w8464 <= not w8462 and w8463;
w8465 <= w8086 and w8410;
w8466 <= pi0039 and not w8465;
w8467 <= not w4989 and not w8309;
w8468 <= not w8466 and w8467;
w8469 <= not w8464 and not w8468;
w8470 <= not pi0072 and w5037;
w8471 <= pi0039 and not w8470;
w8472 <= pi0044 and not pi0072;
w8473 <= not pi0039 and not w8472;
w8474 <= not w8471 and not w8473;
w8475 <= not w183 and w8474;
w8476 <= not w5069 and not w8472;
w8477 <= not pi0039 and not w8476;
w8478 <= not w487 and w8472;
w8479 <= w5069 and not w8478;
w8480 <= w5157 and not w7966;
w8481 <= w5042 and w7879;
w8482 <= w5040 and w8481;
w8483 <= pi0044 and not w7890;
w8484 <= not w8482 and not w8483;
w8485 <= w8480 and not w8484;
w8486 <= w8479 and not w8485;
w8487 <= w8477 and not w8486;
w8488 <= pi0039 and w5037;
w8489 <= not pi0072 and w8488;
w8490 <= not w8487 and not w8489;
w8491 <= w183 and not w8490;
w8492 <= pi0075 and not w8475;
w8493 <= not w8491 and w8492;
w8494 <= pi0228 and w171;
w8495 <= w7879 and w8494;
w8496 <= w7905 and w8494;
w8497 <= w8472 and not w8496;
w8498 <= not pi0039 and not w8497;
w8499 <= not w8495 and w8498;
w8500 <= pi0087 and not w8471;
w8501 <= not w8499 and w8500;
w8502 <= pi0038 and not w8474;
w8503 <= w5042 and w7905;
w8504 <= pi0044 and not w8503;
w8505 <= not w8481 and not w8504;
w8506 <= w8480 and not w8505;
w8507 <= w8479 and not w8506;
w8508 <= w8477 and not w8507;
w8509 <= w3848 and not w8489;
w8510 <= not w8508 and w8509;
w8511 <= pi0287 and w7905;
w8512 <= not pi0072 and not w8511;
w8513 <= w8488 and w8512;
w8514 <= pi0044 and w7970;
w8515 <= not pi0228 and not w8514;
w8516 <= not w7963 and w8515;
w8517 <= pi0044 and w8018;
w8518 <= w487 and not w8013;
w8519 <= not w8517 and w8518;
w8520 <= pi0044 and w7985;
w8521 <= not w487 and not w7995;
w8522 <= not w8520 and w8521;
w8523 <= not w8519 and not w8522;
w8524 <= pi0228 and not w8523;
w8525 <= not pi0039 and not w8516;
w8526 <= not w8524 and w8525;
w8527 <= w171 and not w8513;
w8528 <= not w8526 and w8527;
w8529 <= not pi0087 and not w8502;
w8530 <= not w8510 and w8529;
w8531 <= not w8528 and w8530;
w8532 <= not pi0075 and not w8501;
w8533 <= not w8531 and w8532;
w8534 <= not w8493 and not w8533;
w8535 <= w4992 and not w8534;
w8536 <= not w4992 and not w8474;
w8537 <= w4989 and not w8536;
w8538 <= not w8535 and w8537;
w8539 <= w202 and w5036;
w8540 <= not pi0072 and w8539;
w8541 <= pi0039 and not w8540;
w8542 <= not w4989 and not w8473;
w8543 <= not w8541 and w8542;
w8544 <= not w8538 and not w8543;
w8545 <= not pi0038 and pi0039;
w8546 <= w7760 and w8545;
w8547 <= pi0979 and w8546;
w8548 <= w3943 and w8547;
w8549 <= not pi0102 and not pi0104;
w8550 <= not pi0111 and w8549;
w8551 <= not pi0049 and not pi0076;
w8552 <= w6472 and w8551;
w8553 <= pi0061 and not pi0082;
w8554 <= not pi0083 and not pi0089;
w8555 <= w8553 and w8554;
w8556 <= w5001 and w6478;
w8557 <= w8555 and w8556;
w8558 <= w7735 and w8550;
w8559 <= w8552 and w8558;
w8560 <= w6475 and w8557;
w8561 <= w7810 and w8560;
w8562 <= w8559 and w8561;
w8563 <= w6498 and w8562;
w8564 <= not pi0841 and w8563;
w8565 <= w265 and w451;
w8566 <= pi0024 and w8565;
w8567 <= not w8564 and not w8566;
w8568 <= w7729 and not w8567;
w8569 <= not pi0082 and w37;
w8570 <= not pi0084 and pi0104;
w8571 <= w368 and w8570;
w8572 <= w7734 and w8571;
w8573 <= w8569 and w8572;
w8574 <= not pi0036 and not w8573;
w8575 <= w6479 and w6644;
w8576 <= not pi0067 and not pi0103;
w8577 <= w50 and w8576;
w8578 <= not pi0098 and w8577;
w8579 <= w8575 and w8578;
w8580 <= not w8574 and w8579;
w8581 <= not w366 and w8580;
w8582 <= not pi0088 and not w8581;
w8583 <= not w434 and w5001;
w8584 <= w317 and not w8582;
w8585 <= w8583 and w8584;
w8586 <= w263 and w8585;
w8587 <= not w7722 and not w8586;
w8588 <= w7725 and not w8587;
w8589 <= w5053 and not w8588;
w8590 <= not pi0036 and w8580;
w8591 <= not pi0088 and not w8590;
w8592 <= w8583 and not w8591;
w8593 <= w7749 and w8592;
w8594 <= not pi0824 and w495;
w8595 <= w8593 and w8594;
w8596 <= not w495 and w8588;
w8597 <= pi0829 and not w8595;
w8598 <= not w8596 and w8597;
w8599 <= not w486 and w8598;
w8600 <= not w8589 and not w8599;
w8601 <= pi1091 and not w8600;
w8602 <= not w4980 and w8588;
w8603 <= not pi0829 and not w8602;
w8604 <= not w8598 and not w8603;
w8605 <= not pi1093 and not w8604;
w8606 <= w4980 and w7725;
w8607 <= not w7723 and w8606;
w8608 <= not w3957 and not w5189;
w8609 <= not w8607 and not w8608;
w8610 <= not w8602 and w8609;
w8611 <= w7728 and not w8610;
w8612 <= not w8605 and w8611;
w8613 <= not w8601 and w8612;
w8614 <= not pi0072 and pi0841;
w8615 <= w268 and w8614;
w8616 <= not pi0051 and w8615;
w8617 <= w7819 and w8616;
w8618 <= w7728 and w8617;
w8619 <= w7748 and w8618;
w8620 <= w27 and w50;
w8621 <= not pi0103 and w367;
w8622 <= w7808 and w8621;
w8623 <= w6472 and w6479;
w8624 <= w8622 and w8623;
w8625 <= not pi0045 and pi0049;
w8626 <= w8550 and w8625;
w8627 <= w8620 and w8626;
w8628 <= w8624 and w8627;
w8629 <= w8569 and w8628;
w8630 <= w269 and w6498;
w8631 <= w8629 and w8630;
w8632 <= w7724 and w8615;
w8633 <= w8631 and w8632;
w8634 <= not pi0074 and not w8633;
w8635 <= pi0074 and not w6525;
w8636 <= w4926 and w4989;
w8637 <= not w8634 and w8636;
w8638 <= not w8635 and w8637;
w8639 <= pi0024 and w6460;
w8640 <= not w7937 and not w8639;
w8641 <= not pi0252 and not w6451;
w8642 <= pi0252 and w6468;
w8643 <= not w8641 and not w8642;
w8644 <= pi0024 and not pi0094;
w8645 <= not w6462 and w8644;
w8646 <= w7725 and w8643;
w8647 <= not w8645 and w8646;
w8648 <= not w8640 and w8647;
w8649 <= w525 and w5013;
w8650 <= pi0024 and not pi0090;
w8651 <= w8649 and w8650;
w8652 <= not w8643 and w8651;
w8653 <= w6464 and w8652;
w8654 <= not w8648 and not w8653;
w8655 <= not pi0100 and not w8654;
w8656 <= pi0100 and not w3826;
w8657 <= w3916 and w8656;
w8658 <= not w8655 and not w8657;
w8659 <= w93 and w96;
w8660 <= not w8658 and w8659;
w8661 <= w3845 and w6530;
w8662 <= w6526 and w8661;
w8663 <= not w8660 and not w8662;
w8664 <= w6444 and not w8663;
w8665 <= w6645 and w8620;
w8666 <= w30 and w8665;
w8667 <= not pi0069 and w8666;
w8668 <= w367 and w8667;
w8669 <= w263 and w7729;
w8670 <= w317 and w8669;
w8671 <= w370 and w8668;
w8672 <= w8670 and w8671;
w8673 <= not pi0219 and w8409;
w8674 <= pi0052 and not pi0072;
w8675 <= not pi0039 and not w8674;
w8676 <= not w8088 and not w8675;
w8677 <= not w4992 and not w8676;
w8678 <= not w8164 and w8172;
w8679 <= pi0039 and not w8678;
w8680 <= w3830 and w3833;
w8681 <= not w8674 and not w8680;
w8682 <= not pi0052 and w8121;
w8683 <= pi0052 and w8117;
w8684 <= w8680 and not w8682;
w8685 <= not w8683 and w8684;
w8686 <= not pi0228 and not w8681;
w8687 <= not w8685 and w8686;
w8688 <= not pi0114 and w3830;
w8689 <= not pi0052 and w8136;
w8690 <= pi0052 and w8133;
w8691 <= w8054 and not w8689;
w8692 <= not w8690 and w8691;
w8693 <= not pi0052 and w8143;
w8694 <= pi0052 and w8150;
w8695 <= w8141 and not w8693;
w8696 <= not w8694 and w8695;
w8697 <= not w8692 and not w8696;
w8698 <= w8688 and not w8697;
w8699 <= pi0228 and not w8681;
w8700 <= not w8698 and w8699;
w8701 <= not pi0039 and not w8687;
w8702 <= not w8700 and w8701;
w8703 <= not w8679 and not w8702;
w8704 <= w171 and not w8703;
w8705 <= pi0038 and not w8676;
w8706 <= w5069 and w8054;
w8707 <= w8688 and w8706;
w8708 <= w5042 and w8707;
w8709 <= w8179 and w8708;
w8710 <= w8674 and not w8709;
w8711 <= not pi0039 and not w8710;
w8712 <= not w8088 and not w8711;
w8713 <= w3848 and not w8712;
w8714 <= not w8705 and not w8713;
w8715 <= not w8704 and w8714;
w8716 <= not pi0087 and not w8715;
w8717 <= not w171 and w8676;
w8718 <= pi0087 and not w8717;
w8719 <= pi0228 and w8680;
w8720 <= not pi0052 and w8064;
w8721 <= pi0052 and w8180;
w8722 <= not w8720 and not w8721;
w8723 <= w8719 and not w8722;
w8724 <= w8674 and not w8719;
w8725 <= not w8723 and not w8724;
w8726 <= not pi0039 and w8725;
w8727 <= w171 and not w8088;
w8728 <= not w8726 and w8727;
w8729 <= w8718 and not w8728;
w8730 <= w8050 and not w8729;
w8731 <= not w8716 and w8730;
w8732 <= not w8380 and not w8675;
w8733 <= not w171 and w8732;
w8734 <= w171 and not w8437;
w8735 <= not w8726 and w8734;
w8736 <= w8718 and not w8733;
w8737 <= not w8735 and w8736;
w8738 <= not w8449 and not w8702;
w8739 <= w171 and not w8738;
w8740 <= not w8437 and not w8711;
w8741 <= w3848 and not w8740;
w8742 <= pi0038 and not w8732;
w8743 <= not w8676 and w8742;
w8744 <= not w8741 and not w8743;
w8745 <= not w8739 and w8744;
w8746 <= not pi0087 and not w8745;
w8747 <= not w8050 and not w8737;
w8748 <= not w8746 and w8747;
w8749 <= not w8731 and not w8748;
w8750 <= not pi0075 and not w8749;
w8751 <= w8061 and w8707;
w8752 <= w183 and w8751;
w8753 <= not pi0039 and w8674;
w8754 <= not w8752 and w8753;
w8755 <= not pi0039 and not w8754;
w8756 <= not w8050 and w8437;
w8757 <= w8050 and w8088;
w8758 <= pi0075 and not w8757;
w8759 <= not w8756 and w8758;
w8760 <= not w8755 and w8759;
w8761 <= w4992 and not w8760;
w8762 <= not w8750 and w8761;
w8763 <= w8673 and not w8677;
w8764 <= not w8762 and w8763;
w8765 <= not w4992 and not w8050;
w8766 <= w8732 and w8765;
w8767 <= not w4992 and not w8753;
w8768 <= pi0075 and w8754;
w8769 <= pi0100 and not w8753;
w8770 <= pi0038 and not w8753;
w8771 <= not pi0038 and w8725;
w8772 <= not w8770 and not w8771;
w8773 <= not pi0100 and not w8772;
w8774 <= not pi0100 and w8545;
w8775 <= pi0087 and not w8774;
w8776 <= not w8769 and w8775;
w8777 <= not w8773 and w8776;
w8778 <= pi0100 and not w8710;
w8779 <= not pi0100 and w8702;
w8780 <= not pi0039 and not w8778;
w8781 <= not w8779 and w8780;
w8782 <= not pi0038 and not w8781;
w8783 <= not pi0087 and not w8770;
w8784 <= not w8782 and w8783;
w8785 <= not w8777 and not w8784;
w8786 <= not pi0075 and not w8785;
w8787 <= w4992 and not w8768;
w8788 <= not w8786 and w8787;
w8789 <= w8050 and not w8767;
w8790 <= not w8788 and w8789;
w8791 <= w171 and not w8380;
w8792 <= not w8726 and w8791;
w8793 <= not w8733 and not w8792;
w8794 <= pi0087 and not w8793;
w8795 <= not w8391 and not w8702;
w8796 <= w171 and not w8795;
w8797 <= not w8380 and not w8711;
w8798 <= w3848 and not w8797;
w8799 <= not pi0087 and not w8742;
w8800 <= not w8798 and w8799;
w8801 <= not w8796 and w8800;
w8802 <= not pi0075 and not w8794;
w8803 <= not w8801 and w8802;
w8804 <= not w183 and w8732;
w8805 <= w8674 and not w8751;
w8806 <= not pi0039 and not w8805;
w8807 <= w183 and not w8380;
w8808 <= not w8806 and w8807;
w8809 <= pi0075 and not w8804;
w8810 <= not w8808 and w8809;
w8811 <= w4992 and not w8050;
w8812 <= not w8810 and w8811;
w8813 <= not w8803 and w8812;
w8814 <= not w8790 and not w8813;
w8815 <= not w8673 and not w8814;
w8816 <= w4989 and not w8766;
w8817 <= not w8764 and w8816;
w8818 <= not w8815 and w8817;
w8819 <= pi0039 and w8673;
w8820 <= w8086 and w8819;
w8821 <= not w4989 and not w8753;
w8822 <= not w8820 and w8821;
w8823 <= not w8818 and not w8822;
w8824 <= not pi0287 and not pi0979;
w8825 <= w3744 and w8824;
w8826 <= pi0039 and not w8825;
w8827 <= pi0024 and w7725;
w8828 <= pi0053 and w283;
w8829 <= w280 and w8828;
w8830 <= w284 and w8829;
w8831 <= w8827 and w8830;
w8832 <= not pi0039 and not w8831;
w8833 <= w7763 and not w8826;
w8834 <= not w8832 and w8833;
w8835 <= not w965 and w8834;
w8836 <= w6460 and w6817;
w8837 <= not pi0060 and not pi0085;
w8838 <= pi0106 and w8837;
w8839 <= w42 and w6476;
w8840 <= w8838 and w8839;
w8841 <= w8552 and w8840;
w8842 <= w6482 and w8622;
w8843 <= w8841 and w8842;
w8844 <= w8620 and w8843;
w8845 <= w8836 and w8844;
w8846 <= not pi0841 and w267;
w8847 <= w6523 and w8846;
w8848 <= w174 and w269;
w8849 <= w8847 and w8848;
w8850 <= w8845 and w8849;
w8851 <= not pi0054 and not w8850;
w8852 <= w184 and w7758;
w8853 <= pi0054 and not w8852;
w8854 <= w6443 and not w8851;
w8855 <= not w8853 and w8854;
w8856 <= not pi0054 and w8852;
w8857 <= not pi0074 and w8856;
w8858 <= pi0055 and not w8857;
w8859 <= pi0045 and w42;
w8860 <= w50 and w8859;
w8861 <= w8624 and w8860;
w8862 <= w39 and w8861;
w8863 <= w4042 and w7063;
w8864 <= w28 and w135;
w8865 <= w8863 and w8864;
w8866 <= w8862 and w8865;
w8867 <= not pi0055 and not w8866;
w8868 <= w6441 and not w8867;
w8869 <= not w8858 and w8868;
w8870 <= w81 and w100;
w8871 <= w3735 and w8870;
w8872 <= pi0056 and not w8871;
w8873 <= pi0056 and not pi0062;
w8874 <= pi0055 and w7631;
w8875 <= not w8873 and not w8874;
w8876 <= w891 and not w8872;
w8877 <= not w8875 and w8876;
w8878 <= w3867 and w8857;
w8879 <= pi0057 and not w8878;
w8880 <= w4048 and w8870;
w8881 <= not pi0056 and pi0062;
w8882 <= not pi0924 and w8881;
w8883 <= not w8873 and not w8882;
w8884 <= w8880 and not w8883;
w8885 <= not pi0057 and not w8884;
w8886 <= not pi0059 and not w8879;
w8887 <= not w8885 and w8886;
w8888 <= not pi0093 and w8649;
w8889 <= w7728 and w8888;
w8890 <= w4996 and w8889;
w8891 <= pi0059 and not w8878;
w8892 <= pi0924 and w8881;
w8893 <= w8880 and w8892;
w8894 <= not pi0059 and not w8893;
w8895 <= not pi0057 and not w8891;
w8896 <= not w8894 and w8895;
w8897 <= pi0039 and not pi0979;
w8898 <= not w3744 and w8897;
w8899 <= w3745 and w8898;
w8900 <= w3943 and w8899;
w8901 <= not pi0039 and w8827;
w8902 <= w8836 and w8901;
w8903 <= w281 and w8902;
w8904 <= not w8900 and not w8903;
w8905 <= w7763 and not w8904;
w8906 <= pi0841 and w8563;
w8907 <= not pi0024 and w8836;
w8908 <= w281 and w8907;
w8909 <= not w8906 and not w8908;
w8910 <= w7729 and not w8909;
w8911 <= pi0057 and not w7632;
w8912 <= w8871 and w8881;
w8913 <= not pi0057 and not w8912;
w8914 <= not pi0059 and not w8911;
w8915 <= not w8913 and w8914;
w8916 <= w424 and w6498;
w8917 <= w6663 and w8916;
w8918 <= pi0999 and w8917;
w8919 <= not pi0024 and w8565;
w8920 <= not w8918 and not w8919;
w8921 <= w7729 and not w8920;
w8922 <= not pi0063 and pi0107;
w8923 <= w6663 and w8922;
w8924 <= not pi0841 and not w8923;
w8925 <= w49 and w8922;
w8926 <= not pi0064 and not w8925;
w8927 <= w28 and not w8926;
w8928 <= w7732 and w8927;
w8929 <= pi0841 and not w8928;
w8930 <= w8670 and not w8924;
w8931 <= not w8929 and w8930;
w8932 <= pi0039 and w7764;
w8933 <= w7763 and w8932;
w8934 <= not w7780 and w8933;
w8935 <= not w7786 and w8934;
w8936 <= pi0199 and not pi0299;
w8937 <= w133 and w171;
w8938 <= pi0314 and w27;
w8939 <= w8863 and w8938;
w8940 <= pi0081 and not pi0102;
w8941 <= w8939 and w8940;
w8942 <= w52 and w8941;
w8943 <= w172 and w8936;
w8944 <= w8937 and w8943;
w8945 <= w8942 and w8944;
w8946 <= not pi0219 and not w8945;
w8947 <= not pi0199 and not pi0299;
w8948 <= w135 and w8942;
w8949 <= not w8947 and w8948;
w8950 <= pi0219 and not w8949;
w8951 <= w4989 and not w8946;
w8952 <= not w8950 and w8951;
w8953 <= pi0083 and not pi0103;
w8954 <= w8665 and w8953;
w8955 <= w7728 and w8954;
w8956 <= w8939 and w8955;
w8957 <= w47 and w8956;
w8958 <= not w3807 and w3959;
w8959 <= w873 and w3416;
w8960 <= w8958 and w8959;
w8961 <= not w3770 and w3959;
w8962 <= w914 and w1033;
w8963 <= w8961 and w8962;
w8964 <= not w8960 and not w8963;
w8965 <= w8546 and not w8964;
w8966 <= pi0069 and w8621;
w8967 <= w7716 and w8966;
w8968 <= not pi0071 and not w8967;
w8969 <= not pi0081 and not pi0314;
w8970 <= w28 and w8969;
w8971 <= w4001 and w8970;
w8972 <= not w8968 and w8971;
w8973 <= pi0071 and pi0314;
w8974 <= w5001 and w8973;
w8975 <= w7713 and w8974;
w8976 <= w48 and w8975;
w8977 <= not w8972 and not w8976;
w8978 <= w8670 and not w8977;
w8979 <= w68 and w312;
w8980 <= not pi0096 and w8979;
w8981 <= w7757 and w8980;
w8982 <= pi0198 and pi0589;
w8983 <= w1034 and not w3770;
w8984 <= w8982 and w8983;
w8985 <= pi0210 and pi0589;
w8986 <= not pi0221 and w3416;
w8987 <= not pi0216 and w8986;
w8988 <= not w3807 and w8987;
w8989 <= w8985 and w8988;
w8990 <= not w8984 and not w8989;
w8991 <= not pi0593 and w3944;
w8992 <= not w3952 and w8991;
w8993 <= not w8990 and w8992;
w8994 <= not pi0287 and not w8993;
w8995 <= pi0039 and not w8994;
w8996 <= w84 and w8995;
w8997 <= not w8981 and not w8996;
w8998 <= w7763 and not w8997;
w8999 <= w32 and w44;
w9000 <= w3987 and w8999;
w9001 <= w8577 and w9000;
w9002 <= not pi0064 and w6479;
w9003 <= w9001 and w9002;
w9004 <= not pi0081 and not w9003;
w9005 <= not pi0050 and w6498;
w9006 <= w4007 and w9005;
w9007 <= not pi0199 and pi0200;
w9008 <= not pi0299 and w9007;
w9009 <= pi0211 and not pi0219;
w9010 <= pi0299 and w9009;
w9011 <= not w9008 and not w9010;
w9012 <= pi0314 and not w9011;
w9013 <= w7725 and w9012;
w9014 <= not w9004 and w9013;
w9015 <= w9006 and w9014;
w9016 <= w8575 and w9011;
w9017 <= w8939 and w9016;
w9018 <= w9001 and w9017;
w9019 <= not w9015 and not w9018;
w9020 <= w7728 and not w9019;
w9021 <= pi0024 and w272;
w9022 <= pi0072 and w9021;
w9023 <= pi0088 and w7710;
w9024 <= w3951 and w6704;
w9025 <= w9023 and w9024;
w9026 <= w433 and w9025;
w9027 <= not w9022 and not w9026;
w9028 <= w4042 and not w9027;
w9029 <= not pi0039 and not w9028;
w9030 <= w5167 and w8958;
w9031 <= w5171 and w8961;
w9032 <= pi0039 and not w9030;
w9033 <= not w9031 and w9032;
w9034 <= w7763 and not w9033;
w9035 <= not w9029 and w9034;
w9036 <= not pi0314 and pi1050;
w9037 <= w6653 and w7725;
w9038 <= w9036 and w9037;
w9039 <= not pi0039 and not w9038;
w9040 <= w6614 and w8961;
w9041 <= not pi0299 and not w9040;
w9042 <= w6599 and w8958;
w9043 <= pi0299 and not w9042;
w9044 <= not w9041 and not w9043;
w9045 <= pi0039 and not w9044;
w9046 <= w7763 and not w9039;
w9047 <= not w9045 and w9046;
w9048 <= pi0074 and w8856;
w9049 <= w527 and w5089;
w9050 <= not pi0096 and not w9049;
w9051 <= not pi0096 and not pi1093;
w9052 <= w4980 and w9051;
w9053 <= not pi0096 and not w3732;
w9054 <= pi0479 and not w9053;
w9055 <= w936 and w4992;
w9056 <= not w9052 and w9055;
w9057 <= w6468 and not w9054;
w9058 <= w9056 and w9057;
w9059 <= not w9050 and w9058;
w9060 <= w5019 and w9059;
w9061 <= not w9048 and not w9060;
w9062 <= w4989 and not w9061;
w9063 <= w183 and w7758;
w9064 <= pi0075 and not w9063;
w9065 <= pi0096 and not pi1093;
w9066 <= w494 and not w9050;
w9067 <= not w9065 and not w9066;
w9068 <= w173 and not w9067;
w9069 <= w5097 and w9068;
w9070 <= not pi0075 and not w9069;
w9071 <= w6444 and not w9064;
w9072 <= not w9070 and w9071;
w9073 <= w6493 and w7749;
w9074 <= not w7674 and w9073;
w9075 <= not w3837 and not w9074;
w9076 <= w82 and w7938;
w9077 <= pi0252 and w496;
w9078 <= w9076 and not w9077;
w9079 <= not pi0137 and w9078;
w9080 <= not pi0137 and w487;
w9081 <= not pi0094 and not w6494;
w9082 <= not w6460 and not w7937;
w9083 <= w7725 and not w9081;
w9084 <= not w9082 and w9083;
w9085 <= not w496 and not w9084;
w9086 <= not pi0252 and w9084;
w9087 <= pi0252 and w9073;
w9088 <= w496 and not w9087;
w9089 <= not w9086 and w9088;
w9090 <= not w9085 and not w9089;
w9091 <= pi0122 and not w9090;
w9092 <= w4980 and w9085;
w9093 <= not w3840 and not w9076;
w9094 <= not w9089 and not w9093;
w9095 <= not w9092 and w9094;
w9096 <= not pi0122 and not w9095;
w9097 <= not w9091 and not w9096;
w9098 <= not pi1093 and not w9097;
w9099 <= not pi0122 and not w9078;
w9100 <= not w9091 and not w9099;
w9101 <= pi1093 and not w9100;
w9102 <= not w9098 and not w9101;
w9103 <= w487 and not w9102;
w9104 <= not w9080 and not w9103;
w9105 <= not w9079 and not w9104;
w9106 <= not pi0122 and w9076;
w9107 <= pi1093 and not w9084;
w9108 <= not w4981 and not w9107;
w9109 <= not w9106 and not w9108;
w9110 <= not w9098 and not w9109;
w9111 <= not w487 and not w9110;
w9112 <= not pi0137 and not w487;
w9113 <= not w9111 and not w9112;
w9114 <= pi0252 and pi1092;
w9115 <= not pi1093 and w9114;
w9116 <= w488 and w9115;
w9117 <= not pi0137 and not w9116;
w9118 <= w9076 and w9117;
w9119 <= not w9113 and not w9118;
w9120 <= not w9105 and not w9119;
w9121 <= w3837 and not w9120;
w9122 <= not pi0137 and not w3837;
w9123 <= not w9075 and not w9122;
w9124 <= not w9121 and w9123;
w9125 <= not pi0210 and not w9124;
w9126 <= not w9103 and not w9111;
w9127 <= w3837 and not w9126;
w9128 <= not w9075 and not w9127;
w9129 <= pi0210 and not w9128;
w9130 <= not w9125 and not w9129;
w9131 <= w201 and w7862;
w9132 <= not w9130 and not w9131;
w9133 <= not pi0210 and not w9120;
w9134 <= pi0210 and not w9126;
w9135 <= not w9133 and not w9134;
w9136 <= w9131 and not w9135;
w9137 <= pi0299 and not w9136;
w9138 <= not w9132 and w9137;
w9139 <= not pi0198 and not w9124;
w9140 <= pi0198 and not w9128;
w9141 <= not w9139 and not w9140;
w9142 <= w232 and w3760;
w9143 <= not w9141 and not w9142;
w9144 <= pi0198 and not w9126;
w9145 <= not pi0198 and not w9120;
w9146 <= not w9144 and not w9145;
w9147 <= w9142 and not w9146;
w9148 <= not pi0299 and not w9147;
w9149 <= not w9143 and w9148;
w9150 <= not w9138 and not w9149;
w9151 <= pi0232 and not w9150;
w9152 <= pi0299 and not w9130;
w9153 <= not pi0299 and not w9141;
w9154 <= not pi0232 and not w9152;
w9155 <= not w9153 and w9154;
w9156 <= not w9151 and not w9155;
w9157 <= w4988 and not w9156;
w9158 <= not w487 and w9107;
w9159 <= w496 and not w9076;
w9160 <= not w9077 and not w9085;
w9161 <= not w9159 and w9160;
w9162 <= w4981 and not w9161;
w9163 <= not w9091 and not w9162;
w9164 <= w487 and not w9163;
w9165 <= not pi1093 and not w9090;
w9166 <= not w9158 and not w9165;
w9167 <= not w9164 and w9166;
w9168 <= w3837 and w9167;
w9169 <= not w3837 and w9073;
w9170 <= not w7671 and w9169;
w9171 <= not w9168 and not w9170;
w9172 <= pi0210 and not w9171;
w9173 <= w6467 and w9122;
w9174 <= pi0137 and w9165;
w9175 <= not pi0137 and not w9161;
w9176 <= not pi1093 and w9175;
w9177 <= not w9107 and not w9174;
w9178 <= not w9176 and w9177;
w9179 <= w3837 and w9178;
w9180 <= not w9169 and not w9179;
w9181 <= not w487 and not w9173;
w9182 <= not w9180 and w9181;
w9183 <= pi0137 and not w4981;
w9184 <= w496 and not w9183;
w9185 <= w9073 and not w9184;
w9186 <= not w3837 and not w9185;
w9187 <= pi0137 and not w9163;
w9188 <= not w9174 and not w9175;
w9189 <= not w9187 and w9188;
w9190 <= w3837 and not w9189;
w9191 <= w487 and not w9186;
w9192 <= not w9190 and w9191;
w9193 <= not w9182 and not w9192;
w9194 <= not pi0210 and not w9193;
w9195 <= not w9172 and not w9194;
w9196 <= not w9131 and not w9195;
w9197 <= not w487 and w9178;
w9198 <= w487 and w9189;
w9199 <= not w9197 and not w9198;
w9200 <= not pi0210 and w9199;
w9201 <= pi0210 and not w9167;
w9202 <= w9131 and not w9201;
w9203 <= not w9200 and w9202;
w9204 <= pi0299 and not w9203;
w9205 <= not w9196 and w9204;
w9206 <= pi0198 and not w9171;
w9207 <= not pi0198 and not w9193;
w9208 <= not w9206 and not w9207;
w9209 <= not w9142 and not w9208;
w9210 <= not pi0198 and not w9199;
w9211 <= pi0198 and w9167;
w9212 <= not w9210 and not w9211;
w9213 <= w9142 and not w9212;
w9214 <= not pi0299 and not w9213;
w9215 <= not w9209 and w9214;
w9216 <= not w9205 and not w9215;
w9217 <= pi0232 and not w9216;
w9218 <= not pi0299 and not w9208;
w9219 <= pi0299 and not w9195;
w9220 <= not pi0232 and not w9218;
w9221 <= not w9219 and w9220;
w9222 <= not w4988 and not w9221;
w9223 <= not w9217 and w9222;
w9224 <= not w9157 and not w9223;
w9225 <= w7728 and not w9224;
w9226 <= pi0086 and w6460;
w9227 <= w341 and w9226;
w9228 <= pi0314 and not w9227;
w9229 <= w332 and w347;
w9230 <= not pi0086 and not w9229;
w9231 <= w4015 and not w9230;
w9232 <= w265 and w9231;
w9233 <= not pi0314 and not w9232;
w9234 <= w7729 and not w9228;
w9235 <= not w9233 and w9234;
w9236 <= pi0119 and pi0232;
w9237 <= not pi0468 and w9236;
w9238 <= pi0163 and not w7263;
w9239 <= not pi0163 and not w7259;
w9240 <= not w7261 and w9239;
w9241 <= not w9238 and not w9240;
w9242 <= pi0232 and w9241;
w9243 <= not w6552 and w9242;
w9244 <= pi0074 and not w9243;
w9245 <= pi0075 and not w9242;
w9246 <= pi0100 and not w9242;
w9247 <= not w9245 and not w9246;
w9248 <= pi0147 and w5036;
w9249 <= w6552 and w9248;
w9250 <= w9247 and not w9249;
w9251 <= not w891 and not w9244;
w9252 <= w9250 and w9251;
w9253 <= pi0054 and not w9250;
w9254 <= not pi0038 and not pi0040;
w9255 <= pi0038 and not w9248;
w9256 <= not pi0100 and not w9255;
w9257 <= not w9254 and w9256;
w9258 <= not w9246 and not w9257;
w9259 <= not pi0075 and not w9258;
w9260 <= not w9245 and not w9259;
w9261 <= not pi0054 and not w9260;
w9262 <= not w9253 and not w9261;
w9263 <= not pi0074 and not w9262;
w9264 <= not w9244 and not w9263;
w9265 <= not w92 and not w9264;
w9266 <= w891 and not w9265;
w9267 <= not w7285 and w7287;
w9268 <= not pi0184 and w9267;
w9269 <= pi0184 and w3760;
w9270 <= not w9267 and w9269;
w9271 <= not pi0299 and not w9268;
w9272 <= not w9270 and w9271;
w9273 <= pi0299 and not w9241;
w9274 <= pi0232 and not w9272;
w9275 <= not w9273 and w9274;
w9276 <= not w6552 and w9275;
w9277 <= pi0074 and not w9276;
w9278 <= not pi0055 and not w9277;
w9279 <= not pi0187 and not pi0299;
w9280 <= not pi0147 and pi0299;
w9281 <= not w9279 and not w9280;
w9282 <= w5036 and w9281;
w9283 <= w6552 and not w9282;
w9284 <= pi0054 and not w9283;
w9285 <= not w9276 and w9284;
w9286 <= pi0075 and not w9275;
w9287 <= pi0100 and not w9275;
w9288 <= pi0038 and not w9282;
w9289 <= not pi0100 and not w9288;
w9290 <= not pi0179 and not pi0299;
w9291 <= not pi0156 and pi0299;
w9292 <= not w9290 and not w9291;
w9293 <= w5036 and w9292;
w9294 <= w81 and w172;
w9295 <= w9293 and w9294;
w9296 <= w72 and w9295;
w9297 <= w9254 and not w9296;
w9298 <= w9289 and not w9297;
w9299 <= not w9287 and not w9298;
w9300 <= w6768 and not w9299;
w9301 <= not pi0187 and not w6750;
w9302 <= pi0187 and not w6752;
w9303 <= pi0147 and not w9302;
w9304 <= not w9301 and w9303;
w9305 <= not pi0147 and pi0187;
w9306 <= w6757 and w9305;
w9307 <= not w9304 and not w9306;
w9308 <= pi0038 and not w9307;
w9309 <= w72 and w6656;
w9310 <= not w3805 and w6599;
w9311 <= pi0156 and w3751;
w9312 <= not pi0166 and w6856;
w9313 <= not w9311 and not w9312;
w9314 <= w9310 and not w9313;
w9315 <= w9309 and w9314;
w9316 <= not pi0040 and pi0299;
w9317 <= not w9315 and w9316;
w9318 <= not pi0189 and w6856;
w9319 <= pi0179 and w3751;
w9320 <= not w9318 and not w9319;
w9321 <= not w3768 and w6614;
w9322 <= not w9320 and w9321;
w9323 <= w9309 and w9322;
w9324 <= not pi0040 and not pi0299;
w9325 <= not w9323 and w9324;
w9326 <= pi0039 and not w9317;
w9327 <= not w9325 and w9326;
w9328 <= not pi0175 and not pi0299;
w9329 <= pi0184 and w6710;
w9330 <= not pi0184 and not w6706;
w9331 <= not pi0189 and not w9330;
w9332 <= not w9329 and w9331;
w9333 <= not pi0032 and pi0095;
w9334 <= not pi0479 and w9333;
w9335 <= w72 and w9334;
w9336 <= pi0182 and w9335;
w9337 <= pi0184 and pi0189;
w9338 <= not w6713 and w9337;
w9339 <= not w9336 and not w9338;
w9340 <= not w9332 and w9339;
w9341 <= w3760 and not w9340;
w9342 <= not pi0040 and not w9341;
w9343 <= w9328 and not w9342;
w9344 <= w3760 and w9335;
w9345 <= pi0153 and w6656;
w9346 <= w6696 and w9345;
w9347 <= w6706 and w7862;
w9348 <= not pi0040 and not pi0163;
w9349 <= not w9347 and w9348;
w9350 <= not w9346 and w9349;
w9351 <= not w9344 and w9350;
w9352 <= pi0040 and not w3760;
w9353 <= pi0166 and w3760;
w9354 <= not pi0040 and not w9335;
w9355 <= w6729 and w9354;
w9356 <= w9353 and not w9355;
w9357 <= w6725 and w9354;
w9358 <= w7862 and not w9357;
w9359 <= not pi0153 and not w9356;
w9360 <= not w9358 and w9359;
w9361 <= not pi0210 and not w6683;
w9362 <= not w6681 and w9354;
w9363 <= not w9361 and w9362;
w9364 <= w7862 and not w9363;
w9365 <= not w6692 and w9355;
w9366 <= w9353 and not w9365;
w9367 <= pi0153 and not w9366;
w9368 <= not w9364 and w9367;
w9369 <= not w9360 and not w9368;
w9370 <= pi0163 and not w9352;
w9371 <= not w9369 and w9370;
w9372 <= pi0160 and not w9371;
w9373 <= pi0153 and w6681;
w9374 <= w6725 and not w9373;
w9375 <= w7862 and not w9374;
w9376 <= pi0153 and w6692;
w9377 <= w6729 and not w9376;
w9378 <= w9353 and not w9377;
w9379 <= not pi0040 and pi0163;
w9380 <= not w9378 and w9379;
w9381 <= not w9375 and w9380;
w9382 <= not pi0160 and not w9350;
w9383 <= not w9381 and w9382;
w9384 <= not w9372 and not w9383;
w9385 <= pi0299 and not w9351;
w9386 <= not w9384 and w9385;
w9387 <= not w6684 and w9362;
w9388 <= w7858 and not w9387;
w9389 <= pi0189 and w3760;
w9390 <= w6693 and w9354;
w9391 <= w9389 and not w9390;
w9392 <= pi0182 and pi0184;
w9393 <= not w9352 and w9392;
w9394 <= not w9391 and w9393;
w9395 <= not w9388 and w9394;
w9396 <= pi0175 and not pi0299;
w9397 <= pi0189 and not w6696;
w9398 <= not pi0189 and not w6655;
w9399 <= w81 and not w9397;
w9400 <= not w9398 and w9399;
w9401 <= not w9336 and not w9400;
w9402 <= w3760 and not w9401;
w9403 <= not pi0184 and not w9402;
w9404 <= pi0189 and w6694;
w9405 <= not w6685 and w7858;
w9406 <= not pi0182 and pi0184;
w9407 <= not w9404 and w9406;
w9408 <= not w9405 and w9407;
w9409 <= not w9403 and not w9408;
w9410 <= not pi0040 and not w9409;
w9411 <= not w9395 and w9396;
w9412 <= not w9410 and w9411;
w9413 <= not w9343 and not w9412;
w9414 <= not w9386 and w9413;
w9415 <= not pi0039 and not w9414;
w9416 <= pi0232 and not w9327;
w9417 <= not w9415 and w9416;
w9418 <= not pi0040 and not pi0232;
w9419 <= not pi0038 and not w9418;
w9420 <= not w9417 and w9419;
w9421 <= not w9308 and not w9420;
w9422 <= w131 and not w9421;
w9423 <= pi0087 and not w9254;
w9424 <= w9289 and w9423;
w9425 <= not w9287 and not w9424;
w9426 <= not w9422 and w9425;
w9427 <= w132 and not w9426;
w9428 <= not w9286 and not w9300;
w9429 <= not w9427 and w9428;
w9430 <= not pi0054 and not w9429;
w9431 <= not w9285 and not w9430;
w9432 <= not pi0074 and not w9431;
w9433 <= w9278 and not w9432;
w9434 <= pi0055 and not w9244;
w9435 <= pi0163 and pi0232;
w9436 <= not pi0092 and w172;
w9437 <= w9435 and w9436;
w9438 <= w9309 and w9437;
w9439 <= w9254 and not w9438;
w9440 <= not pi0075 and w9256;
w9441 <= not w9439 and w9440;
w9442 <= w9247 and not w9441;
w9443 <= not pi0054 and not w9442;
w9444 <= not w9253 and not w9443;
w9445 <= not pi0074 and not w9444;
w9446 <= w9434 and not w9445;
w9447 <= w92 and not w9446;
w9448 <= not w9433 and w9447;
w9449 <= w9266 and not w9448;
w9450 <= not w9252 and not w9449;
w9451 <= pi0079 and w9450;
w9452 <= w50 and not w6823;
w9453 <= not pi0040 and not w9452;
w9454 <= not w3760 and w6823;
w9455 <= w6811 and not w9454;
w9456 <= w9435 and w9455;
w9457 <= w9453 and not w9456;
w9458 <= not pi0039 and not w9457;
w9459 <= pi0039 and not w7029;
w9460 <= w6771 and not w9459;
w9461 <= not w9458 and w9460;
w9462 <= pi0087 and not w50;
w9463 <= w9254 and w9462;
w9464 <= w9256 and not w9463;
w9465 <= not w9461 and w9464;
w9466 <= not w9246 and not w9465;
w9467 <= w132 and not w9466;
w9468 <= not w6847 and w9258;
w9469 <= w6768 and not w9468;
w9470 <= not w9245 and not w9469;
w9471 <= not w9467 and w9470;
w9472 <= not pi0054 and not w9471;
w9473 <= not w9253 and not w9472;
w9474 <= not pi0074 and not w9473;
w9475 <= w9434 and not w9474;
w9476 <= w9289 and not w9463;
w9477 <= w50 and w9293;
w9478 <= w9453 and not w9477;
w9479 <= not pi0039 and not w9478;
w9480 <= w9460 and not w9479;
w9481 <= w9476 and not w9480;
w9482 <= not w9287 and not w9481;
w9483 <= w6768 and not w9482;
w9484 <= pi0087 and w9476;
w9485 <= not pi0040 and not w6860;
w9486 <= w3805 and not w9485;
w9487 <= w3790 and w7029;
w9488 <= w50 and not w6858;
w9489 <= not pi0040 and not w9488;
w9490 <= not w3790 and w9489;
w9491 <= not w9487 and not w9490;
w9492 <= not w3805 and w9491;
w9493 <= not w9486 and not w9492;
w9494 <= w6854 and w9493;
w9495 <= w3768 and not w9485;
w9496 <= not w3768 and w9491;
w9497 <= not w9495 and not w9496;
w9498 <= w6614 and not w9497;
w9499 <= not w6614 and not w7029;
w9500 <= not pi0299 and not w9499;
w9501 <= not w9498 and w9500;
w9502 <= not pi0232 and not w9494;
w9503 <= not w9501 and w9502;
w9504 <= not pi0189 and not w9485;
w9505 <= w50 and not w6874;
w9506 <= w6703 and not w9505;
w9507 <= w3761 and w9489;
w9508 <= not w9487 and not w9507;
w9509 <= not w9506 and w9508;
w9510 <= pi0189 and not w3768;
w9511 <= w9509 and w9510;
w9512 <= not w9504 and not w9511;
w9513 <= pi0179 and not w9512;
w9514 <= pi0189 and not w9491;
w9515 <= w6703 and w6887;
w9516 <= not w50 and w6703;
w9517 <= not w9515 and not w9516;
w9518 <= w9508 and w9517;
w9519 <= not pi0189 and not w9518;
w9520 <= not pi0179 and not w3768;
w9521 <= not w9514 and w9520;
w9522 <= not w9519 and w9521;
w9523 <= not w9495 and not w9522;
w9524 <= not w9513 and w9523;
w9525 <= w6614 and not w9524;
w9526 <= not w9499 and not w9525;
w9527 <= not pi0299 and not w9526;
w9528 <= not w6599 and w7029;
w9529 <= pi0299 and not w9528;
w9530 <= not pi0166 and not w3805;
w9531 <= not w9493 and not w9530;
w9532 <= w9518 and w9530;
w9533 <= w6599 and not w9532;
w9534 <= not w9531 and w9533;
w9535 <= w9529 and not w9534;
w9536 <= not w9527 and not w9535;
w9537 <= not pi0156 and pi0232;
w9538 <= not w9536 and w9537;
w9539 <= pi0166 and not w3805;
w9540 <= w9509 and w9539;
w9541 <= not w9485 and not w9539;
w9542 <= w6599 and not w9541;
w9543 <= not w9540 and w9542;
w9544 <= w9529 and not w9543;
w9545 <= not w9527 and not w9544;
w9546 <= pi0156 and pi0232;
w9547 <= not w9545 and w9546;
w9548 <= pi0039 and not w9503;
w9549 <= not w9538 and w9548;
w9550 <= not w9547 and w9549;
w9551 <= not w5 and not w7048;
w9552 <= w6911 and not w6912;
w9553 <= not w9551 and not w9552;
w9554 <= not pi0040 and not w7019;
w9555 <= not pi0095 and not w9554;
w9556 <= not w9553 and not w9555;
w9557 <= not pi0299 and w9556;
w9558 <= not pi0040 and not w7144;
w9559 <= not pi0095 and not w9558;
w9560 <= not w9553 and not w9559;
w9561 <= pi0299 and w9560;
w9562 <= not pi0232 and not w9557;
w9563 <= not w9561 and w9562;
w9564 <= not w3760 and w9556;
w9565 <= not pi0040 and not w6990;
w9566 <= not pi0095 and not w9565;
w9567 <= not pi0040 and not w7005;
w9568 <= pi0189 and w9567;
w9569 <= w9566 and not w9568;
w9570 <= not pi0182 and w9553;
w9571 <= pi0182 and w7048;
w9572 <= w3760 and not w9571;
w9573 <= not w9570 and w9572;
w9574 <= not w9569 and w9573;
w9575 <= pi0184 and not w9574;
w9576 <= not pi0040 and w6966;
w9577 <= not pi0032 and not w9576;
w9578 <= not w7050 and not w9577;
w9579 <= not pi0095 and not w9578;
w9580 <= not w7048 and not w9579;
w9581 <= not pi0198 and not w9580;
w9582 <= not w7030 and not w9577;
w9583 <= not pi0095 and not w9582;
w9584 <= not w7048 and not w9583;
w9585 <= pi0198 and not w9584;
w9586 <= w7858 and not w9581;
w9587 <= not w9585 and w9586;
w9588 <= w9389 and w9554;
w9589 <= pi0182 and not pi0184;
w9590 <= not w9587 and w9589;
w9591 <= not w9588 and w9590;
w9592 <= not w9575 and not w9591;
w9593 <= w9328 and not w9592;
w9594 <= pi0095 and not pi0182;
w9595 <= not pi0040 and not w7066;
w9596 <= not pi0095 and pi0189;
w9597 <= w50 and not w9596;
w9598 <= w9595 and not w9597;
w9599 <= not w9594 and not w9598;
w9600 <= w9269 and not w9599;
w9601 <= not w9570 and w9600;
w9602 <= w7123 and w7858;
w9603 <= not pi0198 and not w7053;
w9604 <= not pi0095 and not w7042;
w9605 <= not w7048 and not w9604;
w9606 <= pi0198 and not w9605;
w9607 <= w9389 and not w9603;
w9608 <= not w9606 and w9607;
w9609 <= pi0182 and not w9602;
w9610 <= not w9608 and w9609;
w9611 <= not w7052 and not w9553;
w9612 <= not pi0198 and not w9611;
w9613 <= not w9553 and not w9604;
w9614 <= pi0198 and not w9613;
w9615 <= w9389 and not w9612;
w9616 <= not w9614 and w9615;
w9617 <= not pi0182 and not w9616;
w9618 <= not w9610 and not w9617;
w9619 <= not w7123 and not w9594;
w9620 <= w7858 and not w9553;
w9621 <= not w9619 and w9620;
w9622 <= not w9618 and not w9621;
w9623 <= not pi0184 and not w9622;
w9624 <= w9396 and not w9601;
w9625 <= not w9623 and w9624;
w9626 <= not w9593 and not w9625;
w9627 <= not w9564 and not w9626;
w9628 <= not w3760 and w9560;
w9629 <= not pi0095 and not w9595;
w9630 <= pi0166 and not w9629;
w9631 <= not w9037 and not w9629;
w9632 <= pi0153 and not w9630;
w9633 <= not w9631 and w9632;
w9634 <= pi0166 and w9567;
w9635 <= w9566 and not w9634;
w9636 <= not pi0153 and w9635;
w9637 <= not pi0160 and w3760;
w9638 <= not w9633 and w9637;
w9639 <= not w9553 and w9638;
w9640 <= not w9636 and w9639;
w9641 <= w3760 and not w7048;
w9642 <= w9630 and w9641;
w9643 <= w7029 and w7862;
w9644 <= pi0153 and not w9643;
w9645 <= not w9642 and w9644;
w9646 <= not w9635 and w9641;
w9647 <= not pi0153 and not w9646;
w9648 <= pi0160 and not w9645;
w9649 <= not w9647 and w9648;
w9650 <= pi0163 and not w9640;
w9651 <= not w9649 and w9650;
w9652 <= pi0210 and not w9613;
w9653 <= not pi0210 and not w9611;
w9654 <= w9353 and not w9652;
w9655 <= not w9653 and w9654;
w9656 <= not w7120 and not w9553;
w9657 <= not pi0210 and not w9656;
w9658 <= not w7116 and not w9553;
w9659 <= pi0210 and not w9658;
w9660 <= w7862 and not w9657;
w9661 <= not w9659 and w9660;
w9662 <= pi0153 and not w9655;
w9663 <= not w9661 and w9662;
w9664 <= pi0166 and w9560;
w9665 <= not w9553 and not w9583;
w9666 <= pi0210 and not w9665;
w9667 <= not w9553 and not w9579;
w9668 <= not pi0210 and not w9667;
w9669 <= w7862 and not w9666;
w9670 <= not w9668 and w9669;
w9671 <= not pi0153 and not w9670;
w9672 <= not w9664 and w9671;
w9673 <= not pi0160 and not w9663;
w9674 <= not w9672 and w9673;
w9675 <= pi0210 and not w7117;
w9676 <= not pi0210 and not w7121;
w9677 <= w7862 and not w9675;
w9678 <= not w9676 and w9677;
w9679 <= not pi0210 and not w7053;
w9680 <= pi0210 and not w9605;
w9681 <= w9353 and not w9679;
w9682 <= not w9680 and w9681;
w9683 <= pi0153 and not w9678;
w9684 <= not w9682 and w9683;
w9685 <= w9353 and w9558;
w9686 <= not pi0210 and not w9580;
w9687 <= pi0210 and not w9584;
w9688 <= w7862 and not w9686;
w9689 <= not w9687 and w9688;
w9690 <= not pi0153 and not w9689;
w9691 <= not w9685 and w9690;
w9692 <= pi0160 and not w9684;
w9693 <= not w9691 and w9692;
w9694 <= not pi0163 and not w9693;
w9695 <= not w9674 and w9694;
w9696 <= not w9651 and not w9695;
w9697 <= pi0299 and not w9628;
w9698 <= not w9696 and w9697;
w9699 <= not w7858 and w9556;
w9700 <= pi0198 and not w9665;
w9701 <= not pi0198 and not w9667;
w9702 <= w7858 and not w9700;
w9703 <= not w9701 and w9702;
w9704 <= not pi0182 and not pi0184;
w9705 <= w9328 and w9704;
w9706 <= not w9703 and w9705;
w9707 <= not w9699 and w9706;
w9708 <= not w9627 and not w9707;
w9709 <= not w9698 and w9708;
w9710 <= pi0232 and not w9709;
w9711 <= not pi0039 and not w9563;
w9712 <= not w9710 and w9711;
w9713 <= not pi0038 and not w9550;
w9714 <= not w9712 and w9713;
w9715 <= not w9308 and not w9714;
w9716 <= w131 and not w9715;
w9717 <= not w9287 and not w9484;
w9718 <= not w9716 and w9717;
w9719 <= w132 and not w9718;
w9720 <= not w9286 and not w9483;
w9721 <= not w9719 and w9720;
w9722 <= not pi0054 and not w9721;
w9723 <= not w9285 and not w9722;
w9724 <= not pi0074 and not w9723;
w9725 <= w9278 and not w9724;
w9726 <= w92 and not w9475;
w9727 <= not w9725 and w9726;
w9728 <= not w6815 and w9266;
w9729 <= not w9727 and w9728;
w9730 <= not w9252 and not w9729;
w9731 <= not pi0079 and w9730;
w9732 <= not pi0034 and w7621;
w9733 <= not w9451 and not w9732;
w9734 <= not w9731 and w9733;
w9735 <= not pi0079 and not w6540;
w9736 <= w9450 and w9735;
w9737 <= w9730 and not w9735;
w9738 <= w9732 and not w9736;
w9739 <= not w9737 and w9738;
w9740 <= not w9734 and not w9739;
w9741 <= pi0098 and pi1092;
w9742 <= pi1093 and w9741;
w9743 <= not pi0567 and w489;
w9744 <= not w9742 and not w9743;
w9745 <= not pi0080 and not w9744;
w9746 <= pi0217 and not w9745;
w9747 <= w4988 and w9744;
w9748 <= not w5604 and w9744;
w9749 <= pi0588 and not w9748;
w9750 <= pi0592 and not w5656;
w9751 <= w4985 and not w5682;
w9752 <= not w9750 and w9751;
w9753 <= w9744 and not w9752;
w9754 <= not pi1199 and not w9753;
w9755 <= pi0428 and not w9753;
w9756 <= not w5207 and w9744;
w9757 <= not pi0428 and not w9756;
w9758 <= not w9755 and not w9757;
w9759 <= not pi0427 and not w9758;
w9760 <= not pi0428 and not w9753;
w9761 <= pi0428 and not w9756;
w9762 <= not w9760 and not w9761;
w9763 <= pi0427 and not w9762;
w9764 <= not w9759 and not w9763;
w9765 <= not pi0430 and not w9764;
w9766 <= not pi0427 and not w9762;
w9767 <= pi0427 and not w9758;
w9768 <= not w9766 and not w9767;
w9769 <= pi0430 and not w9768;
w9770 <= not w9765 and not w9769;
w9771 <= not pi0426 and not w9770;
w9772 <= not pi0430 and not w9768;
w9773 <= pi0430 and not w9764;
w9774 <= not w9772 and not w9773;
w9775 <= pi0426 and not w9774;
w9776 <= not w9771 and not w9775;
w9777 <= not pi0445 and not w9776;
w9778 <= not pi0426 and not w9774;
w9779 <= pi0426 and not w9770;
w9780 <= not w9778 and not w9779;
w9781 <= pi0445 and not w9780;
w9782 <= not w9777 and not w9781;
w9783 <= pi0448 and not w9782;
w9784 <= not pi0445 and not w9780;
w9785 <= pi0445 and not w9776;
w9786 <= not w9784 and not w9785;
w9787 <= not pi0448 and not w9786;
w9788 <= w5691 and not w9783;
w9789 <= not w9787 and w9788;
w9790 <= not pi0448 and not w9782;
w9791 <= pi0448 and not w9786;
w9792 <= not w5691 and not w9790;
w9793 <= not w9791 and w9792;
w9794 <= pi1199 and not w9789;
w9795 <= not w9793 and w9794;
w9796 <= w5604 and not w9754;
w9797 <= not w9795 and w9796;
w9798 <= w9749 and not w9797;
w9799 <= pi0591 and not w9744;
w9800 <= pi0590 and not w9799;
w9801 <= not w5208 and w9744;
w9802 <= w5417 and w9801;
w9803 <= not w5320 and w9802;
w9804 <= not w9756 and not w9803;
w9805 <= pi0461 and not w9804;
w9806 <= not w5425 and w9802;
w9807 <= not w9756 and not w9806;
w9808 <= not pi0461 and not w9807;
w9809 <= not w9805 and not w9808;
w9810 <= pi0357 and not w9809;
w9811 <= pi0461 and not w9807;
w9812 <= not pi0461 and not w9804;
w9813 <= not w9811 and not w9812;
w9814 <= not pi0357 and not w9813;
w9815 <= not w9810 and not w9814;
w9816 <= pi0356 and not w9815;
w9817 <= pi0357 and not w9813;
w9818 <= not pi0357 and not w9809;
w9819 <= not w9817 and not w9818;
w9820 <= not pi0356 and not w9819;
w9821 <= not w9816 and not w9820;
w9822 <= pi0354 and w9821;
w9823 <= pi0356 and not w9819;
w9824 <= not pi0356 and not w9815;
w9825 <= not w9823 and not w9824;
w9826 <= not pi0354 and w9825;
w9827 <= not w5450 and not w9822;
w9828 <= not w9826 and w9827;
w9829 <= pi0354 and w9825;
w9830 <= not pi0354 and w9821;
w9831 <= w5450 and not w9829;
w9832 <= not w9830 and w9831;
w9833 <= not pi0591 and not w9828;
w9834 <= not w9832 and w9833;
w9835 <= w9800 and not w9834;
w9836 <= not pi1197 and not w5958;
w9837 <= not w9756 and not w9836;
w9838 <= pi0592 and not w9744;
w9839 <= not pi1196 and not w9744;
w9840 <= not w9838 and not w9839;
w9841 <= pi0397 and not pi0404;
w9842 <= not pi0397 and pi0404;
w9843 <= not w9841 and not w9842;
w9844 <= pi0411 and not w9843;
w9845 <= not pi0411 and w9843;
w9846 <= not w9844 and not w9845;
w9847 <= not w5495 and w9846;
w9848 <= w5495 and not w9846;
w9849 <= not w9847 and not w9848;
w9850 <= w4980 and not w9849;
w9851 <= not w9741 and not w9850;
w9852 <= not pi0412 and not w9851;
w9853 <= w4980 and w9849;
w9854 <= not w9741 and not w9853;
w9855 <= pi0412 and not w9854;
w9856 <= w5507 and not w9852;
w9857 <= not w9855 and w9856;
w9858 <= pi0412 and not w9851;
w9859 <= not pi0412 and not w9854;
w9860 <= not w5507 and not w9858;
w9861 <= not w9859 and w9860;
w9862 <= not pi0122 and not w9857;
w9863 <= not w9861 and w9862;
w9864 <= not w9741 and not w9863;
w9865 <= w5189 and not w9864;
w9866 <= pi1091 and w9742;
w9867 <= not w9865 and not w9866;
w9868 <= pi0567 and not w9867;
w9869 <= not w9743 and not w9868;
w9870 <= w5521 and not w9869;
w9871 <= w9840 and not w9870;
w9872 <= not pi1199 and not w9871;
w9873 <= not pi0122 and w4980;
w9874 <= not w9741 and not w9873;
w9875 <= not w5189 and not w9866;
w9876 <= w4980 and w5489;
w9877 <= not pi0122 and not w9741;
w9878 <= not w9876 and w9877;
w9879 <= not w9875 and not w9878;
w9880 <= not w9874 and w9879;
w9881 <= pi0567 and w9880;
w9882 <= not w9743 and not w9881;
w9883 <= not w9868 and w9882;
w9884 <= w5521 and not w9883;
w9885 <= w6231 and not w9882;
w9886 <= not w9838 and not w9885;
w9887 <= not w9884 and w9886;
w9888 <= pi1199 and not w9887;
w9889 <= not w9872 and not w9888;
w9890 <= w9836 and not w9889;
w9891 <= not w9837 and not w9890;
w9892 <= pi0333 and not w9891;
w9893 <= w5958 and not w9756;
w9894 <= not w5958 and not w9889;
w9895 <= not w9893 and not w9894;
w9896 <= not pi0333 and not w9895;
w9897 <= not w9892 and not w9896;
w9898 <= pi0391 and not w9897;
w9899 <= not pi0333 and not w9891;
w9900 <= pi0333 and not w9895;
w9901 <= not w9899 and not w9900;
w9902 <= not pi0391 and not w9901;
w9903 <= pi0392 and w6364;
w9904 <= not pi0392 and not w6364;
w9905 <= not w9903 and not w9904;
w9906 <= not w9898 and not w9905;
w9907 <= not w9902 and w9906;
w9908 <= pi0391 and not w9901;
w9909 <= not pi0391 and not w9897;
w9910 <= w9905 and not w9908;
w9911 <= not w9909 and w9910;
w9912 <= pi0591 and not w9907;
w9913 <= not w9911 and w9912;
w9914 <= not w5207 and not w5318;
w9915 <= w4985 and not w5289;
w9916 <= not pi1198 and not w9915;
w9917 <= not w5533 and not w9916;
w9918 <= not w9914 and w9917;
w9919 <= w9744 and not w9918;
w9920 <= not pi0591 and not w9919;
w9921 <= not pi0590 and not w9920;
w9922 <= not w9913 and w9921;
w9923 <= not pi0588 and not w9835;
w9924 <= not w9922 and w9923;
w9925 <= not w4988 and not w9798;
w9926 <= not w9924 and w9925;
w9927 <= not pi0080 and not w4989;
w9928 <= not w9747 and w9927;
w9929 <= not w9926 and w9928;
w9930 <= pi0567 and w4992;
w9931 <= not w4983 and not w9742;
w9932 <= not pi0122 and w9931;
w9933 <= w5189 and not w9932;
w9934 <= w188 and not w9866;
w9935 <= not w9933 and w9934;
w9936 <= pi0824 and pi0950;
w9937 <= not pi0110 and w264;
w9938 <= not pi0088 and w58;
w9939 <= w7942 and w9938;
w9940 <= w9937 and w9939;
w9941 <= w5003 and w9940;
w9942 <= w5009 and w9941;
w9943 <= pi0051 and w9942;
w9944 <= pi0090 and pi0093;
w9945 <= not pi0841 and not w267;
w9946 <= not w9944 and w9945;
w9947 <= w525 and w9946;
w9948 <= w9941 and w9947;
w9949 <= not w9943 and not w9948;
w9950 <= w5013 and w9936;
w9951 <= not w9949 and w9950;
w9952 <= not pi0098 and not w9951;
w9953 <= pi1092 and not w9952;
w9954 <= not pi0087 and w9934;
w9955 <= not w9953 and w9954;
w9956 <= w83 and w9936;
w9957 <= w9942 and w9956;
w9958 <= not pi0098 and not w9957;
w9959 <= pi1092 and not w9958;
w9960 <= pi0087 and w9934;
w9961 <= not w9959 and w9960;
w9962 <= not w9955 and not w9961;
w9963 <= pi0122 and not w9962;
w9964 <= not w9935 and not w9963;
w9965 <= not pi0075 and not w9964;
w9966 <= not w5028 and w9931;
w9967 <= w9930 and not w9966;
w9968 <= not w9965 and w9967;
w9969 <= not w4992 and not w9931;
w9970 <= not w9743 and not w9969;
w9971 <= not w9968 and w9970;
w9972 <= not pi0592 and not w9971;
w9973 <= not w9838 and not w9972;
w9974 <= not w5656 and w9973;
w9975 <= w5656 and not w9839;
w9976 <= not pi0443 and not w9744;
w9977 <= pi0443 and not w9973;
w9978 <= not w9976 and not w9977;
w9979 <= w5812 and w9978;
w9980 <= pi0443 and not w9744;
w9981 <= not pi0443 and not w9973;
w9982 <= not w9980 and not w9981;
w9983 <= not w5812 and w9982;
w9984 <= not w9979 and not w9983;
w9985 <= pi0435 and not w9984;
w9986 <= not pi0444 and w9982;
w9987 <= pi0444 and w9978;
w9988 <= not pi0436 and not w9986;
w9989 <= not w9987 and w9988;
w9990 <= not pi0444 and w9978;
w9991 <= pi0444 and w9982;
w9992 <= pi0436 and not w9990;
w9993 <= not w9991 and w9992;
w9994 <= not w9989 and not w9993;
w9995 <= not pi0435 and w9994;
w9996 <= not w9985 and not w9995;
w9997 <= not pi0429 and w9996;
w9998 <= not pi0435 and not w9984;
w9999 <= pi0435 and w9994;
w10000 <= not w9998 and not w9999;
w10001 <= pi0429 and w10000;
w10002 <= w5668 and not w9997;
w10003 <= not w10001 and w10002;
w10004 <= not pi0429 and w10000;
w10005 <= pi0429 and w9996;
w10006 <= not w5668 and not w10004;
w10007 <= not w10005 and w10006;
w10008 <= pi1196 and not w10003;
w10009 <= not w10007 and w10008;
w10010 <= w9975 and not w10009;
w10011 <= not w9974 and not w10010;
w10012 <= not pi1199 and w10011;
w10013 <= pi0428 and not w10011;
w10014 <= not pi0428 and w9973;
w10015 <= not w10013 and not w10014;
w10016 <= not pi0427 and not w10015;
w10017 <= not pi0428 and not w10011;
w10018 <= pi0428 and w9973;
w10019 <= not w10017 and not w10018;
w10020 <= pi0427 and not w10019;
w10021 <= not w10016 and not w10020;
w10022 <= pi0430 and not w10021;
w10023 <= not pi0427 and not w10019;
w10024 <= pi0427 and not w10015;
w10025 <= not w10023 and not w10024;
w10026 <= not pi0430 and not w10025;
w10027 <= not w10022 and not w10026;
w10028 <= pi0426 and not w10027;
w10029 <= pi0430 and not w10025;
w10030 <= not pi0430 and not w10021;
w10031 <= not w10029 and not w10030;
w10032 <= not pi0426 and not w10031;
w10033 <= not w10028 and not w10032;
w10034 <= pi0445 and not w10033;
w10035 <= pi0426 and not w10031;
w10036 <= not pi0426 and not w10027;
w10037 <= not w10035 and not w10036;
w10038 <= not pi0445 and not w10037;
w10039 <= not w10034 and not w10038;
w10040 <= pi0448 and w10039;
w10041 <= pi0445 and not w10037;
w10042 <= not pi0445 and not w10033;
w10043 <= not w10041 and not w10042;
w10044 <= not pi0448 and w10043;
w10045 <= not w5691 and not w10040;
w10046 <= not w10044 and w10045;
w10047 <= not pi0448 and w10039;
w10048 <= pi0448 and w10043;
w10049 <= w5691 and not w10047;
w10050 <= not w10048 and w10049;
w10051 <= pi1199 and not w10046;
w10052 <= not w10050 and w10051;
w10053 <= w5604 and not w10012;
w10054 <= not w10052 and w10053;
w10055 <= w9749 and not w10054;
w10056 <= w5413 and w9744;
w10057 <= not w5413 and w9973;
w10058 <= not w10056 and not w10057;
w10059 <= pi1198 and not w10058;
w10060 <= not pi1198 and not w9839;
w10061 <= w5354 and w9744;
w10062 <= not w5354 and w9973;
w10063 <= not w10061 and not w10062;
w10064 <= not pi0355 and not w10063;
w10065 <= pi0455 and not w9744;
w10066 <= not pi0455 and not w9973;
w10067 <= not w10065 and not w10066;
w10068 <= not pi0452 and not w10067;
w10069 <= not pi0455 and not w9744;
w10070 <= pi0455 and not w9973;
w10071 <= not w10069 and not w10070;
w10072 <= pi0452 and not w10071;
w10073 <= not w10068 and not w10072;
w10074 <= pi0355 and w10073;
w10075 <= not w10064 and not w10074;
w10076 <= not pi0458 and w10075;
w10077 <= pi0355 and not w10063;
w10078 <= not pi0355 and w10073;
w10079 <= not w10077 and not w10078;
w10080 <= pi0458 and w10079;
w10081 <= w5375 and not w10076;
w10082 <= not w10080 and w10081;
w10083 <= not pi0458 and w10079;
w10084 <= pi0458 and w10075;
w10085 <= not w5375 and not w10083;
w10086 <= not w10084 and w10085;
w10087 <= pi1196 and not w10082;
w10088 <= not w10086 and w10087;
w10089 <= w10060 and not w10088;
w10090 <= not w10059 and not w10089;
w10091 <= not w5345 and not w10090;
w10092 <= w5345 and w9973;
w10093 <= not w10091 and not w10092;
w10094 <= not w5320 and w10093;
w10095 <= pi1199 and not w9973;
w10096 <= pi0351 and w10095;
w10097 <= not w10094 and not w10096;
w10098 <= not pi0461 and not w10097;
w10099 <= not w5425 and w10093;
w10100 <= not pi0351 and w10095;
w10101 <= not w10099 and not w10100;
w10102 <= pi0461 and not w10101;
w10103 <= not w10098 and not w10102;
w10104 <= not pi0357 and not w10103;
w10105 <= not pi0461 and not w10101;
w10106 <= pi0461 and not w10097;
w10107 <= not w10105 and not w10106;
w10108 <= pi0357 and not w10107;
w10109 <= not w10104 and not w10108;
w10110 <= not pi0356 and not w10109;
w10111 <= not pi0357 and not w10107;
w10112 <= pi0357 and not w10103;
w10113 <= not w10111 and not w10112;
w10114 <= pi0356 and not w10113;
w10115 <= not w10110 and not w10114;
w10116 <= not pi0354 and not w10115;
w10117 <= not pi0356 and not w10113;
w10118 <= pi0356 and not w10109;
w10119 <= not w10117 and not w10118;
w10120 <= pi0354 and not w10119;
w10121 <= not w5450 and not w10116;
w10122 <= not w10120 and w10121;
w10123 <= not pi0354 and not w10119;
w10124 <= pi0354 and not w10115;
w10125 <= w5450 and not w10123;
w10126 <= not w10124 and w10125;
w10127 <= not pi0591 and not w10122;
w10128 <= not w10126 and w10127;
w10129 <= w9800 and not w10128;
w10130 <= not w9836 and w9973;
w10131 <= w4992 and not w9743;
w10132 <= not w9869 and not w10131;
w10133 <= pi0075 and w9867;
w10134 <= not pi0411 and w9741;
w10135 <= w5513 and not w10134;
w10136 <= pi0411 and w9959;
w10137 <= w10135 and not w10136;
w10138 <= not pi0411 and w9959;
w10139 <= not w5513 and not w9741;
w10140 <= not w5515 and not w10139;
w10141 <= not w10138 and not w10140;
w10142 <= not w10137 and not w10141;
w10143 <= pi0122 and w10142;
w10144 <= not w9863 and not w10143;
w10145 <= w5189 and not w10144;
w10146 <= w9960 and not w10145;
w10147 <= pi0411 and w9953;
w10148 <= w10135 and not w10147;
w10149 <= not pi0411 and w9953;
w10150 <= not w10140 and not w10149;
w10151 <= not w10148 and not w10150;
w10152 <= pi0122 and w10151;
w10153 <= not w9863 and not w10152;
w10154 <= w5189 and not w10153;
w10155 <= w9954 and not w10154;
w10156 <= not w188 and w9867;
w10157 <= not w10146 and not w10156;
w10158 <= not w10155 and w10157;
w10159 <= not pi0075 and not w10158;
w10160 <= w9930 and not w10133;
w10161 <= not w10159 and w10160;
w10162 <= not w10132 and not w10161;
w10163 <= w5521 and not w10162;
w10164 <= not w9839 and not w10163;
w10165 <= not pi1199 and not w10164;
w10166 <= not w9883 and not w10131;
w10167 <= not w5028 and not w9880;
w10168 <= not w9865 and w10167;
w10169 <= w188 and not w9879;
w10170 <= not w9865 and w10169;
w10171 <= not pi0122 and w9876;
w10172 <= w5489 and w9953;
w10173 <= not w5489 and w9741;
w10174 <= not w10172 and not w10173;
w10175 <= w9954 and w10174;
w10176 <= not w5513 and not w10149;
w10177 <= not w10148 and not w10176;
w10178 <= w10175 and not w10177;
w10179 <= w5489 and w9959;
w10180 <= w9960 and not w10179;
w10181 <= not w10142 and w10180;
w10182 <= not w10178 and not w10181;
w10183 <= not w9863 and not w10171;
w10184 <= not w10182 and w10183;
w10185 <= not w10170 and not w10184;
w10186 <= not pi0075 and not w10185;
w10187 <= w9930 and not w10168;
w10188 <= not w10186 and w10187;
w10189 <= not w10166 and not w10188;
w10190 <= w5521 and not w10189;
w10191 <= not w9882 and not w10131;
w10192 <= not w10173 and not w10179;
w10193 <= w9960 and w10192;
w10194 <= not w10175 and not w10193;
w10195 <= pi0122 and not w10194;
w10196 <= not w10169 and not w10195;
w10197 <= not pi0075 and not w10196;
w10198 <= w9930 and not w10167;
w10199 <= not w10197 and w10198;
w10200 <= not w10191 and not w10199;
w10201 <= w6231 and not w10200;
w10202 <= not w10190 and not w10201;
w10203 <= pi1199 and not w10202;
w10204 <= not w9838 and not w10203;
w10205 <= not w10165 and w10204;
w10206 <= w9836 and w10205;
w10207 <= not w10130 and not w10206;
w10208 <= pi0333 and not w10207;
w10209 <= w5958 and not w9973;
w10210 <= not w5958 and not w10205;
w10211 <= not w10209 and not w10210;
w10212 <= not pi0333 and w10211;
w10213 <= not w10208 and not w10212;
w10214 <= pi0391 and not w10213;
w10215 <= pi0333 and not w10211;
w10216 <= not pi0333 and w10207;
w10217 <= not w10215 and not w10216;
w10218 <= not pi0391 and w10217;
w10219 <= not w10214 and not w10218;
w10220 <= pi0392 and not w10219;
w10221 <= not pi0391 and w10213;
w10222 <= pi0391 and not w10217;
w10223 <= not w10221 and not w10222;
w10224 <= not pi0392 and w10223;
w10225 <= not w10220 and not w10224;
w10226 <= pi0393 and not w10225;
w10227 <= not pi0392 and not w10219;
w10228 <= pi0392 and w10223;
w10229 <= not w10227 and not w10228;
w10230 <= not pi0393 and not w10229;
w10231 <= not w10226 and not w10230;
w10232 <= not w5591 and not w10231;
w10233 <= pi0393 and not w10229;
w10234 <= not pi0393 and not w10225;
w10235 <= not w10233 and not w10234;
w10236 <= w5591 and not w10235;
w10237 <= pi0591 and not w10232;
w10238 <= not w10236 and w10237;
w10239 <= not pi0592 and not w9744;
w10240 <= pi0592 and not w9971;
w10241 <= not w10239 and not w10240;
w10242 <= not w5285 and w10241;
w10243 <= w5285 and w9744;
w10244 <= not w10242 and not w10243;
w10245 <= pi1199 and w10244;
w10246 <= w5233 and w10241;
w10247 <= not pi1197 and not w9744;
w10248 <= not w5233 and not w10247;
w10249 <= pi0367 and not w9744;
w10250 <= not pi0367 and not w10241;
w10251 <= not w10249 and not w10250;
w10252 <= w5236 and not w10251;
w10253 <= not pi0367 and not w9744;
w10254 <= pi0367 and not w10241;
w10255 <= not w10253 and not w10254;
w10256 <= not w5236 and not w10255;
w10257 <= not w10252 and not w10256;
w10258 <= w5239 and not w10257;
w10259 <= not w5236 and w10251;
w10260 <= w5236 and w10255;
w10261 <= not w10259 and not w10260;
w10262 <= not w5239 and w10261;
w10263 <= not w5248 and not w10258;
w10264 <= not w10262 and w10263;
w10265 <= not w5239 and not w10257;
w10266 <= w5239 and w10261;
w10267 <= w5248 and not w10265;
w10268 <= not w10266 and w10267;
w10269 <= pi1197 and not w10264;
w10270 <= not w10268 and w10269;
w10271 <= w10248 and not w10270;
w10272 <= not pi1199 and not w10246;
w10273 <= not w10271 and w10272;
w10274 <= not w10245 and not w10273;
w10275 <= not pi0374 and not w10274;
w10276 <= w6062 and w10244;
w10277 <= not pi1198 and w10273;
w10278 <= pi1198 and not w10241;
w10279 <= not w10276 and not w10278;
w10280 <= not w10277 and w10279;
w10281 <= pi0374 and not w10280;
w10282 <= not w10275 and not w10281;
w10283 <= pi0369 and not w10282;
w10284 <= not pi0374 and not w10280;
w10285 <= pi0374 and not w10274;
w10286 <= not w10284 and not w10285;
w10287 <= not pi0369 and not w10286;
w10288 <= pi0371 and w6416;
w10289 <= not pi0371 and not w6416;
w10290 <= not w10288 and not w10289;
w10291 <= pi0370 and not w10290;
w10292 <= not pi0370 and w10290;
w10293 <= not w10291 and not w10292;
w10294 <= not w10283 and w10293;
w10295 <= not w10287 and w10294;
w10296 <= not pi0369 and not w10282;
w10297 <= pi0369 and not w10286;
w10298 <= not w10293 and not w10296;
w10299 <= not w10297 and w10298;
w10300 <= not pi0591 and not w10295;
w10301 <= not w10299 and w10300;
w10302 <= not pi0590 and not w10238;
w10303 <= not w10301 and w10302;
w10304 <= not pi0588 and not w10303;
w10305 <= not w10129 and w10304;
w10306 <= not w4988 and not w10305;
w10307 <= not w10055 and w10306;
w10308 <= not w4992 and w9744;
w10309 <= pi0075 and w9742;
w10310 <= not w9866 and not w9959;
w10311 <= w5725 and not w9875;
w10312 <= not w10310 and w10311;
w10313 <= not w9866 and not w9953;
w10314 <= w173 and not w9875;
w10315 <= not w10313 and w10314;
w10316 <= not w188 and w9742;
w10317 <= not w10312 and not w10316;
w10318 <= not w10315 and w10317;
w10319 <= not pi0075 and not w10318;
w10320 <= not w10309 and not w10319;
w10321 <= pi0567 and not w10320;
w10322 <= w10131 and not w10321;
w10323 <= not w10308 and not w10322;
w10324 <= not pi0592 and w10323;
w10325 <= not w9838 and not w10324;
w10326 <= not w5656 and w10325;
w10327 <= pi0443 and not w10325;
w10328 <= not w9976 and not w10327;
w10329 <= w5812 and w10328;
w10330 <= not pi0443 and not w10325;
w10331 <= not w9980 and not w10330;
w10332 <= not w5812 and w10331;
w10333 <= not w10329 and not w10332;
w10334 <= pi0435 and not w10333;
w10335 <= not pi0444 and w10331;
w10336 <= pi0444 and w10328;
w10337 <= not pi0436 and not w10335;
w10338 <= not w10336 and w10337;
w10339 <= not pi0444 and w10328;
w10340 <= pi0444 and w10331;
w10341 <= pi0436 and not w10339;
w10342 <= not w10340 and w10341;
w10343 <= not w10338 and not w10342;
w10344 <= not pi0435 and w10343;
w10345 <= not w10334 and not w10344;
w10346 <= not pi0429 and w10345;
w10347 <= not pi0435 and not w10333;
w10348 <= pi0435 and w10343;
w10349 <= not w10347 and not w10348;
w10350 <= pi0429 and w10349;
w10351 <= w5668 and not w10346;
w10352 <= not w10350 and w10351;
w10353 <= not pi0429 and w10349;
w10354 <= pi0429 and w10345;
w10355 <= not w5668 and not w10353;
w10356 <= not w10354 and w10355;
w10357 <= pi1196 and not w10352;
w10358 <= not w10356 and w10357;
w10359 <= w9975 and not w10358;
w10360 <= not w10326 and not w10359;
w10361 <= not pi1199 and w10360;
w10362 <= not pi0428 and not w10360;
w10363 <= pi0428 and w10325;
w10364 <= not w10362 and not w10363;
w10365 <= not pi0427 and not w10364;
w10366 <= pi0428 and not w10360;
w10367 <= not pi0428 and w10325;
w10368 <= not w10366 and not w10367;
w10369 <= pi0427 and not w10368;
w10370 <= not w10365 and not w10369;
w10371 <= pi0430 and not w10370;
w10372 <= not pi0427 and not w10368;
w10373 <= pi0427 and not w10364;
w10374 <= not w10372 and not w10373;
w10375 <= not pi0430 and not w10374;
w10376 <= not w10371 and not w10375;
w10377 <= pi0426 and not w10376;
w10378 <= pi0430 and not w10374;
w10379 <= not pi0430 and not w10370;
w10380 <= not w10378 and not w10379;
w10381 <= not pi0426 and not w10380;
w10382 <= not w10377 and not w10381;
w10383 <= pi0445 and not w10382;
w10384 <= pi0426 and not w10380;
w10385 <= not pi0426 and not w10376;
w10386 <= not w10384 and not w10385;
w10387 <= not pi0445 and not w10386;
w10388 <= not w10383 and not w10387;
w10389 <= pi0448 and w10388;
w10390 <= pi0445 and not w10386;
w10391 <= not pi0445 and not w10382;
w10392 <= not w10390 and not w10391;
w10393 <= not pi0448 and w10392;
w10394 <= w5691 and not w10389;
w10395 <= not w10393 and w10394;
w10396 <= pi0448 and w10392;
w10397 <= not pi0448 and w10388;
w10398 <= not w5691 and not w10396;
w10399 <= not w10397 and w10398;
w10400 <= pi1199 and not w10395;
w10401 <= not w10399 and w10400;
w10402 <= w5604 and not w10361;
w10403 <= not w10401 and w10402;
w10404 <= w9749 and not w10403;
w10405 <= not w9836 and not w10325;
w10406 <= w5973 and w10131;
w10407 <= not w9744 and not w10406;
w10408 <= w5521 and not w10308;
w10409 <= not w9866 and not w10142;
w10410 <= w10311 and not w10409;
w10411 <= not w9866 and not w10151;
w10412 <= w10314 and not w10411;
w10413 <= not w10316 and not w10410;
w10414 <= not w10412 and w10413;
w10415 <= w5489 and w10312;
w10416 <= not w10174 and w10315;
w10417 <= not w10415 and not w10416;
w10418 <= w10414 and w10417;
w10419 <= w10408 and not w10418;
w10420 <= not w10192 and w10312;
w10421 <= not w10316 and not w10420;
w10422 <= not w10416 and w10421;
w10423 <= w6231 and not w10308;
w10424 <= not w10422 and w10423;
w10425 <= not w10419 and not w10424;
w10426 <= not pi0075 and pi0567;
w10427 <= not w10425 and w10426;
w10428 <= pi1199 and not w10407;
w10429 <= not w10427 and w10428;
w10430 <= not pi0075 and not w10414;
w10431 <= not w10309 and not w10430;
w10432 <= pi0567 and not w10431;
w10433 <= w10131 and not w10432;
w10434 <= w10408 and not w10433;
w10435 <= not pi1199 and w9840;
w10436 <= not w10434 and w10435;
w10437 <= not w5958 and not w10429;
w10438 <= not w10436 and w10437;
w10439 <= not pi1197 and w10438;
w10440 <= not w10405 and not w10439;
w10441 <= not pi0333 and not w10440;
w10442 <= w5958 and not w10325;
w10443 <= not w10438 and not w10442;
w10444 <= pi0333 and not w10443;
w10445 <= not w10441 and not w10444;
w10446 <= not pi0391 and not w10445;
w10447 <= pi0333 and not w10440;
w10448 <= not pi0333 and not w10443;
w10449 <= not w10447 and not w10448;
w10450 <= pi0391 and not w10449;
w10451 <= not w10446 and not w10450;
w10452 <= not pi0392 and not w10451;
w10453 <= not pi0391 and not w10449;
w10454 <= pi0391 and not w10445;
w10455 <= not w10453 and not w10454;
w10456 <= pi0392 and not w10455;
w10457 <= not w10452 and not w10456;
w10458 <= not pi0393 and not w10457;
w10459 <= not pi0392 and not w10455;
w10460 <= pi0392 and not w10451;
w10461 <= not w10459 and not w10460;
w10462 <= pi0393 and not w10461;
w10463 <= not w5591 and not w10458;
w10464 <= not w10462 and w10463;
w10465 <= not pi0393 and not w10461;
w10466 <= pi0393 and not w10457;
w10467 <= w5591 and not w10465;
w10468 <= not w10466 and w10467;
w10469 <= pi0591 and not w10464;
w10470 <= not w10468 and w10469;
w10471 <= pi0592 and w10323;
w10472 <= not w10239 and not w10471;
w10473 <= not w5285 and w10472;
w10474 <= pi1199 and not w10243;
w10475 <= not w10473 and w10474;
w10476 <= w5236 and w5251;
w10477 <= not w5236 and not w5251;
w10478 <= not w10476 and not w10477;
w10479 <= pi0367 and not w10478;
w10480 <= not pi0367 and w10478;
w10481 <= not w10479 and not w10480;
w10482 <= w9744 and not w10481;
w10483 <= w10472 and w10481;
w10484 <= pi1197 and not w10482;
w10485 <= not w10483 and w10484;
w10486 <= w10248 and not w10485;
w10487 <= w5233 and w10472;
w10488 <= not pi1199 and not w10487;
w10489 <= not w10486 and w10488;
w10490 <= not w10475 and not w10489;
w10491 <= not pi0374 and not w10490;
w10492 <= not pi1198 and not w10490;
w10493 <= pi1198 and not w10472;
w10494 <= not w10492 and not w10493;
w10495 <= pi0374 and not w10494;
w10496 <= not w10491 and not w10495;
w10497 <= not pi0369 and not w10496;
w10498 <= not pi0374 and not w10494;
w10499 <= pi0374 and not w10490;
w10500 <= not w10498 and not w10499;
w10501 <= pi0369 and not w10500;
w10502 <= not w10293 and not w10497;
w10503 <= not w10501 and w10502;
w10504 <= pi0369 and not w10496;
w10505 <= not pi0369 and not w10500;
w10506 <= w10293 and not w10504;
w10507 <= not w10505 and w10506;
w10508 <= not pi0591 and not w10503;
w10509 <= not w10507 and w10508;
w10510 <= not pi0590 and not w10509;
w10511 <= not w10470 and w10510;
w10512 <= not w5413 and w10325;
w10513 <= not w10056 and not w10512;
w10514 <= pi1198 and not w10513;
w10515 <= not w5354 and w10325;
w10516 <= not w10061 and not w10515;
w10517 <= pi0355 and not w10516;
w10518 <= not pi0455 and not w10325;
w10519 <= not w10065 and not w10518;
w10520 <= not pi0452 and not w10519;
w10521 <= pi0455 and not w10325;
w10522 <= not w10069 and not w10521;
w10523 <= pi0452 and not w10522;
w10524 <= not w10520 and not w10523;
w10525 <= not pi0355 and w10524;
w10526 <= not w10517 and not w10525;
w10527 <= not pi0458 and w10526;
w10528 <= not pi0355 and not w10516;
w10529 <= pi0355 and w10524;
w10530 <= not w10528 and not w10529;
w10531 <= pi0458 and w10530;
w10532 <= not w5375 and not w10527;
w10533 <= not w10531 and w10532;
w10534 <= not pi0458 and w10530;
w10535 <= pi0458 and w10526;
w10536 <= w5375 and not w10534;
w10537 <= not w10535 and w10536;
w10538 <= pi1196 and not w10533;
w10539 <= not w10537 and w10538;
w10540 <= w10060 and not w10539;
w10541 <= not w10514 and not w10540;
w10542 <= not w5345 and not w10541;
w10543 <= w5345 and w10325;
w10544 <= not w10542 and not w10543;
w10545 <= not w5320 and w10544;
w10546 <= pi1199 and not w10325;
w10547 <= pi0351 and w10546;
w10548 <= not w10545 and not w10547;
w10549 <= not pi0461 and not w10548;
w10550 <= not w5425 and w10544;
w10551 <= not pi0351 and w10546;
w10552 <= not w10550 and not w10551;
w10553 <= pi0461 and not w10552;
w10554 <= not w10549 and not w10553;
w10555 <= not pi0357 and not w10554;
w10556 <= not pi0461 and not w10552;
w10557 <= pi0461 and not w10548;
w10558 <= not w10556 and not w10557;
w10559 <= pi0357 and not w10558;
w10560 <= not w10555 and not w10559;
w10561 <= not pi0356 and not w10560;
w10562 <= not pi0357 and not w10558;
w10563 <= pi0357 and not w10554;
w10564 <= not w10562 and not w10563;
w10565 <= pi0356 and not w10564;
w10566 <= not w10561 and not w10565;
w10567 <= not pi0354 and not w10566;
w10568 <= not pi0356 and not w10564;
w10569 <= pi0356 and not w10560;
w10570 <= not w10568 and not w10569;
w10571 <= pi0354 and not w10570;
w10572 <= not w5450 and not w10567;
w10573 <= not w10571 and w10572;
w10574 <= not pi0354 and not w10570;
w10575 <= pi0354 and not w10566;
w10576 <= w5450 and not w10574;
w10577 <= not w10575 and w10576;
w10578 <= not pi0591 and not w10573;
w10579 <= not w10577 and w10578;
w10580 <= w9800 and not w10579;
w10581 <= not pi0588 and not w10511;
w10582 <= not w10580 and w10581;
w10583 <= w4988 and not w10582;
w10584 <= not w10404 and w10583;
w10585 <= not pi0080 and w4989;
w10586 <= not w10307 and w10585;
w10587 <= not w10584 and w10586;
w10588 <= not pi0217 and not w9929;
w10589 <= not w10587 and w10588;
w10590 <= w5206 and not w9746;
w10591 <= not w10589 and w10590;
w10592 <= w4989 and w8865;
w10593 <= pi0081 and not pi0314;
w10594 <= w52 and w10593;
w10595 <= pi0068 and not pi0081;
w10596 <= w43 and w10595;
w10597 <= w8577 and w10596;
w10598 <= w9002 and w10597;
w10599 <= w363 and w10598;
w10600 <= not w10594 and not w10599;
w10601 <= w10592 and not w10600;
w10602 <= pi0069 and pi0314;
w10603 <= w355 and w10602;
w10604 <= pi0066 and not pi0073;
w10605 <= w31 and w10604;
w10606 <= w45 and w10605;
w10607 <= not w10603 and not w10606;
w10608 <= w8666 and w8670;
w10609 <= not w10607 and w10608;
w10610 <= w43 and w362;
w10611 <= pi0084 and w6640;
w10612 <= w10610 and w10611;
w10613 <= w30 and w10612;
w10614 <= w62 and w8665;
w10615 <= w265 and w10614;
w10616 <= w10613 and w10615;
w10617 <= pi0314 and not w10616;
w10618 <= not pi0083 and not w10612;
w10619 <= w10615 and not w10618;
w10620 <= w358 and w10619;
w10621 <= not pi0314 and not w10620;
w10622 <= w7729 and not w10617;
w10623 <= not w10621 and w10622;
w10624 <= pi0211 and pi0299;
w10625 <= pi0219 and pi0299;
w10626 <= not w10624 and not w10625;
w10627 <= not w8373 and w10626;
w10628 <= w4989 and w10627;
w10629 <= w8948 and w10628;
w10630 <= w3986 and w8667;
w10631 <= not pi0314 and w8668;
w10632 <= w9000 and w10631;
w10633 <= not w10630 and not w10632;
w10634 <= w8670 and not w10633;
w10635 <= w5166 and w8959;
w10636 <= w5169 and w8962;
w10637 <= not w10635 and not w10636;
w10638 <= w8546 and not w10637;
w10639 <= w408 and w10614;
w10640 <= pi0314 and w7729;
w10641 <= w265 and w10640;
w10642 <= w10639 and w10641;
w10643 <= w271 and w4980;
w10644 <= not pi1093 and w82;
w10645 <= w135 and w10644;
w10646 <= w10643 and w10645;
w10647 <= w9023 and w10646;
w10648 <= w433 and w10647;
w10649 <= not w4988 and not w10648;
w10650 <= w4980 and w8593;
w10651 <= not pi1093 and not w10650;
w10652 <= w5002 and w9939;
w10653 <= w8590 and w10652;
w10654 <= w8606 and w9937;
w10655 <= w10653 and w10654;
w10656 <= pi1093 and not w10655;
w10657 <= w135 and not w7637;
w10658 <= not w10656 and w10657;
w10659 <= not w10651 and w10658;
w10660 <= w4988 and not w10659;
w10661 <= w4989 and not w10649;
w10662 <= not w10660 and w10661;
w10663 <= w28 and w6484;
w10664 <= w6498 and w10663;
w10665 <= w7744 and w10664;
w10666 <= pi0841 and w5008;
w10667 <= w10665 and w10666;
w10668 <= not pi0070 and not w10667;
w10669 <= pi0070 and not w6522;
w10670 <= w83 and w7728;
w10671 <= not w10668 and w10670;
w10672 <= not w10669 and w10671;
w10673 <= not pi1050 and w6653;
w10674 <= not pi0090 and not w10673;
w10675 <= w8889 and not w10674;
w10676 <= not w459 and w10675;
w10677 <= not w4996 and w10676;
w10678 <= not pi0058 and w319;
w10679 <= not w7721 and not w10678;
w10680 <= w491 and w7725;
w10681 <= not w10679 and w10680;
w10682 <= pi0024 and w501;
w10683 <= not w491 and w10682;
w10684 <= w8649 and w10683;
w10685 <= w319 and w10684;
w10686 <= not pi0039 and not w10685;
w10687 <= not w10681 and w10686;
w10688 <= w7760 and not w10687;
w10689 <= w5175 and w10688;
w10690 <= pi0092 and w84;
w10691 <= w936 and w9036;
w10692 <= w10690 and w10691;
w10693 <= w3416 and w3798;
w10694 <= w5166 and w10693;
w10695 <= w1033 and w3752;
w10696 <= w5169 and w10695;
w10697 <= not w10694 and not w10696;
w10698 <= w97 and w8774;
w10699 <= not w10697 and w10698;
w10700 <= not w10692 and not w10699;
w10701 <= w7726 and not w10700;
w10702 <= pi0093 and w8649;
w10703 <= w477 and w10702;
w10704 <= not pi0092 and not w10703;
w10705 <= not pi1050 and w84;
w10706 <= pi0092 and not w10705;
w10707 <= w7727 and not w10704;
w10708 <= not w10706 and w10707;
w10709 <= w8631 and w8847;
w10710 <= not w6451 and not w10709;
w10711 <= w487 and w10709;
w10712 <= pi1093 and not w10711;
w10713 <= w496 and not w10712;
w10714 <= w7806 and w8629;
w10715 <= not w343 and not w10714;
w10716 <= w280 and w7725;
w10717 <= pi0252 and w10716;
w10718 <= not w10715 and w10717;
w10719 <= not w10713 and not w10718;
w10720 <= w6468 and not w10719;
w10721 <= not w10709 and not w10720;
w10722 <= pi0252 and w10719;
w10723 <= not w10721 and not w10722;
w10724 <= w6451 and not w10723;
w10725 <= w7728 and not w10710;
w10726 <= not w10724 and w10725;
w10727 <= w80 and w9333;
w10728 <= w9021 and w10727;
w10729 <= not pi0332 and w7725;
w10730 <= w8846 and w10729;
w10731 <= w10665 and w10730;
w10732 <= not pi0039 and not w10731;
w10733 <= not w10728 and w10732;
w10734 <= not w8985 and w8988;
w10735 <= not w3955 and w10734;
w10736 <= not w3770 and not w3955;
w10737 <= w1034 and not w8982;
w10738 <= w10736 and w10737;
w10739 <= pi0039 and not w10735;
w10740 <= not w10738 and w10739;
w10741 <= w7763 and not w10733;
w10742 <= not w10740 and w10741;
w10743 <= w7888 and w10727;
w10744 <= pi0479 and w6468;
w10745 <= w746 and w10744;
w10746 <= pi0096 and w73;
w10747 <= w524 and w10746;
w10748 <= not w10744 and w10747;
w10749 <= w479 and w10748;
w10750 <= not w10745 and not w10749;
w10751 <= not pi0095 and not w10750;
w10752 <= not w10743 and not w10751;
w10753 <= w7728 and not w10752;
w10754 <= pi0039 and pi0593;
w10755 <= not w8990 and w10754;
w10756 <= not w3955 and w10755;
w10757 <= w3732 and w10744;
w10758 <= not w3841 and not w10757;
w10759 <= not pi0096 and w7756;
w10760 <= not w10758 and w10759;
w10761 <= w9049 and w10760;
w10762 <= not w10756 and not w10761;
w10763 <= w7763 and not w10762;
w10764 <= not pi0092 and w9037;
w10765 <= not w10690 and not w10764;
w10766 <= pi0314 and pi1050;
w10767 <= w7727 and w10766;
w10768 <= not w10765 and w10767;
w10769 <= not pi0072 and pi0152;
w10770 <= w7863 and w10769;
w10771 <= pi0299 and w10770;
w10772 <= not pi0072 and pi0174;
w10773 <= not pi0299 and w10772;
w10774 <= w7859 and w10773;
w10775 <= not w10771 and not w10774;
w10776 <= pi0232 and not w10775;
w10777 <= pi0039 and not w10776;
w10778 <= not pi0072 and pi0099;
w10779 <= not pi0039 and not w10778;
w10780 <= not w10777 and not w10779;
w10781 <= not w183 and w10780;
w10782 <= not w5069 and not w10778;
w10783 <= not w487 and w10778;
w10784 <= w5069 and not w10783;
w10785 <= not w7892 and w10778;
w10786 <= w3829 and w8482;
w10787 <= not w10785 and not w10786;
w10788 <= w7919 and not w10787;
w10789 <= w10784 and not w10788;
w10790 <= not w10782 and not w10789;
w10791 <= not pi0039 and not w10790;
w10792 <= w183 and not w10777;
w10793 <= not w10791 and w10792;
w10794 <= pi0075 and not w10781;
w10795 <= not w10793 and w10794;
w10796 <= pi0228 and w8063;
w10797 <= pi0228 and w7907;
w10798 <= w10778 and not w10797;
w10799 <= w94 and not w10798;
w10800 <= not w10796 and w10799;
w10801 <= not w94 and not w10780;
w10802 <= pi0087 and not w10801;
w10803 <= not w10800 and w10802;
w10804 <= pi0038 and not w10780;
w10805 <= w8041 and not w10775;
w10806 <= not w8511 and w10805;
w10807 <= pi0041 and pi0072;
w10808 <= pi0099 and not w10807;
w10809 <= not w7974 and w10808;
w10810 <= not pi0228 and not w8119;
w10811 <= not w10809 and w10810;
w10812 <= not w8022 and w10808;
w10813 <= w8342 and not w10812;
w10814 <= not w7989 and w10808;
w10815 <= w8341 and not w10814;
w10816 <= not w10813 and not w10815;
w10817 <= pi0228 and not w10816;
w10818 <= not pi0039 and not w10811;
w10819 <= not w10817 and w10818;
w10820 <= w171 and not w10806;
w10821 <= not w10819 and w10820;
w10822 <= not w7922 and w10778;
w10823 <= w3828 and w7881;
w10824 <= not w10822 and not w10823;
w10825 <= w7919 and not w10824;
w10826 <= w10784 and not w10825;
w10827 <= not w10782 and not w10826;
w10828 <= not pi0039 and not w10827;
w10829 <= not w10777 and not w10828;
w10830 <= w3848 and not w10829;
w10831 <= not pi0087 and not w10804;
w10832 <= not w10830 and w10831;
w10833 <= not w10821 and w10832;
w10834 <= not pi0075 and not w10803;
w10835 <= not w10833 and w10834;
w10836 <= not w10795 and not w10835;
w10837 <= w4992 and not w10836;
w10838 <= not w4992 and not w10780;
w10839 <= w4989 and not w10838;
w10840 <= not w10837 and w10839;
w10841 <= pi0232 and w10770;
w10842 <= pi0039 and not w10841;
w10843 <= not w4989 and not w10779;
w10844 <= not w10842 and w10843;
w10845 <= not w10840 and not w10844;
w10846 <= not w3826 and not w3844;
w10847 <= not w5036 and w7641;
w10848 <= pi0129 and not w10847;
w10849 <= w5035 and not w10848;
w10850 <= pi0129 and not w7641;
w10851 <= not w7644 and not w10850;
w10852 <= not w10846 and not w10851;
w10853 <= not w10849 and w10852;
w10854 <= not pi0075 and w172;
w10855 <= w3848 and w10854;
w10856 <= not w10853 and w10855;
w10857 <= not pi0024 and w6530;
w10858 <= not w6468 and w10857;
w10859 <= not w6527 and w10858;
w10860 <= not w10856 and not w10859;
w10861 <= w6444 and not w10860;
w10862 <= w84 and w10861;
w10863 <= not pi0039 and not w7885;
w10864 <= pi0152 and w952;
w10865 <= w3760 and w10864;
w10866 <= not pi0072 and w10865;
w10867 <= pi0299 and not w10866;
w10868 <= not pi0144 and pi0174;
w10869 <= w7858 and w10868;
w10870 <= not pi0072 and w10869;
w10871 <= not pi0299 and not w10870;
w10872 <= pi0232 and not w10867;
w10873 <= not w10871 and w10872;
w10874 <= pi0039 and not w10873;
w10875 <= not w10863 and not w10874;
w10876 <= not w183 and w10875;
w10877 <= not w5069 and not w7885;
w10878 <= not w487 and w7885;
w10879 <= w5069 and not w10878;
w10880 <= w487 and not w3836;
w10881 <= w7885 and not w7891;
w10882 <= not w7882 and not w10881;
w10883 <= w10880 and not w10882;
w10884 <= w10879 and not w10883;
w10885 <= not w10877 and not w10884;
w10886 <= not pi0039 and not w10885;
w10887 <= w183 and not w10874;
w10888 <= not w10886 and w10887;
w10889 <= pi0075 and not w10876;
w10890 <= not w10888 and w10889;
w10891 <= w7906 and w8494;
w10892 <= w7885 and not w10891;
w10893 <= not pi0101 and w8495;
w10894 <= not pi0039 and not w10892;
w10895 <= not w10893 and w10894;
w10896 <= pi0087 and not w10874;
w10897 <= not w10895 and w10896;
w10898 <= pi0038 and not w10875;
w10899 <= w8512 and w10865;
w10900 <= pi0299 and not w10899;
w10901 <= w8512 and w10869;
w10902 <= not pi0299 and not w10901;
w10903 <= w8041 and not w10900;
w10904 <= not w10902 and w10903;
w10905 <= pi0101 and w7972;
w10906 <= not pi0228 and not w7964;
w10907 <= not w10905 and w10906;
w10908 <= pi0101 and w8020;
w10909 <= w487 and not w8014;
w10910 <= not w10908 and w10909;
w10911 <= pi0101 and w7987;
w10912 <= not w487 and not w7996;
w10913 <= not w10911 and w10912;
w10914 <= not w10910 and not w10913;
w10915 <= pi0228 and not w10914;
w10916 <= not pi0039 and not w10907;
w10917 <= not w10915 and w10916;
w10918 <= w171 and not w10904;
w10919 <= not w10917 and w10918;
w10920 <= not pi0044 and w8503;
w10921 <= w7885 and not w10920;
w10922 <= not w7881 and not w10921;
w10923 <= w10880 and not w10922;
w10924 <= w10879 and not w10923;
w10925 <= not w10877 and not w10924;
w10926 <= not pi0039 and not w10925;
w10927 <= not w10874 and not w10926;
w10928 <= w3848 and not w10927;
w10929 <= not pi0087 and not w10898;
w10930 <= not w10928 and w10929;
w10931 <= not w10919 and w10930;
w10932 <= not pi0075 and not w10897;
w10933 <= not w10931 and w10932;
w10934 <= not w10890 and not w10933;
w10935 <= w4992 and not w10934;
w10936 <= not w4992 and not w10875;
w10937 <= w4989 and not w10936;
w10938 <= not w10935 and w10937;
w10939 <= pi0232 and w10866;
w10940 <= pi0039 and not w10939;
w10941 <= not w4989 and not w10863;
w10942 <= not w10940 and w10941;
w10943 <= not w10938 and not w10942;
w10944 <= w414 and w6485;
w10945 <= w10592 and w10944;
w10946 <= pi0109 and w328;
w10947 <= w262 and w10946;
w10948 <= pi0314 and not w10947;
w10949 <= not pi0109 and not w10639;
w10950 <= w3985 and not w10949;
w10951 <= not pi0314 and not w10950;
w10952 <= w8669 and not w10948;
w10953 <= not w10951 and w10952;
w10954 <= w4988 and not w6451;
w10955 <= w7638 and not w10954;
w10956 <= w7959 and not w10955;
w10957 <= not w3837 and not w10655;
w10958 <= not pi0110 and not w10653;
w10959 <= not pi0047 and w8606;
w10960 <= not w10958 and w10959;
w10961 <= w7941 and w10960;
w10962 <= w3837 and not w10961;
w10963 <= not w5037 and not w7637;
w10964 <= not w10957 and w10963;
w10965 <= not w10962 and w10964;
w10966 <= w5037 and not w7637;
w10967 <= w10961 and w10966;
w10968 <= not w10965 and not w10967;
w10969 <= not w4988 and not w10968;
w10970 <= not w10956 and not w10969;
w10971 <= w7728 and not w10970;
w10972 <= pi0024 and w8845;
w10973 <= not pi0053 and not w8844;
w10974 <= w286 and not w10973;
w10975 <= not pi0024 and w280;
w10976 <= w10974 and w10975;
w10977 <= not w10972 and not w10976;
w10978 <= pi0841 and not w10977;
w10979 <= w6509 and w8830;
w10980 <= not w10978 and not w10979;
w10981 <= w7729 and not w10980;
w10982 <= not pi0999 and w7729;
w10983 <= w8917 and w10982;
w10984 <= not pi0097 and w5005;
w10985 <= not pi0108 and not w10984;
w10986 <= w264 and not w10985;
w10987 <= w7807 and w10986;
w10988 <= not pi0314 and not w10987;
w10989 <= pi0314 and not w5007;
w10990 <= w5009 and not w7801;
w10991 <= not w10989 and w10990;
w10992 <= not w10988 and w10991;
w10993 <= w5009 and w7801;
w10994 <= w10987 and w10993;
w10995 <= not pi0051 and not w10994;
w10996 <= not w10992 and w10995;
w10997 <= w188 and w5081;
w10998 <= not w10996 and w10997;
w10999 <= not pi0087 and not w10998;
w11000 <= w3696 and w6444;
w11001 <= not w10999 and w11000;
w11002 <= w347 and w9005;
w11003 <= w10640 and w11002;
w11004 <= not pi0082 and not pi0109;
w11005 <= pi0111 and w11004;
w11006 <= w9937 and w11005;
w11007 <= w62 and w11006;
w11008 <= w8668 and w11007;
w11009 <= w364 and w11008;
w11010 <= pi0314 and w11009;
w11011 <= w6451 and w7638;
w11012 <= w7951 and w11011;
w11013 <= not w11010 and not w11012;
w11014 <= w7729 and not w11013;
w11015 <= pi0072 and w7888;
w11016 <= not pi0314 and w11009;
w11017 <= w6704 and w11016;
w11018 <= not w11015 and not w11017;
w11019 <= w4042 and w7728;
w11020 <= not w11018 and w11019;
w11021 <= pi0124 and not pi0468;
w11022 <= not pi0072 and pi0113;
w11023 <= not pi0039 and w11022;
w11024 <= pi0038 and not w11023;
w11025 <= w487 and w5069;
w11026 <= w5042 and w8094;
w11027 <= not w3835 and not w11026;
w11028 <= w11025 and not w11027;
w11029 <= w11022 and not w11028;
w11030 <= not w3835 and w11025;
w11031 <= not pi0113 and w11030;
w11032 <= w10823 and w11031;
w11033 <= not w11029 and not w11032;
w11034 <= not pi0039 and not w11033;
w11035 <= w3848 and not w11034;
w11036 <= pi0113 and w8113;
w11037 <= not pi0228 and not w8120;
w11038 <= not w11036 and w11037;
w11039 <= not pi0113 and w8343;
w11040 <= not w487 and not w7989;
w11041 <= not pi0099 and not w11040;
w11042 <= not w8023 and w11041;
w11043 <= pi0113 and not w8111;
w11044 <= not w11042 and w11043;
w11045 <= pi0228 and not w11039;
w11046 <= not w11044 and w11045;
w11047 <= not pi0039 and not w11038;
w11048 <= not w11046 and w11047;
w11049 <= w171 and not w11048;
w11050 <= not w11024 and not w11035;
w11051 <= not w11049 and w11050;
w11052 <= not pi0087 and not w11051;
w11053 <= not w171 and w11023;
w11054 <= not w8095 and w11022;
w11055 <= not pi0113 and w10796;
w11056 <= not w11054 and not w11055;
w11057 <= w94 and not w11056;
w11058 <= pi0087 and not w11053;
w11059 <= not w11057 and w11058;
w11060 <= not w11052 and not w11059;
w11061 <= not pi0075 and not w11060;
w11062 <= w5040 and w11032;
w11063 <= not w3835 and not w8059;
w11064 <= w11025 and not w11063;
w11065 <= w11022 and not w11064;
w11066 <= not w11062 and not w11065;
w11067 <= w173 and not w11066;
w11068 <= not w183 and w11023;
w11069 <= pi0075 and not w11068;
w11070 <= not w11067 and w11069;
w11071 <= not w11061 and not w11070;
w11072 <= w6444 and not w11071;
w11073 <= not w6444 and not w11023;
w11074 <= not w11072 and not w11073;
w11075 <= not pi0072 and pi0114;
w11076 <= not pi0039 and w11075;
w11077 <= not w183 and w11076;
w11078 <= not w8706 and not w11075;
w11079 <= pi0114 and w8298;
w11080 <= w8706 and not w11079;
w11081 <= not w8068 and w11080;
w11082 <= w173 and not w11078;
w11083 <= not w11081 and w11082;
w11084 <= pi0075 and not w11077;
w11085 <= not w11083 and w11084;
w11086 <= not w171 and not w11076;
w11087 <= pi0228 and w8179;
w11088 <= not pi0115 and w11087;
w11089 <= w11075 and not w11088;
w11090 <= w171 and not w11089;
w11091 <= not w8100 and w11090;
w11092 <= w8775 and not w11086;
w11093 <= not w11091 and w11092;
w11094 <= pi0038 and not w11076;
w11095 <= pi0114 and not w8181;
w11096 <= w8706 and not w11095;
w11097 <= not w8067 and w11096;
w11098 <= not pi0039 and not w11078;
w11099 <= not w11097 and w11098;
w11100 <= w3848 and not w11099;
w11101 <= not pi0114 and not w8346;
w11102 <= pi0114 and not w8354;
w11103 <= not w11101 and not w11102;
w11104 <= not pi0115 and not w11103;
w11105 <= pi0115 and not w11075;
w11106 <= not pi0039 and not w11105;
w11107 <= not w11104 and w11106;
w11108 <= w171 and not w11107;
w11109 <= not pi0087 and not w11094;
w11110 <= not w11100 and w11109;
w11111 <= not w11108 and w11110;
w11112 <= not pi0075 and not w11093;
w11113 <= not w11111 and w11112;
w11114 <= not w11085 and not w11113;
w11115 <= w6444 and not w11114;
w11116 <= not w6444 and not w11076;
w11117 <= not w11115 and not w11116;
w11118 <= not pi0072 and pi0115;
w11119 <= not pi0039 and w11118;
w11120 <= not w183 and w11119;
w11121 <= not w11025 and not w11118;
w11122 <= pi0115 and w8298;
w11123 <= not pi0052 and w8688;
w11124 <= not pi0115 and not w11123;
w11125 <= w8065 and w11124;
w11126 <= w5040 and w11125;
w11127 <= w11025 and not w11122;
w11128 <= not w11126 and w11127;
w11129 <= w173 and not w11121;
w11130 <= not w11128 and w11129;
w11131 <= pi0075 and not w11120;
w11132 <= not w11130 and w11131;
w11133 <= not w171 and not w11119;
w11134 <= not w11087 and w11118;
w11135 <= w171 and not w11134;
w11136 <= not w8099 and w11135;
w11137 <= w8775 and not w11133;
w11138 <= not w11136 and w11137;
w11139 <= pi0038 and not w11119;
w11140 <= pi0115 and not w8181;
w11141 <= w11025 and not w11140;
w11142 <= not w11125 and w11141;
w11143 <= not pi0039 and not w11121;
w11144 <= not w11142 and w11143;
w11145 <= w3848 and not w11144;
w11146 <= not pi0115 and not w8346;
w11147 <= pi0115 and not w8354;
w11148 <= not pi0039 and not w11146;
w11149 <= not w11147 and w11148;
w11150 <= w171 and not w11149;
w11151 <= not pi0087 and not w11139;
w11152 <= not w11145 and w11151;
w11153 <= not w11150 and w11152;
w11154 <= not pi0075 and not w11138;
w11155 <= not w11153 and w11154;
w11156 <= not w11132 and not w11155;
w11157 <= w6444 and not w11156;
w11158 <= not w6444 and not w11119;
w11159 <= not w11157 and not w11158;
w11160 <= not pi0072 and pi0116;
w11161 <= not pi0039 and w11160;
w11162 <= pi0038 and not w11161;
w11163 <= not pi0113 and w8095;
w11164 <= w11160 and not w11163;
w11165 <= not pi0038 and not w11164;
w11166 <= not w8098 and w11165;
w11167 <= not w11162 and not w11166;
w11168 <= not pi0100 and not w11167;
w11169 <= pi0100 and not w11161;
w11170 <= w8775 and not w11169;
w11171 <= not w11168 and w11170;
w11172 <= not w487 and w8143;
w11173 <= pi0116 and w8148;
w11174 <= not w487 and not w11173;
w11175 <= w487 and not w8131;
w11176 <= pi0116 and not w11175;
w11177 <= not w8136 and not w11176;
w11178 <= not w11174 and not w11177;
w11179 <= pi0228 and not w11172;
w11180 <= not w11178 and w11179;
w11181 <= pi0116 and w8115;
w11182 <= w8340 and not w11181;
w11183 <= not pi0039 and not w11182;
w11184 <= not w11180 and w11183;
w11185 <= w171 and not w11184;
w11186 <= not w11025 and w11160;
w11187 <= not pi0113 and w11026;
w11188 <= w11160 and not w11187;
w11189 <= not w8065 and not w11188;
w11190 <= w11030 and not w11189;
w11191 <= not w11186 and not w11190;
w11192 <= not pi0039 and not w11191;
w11193 <= w3848 and not w11192;
w11194 <= not pi0087 and not w11162;
w11195 <= not w11193 and w11194;
w11196 <= not w11185 and w11195;
w11197 <= not pi0075 and not w11171;
w11198 <= not w11196 and w11197;
w11199 <= not w8060 and w11160;
w11200 <= not w8301 and not w11199;
w11201 <= w11030 and not w11200;
w11202 <= not w11186 and not w11201;
w11203 <= w173 and not w11202;
w11204 <= not w183 and w11161;
w11205 <= pi0075 and not w11204;
w11206 <= not w11203 and w11205;
w11207 <= not w11198 and not w11206;
w11208 <= w6444 and not w11207;
w11209 <= not w6444 and not w11161;
w11210 <= not w11208 and not w11209;
w11211 <= w1249 and w4942;
w11212 <= not w1248 and not w11211;
w11213 <= not pi0038 and not w11212;
w11214 <= not pi0087 and not w11213;
w11215 <= w3696 and not w11214;
w11216 <= not pi0092 and not w11215;
w11217 <= not pi0054 and not w4868;
w11218 <= not pi0074 and w11217;
w11219 <= not w11216 and w11218;
w11220 <= not pi0055 and not w11219;
w11221 <= not w4910 and not w11220;
w11222 <= not pi0056 and not w11221;
w11223 <= not w3690 and not w11222;
w11224 <= not pi0062 and not w11223;
w11225 <= not pi0057 and w3863;
w11226 <= not w11224 and w11225;
w11227 <= not pi0079 and w9732;
w11228 <= pi0163 and w3760;
w11229 <= not w9241 and not w11228;
w11230 <= not pi0150 and not w11229;
w11231 <= pi0150 and w7262;
w11232 <= w9239 and w11231;
w11233 <= not w11230 and not w11232;
w11234 <= pi0232 and not w11233;
w11235 <= not w6552 and w11234;
w11236 <= pi0074 and not w11235;
w11237 <= pi0165 and w5036;
w11238 <= not pi0038 and not pi0054;
w11239 <= not w11237 and not w11238;
w11240 <= w6552 and w11239;
w11241 <= not pi0074 and not w11235;
w11242 <= not w11240 and w11241;
w11243 <= not w11236 and not w11242;
w11244 <= not w92 and not w11243;
w11245 <= w891 and not w11244;
w11246 <= not w7446 and not w11245;
w11247 <= pi0055 and not w11236;
w11248 <= pi0150 and w5036;
w11249 <= not pi0092 and w6845;
w11250 <= w11248 and w11249;
w11251 <= w6811 and w11238;
w11252 <= not w11250 and w11251;
w11253 <= not w11239 and not w11252;
w11254 <= w6552 and not w11253;
w11255 <= w11241 and not w11254;
w11256 <= w11247 and not w11255;
w11257 <= not pi0184 and not w9267;
w11258 <= pi0185 and not w11257;
w11259 <= not pi0185 and w11257;
w11260 <= w3760 and not w11258;
w11261 <= not w11259 and w11260;
w11262 <= not pi0299 and not w11261;
w11263 <= pi0299 and w11233;
w11264 <= pi0232 and not w11262;
w11265 <= not w11263 and w11264;
w11266 <= not w6552 and w11265;
w11267 <= pi0074 and not w11266;
w11268 <= not pi0055 and not w11267;
w11269 <= not pi0143 and not pi0299;
w11270 <= not pi0165 and pi0299;
w11271 <= not w11269 and not w11270;
w11272 <= w5036 and w11271;
w11273 <= w6552 and not w11272;
w11274 <= pi0054 and not w11273;
w11275 <= not w11266 and w11274;
w11276 <= pi0075 and not w11265;
w11277 <= pi0100 and not w11265;
w11278 <= pi0038 and not w11272;
w11279 <= not pi0100 and not w11278;
w11280 <= not pi0157 and pi0299;
w11281 <= not pi0178 and not pi0299;
w11282 <= not w11280 and not w11281;
w11283 <= w5036 and w11282;
w11284 <= w6845 and w11283;
w11285 <= w6812 and not w11284;
w11286 <= w11279 and not w11285;
w11287 <= not w11277 and not w11286;
w11288 <= w6768 and not w11287;
w11289 <= not pi0143 and not w6750;
w11290 <= pi0143 and not w6752;
w11291 <= pi0165 and not w11290;
w11292 <= not w11289 and w11291;
w11293 <= pi0143 and not pi0165;
w11294 <= w6757 and w11293;
w11295 <= pi0038 and not w11294;
w11296 <= not w11292 and w11295;
w11297 <= w131 and not w11296;
w11298 <= not pi0232 and w7095;
w11299 <= not w3760 and not w7095;
w11300 <= w3760 and not w7137;
w11301 <= not w11299 and not w11300;
w11302 <= pi0151 and pi0168;
w11303 <= not w11301 and w11302;
w11304 <= not w3760 and w7095;
w11305 <= pi0151 and not pi0168;
w11306 <= not w7169 and w11305;
w11307 <= not pi0168 and w7178;
w11308 <= pi0168 and w7175;
w11309 <= not pi0151 and not w11307;
w11310 <= not w11308 and w11309;
w11311 <= not w11306 and not w11310;
w11312 <= not w11304 and not w11311;
w11313 <= pi0150 and not w11303;
w11314 <= not w11312 and w11313;
w11315 <= pi0168 and w3760;
w11316 <= w7095 and not w11315;
w11317 <= pi0168 and w7069;
w11318 <= not pi0151 and not w11316;
w11319 <= not w11317 and w11318;
w11320 <= not w7208 and not w11299;
w11321 <= not pi0168 and w11320;
w11322 <= not w7008 and not w11299;
w11323 <= pi0168 and w11322;
w11324 <= pi0151 and not w11321;
w11325 <= not w11323 and w11324;
w11326 <= not pi0150 and not w11319;
w11327 <= not w11325 and w11326;
w11328 <= pi0299 and not w11327;
w11329 <= not w11314 and w11328;
w11330 <= not w7069 and not w11304;
w11331 <= not pi0173 and not w11330;
w11332 <= pi0173 and w11322;
w11333 <= not pi0185 and not w11331;
w11334 <= not w11332 and w11333;
w11335 <= w3760 and not w6954;
w11336 <= pi0173 and not w11299;
w11337 <= not w11335 and w11336;
w11338 <= not w7059 and not w11304;
w11339 <= not pi0173 and not w11338;
w11340 <= pi0185 and not w11337;
w11341 <= not w11339 and w11340;
w11342 <= pi0190 and not w11334;
w11343 <= not w11341 and w11342;
w11344 <= not pi0173 and not w7090;
w11345 <= pi0173 and not w7512;
w11346 <= w3760 and not w11344;
w11347 <= not w11345 and w11346;
w11348 <= pi0185 and not w11304;
w11349 <= not w11347 and w11348;
w11350 <= pi0173 and w11320;
w11351 <= not pi0173 and w7095;
w11352 <= not pi0185 and not w11351;
w11353 <= not w11350 and w11352;
w11354 <= not pi0190 and not w11353;
w11355 <= not w11349 and w11354;
w11356 <= not pi0299 and not w11355;
w11357 <= not w11343 and w11356;
w11358 <= pi0232 and not w11357;
w11359 <= not w11329 and w11358;
w11360 <= not pi0039 and not w11298;
w11361 <= not w11359 and w11360;
w11362 <= pi0168 and w6874;
w11363 <= pi0157 and w6887;
w11364 <= not w11362 and not w11363;
w11365 <= w3760 and w9310;
w11366 <= not w11364 and w11365;
w11367 <= pi0299 and not w11366;
w11368 <= not w11281 and not w11367;
w11369 <= w6811 and not w11368;
w11370 <= pi0178 and not w6901;
w11371 <= not pi0190 and not w11370;
w11372 <= not pi0299 and not w11371;
w11373 <= not w11369 and not w11372;
w11374 <= w3768 and not w6811;
w11375 <= w6614 and not w11374;
w11376 <= not pi0178 and w11375;
w11377 <= not w6877 and w11376;
w11378 <= not pi0299 and not w6866;
w11379 <= pi0178 and w11375;
w11380 <= not w6868 and w11379;
w11381 <= pi0190 and w11378;
w11382 <= not w11377 and w11381;
w11383 <= not w11380 and w11382;
w11384 <= pi0232 and not w11383;
w11385 <= not w11373 and w11384;
w11386 <= not pi0232 and w6811;
w11387 <= pi0039 and not w11386;
w11388 <= not w11385 and w11387;
w11389 <= not pi0038 and not w11388;
w11390 <= not w11361 and w11389;
w11391 <= w11297 and not w11390;
w11392 <= w5724 and not w11278;
w11393 <= not w6812 and w11392;
w11394 <= not w11277 and not w11393;
w11395 <= not w11391 and w11394;
w11396 <= w132 and not w11395;
w11397 <= not w11276 and not w11288;
w11398 <= not w11396 and w11397;
w11399 <= not pi0054 and not w11398;
w11400 <= not w11275 and not w11399;
w11401 <= not pi0074 and not w11400;
w11402 <= w11268 and not w11401;
w11403 <= w92 and not w11256;
w11404 <= not w11402 and w11403;
w11405 <= not w11246 and not w11404;
w11406 <= w6552 and w11237;
w11407 <= not w6552 and not w11234;
w11408 <= not w891 and not w11406;
w11409 <= not w11407 and w11408;
w11410 <= not w11236 and w11409;
w11411 <= not w11405 and not w11410;
w11412 <= pi0118 and w11411;
w11413 <= w6528 and not w11283;
w11414 <= w84 and w11413;
w11415 <= w11279 and not w11414;
w11416 <= not w11277 and not w11415;
w11417 <= w6768 and not w11416;
w11418 <= w4872 and w6624;
w11419 <= not w3807 and w10693;
w11420 <= not w3955 and w11419;
w11421 <= not pi0232 and not w11420;
w11422 <= not w11418 and w11421;
w11423 <= w3761 and not w3955;
w11424 <= pi0157 and not w6602;
w11425 <= not pi0157 and w6607;
w11426 <= pi0168 and not w11425;
w11427 <= not pi0157 and not pi0168;
w11428 <= not w6600 and w11427;
w11429 <= not w11424 and not w11428;
w11430 <= not w11426 and w11429;
w11431 <= not w11423 and not w11430;
w11432 <= w10693 and not w11431;
w11433 <= not pi0178 and not w3768;
w11434 <= w6606 and w11433;
w11435 <= not w11423 and not w11434;
w11436 <= pi0190 and not w11435;
w11437 <= pi0178 and not w6615;
w11438 <= not w11423 and w11437;
w11439 <= not pi0178 and not w10736;
w11440 <= not pi0190 and not w11438;
w11441 <= not w11439 and w11440;
w11442 <= not w11436 and not w11441;
w11443 <= w10695 and not w11442;
w11444 <= pi0232 and not w11443;
w11445 <= not w11432 and w11444;
w11446 <= pi0039 and not w11422;
w11447 <= not w11445 and w11446;
w11448 <= not w3732 and not w6683;
w11449 <= not pi0232 and not w6681;
w11450 <= not w11448 and w11449;
w11451 <= not w6681 and not w9361;
w11452 <= not w3760 and not w11451;
w11453 <= w6705 and w11305;
w11454 <= pi0168 and not w6696;
w11455 <= not pi0168 and not w6655;
w11456 <= not pi0151 and not w11454;
w11457 <= not w11455 and w11456;
w11458 <= not w11453 and not w11457;
w11459 <= w6657 and not w11458;
w11460 <= pi0150 and not w11459;
w11461 <= not pi0151 and w6692;
w11462 <= w6729 and not w11461;
w11463 <= w11315 and not w11462;
w11464 <= not pi0151 and w6681;
w11465 <= w6725 and not w11464;
w11466 <= not pi0168 and not w11465;
w11467 <= not pi0150 and not w11463;
w11468 <= not w11466 and w11467;
w11469 <= not w11460 and not w11468;
w11470 <= pi0299 and not w11452;
w11471 <= not w11469 and w11470;
w11472 <= not w3760 and not w6685;
w11473 <= w4042 and w6705;
w11474 <= pi0173 and w11473;
w11475 <= not pi0173 and w4042;
w11476 <= w6655 and w11475;
w11477 <= not w11474 and not w11476;
w11478 <= not pi0190 and w3760;
w11479 <= not w11477 and w11478;
w11480 <= not pi0173 and pi0190;
w11481 <= w6697 and w11480;
w11482 <= pi0185 and not w11481;
w11483 <= not w11479 and w11482;
w11484 <= pi0173 and w6713;
w11485 <= pi0190 and w6694;
w11486 <= not w11484 and w11485;
w11487 <= not pi0173 and w6681;
w11488 <= w6710 and not w11487;
w11489 <= not pi0190 and not w11488;
w11490 <= not pi0185 and not w11486;
w11491 <= not w11489 and w11490;
w11492 <= not w11483 and not w11491;
w11493 <= not pi0299 and not w11472;
w11494 <= not w11492 and w11493;
w11495 <= not w11471 and not w11494;
w11496 <= pi0232 and not w11495;
w11497 <= not pi0039 and not w11450;
w11498 <= not w11496 and w11497;
w11499 <= not w11447 and not w11498;
w11500 <= not pi0038 and not w11499;
w11501 <= w11297 and not w11500;
w11502 <= not w11277 and not w11392;
w11503 <= not w11501 and w11502;
w11504 <= w132 and not w11503;
w11505 <= not w11276 and not w11417;
w11506 <= not w11504 and w11505;
w11507 <= not pi0054 and not w11506;
w11508 <= not w11275 and not w11507;
w11509 <= not pi0074 and not w11508;
w11510 <= w11268 and not w11509;
w11511 <= pi0054 and w11237;
w11512 <= not pi0092 and w6552;
w11513 <= w6528 and w11512;
w11514 <= not w11248 and w11513;
w11515 <= not w11511 and w11514;
w11516 <= w84 and w11515;
w11517 <= w11242 and not w11516;
w11518 <= w11247 and not w11517;
w11519 <= w92 and not w11518;
w11520 <= not w11510 and w11519;
w11521 <= w11245 and not w11520;
w11522 <= not w11410 and not w11521;
w11523 <= not pi0118 and w11522;
w11524 <= not w11227 and not w11523;
w11525 <= not w11412 and w11524;
w11526 <= not pi0118 and not w6539;
w11527 <= w11522 and not w11526;
w11528 <= w11411 and w11526;
w11529 <= w11227 and not w11527;
w11530 <= not w11528 and w11529;
w11531 <= not w11525 and not w11530;
w11532 <= pi0128 and pi0228;
w11533 <= not w7726 and w11532;
w11534 <= w4947 and w6528;
w11535 <= not w11532 and not w11534;
w11536 <= pi0075 and not w11535;
w11537 <= pi0087 and not w11532;
w11538 <= w93 and w898;
w11539 <= not w11532 and not w11538;
w11540 <= pi0100 and not w11539;
w11541 <= not w166 and w1033;
w11542 <= w5169 and w11541;
w11543 <= not w1011 and w3416;
w11544 <= w5166 and w11543;
w11545 <= not w11542 and not w11544;
w11546 <= pi0039 and not w11545;
w11547 <= pi0299 and w3981;
w11548 <= not w4091 and not w11547;
w11549 <= w5036 and not w11548;
w11550 <= pi0109 and not w11549;
w11551 <= not w491 and w9231;
w11552 <= w333 and w7720;
w11553 <= w9230 and not w11552;
w11554 <= w346 and not w11553;
w11555 <= not pi0097 and not w11554;
w11556 <= not pi0046 and w491;
w11557 <= w499 and w11556;
w11558 <= not w11555 and w11557;
w11559 <= not w11550 and not w11551;
w11560 <= not w11558 and w11559;
w11561 <= not w3985 and not w11549;
w11562 <= not w4054 and w11549;
w11563 <= not w11561 and not w11562;
w11564 <= not w11560 and w11563;
w11565 <= not pi0091 and not w11564;
w11566 <= w501 and not w3982;
w11567 <= not w11565 and w11566;
w11568 <= not w315 and not w11567;
w11569 <= not pi0039 and w8649;
w11570 <= not w11568 and w11569;
w11571 <= not w11546 and not w11570;
w11572 <= not pi0038 and not w11571;
w11573 <= not pi0228 and w11572;
w11574 <= not w11532 and not w11573;
w11575 <= not pi0100 and not w11574;
w11576 <= not pi0087 and not w11540;
w11577 <= not w11575 and w11576;
w11578 <= not pi0075 and not w11537;
w11579 <= not w11577 and w11578;
w11580 <= not pi0092 and not w11536;
w11581 <= not w11579 and w11580;
w11582 <= pi0092 and not w11532;
w11583 <= not w4932 and w11582;
w11584 <= w7726 and not w11583;
w11585 <= not w11581 and w11584;
w11586 <= not w11533 and not w11585;
w11587 <= not pi0031 and not pi0080;
w11588 <= pi0818 and w11587;
w11589 <= w4983 and not w4992;
w11590 <= not w4988 and not w11589;
w11591 <= not pi0120 and not w4992;
w11592 <= not pi1093 and w11591;
w11593 <= w11590 and not w11592;
w11594 <= pi0120 and not w4983;
w11595 <= not pi0120 and pi1093;
w11596 <= not pi1091 and w9873;
w11597 <= w11595 and not w11596;
w11598 <= not w11594 and not w11597;
w11599 <= w84 and w5158;
w11600 <= not w5182 and w11594;
w11601 <= w11599 and not w11600;
w11602 <= w5182 and not w11595;
w11603 <= not w11601 and not w11602;
w11604 <= w93 and w5069;
w11605 <= not w11603 and w11604;
w11606 <= pi0100 and not w11598;
w11607 <= not w11605 and w11606;
w11608 <= pi0038 and w4983;
w11609 <= not pi1093 and w5023;
w11610 <= pi0120 and w11609;
w11611 <= not pi0039 and not w11610;
w11612 <= pi0122 and not w5015;
w11613 <= w5097 and not w8008;
w11614 <= w4980 and w5014;
w11615 <= not pi0829 and w11614;
w11616 <= not pi0122 and not w11615;
w11617 <= not w11613 and w11616;
w11618 <= not w486 and not w11612;
w11619 <= not w11617 and w11618;
w11620 <= w493 and not w11619;
w11621 <= w5189 and not w11614;
w11622 <= not w9873 and w11621;
w11623 <= not w11620 and not w11622;
w11624 <= w11611 and w11623;
w11625 <= not w5133 and w11598;
w11626 <= not w3761 and w11598;
w11627 <= not w5165 and w11594;
w11628 <= pi1091 and pi1092;
w11629 <= w5117 and w11628;
w11630 <= w11597 and not w11629;
w11631 <= not w11627 and not w11630;
w11632 <= w3761 and w11631;
w11633 <= not w11626 and not w11632;
w11634 <= w3805 and w11633;
w11635 <= w3790 and not w11598;
w11636 <= not w3790 and not w11631;
w11637 <= not w11635 and not w11636;
w11638 <= not w3805 and not w11637;
w11639 <= w5133 and not w11634;
w11640 <= not w11638 and w11639;
w11641 <= pi0299 and not w11625;
w11642 <= not w11640 and w11641;
w11643 <= w3768 and w11633;
w11644 <= not w3768 and not w11637;
w11645 <= w5114 and not w11643;
w11646 <= not w11644 and w11645;
w11647 <= not w5114 and w11598;
w11648 <= not pi0299 and not w11647;
w11649 <= not w11646 and w11648;
w11650 <= pi0039 and not w11642;
w11651 <= not w11649 and w11650;
w11652 <= not w11624 and not w11651;
w11653 <= not pi0038 and not w11652;
w11654 <= not pi0120 and not pi1093;
w11655 <= pi0038 and w11654;
w11656 <= not pi0100 and not w11655;
w11657 <= not w11608 and w11656;
w11658 <= not w11653 and w11657;
w11659 <= not w11607 and not w11658;
w11660 <= not pi0087 and not w11659;
w11661 <= w5194 and not w11654;
w11662 <= not w188 and w4983;
w11663 <= w5189 and not w9873;
w11664 <= not w5059 and w11663;
w11665 <= w5192 and not w11664;
w11666 <= pi0087 and not w11662;
w11667 <= not w11665 and w11666;
w11668 <= w11661 and w11667;
w11669 <= not w11660 and not w11668;
w11670 <= not pi0075 and not w11669;
w11671 <= w5037 and w11598;
w11672 <= not w5159 and w11597;
w11673 <= not pi1091 and not w4982;
w11674 <= not w5045 and not w11673;
w11675 <= pi0120 and not w11674;
w11676 <= not w5037 and not w11675;
w11677 <= not w11672 and w11676;
w11678 <= not w11671 and not w11677;
w11679 <= w173 and not w11678;
w11680 <= not w173 and w11598;
w11681 <= pi0075 and not w11680;
w11682 <= not w11679 and w11681;
w11683 <= w4992 and not w11682;
w11684 <= not w11670 and w11683;
w11685 <= w11593 and not w11684;
w11686 <= w5162 and not w11654;
w11687 <= not w11620 and not w11621;
w11688 <= w11611 and w11687;
w11689 <= pi1093 and not w3761;
w11690 <= w3805 and w11689;
w11691 <= w3790 and not w3805;
w11692 <= w5133 and not w11691;
w11693 <= not w11690 and w11692;
w11694 <= w5165 and w11693;
w11695 <= pi0299 and not w11654;
w11696 <= not w11694 and w11695;
w11697 <= w3768 and w11689;
w11698 <= not w3768 and w3790;
w11699 <= w5114 and not w11698;
w11700 <= not w11697 and w11699;
w11701 <= w5165 and w11700;
w11702 <= not pi0299 and not w11654;
w11703 <= not w11701 and w11702;
w11704 <= pi0039 and not w11696;
w11705 <= not w11703 and w11704;
w11706 <= not w11688 and not w11705;
w11707 <= not pi0038 and not w11706;
w11708 <= w11656 and not w11707;
w11709 <= pi0120 and w5182;
w11710 <= not pi0120 and w11599;
w11711 <= not w11709 and not w11710;
w11712 <= w11604 and not w11711;
w11713 <= pi0100 and not w11654;
w11714 <= not w11712 and w11713;
w11715 <= not w11708 and not w11714;
w11716 <= not pi0087 and not w11715;
w11717 <= not w11661 and not w11716;
w11718 <= not pi0075 and not w11717;
w11719 <= w4992 and not w11686;
w11720 <= not w11718 and w11719;
w11721 <= w4988 and not w11592;
w11722 <= not w11720 and w11721;
w11723 <= not w11685 and not w11722;
w11724 <= w11588 and not w11723;
w11725 <= w4989 and not w11724;
w11726 <= not w4988 and w11598;
w11727 <= pi0120 and not w11726;
w11728 <= w11588 and not w11654;
w11729 <= not w11726 and w11728;
w11730 <= not w4989 and not w11729;
w11731 <= not w11727 and w11730;
w11732 <= not w5206 and not w11731;
w11733 <= pi0951 and pi0982;
w11734 <= pi1092 and w11733;
w11735 <= pi1093 and w11734;
w11736 <= not pi0120 and not w11735;
w11737 <= not w11726 and not w11736;
w11738 <= w11730 and not w11737;
w11739 <= w5206 and not w11738;
w11740 <= not w11732 and not w11739;
w11741 <= not w11725 and not w11740;
w11742 <= w11591 and not w11735;
w11743 <= not w173 and not w11736;
w11744 <= pi0120 and w5160;
w11745 <= not pi1091 and w11735;
w11746 <= not pi0120 and not w11745;
w11747 <= w493 and w11734;
w11748 <= not pi0093 and not pi0122;
w11749 <= w69 and w11748;
w11750 <= w488 and w6457;
w11751 <= w11749 and w11750;
w11752 <= w525 and w11751;
w11753 <= w7887 and w11752;
w11754 <= w5041 and w11753;
w11755 <= w266 and w11754;
w11756 <= w11747 and not w11755;
w11757 <= w11746 and not w11756;
w11758 <= not w11744 and not w11757;
w11759 <= not w5037 and not w11758;
w11760 <= w5037 and w11736;
w11761 <= w173 and not w11760;
w11762 <= not w11759 and w11761;
w11763 <= pi0075 and not w11743;
w11764 <= not w11762 and w11763;
w11765 <= not w188 and w11736;
w11766 <= pi0087 and not w11765;
w11767 <= pi0950 and w84;
w11768 <= not w486 and not w3776;
w11769 <= w11767 and w11768;
w11770 <= w11747 and not w11769;
w11771 <= pi0824 and w11767;
w11772 <= w11745 and not w11771;
w11773 <= not w11770 and not w11772;
w11774 <= not pi0120 and not w11773;
w11775 <= not w5190 and not w5191;
w11776 <= pi0120 and not w11775;
w11777 <= w188 and not w11776;
w11778 <= not w11774 and w11777;
w11779 <= w11766 and not w11778;
w11780 <= w4993 and w5041;
w11781 <= w11767 and w11780;
w11782 <= w11747 and not w11781;
w11783 <= w11746 and not w11782;
w11784 <= not w11709 and not w11783;
w11785 <= not pi0039 and w5069;
w11786 <= not w11784 and w11785;
w11787 <= pi0100 and not w11786;
w11788 <= not pi0038 and not w11787;
w11789 <= not w11604 and w11736;
w11790 <= not w11788 and not w11789;
w11791 <= not w5114 and w11736;
w11792 <= not pi0299 and not w11791;
w11793 <= not w6184 and not w11736;
w11794 <= not w3768 and w11793;
w11795 <= not w6187 and not w11736;
w11796 <= w3768 and w11795;
w11797 <= w5114 and not w11794;
w11798 <= not w11796 and w11797;
w11799 <= w11792 and not w11798;
w11800 <= not w5133 and w11736;
w11801 <= pi0299 and not w11800;
w11802 <= not w3805 and w11793;
w11803 <= w3805 and w11795;
w11804 <= w5133 and not w11802;
w11805 <= not w11803 and w11804;
w11806 <= w11801 and not w11805;
w11807 <= not w11799 and not w11806;
w11808 <= pi0039 and not w11807;
w11809 <= w334 and w5000;
w11810 <= w330 and w11809;
w11811 <= w6673 and w11810;
w11812 <= w4994 and w11811;
w11813 <= w4999 and not w11812;
w11814 <= pi0950 and w5081;
w11815 <= not w11813 and w11814;
w11816 <= pi0824 and w11815;
w11817 <= w11734 and not w11816;
w11818 <= not pi0829 and w11817;
w11819 <= not pi0097 and not w11810;
w11820 <= w498 and not w11819;
w11821 <= w500 and w11820;
w11822 <= not w5085 and not w11821;
w11823 <= w24 and not w11822;
w11824 <= w4997 and not w11823;
w11825 <= w4994 and not w11824;
w11826 <= not pi0051 and not w11825;
w11827 <= not w310 and not w11826;
w11828 <= not pi0096 and not w11827;
w11829 <= not pi0072 and pi0950;
w11830 <= w7979 and w11829;
w11831 <= not w11828 and w11830;
w11832 <= w4993 and w11734;
w11833 <= not w11831 and w11832;
w11834 <= pi0829 and pi1092;
w11835 <= pi0122 and w11733;
w11836 <= w11834 and w11835;
w11837 <= not w11815 and w11836;
w11838 <= not w11818 and not w11837;
w11839 <= not w11833 and w11838;
w11840 <= w5080 and not w11839;
w11841 <= w486 and w11735;
w11842 <= not w11840 and not w11841;
w11843 <= pi1091 and not w11842;
w11844 <= w11745 and not w11816;
w11845 <= not pi0120 and not w11844;
w11846 <= not w11843 and w11845;
w11847 <= not w11609 and w11687;
w11848 <= pi0120 and w11847;
w11849 <= not pi0039 and not w11846;
w11850 <= not w11848 and w11849;
w11851 <= not w11808 and not w11850;
w11852 <= w171 and not w11851;
w11853 <= not w11790 and not w11852;
w11854 <= not pi0087 and not w11853;
w11855 <= not pi0075 and not w11779;
w11856 <= not w11854 and w11855;
w11857 <= not w11764 and not w11856;
w11858 <= w4992 and not w11857;
w11859 <= w4988 and not w11858;
w11860 <= not w11598 and not w11736;
w11861 <= not w93 and not w11860;
w11862 <= not w5069 and w11860;
w11863 <= not w9873 and w11745;
w11864 <= not w11782 and not w11863;
w11865 <= not pi0120 and not w11864;
w11866 <= not w11600 and not w11865;
w11867 <= w5069 and not w11866;
w11868 <= w93 and not w11862;
w11869 <= not w11867 and w11868;
w11870 <= pi0100 and not w11861;
w11871 <= not w11869 and w11870;
w11872 <= pi0038 and not w11860;
w11873 <= not w11609 and w11623;
w11874 <= pi0120 and w11873;
w11875 <= w11663 and w11817;
w11876 <= not pi0120 and not w11875;
w11877 <= not w11843 and w11876;
w11878 <= not w11874 and not w11877;
w11879 <= not pi0039 and not w11878;
w11880 <= not w5117 and w11747;
w11881 <= not w11863 and not w11880;
w11882 <= not pi0120 and not w11881;
w11883 <= not w11627 and not w11882;
w11884 <= w3761 and not w11883;
w11885 <= not w3761 and w11860;
w11886 <= not w11884 and not w11885;
w11887 <= w3768 and not w11886;
w11888 <= not w3790 and not w11883;
w11889 <= w3790 and w11860;
w11890 <= not w11888 and not w11889;
w11891 <= not w3768 and not w11890;
w11892 <= w5114 and not w11887;
w11893 <= not w11891 and w11892;
w11894 <= not w11647 and w11792;
w11895 <= not w11893 and w11894;
w11896 <= w3805 and not w11886;
w11897 <= not w3805 and not w11890;
w11898 <= w5133 and not w11896;
w11899 <= not w11897 and w11898;
w11900 <= w4983 and not w5133;
w11901 <= w11801 and not w11900;
w11902 <= not w11899 and w11901;
w11903 <= pi0039 and not w11895;
w11904 <= not w11902 and w11903;
w11905 <= not w11879 and not w11904;
w11906 <= not pi0038 and not w11905;
w11907 <= not pi0100 and not w11872;
w11908 <= not w11906 and w11907;
w11909 <= not w11871 and not w11908;
w11910 <= not pi0087 and not w11909;
w11911 <= not w11665 and not w11777;
w11912 <= not w11770 and not w11863;
w11913 <= w11774 and not w11912;
w11914 <= not w11911 and not w11913;
w11915 <= not w11662 and w11766;
w11916 <= not w11914 and w11915;
w11917 <= not w11910 and not w11916;
w11918 <= not pi0075 and not w11917;
w11919 <= w5037 and not w11860;
w11920 <= not w11756 and not w11863;
w11921 <= not pi0120 and not w11920;
w11922 <= w11676 and not w11921;
w11923 <= not w11919 and not w11922;
w11924 <= w173 and not w11923;
w11925 <= not w173 and not w11860;
w11926 <= pi0075 and not w11925;
w11927 <= not w11924 and w11926;
w11928 <= w4992 and not w11927;
w11929 <= not w11918 and w11928;
w11930 <= w11593 and not w11929;
w11931 <= not w11859 and not w11930;
w11932 <= w11739 and not w11742;
w11933 <= not w11931 and w11932;
w11934 <= not w4983 and w5186;
w11935 <= not pi0039 and not w11873;
w11936 <= w4983 and not w5114;
w11937 <= not w5119 and not w11673;
w11938 <= w3761 and not w11937;
w11939 <= not w3761 and not w4983;
w11940 <= not w11938 and not w11939;
w11941 <= w3768 and not w11940;
w11942 <= not w3790 and not w11937;
w11943 <= w3790 and not w4983;
w11944 <= not w11942 and not w11943;
w11945 <= not w3768 and not w11944;
w11946 <= w5114 and not w11941;
w11947 <= not w11945 and w11946;
w11948 <= not pi0299 and not w11936;
w11949 <= not w11947 and w11948;
w11950 <= w3805 and not w11940;
w11951 <= not w3805 and not w11944;
w11952 <= w5133 and not w11950;
w11953 <= not w11951 and w11952;
w11954 <= pi0299 and not w11900;
w11955 <= not w11953 and w11954;
w11956 <= not w11949 and not w11955;
w11957 <= pi0039 and not w11956;
w11958 <= not pi0038 and not w11957;
w11959 <= not w11935 and w11958;
w11960 <= not pi0100 and not w11608;
w11961 <= not w11959 and w11960;
w11962 <= not w11934 and not w11961;
w11963 <= not pi0087 and not w11962;
w11964 <= not w11667 and not w11963;
w11965 <= not pi0075 and not w11964;
w11966 <= w4983 and not w5038;
w11967 <= w5038 and w11674;
w11968 <= pi0075 and not w11966;
w11969 <= not w11967 and w11968;
w11970 <= not w11965 and not w11969;
w11971 <= w11590 and not w11970;
w11972 <= not w4992 and not w11726;
w11973 <= not pi0039 and not w11847;
w11974 <= w5175 and not w11973;
w11975 <= not pi0100 and not w11974;
w11976 <= not w5186 and not w11975;
w11977 <= not pi0087 and not w11976;
w11978 <= not w5194 and not w11977;
w11979 <= not pi0075 and not w11978;
w11980 <= not w5162 and not w11979;
w11981 <= w4988 and not w11591;
w11982 <= not w11980 and w11981;
w11983 <= not w11971 and not w11972;
w11984 <= not w11982 and w11983;
w11985 <= pi0120 and w11732;
w11986 <= not w11984 and w11985;
w11987 <= not w11933 and not w11986;
w11988 <= not w11588 and not w11987;
w11989 <= not w11741 and not w11988;
w11990 <= not pi0134 and not pi0135;
w11991 <= not pi0136 and w11990;
w11992 <= not pi0130 and w11991;
w11993 <= not pi0132 and w11992;
w11994 <= not pi0126 and w11993;
w11995 <= not pi0121 and w11994;
w11996 <= not pi0125 and not pi0133;
w11997 <= pi0121 and not w11996;
w11998 <= not pi0121 and w11996;
w11999 <= not w11997 and not w11998;
w12000 <= not w11995 and not w11999;
w12001 <= w41 and w7715;
w12002 <= not pi0051 and w12001;
w12003 <= not pi0087 and w12002;
w12004 <= not w12000 and w12003;
w12005 <= pi0051 and pi0146;
w12006 <= pi0051 and w3760;
w12007 <= not pi0146 and w12006;
w12008 <= pi0161 and not w12007;
w12009 <= w3760 and not w12002;
w12010 <= not w12005 and not w12008;
w12011 <= w12009 and w12010;
w12012 <= not pi0087 and not w12011;
w12013 <= pi0087 and not w11228;
w12014 <= pi0232 and not w12013;
w12015 <= not w12012 and w12014;
w12016 <= not w4989 and not w12004;
w12017 <= not w12015 and w12016;
w12018 <= not pi0087 and not w133;
w12019 <= not w12002 and w12018;
w12020 <= not pi0142 and w12006;
w12021 <= pi0144 and not w12020;
w12022 <= pi0051 and pi0142;
w12023 <= w12009 and not w12022;
w12024 <= not w12021 and w12023;
w12025 <= not pi0299 and not w12024;
w12026 <= pi0299 and not w12011;
w12027 <= pi0232 and not w12025;
w12028 <= not w12026 and w12027;
w12029 <= w12019 and not w12028;
w12030 <= pi0100 and w12002;
w12031 <= w98 and not w12030;
w12032 <= pi0100 and w12028;
w12033 <= pi0038 and not w12028;
w12034 <= not pi0100 and not w12033;
w12035 <= pi0038 and not w12002;
w12036 <= not pi0100 and not w12035;
w12037 <= not w12034 and not w12036;
w12038 <= not pi0161 and not w12007;
w12039 <= w268 and w5008;
w12040 <= not pi0024 and pi0314;
w12041 <= w12039 and w12040;
w12042 <= w30 and w7714;
w12043 <= w10610 and w12042;
w12044 <= not pi0050 and pi0077;
w12045 <= w58 and w12044;
w12046 <= w12043 and w12045;
w12047 <= w6460 and w12041;
w12048 <= w12046 and w12047;
w12049 <= w82 and w12048;
w12050 <= w333 and w12043;
w12051 <= not pi0058 and w12039;
w12052 <= w6816 and w12051;
w12053 <= w12050 and w12052;
w12054 <= pi0072 and w4042;
w12055 <= w12053 and w12054;
w12056 <= w12001 and not w12039;
w12057 <= not pi0051 and not w12056;
w12058 <= not pi0024 and w9226;
w12059 <= w12050 and w12058;
w12060 <= pi0086 and w12050;
w12061 <= not w12046 and not w12060;
w12062 <= w8639 and not w12061;
w12063 <= w12001 and not w12059;
w12064 <= not w12062 and w12063;
w12065 <= w12057 and not w12064;
w12066 <= w82 and w12065;
w12067 <= w12002 and not w12066;
w12068 <= not w12055 and w12067;
w12069 <= not w12049 and w12068;
w12070 <= not w3760 and not w12069;
w12071 <= pi0072 and w7905;
w12072 <= not w12006 and not w12071;
w12073 <= w3760 and not w12072;
w12074 <= not w12070 and not w12073;
w12075 <= w12038 and not w12074;
w12076 <= w12002 and not w12049;
w12077 <= not w12066 and w12076;
w12078 <= not w3760 and not w12077;
w12079 <= not w12009 and not w12078;
w12080 <= not w12055 and w12079;
w12081 <= pi0146 and w12080;
w12082 <= not pi0051 and w3760;
w12083 <= w12001 and not w12055;
w12084 <= w12082 and not w12083;
w12085 <= not pi0146 and not w12084;
w12086 <= not w12070 and w12085;
w12087 <= pi0161 and not w12081;
w12088 <= not w12086 and w12087;
w12089 <= not w12075 and not w12088;
w12090 <= w7135 and not w12089;
w12091 <= not w3760 and w12069;
w12092 <= not pi0051 and w12041;
w12093 <= w11002 and w12092;
w12094 <= not pi0072 and not w12093;
w12095 <= w4043 and not w12094;
w12096 <= w3760 and not w12095;
w12097 <= not w12091 and not w12096;
w12098 <= not pi0146 and not w12097;
w12099 <= w82 and w3760;
w12100 <= w12093 and w12099;
w12101 <= w12074 and not w12100;
w12102 <= pi0146 and w12101;
w12103 <= not pi0161 and not w12098;
w12104 <= not w12102 and w12103;
w12105 <= w12082 and w12083;
w12106 <= not w12049 and w12105;
w12107 <= not w12006 and not w12106;
w12108 <= pi0146 and not w12002;
w12109 <= not w12107 and not w12108;
w12110 <= pi0161 and not w12109;
w12111 <= not w12091 and w12110;
w12112 <= not w12104 and not w12111;
w12113 <= w7166 and not w12112;
w12114 <= not w12090 and not w12113;
w12115 <= pi0156 and not w12114;
w12116 <= pi0144 and not w12080;
w12117 <= not pi0144 and not w12074;
w12118 <= not w12116 and not w12117;
w12119 <= not w12020 and not w12118;
w12120 <= pi0180 and not w12119;
w12121 <= not pi0142 and not w12097;
w12122 <= pi0142 and w12101;
w12123 <= not pi0144 and not w12121;
w12124 <= not w12122 and w12123;
w12125 <= not w12049 and w12080;
w12126 <= w12021 and not w12125;
w12127 <= not pi0180 and not w12126;
w12128 <= not w12124 and w12127;
w12129 <= pi0179 and not w12120;
w12130 <= not w12128 and w12129;
w12131 <= w12021 and not w12069;
w12132 <= not pi0024 and not w9227;
w12133 <= pi0024 and not w9232;
w12134 <= not w12132 and not w12133;
w12135 <= not pi0314 and not w12134;
w12136 <= pi0314 and not w9232;
w12137 <= not w12135 and not w12136;
w12138 <= w5008 and w6523;
w12139 <= w12137 and w12138;
w12140 <= not pi0051 and not w12139;
w12141 <= not w12071 and w12140;
w12142 <= w3760 and not w12141;
w12143 <= not w12070 and not w12142;
w12144 <= pi0142 and w12143;
w12145 <= w271 and w12137;
w12146 <= not pi0072 and not w12145;
w12147 <= w4043 and not w12146;
w12148 <= w3760 and not w12147;
w12149 <= not w12091 and not w12148;
w12150 <= not pi0142 and not w12149;
w12151 <= not pi0144 and not w12144;
w12152 <= not w12150 and w12151;
w12153 <= not pi0180 and not w12131;
w12154 <= not w12152 and w12153;
w12155 <= not w12068 and w12082;
w12156 <= not w12070 and not w12155;
w12157 <= w3760 and not w12067;
w12158 <= not pi0142 and not w12157;
w12159 <= not pi0051 and not w12001;
w12160 <= w3760 and w12159;
w12161 <= not w12099 and not w12160;
w12162 <= w82 and not w12065;
w12163 <= not w12161 and not w12162;
w12164 <= pi0142 and not w12163;
w12165 <= not w12158 and not w12164;
w12166 <= not w12079 and not w12165;
w12167 <= w12156 and not w12166;
w12168 <= pi0144 and not w12167;
w12169 <= w271 and w12134;
w12170 <= not pi0072 and not w12169;
w12171 <= w4043 and not w12170;
w12172 <= w3760 and not w12171;
w12173 <= not w12091 and not w12172;
w12174 <= not pi0142 and not w12173;
w12175 <= w12099 and w12169;
w12176 <= not w12073 and not w12175;
w12177 <= not w12070 and w12176;
w12178 <= pi0142 and w12177;
w12179 <= not pi0144 and not w12178;
w12180 <= not w12174 and w12179;
w12181 <= pi0180 and not w12168;
w12182 <= not w12180 and w12181;
w12183 <= not pi0179 and not w12182;
w12184 <= not w12154 and w12183;
w12185 <= not w12130 and not w12184;
w12186 <= not pi0299 and not w12185;
w12187 <= pi0146 and w12177;
w12188 <= not pi0146 and not w12173;
w12189 <= w7135 and not w12187;
w12190 <= not w12188 and w12189;
w12191 <= not pi0146 and not w12149;
w12192 <= pi0146 and w12143;
w12193 <= w7166 and not w12191;
w12194 <= not w12192 and w12193;
w12195 <= not pi0161 and not w12190;
w12196 <= not w12194 and w12195;
w12197 <= not pi0146 and not w12157;
w12198 <= pi0146 and not w12163;
w12199 <= not w12197 and not w12198;
w12200 <= not w12079 and not w12199;
w12201 <= w12156 and not w12200;
w12202 <= w7135 and not w12201;
w12203 <= w7166 and not w12007;
w12204 <= not w12069 and w12203;
w12205 <= pi0161 and not w12204;
w12206 <= not w12202 and w12205;
w12207 <= not pi0156 and not w12206;
w12208 <= not w12196 and w12207;
w12209 <= not w12115 and not w12208;
w12210 <= not w12186 and w12209;
w12211 <= w6722 and not w12210;
w12212 <= w82 and w12053;
w12213 <= not w4203 and not w5170;
w12214 <= w12212 and not w12213;
w12215 <= not pi0232 and w12002;
w12216 <= not w12214 and w12215;
w12217 <= w12002 and not w12212;
w12218 <= not pi0051 and not w12217;
w12219 <= not pi0287 and not w12218;
w12220 <= not pi0287 and w3760;
w12221 <= not w12160 and not w12220;
w12222 <= not w12219 and not w12221;
w12223 <= not w12023 and not w12222;
w12224 <= w6614 and not w12223;
w12225 <= w12001 and w12224;
w12226 <= not w12002 and not w12020;
w12227 <= not w3968 and not w12226;
w12228 <= pi0144 and not w12227;
w12229 <= pi0051 and not w3760;
w12230 <= not w12218 and not w12229;
w12231 <= w3968 and not w12022;
w12232 <= w12230 and w12231;
w12233 <= w12228 and not w12232;
w12234 <= not w12225 and w12233;
w12235 <= not w3760 and not w12217;
w12236 <= not w3785 and not w12235;
w12237 <= not pi0142 and not w12236;
w12238 <= w78 and w5013;
w12239 <= not pi0051 and not w12238;
w12240 <= w3760 and not w12239;
w12241 <= not w12235 and not w12240;
w12242 <= pi0142 and not w12241;
w12243 <= w3968 and not w12237;
w12244 <= not w12242 and w12243;
w12245 <= not w6614 and not w12244;
w12246 <= not pi0051 and w12220;
w12247 <= not w12241 and not w12246;
w12248 <= pi0224 and not w12020;
w12249 <= w12247 and w12248;
w12250 <= not w12245 and not w12249;
w12251 <= not w3968 and w12160;
w12252 <= not w12227 and not w12251;
w12253 <= not w12228 and w12252;
w12254 <= not w12250 and w12253;
w12255 <= pi0181 and not w12234;
w12256 <= not w12254 and w12255;
w12257 <= not w12244 and w12253;
w12258 <= not pi0181 and not w12233;
w12259 <= not w12257 and w12258;
w12260 <= not pi0299 and not w12259;
w12261 <= not w12256 and w12260;
w12262 <= not w12007 and not w12217;
w12263 <= pi0161 and not w12262;
w12264 <= not pi0146 and not w12236;
w12265 <= pi0146 and not w12241;
w12266 <= not pi0161 and not w12264;
w12267 <= not w12265 and w12266;
w12268 <= not w12263 and not w12267;
w12269 <= w3942 and not w12268;
w12270 <= not w12002 and not w12011;
w12271 <= not w3942 and not w12270;
w12272 <= w7356 and not w12271;
w12273 <= not w12269 and w12272;
w12274 <= not w6599 and not w12269;
w12275 <= w12038 and w12247;
w12276 <= w12212 and not w12220;
w12277 <= w12002 and not w12276;
w12278 <= w12008 and not w12277;
w12279 <= not w12275 and not w12278;
w12280 <= pi0216 and not w12279;
w12281 <= not w12274 and not w12280;
w12282 <= w7357 and not w12271;
w12283 <= not w12281 and w12282;
w12284 <= pi0232 and not w12273;
w12285 <= not w12261 and w12284;
w12286 <= not w12283 and w12285;
w12287 <= pi0039 and not w12216;
w12288 <= not w12286 and w12287;
w12289 <= not pi0039 and not pi0232;
w12290 <= not w12069 and w12289;
w12291 <= not w12288 and not w12290;
w12292 <= not w12211 and w12291;
w12293 <= not pi0038 and not w12292;
w12294 <= not w12037 and not w12293;
w12295 <= w12031 and not w12032;
w12296 <= not w12294 and w12295;
w12297 <= not pi0184 and not pi0299;
w12298 <= not pi0163 and pi0299;
w12299 <= not w12297 and not w12298;
w12300 <= w5036 and w12299;
w12301 <= pi0087 and not w12300;
w12302 <= not w12000 and not w12301;
w12303 <= not w12029 and w12302;
w12304 <= not w12296 and w12303;
w12305 <= w12018 and not w12028;
w12306 <= not pi0158 and w12026;
w12307 <= w12008 and not w12100;
w12308 <= w3760 and not w12076;
w12309 <= not pi0146 and w12308;
w12310 <= w12001 and not w12048;
w12311 <= not pi0051 and not w12310;
w12312 <= w82 and not w12311;
w12313 <= not w12161 and not w12312;
w12314 <= pi0146 and w12313;
w12315 <= not pi0161 and not w12309;
w12316 <= not w12314 and w12315;
w12317 <= not w12307 and not w12316;
w12318 <= w7135 and not w12317;
w12319 <= pi0232 and not w12306;
w12320 <= not w12318 and w12319;
w12321 <= not pi0156 and w93;
w12322 <= not w12320 and w12321;
w12323 <= not pi0159 and w12026;
w12324 <= not pi0181 and w12024;
w12325 <= not pi0144 and not w12023;
w12326 <= not w12224 and w12325;
w12327 <= w6614 and w12220;
w12328 <= pi0142 and not w84;
w12329 <= not pi0142 and not w12238;
w12330 <= w12327 and not w12328;
w12331 <= not w12329 and w12330;
w12332 <= w12021 and not w12331;
w12333 <= pi0181 and not w12326;
w12334 <= not w12332 and w12333;
w12335 <= not pi0299 and not w12324;
w12336 <= not w12334 and w12335;
w12337 <= not w6599 and w12011;
w12338 <= w12038 and not w12222;
w12339 <= w3760 and w3943;
w12340 <= w12008 and not w12339;
w12341 <= w6599 and not w12338;
w12342 <= not w12340 and w12341;
w12343 <= w7357 and not w12337;
w12344 <= not w12342 and w12343;
w12345 <= w8041 and not w12323;
w12346 <= not w12344 and w12345;
w12347 <= not w12336 and w12346;
w12348 <= w3760 and not w12140;
w12349 <= not w12005 and w12348;
w12350 <= pi0161 and not w12349;
w12351 <= w3760 and not w12077;
w12352 <= not pi0146 and w12351;
w12353 <= w12039 and w12310;
w12354 <= w12064 and w12353;
w12355 <= w12057 and not w12354;
w12356 <= w82 and not w12355;
w12357 <= not w12161 and not w12356;
w12358 <= pi0146 and w12357;
w12359 <= not pi0161 and not w12352;
w12360 <= not w12358 and w12359;
w12361 <= not w12350 and not w12360;
w12362 <= w7135 and not w12361;
w12363 <= w12008 and not w12175;
w12364 <= not pi0161 and not w12199;
w12365 <= not w12363 and not w12364;
w12366 <= w7166 and not w12365;
w12367 <= pi0232 and not w12366;
w12368 <= not w12362 and w12367;
w12369 <= pi0156 and not w12368;
w12370 <= not pi0142 and w12351;
w12371 <= pi0142 and w12357;
w12372 <= not pi0144 and not w12370;
w12373 <= not w12371 and w12372;
w12374 <= not w12022 and w12348;
w12375 <= pi0144 and not w12374;
w12376 <= pi0180 and not w12373;
w12377 <= not w12375 and w12376;
w12378 <= w12021 and not w12175;
w12379 <= not pi0144 and not w12165;
w12380 <= not pi0180 and not w12379;
w12381 <= not w12378 and w12380;
w12382 <= pi0179 and not w12381;
w12383 <= not w12377 and w12382;
w12384 <= not pi0180 and w12024;
w12385 <= not pi0142 and w12308;
w12386 <= pi0142 and w12313;
w12387 <= not pi0144 and not w12385;
w12388 <= not w12386 and w12387;
w12389 <= w12021 and not w12100;
w12390 <= pi0180 and not w12388;
w12391 <= not w12389 and w12390;
w12392 <= not pi0179 and not w12384;
w12393 <= not w12391 and w12392;
w12394 <= not w12383 and not w12393;
w12395 <= not pi0299 and not w12394;
w12396 <= not pi0039 and not w12369;
w12397 <= not w12395 and w12396;
w12398 <= not pi0038 and not w12347;
w12399 <= not w12397 and w12398;
w12400 <= w12034 and not w12322;
w12401 <= not w12399 and w12400;
w12402 <= w98 and not w12032;
w12403 <= not w12401 and w12402;
w12404 <= w12000 and not w12301;
w12405 <= not w12305 and w12404;
w12406 <= not w12403 and w12405;
w12407 <= w4989 and not w12406;
w12408 <= not w12304 and w12407;
w12409 <= not w12017 and not w12408;
w12410 <= w4983 and w4990;
w12411 <= w4992 and w11970;
w12412 <= w11590 and not w12411;
w12413 <= w4992 and w11980;
w12414 <= w4988 and not w12413;
w12415 <= w4989 and not w12412;
w12416 <= not w12414 and w12415;
w12417 <= not w12410 and not w12416;
w12418 <= pi0110 and w7638;
w12419 <= not w8539 and w12418;
w12420 <= not w3837 and w12419;
w12421 <= not pi0039 and not w12420;
w12422 <= not pi0110 and w6856;
w12423 <= not w3807 and w3942;
w12424 <= w12422 and w12423;
w12425 <= pi0039 and not w12424;
w12426 <= not w4989 and not w12421;
w12427 <= not w12425 and w12426;
w12428 <= pi0110 and w11011;
w12429 <= not pi0039 and not w12428;
w12430 <= not w3770 and w5170;
w12431 <= w12422 and w12430;
w12432 <= pi0299 and w12424;
w12433 <= pi0039 and not w12431;
w12434 <= not w12432 and w12433;
w12435 <= not w12429 and not w12434;
w12436 <= not pi0038 and w134;
w12437 <= not w12435 and not w12436;
w12438 <= pi0090 and not w7950;
w12439 <= not pi0111 and not w3992;
w12440 <= not pi0036 and w372;
w12441 <= not w12439 and w12440;
w12442 <= w31 and not w12441;
w12443 <= not w356 and not w361;
w12444 <= not w12442 and w12443;
w12445 <= not pi0083 and not w12444;
w12446 <= w358 and not w12445;
w12447 <= not pi0071 and not w12446;
w12448 <= w4001 and not w12447;
w12449 <= not pi0081 and not w12448;
w12450 <= w9006 and not w12449;
w12451 <= not pi0090 and not w12450;
w12452 <= w270 and not w12451;
w12453 <= w6636 and not w12438;
w12454 <= w12452 and w12453;
w12455 <= pi0072 and w271;
w12456 <= w7950 and w12455;
w12457 <= not w12454 and not w12456;
w12458 <= w4042 and not w12457;
w12459 <= not pi0110 and not w12458;
w12460 <= w11011 and not w12459;
w12461 <= w460 and w12452;
w12462 <= not pi0072 and not w12461;
w12463 <= w4043 and not w11011;
w12464 <= not w12462 and w12463;
w12465 <= not pi0039 and not w12464;
w12466 <= not w12460 and w12465;
w12467 <= not w12434 and not w12466;
w12468 <= w12436 and not w12467;
w12469 <= w4989 and not w12437;
w12470 <= not w12468 and w12469;
w12471 <= not w12427 and not w12470;
w12472 <= not pi0125 and w11995;
w12473 <= pi0125 and pi0133;
w12474 <= not w11996 and not w12473;
w12475 <= not w12472 and not w12474;
w12476 <= w12002 and not w12475;
w12477 <= pi0172 and w12006;
w12478 <= not pi0152 and w12160;
w12479 <= not w12477 and not w12478;
w12480 <= pi0232 and not w12479;
w12481 <= not w12476 and not w12480;
w12482 <= not pi0087 and not w12481;
w12483 <= pi0087 and w5036;
w12484 <= pi0162 and w12483;
w12485 <= not w4989 and not w12484;
w12486 <= not w12482 and w12485;
w12487 <= pi0193 and w12006;
w12488 <= not pi0174 and w12160;
w12489 <= not pi0299 and not w12487;
w12490 <= not w12488 and w12489;
w12491 <= pi0299 and w12479;
w12492 <= pi0232 and not w12490;
w12493 <= not w12491 and w12492;
w12494 <= w12018 and not w12493;
w12495 <= pi0140 and not pi0299;
w12496 <= pi0162 and pi0299;
w12497 <= not w12495 and not w12496;
w12498 <= w5036 and not w12497;
w12499 <= pi0087 and not w12498;
w12500 <= pi0100 and w12493;
w12501 <= not pi0232 and not w12071;
w12502 <= not pi0039 and not w12501;
w12503 <= not pi0299 and not w5114;
w12504 <= pi0299 and not w5133;
w12505 <= not w12503 and not w12504;
w12506 <= w84 and w12505;
w12507 <= not pi0232 and not w12506;
w12508 <= pi0039 and not w12507;
w12509 <= not w5133 and w12479;
w12510 <= w84 and not w3760;
w12511 <= w3760 and not w12217;
w12512 <= not w12510 and not w12511;
w12513 <= not pi0152 and not w12512;
w12514 <= not w12240 and not w12510;
w12515 <= pi0152 and not w12514;
w12516 <= not w12513 and not w12515;
w12517 <= pi0051 and not pi0172;
w12518 <= not w12516 and not w12517;
w12519 <= not pi0216 and not w12518;
w12520 <= w3942 and w12519;
w12521 <= not w12509 and not w12520;
w12522 <= w7166 and not w12521;
w12523 <= not w3942 and not w12479;
w12524 <= w12212 and w12220;
w12525 <= not w12009 and not w12524;
w12526 <= not pi0152 and w12525;
w12527 <= w12220 and w12238;
w12528 <= not w12006 and not w12527;
w12529 <= pi0152 and w12528;
w12530 <= pi0172 and not w12526;
w12531 <= not w12529 and w12530;
w12532 <= not pi0152 and not w12222;
w12533 <= pi0152 and not w12339;
w12534 <= not pi0172 and not w12532;
w12535 <= not w12533 and w12534;
w12536 <= pi0216 and not w12531;
w12537 <= not w12535 and w12536;
w12538 <= w3942 and not w12537;
w12539 <= not w12519 and w12538;
w12540 <= w7135 and not w12523;
w12541 <= not w12539 and w12540;
w12542 <= not w5114 and not w12009;
w12543 <= w3760 and w12218;
w12544 <= not w12510 and not w12543;
w12545 <= not w12542 and not w12544;
w12546 <= not pi0174 and w12545;
w12547 <= w84 and w5114;
w12548 <= pi0174 and w12547;
w12549 <= not w12487 and not w12548;
w12550 <= not w12546 and w12549;
w12551 <= not pi0180 and not w12550;
w12552 <= w5114 and w12512;
w12553 <= pi0224 and not w12524;
w12554 <= w3968 and not w12553;
w12555 <= not w12009 and not w12554;
w12556 <= not w12552 and not w12555;
w12557 <= not pi0174 and w12556;
w12558 <= pi0224 and w12528;
w12559 <= w3968 and not w12558;
w12560 <= w5114 and w12514;
w12561 <= w12559 and not w12560;
w12562 <= not w12006 and not w12561;
w12563 <= pi0174 and not w12562;
w12564 <= pi0193 and not w12557;
w12565 <= not w12563 and w12564;
w12566 <= not w5114 and not w12327;
w12567 <= w84 and not w12566;
w12568 <= pi0174 and w12567;
w12569 <= pi0224 and not w12222;
w12570 <= not pi0224 and w12544;
w12571 <= w3968 and not w12569;
w12572 <= not w12570 and w12571;
w12573 <= not w12251 and not w12572;
w12574 <= not pi0174 and not w12573;
w12575 <= not pi0193 and not w12568;
w12576 <= not w12574 and w12575;
w12577 <= pi0180 and not w12576;
w12578 <= not w12565 and w12577;
w12579 <= not pi0299 and not w12551;
w12580 <= not w12578 and w12579;
w12581 <= not w12522 and not w12541;
w12582 <= not w12580 and w12581;
w12583 <= pi0232 and not w12582;
w12584 <= w12508 and not w12583;
w12585 <= not pi0038 and not w12502;
w12586 <= not w12584 and w12585;
w12587 <= pi0038 and not w12493;
w12588 <= not pi0100 and not w12587;
w12589 <= not pi0152 and w12084;
w12590 <= not pi0152 and w3760;
w12591 <= w12071 and not w12590;
w12592 <= not pi0197 and not w12589;
w12593 <= not w12591 and w12592;
w12594 <= not w3760 and w12071;
w12595 <= not w12082 and not w12594;
w12596 <= not w12106 and not w12595;
w12597 <= not pi0152 and pi0197;
w12598 <= not w12596 and w12597;
w12599 <= not w12593 and not w12598;
w12600 <= not w12477 and not w12599;
w12601 <= not w3760 and not w12071;
w12602 <= not w12096 and not w12601;
w12603 <= not pi0172 and w12602;
w12604 <= not w12006 and not w12100;
w12605 <= not w12071 and w12604;
w12606 <= pi0172 and not w12605;
w12607 <= pi0152 and pi0197;
w12608 <= not w12606 and w12607;
w12609 <= not w12603 and w12608;
w12610 <= not w12600 and not w12609;
w12611 <= w7329 and not w12610;
w12612 <= w12068 and w12105;
w12613 <= not w12601 and not w12612;
w12614 <= not pi0152 and w12613;
w12615 <= w12072 and not w12175;
w12616 <= pi0152 and not w12615;
w12617 <= pi0172 and not w12614;
w12618 <= not w12616 and w12617;
w12619 <= not w12172 and not w12601;
w12620 <= pi0152 and w12619;
w12621 <= not w12155 and not w12594;
w12622 <= not pi0152 and not w12621;
w12623 <= not pi0172 and not w12622;
w12624 <= not w12620 and w12623;
w12625 <= not pi0197 and not w12618;
w12626 <= not w12624 and w12625;
w12627 <= not w12148 and not w12601;
w12628 <= not pi0172 and w12627;
w12629 <= not w12141 and not w12601;
w12630 <= pi0172 and w12629;
w12631 <= pi0152 and not w12630;
w12632 <= not w12628 and w12631;
w12633 <= w3760 and w12069;
w12634 <= not w12595 and not w12633;
w12635 <= not pi0152 and not w12477;
w12636 <= not w12634 and w12635;
w12637 <= pi0197 and not w12636;
w12638 <= not w12632 and w12637;
w12639 <= w7323 and not w12626;
w12640 <= not w12638 and w12639;
w12641 <= not w12611 and not w12640;
w12642 <= pi0299 and not w12641;
w12643 <= not pi0145 and w12071;
w12644 <= pi0145 and w12602;
w12645 <= pi0174 and not w12643;
w12646 <= not w12644 and w12645;
w12647 <= not w12084 and not w12594;
w12648 <= not pi0145 and not w12647;
w12649 <= pi0145 and w12596;
w12650 <= not pi0174 and not w12648;
w12651 <= not w12649 and w12650;
w12652 <= not w12646 and not w12651;
w12653 <= not pi0193 and not w12652;
w12654 <= not pi0145 and w12100;
w12655 <= not w12604 and not w12654;
w12656 <= not w12071 and not w12655;
w12657 <= pi0174 and not w12656;
w12658 <= not w12006 and not w12049;
w12659 <= pi0145 and not w12658;
w12660 <= w12105 and not w12659;
w12661 <= not pi0174 and not w12660;
w12662 <= not w12601 and w12661;
w12663 <= pi0193 and not w12662;
w12664 <= not w12657 and w12663;
w12665 <= not w12653 and not w12664;
w12666 <= w7335 and not w12665;
w12667 <= pi0193 and w12613;
w12668 <= not pi0193 and not w12621;
w12669 <= not pi0145 and not w12667;
w12670 <= not w12668 and w12669;
w12671 <= pi0145 and not w12487;
w12672 <= not w12634 and w12671;
w12673 <= not pi0174 and not w12672;
w12674 <= not w12670 and w12673;
w12675 <= pi0145 and w12629;
w12676 <= not pi0145 and not w12615;
w12677 <= pi0193 and not w12676;
w12678 <= not w12675 and w12677;
w12679 <= not pi0145 and w12619;
w12680 <= pi0145 and w12627;
w12681 <= not pi0193 and not w12679;
w12682 <= not w12680 and w12681;
w12683 <= pi0174 and not w12678;
w12684 <= not w12682 and w12683;
w12685 <= w7339 and not w12674;
w12686 <= not w12684 and w12685;
w12687 <= not w12666 and not w12686;
w12688 <= not pi0038 and not w12687;
w12689 <= not w12642 and not w12688;
w12690 <= w6722 and not w12689;
w12691 <= not w12586 and w12588;
w12692 <= not w12690 and w12691;
w12693 <= w98 and not w12500;
w12694 <= not w12692 and w12693;
w12695 <= w12475 and not w12499;
w12696 <= not w12494 and w12695;
w12697 <= not w12694 and w12696;
w12698 <= w12019 and not w12493;
w12699 <= not w12036 and not w12588;
w12700 <= not w12078 and not w12175;
w12701 <= pi0145 and w12700;
w12702 <= w12099 and w12145;
w12703 <= not w12078 and not w12702;
w12704 <= not pi0145 and w12703;
w12705 <= not pi0174 and not w12701;
w12706 <= not w12704 and w12705;
w12707 <= not w12078 and not w12357;
w12708 <= not pi0145 and not w12076;
w12709 <= not w3760 and not w12076;
w12710 <= not w12009 and not w12709;
w12711 <= not w12066 and w12710;
w12712 <= not w12708 and w12711;
w12713 <= w82 and w12712;
w12714 <= pi0174 and not w12707;
w12715 <= not w12713 and w12714;
w12716 <= pi0193 and not w12715;
w12717 <= not w12706 and w12716;
w12718 <= pi0174 and not w12712;
w12719 <= not pi0051 and w12701;
w12720 <= not pi0145 and not w12078;
w12721 <= not w12348 and w12720;
w12722 <= not pi0174 and not w12719;
w12723 <= not w12721 and w12722;
w12724 <= not pi0193 and not w12718;
w12725 <= not w12723 and w12724;
w12726 <= w7335 and not w12717;
w12727 <= not w12725 and w12726;
w12728 <= pi0145 and not w12160;
w12729 <= not pi0174 and not w12654;
w12730 <= not pi0145 and pi0174;
w12731 <= not w12313 and w12730;
w12732 <= not w12728 and not w12731;
w12733 <= not w12729 and w12732;
w12734 <= pi0193 and not w12078;
w12735 <= not w12733 and w12734;
w12736 <= not w12006 and not w12078;
w12737 <= pi0145 and w12001;
w12738 <= not w12729 and not w12737;
w12739 <= w12736 and not w12738;
w12740 <= not w12078 and not w12308;
w12741 <= pi0174 and w12740;
w12742 <= not w12739 and not w12741;
w12743 <= not pi0193 and not w12742;
w12744 <= w7339 and not w12735;
w12745 <= not w12743 and w12744;
w12746 <= not w12727 and not w12745;
w12747 <= not pi0038 and not w12746;
w12748 <= not pi0172 and w12006;
w12749 <= not pi0172 and w12711;
w12750 <= not w12078 and not w12163;
w12751 <= pi0172 and w12750;
w12752 <= pi0152 and not w12749;
w12753 <= not w12751 and w12752;
w12754 <= not pi0152 and not w12700;
w12755 <= pi0197 and not w12748;
w12756 <= not w12753 and w12755;
w12757 <= not w12754 and w12756;
w12758 <= not pi0152 and not w12703;
w12759 <= pi0152 and not w12707;
w12760 <= pi0172 and not w12759;
w12761 <= not w12758 and w12760;
w12762 <= not pi0152 and w12348;
w12763 <= not w12077 and not w12590;
w12764 <= not pi0172 and not w12763;
w12765 <= not w12762 and w12764;
w12766 <= not w12761 and not w12765;
w12767 <= not pi0197 and not w12766;
w12768 <= pi0299 and w7329;
w12769 <= not w12757 and w12768;
w12770 <= not w12767 and w12769;
w12771 <= pi0152 and w12160;
w12772 <= not w12078 and not w12771;
w12773 <= pi0172 and not w12772;
w12774 <= not pi0172 and not w12478;
w12775 <= not w12079 and w12774;
w12776 <= pi0197 and not w12773;
w12777 <= not w12775 and w12776;
w12778 <= pi0152 and w12740;
w12779 <= not w12078 and not w12100;
w12780 <= not pi0152 and w12779;
w12781 <= not w12006 and w12780;
w12782 <= not pi0172 and not w12778;
w12783 <= not w12781 and w12782;
w12784 <= not w12078 and not w12313;
w12785 <= pi0152 and w12784;
w12786 <= pi0172 and not w12785;
w12787 <= not w12780 and w12786;
w12788 <= not pi0197 and not w12787;
w12789 <= not w12783 and w12788;
w12790 <= pi0299 and w7323;
w12791 <= not w12777 and w12790;
w12792 <= not w12789 and w12791;
w12793 <= not w12770 and not w12792;
w12794 <= not w12747 and w12793;
w12795 <= w6722 and not w12794;
w12796 <= not w12002 and w12479;
w12797 <= not w6599 and not w12796;
w12798 <= not w12217 and not w12590;
w12799 <= not pi0152 and w12240;
w12800 <= not w12798 and not w12799;
w12801 <= not pi0172 and not w12800;
w12802 <= not pi0152 and w12236;
w12803 <= pi0152 and w12230;
w12804 <= pi0172 and not w12803;
w12805 <= not w12802 and w12804;
w12806 <= w6599 and not w12801;
w12807 <= not w12805 and w12806;
w12808 <= w7166 and not w12807;
w12809 <= pi0152 and not w12477;
w12810 <= not w12277 and w12809;
w12811 <= w12247 and w12635;
w12812 <= w6599 and not w12810;
w12813 <= not w12811 and w12812;
w12814 <= w7135 and not w12813;
w12815 <= not w12808 and not w12814;
w12816 <= not w12797 and not w12815;
w12817 <= pi0180 and w12277;
w12818 <= w6614 and w12212;
w12819 <= w12002 and not w12818;
w12820 <= pi0174 and not w12819;
w12821 <= not w12817 and w12820;
w12822 <= w6614 and w12241;
w12823 <= not w3760 and not w12001;
w12824 <= not w6614 and not w12823;
w12825 <= not pi0051 and w12824;
w12826 <= not w12822 and not w12825;
w12827 <= pi0180 and w12246;
w12828 <= not pi0174 and not w12827;
w12829 <= w12826 and w12828;
w12830 <= not pi0193 and not w12821;
w12831 <= not w12829 and w12830;
w12832 <= not w12229 and w12824;
w12833 <= w6614 and w12236;
w12834 <= not w12832 and not w12833;
w12835 <= not pi0174 and not w12834;
w12836 <= not w12006 and not w12819;
w12837 <= pi0174 and not w12836;
w12838 <= not pi0180 and not w12837;
w12839 <= not w12835 and w12838;
w12840 <= w6614 and not w12235;
w12841 <= not w8166 and w12840;
w12842 <= not w12832 and not w12841;
w12843 <= not pi0174 and not w12842;
w12844 <= not pi0051 and not w12277;
w12845 <= w3760 and not w12844;
w12846 <= not w12819 and not w12845;
w12847 <= pi0174 and not w12846;
w12848 <= pi0180 and not w12847;
w12849 <= not w12843 and w12848;
w12850 <= pi0193 and not w12849;
w12851 <= not w12839 and w12850;
w12852 <= not pi0299 and not w12831;
w12853 <= not w12851 and w12852;
w12854 <= not w12816 and not w12853;
w12855 <= pi0232 and not w12854;
w12856 <= not pi0299 and not w12819;
w12857 <= w6599 and w12212;
w12858 <= w12002 and not w12857;
w12859 <= pi0299 and not w12858;
w12860 <= not w12856 and not w12859;
w12861 <= not pi0232 and not w12860;
w12862 <= pi0039 and not w12861;
w12863 <= not w12855 and w12862;
w12864 <= not pi0232 and not w12077;
w12865 <= not pi0039 and not w12864;
w12866 <= not pi0038 and not w12865;
w12867 <= not w12863 and w12866;
w12868 <= not w12699 and not w12867;
w12869 <= not w12795 and w12868;
w12870 <= w12031 and not w12500;
w12871 <= not w12869 and w12870;
w12872 <= not w12475 and not w12499;
w12873 <= not w12698 and w12872;
w12874 <= not w12871 and w12873;
w12875 <= w4989 and not w12874;
w12876 <= not w12697 and w12875;
w12877 <= not w12486 and not w12876;
w12878 <= pi0175 and w12006;
w12879 <= not pi0189 and w12160;
w12880 <= not pi0299 and not w12878;
w12881 <= not w12879 and w12880;
w12882 <= not pi0051 and not w12160;
w12883 <= not w7862 and not w12001;
w12884 <= not pi0051 and not w12883;
w12885 <= pi0153 and w12006;
w12886 <= not w12884 and not w12885;
w12887 <= not w12882 and not w12886;
w12888 <= pi0299 and not w12887;
w12889 <= pi0232 and not w12881;
w12890 <= not w12888 and w12889;
w12891 <= not w171 and w12890;
w12892 <= not pi0126 and w11998;
w12893 <= pi0126 and not w11998;
w12894 <= not w12892 and not w12893;
w12895 <= not w11994 and not w12894;
w12896 <= not w171 and w12002;
w12897 <= not w12895 and w12896;
w12898 <= pi0182 and w12277;
w12899 <= pi0189 and not w12819;
w12900 <= not w12898 and w12899;
w12901 <= pi0182 and w12246;
w12902 <= not pi0189 and not w12901;
w12903 <= w12826 and w12902;
w12904 <= not w12900 and not w12903;
w12905 <= w9328 and not w12904;
w12906 <= not pi0189 and not w12834;
w12907 <= pi0189 and not w12836;
w12908 <= not pi0182 and not w12907;
w12909 <= not w12906 and w12908;
w12910 <= not pi0189 and not w12842;
w12911 <= pi0189 and not w12846;
w12912 <= pi0182 and not w12911;
w12913 <= not w12910 and w12912;
w12914 <= not w12909 and not w12913;
w12915 <= w9396 and not w12914;
w12916 <= not w6599 and not w12886;
w12917 <= not pi0166 and w12247;
w12918 <= pi0166 and not w12277;
w12919 <= not w12917 and not w12918;
w12920 <= pi0160 and not w12885;
w12921 <= not w12919 and w12920;
w12922 <= not w7862 and not w12217;
w12923 <= not pi0166 and w12240;
w12924 <= not w12922 and not w12923;
w12925 <= not pi0153 and not w12924;
w12926 <= not pi0166 and w12236;
w12927 <= pi0166 and w12230;
w12928 <= pi0153 and not w12927;
w12929 <= not w12926 and w12928;
w12930 <= not w12925 and not w12929;
w12931 <= not pi0160 and not w12930;
w12932 <= w6599 and not w12921;
w12933 <= not w12931 and w12932;
w12934 <= pi0299 and not w12916;
w12935 <= not w12933 and w12934;
w12936 <= not w12905 and not w12915;
w12937 <= not w12935 and w12936;
w12938 <= pi0232 and not w12937;
w12939 <= w12862 and not w12938;
w12940 <= not pi0189 and w12736;
w12941 <= pi0178 and not w12940;
w12942 <= pi0189 and w12079;
w12943 <= w12941 and not w12942;
w12944 <= pi0189 and w12711;
w12945 <= not w12175 and w12940;
w12946 <= not pi0178 and not w12944;
w12947 <= not w12945 and w12946;
w12948 <= pi0181 and not w12943;
w12949 <= not w12947 and w12948;
w12950 <= pi0189 and w12740;
w12951 <= not pi0189 and w12779;
w12952 <= pi0178 and not w12951;
w12953 <= not w12941 and not w12952;
w12954 <= not w12950 and not w12953;
w12955 <= not w7858 and not w12077;
w12956 <= not pi0189 and w12348;
w12957 <= not w12955 and not w12956;
w12958 <= not pi0178 and not w12957;
w12959 <= not pi0181 and not w12954;
w12960 <= not w12958 and w12959;
w12961 <= w9328 and not w12949;
w12962 <= not w12960 and w12961;
w12963 <= not pi0189 and not w12175;
w12964 <= pi0189 and not w12163;
w12965 <= not pi0178 and not w12964;
w12966 <= not w12963 and w12965;
w12967 <= pi0178 and w9389;
w12968 <= w12159 and w12967;
w12969 <= pi0181 and not w12968;
w12970 <= not w12078 and w12969;
w12971 <= not w12966 and w12970;
w12972 <= pi0189 and w12784;
w12973 <= w12952 and not w12972;
w12974 <= not pi0189 and w12703;
w12975 <= pi0189 and w12707;
w12976 <= not pi0178 and not w12975;
w12977 <= not w12974 and w12976;
w12978 <= not pi0181 and not w12973;
w12979 <= not w12977 and w12978;
w12980 <= w9396 and not w12971;
w12981 <= not w12979 and w12980;
w12982 <= pi0166 and w12160;
w12983 <= not w12078 and not w12982;
w12984 <= pi0153 and not w12983;
w12985 <= not pi0153 and not w12887;
w12986 <= not w12079 and w12985;
w12987 <= pi0157 and not w12984;
w12988 <= not w12986 and w12987;
w12989 <= pi0153 and pi0166;
w12990 <= not w12750 and w12989;
w12991 <= not pi0166 and not w12700;
w12992 <= pi0166 and not w12711;
w12993 <= pi0051 and w7862;
w12994 <= not w12992 and not w12993;
w12995 <= not pi0153 and not w12994;
w12996 <= not pi0157 and not w12990;
w12997 <= not w12995 and w12996;
w12998 <= not w12991 and w12997;
w12999 <= w7357 and not w12988;
w13000 <= not w12998 and w12999;
w13001 <= not pi0166 and not w12779;
w13002 <= pi0166 and not w12740;
w13003 <= not w12993 and not w13002;
w13004 <= not pi0153 and not w13003;
w13005 <= not w12784 and w12989;
w13006 <= pi0157 and not w13005;
w13007 <= not w13001 and w13006;
w13008 <= not w13004 and w13007;
w13009 <= not pi0166 and not w12703;
w13010 <= pi0166 and not w12707;
w13011 <= pi0153 and not w13010;
w13012 <= not w13009 and w13011;
w13013 <= not pi0166 and w12348;
w13014 <= not w7862 and not w12077;
w13015 <= not pi0153 and not w13014;
w13016 <= not w13013 and w13015;
w13017 <= not w13012 and not w13016;
w13018 <= not pi0157 and not w13017;
w13019 <= w7356 and not w13008;
w13020 <= not w13018 and w13019;
w13021 <= not w12981 and not w13000;
w13022 <= not w12962 and w13021;
w13023 <= not w13020 and w13022;
w13024 <= pi0232 and not w13023;
w13025 <= w12865 and not w13024;
w13026 <= not w12895 and not w12939;
w13027 <= not w13025 and w13026;
w13028 <= not pi0189 and w12545;
w13029 <= pi0189 and w12547;
w13030 <= not pi0182 and not w13029;
w13031 <= not w13028 and w13030;
w13032 <= not w12006 and w13031;
w13033 <= not pi0189 and w12556;
w13034 <= pi0189 and not w12562;
w13035 <= pi0182 and not w13033;
w13036 <= not w13034 and w13035;
w13037 <= not w13032 and not w13036;
w13038 <= w9396 and not w13037;
w13039 <= not pi0189 and not w12573;
w13040 <= pi0189 and w12567;
w13041 <= pi0182 and not w13040;
w13042 <= not w13039 and w13041;
w13043 <= not w13031 and not w13042;
w13044 <= w9328 and not w13043;
w13045 <= not pi0160 and pi0216;
w13046 <= w3942 and not w13045;
w13047 <= w12887 and not w13046;
w13048 <= not pi0166 and w12222;
w13049 <= pi0166 and w12339;
w13050 <= not pi0153 and not w13048;
w13051 <= not w13049 and w13050;
w13052 <= pi0166 and not w12528;
w13053 <= not pi0166 and not w12525;
w13054 <= pi0153 and not w13053;
w13055 <= not w13052 and w13054;
w13056 <= pi0160 and not w13051;
w13057 <= not w13055 and w13056;
w13058 <= pi0216 and not w13057;
w13059 <= not pi0166 and not w12512;
w13060 <= pi0166 and not w12514;
w13061 <= not w13059 and not w13060;
w13062 <= pi0051 and not pi0153;
w13063 <= not w13061 and not w13062;
w13064 <= not pi0216 and not w13063;
w13065 <= w3942 and not w13058;
w13066 <= not w13064 and w13065;
w13067 <= pi0299 and not w13047;
w13068 <= not w13066 and w13067;
w13069 <= not w13038 and not w13044;
w13070 <= not w13068 and w13069;
w13071 <= pi0232 and not w13070;
w13072 <= w12508 and not w13071;
w13073 <= not pi0153 and w12627;
w13074 <= pi0153 and w12629;
w13075 <= pi0157 and not w13074;
w13076 <= not w13073 and w13075;
w13077 <= not pi0153 and w12602;
w13078 <= pi0153 and not w12605;
w13079 <= not pi0157 and not w13078;
w13080 <= not w13077 and w13079;
w13081 <= not w13076 and not w13080;
w13082 <= pi0166 and not w13081;
w13083 <= pi0157 and w12634;
w13084 <= not pi0157 and w12596;
w13085 <= not pi0166 and not w12885;
w13086 <= not w13083 and w13085;
w13087 <= not w13084 and w13086;
w13088 <= not w13082 and not w13087;
w13089 <= w7357 and not w13088;
w13090 <= not pi0166 and w12613;
w13091 <= pi0166 and not w12615;
w13092 <= pi0153 and not w13090;
w13093 <= not w13091 and w13092;
w13094 <= pi0166 and w12619;
w13095 <= not pi0166 and not w12621;
w13096 <= not pi0153 and not w13095;
w13097 <= not w13094 and w13096;
w13098 <= not w13093 and not w13097;
w13099 <= pi0157 and not w13098;
w13100 <= pi0166 and w12071;
w13101 <= not pi0166 and not w12647;
w13102 <= not pi0157 and not w12885;
w13103 <= not w13100 and w13102;
w13104 <= not w13101 and w13103;
w13105 <= not w13099 and not w13104;
w13106 <= w7356 and not w13105;
w13107 <= not pi0189 and not w12647;
w13108 <= pi0189 and w12071;
w13109 <= not pi0178 and not w13108;
w13110 <= not w12006 and w13109;
w13111 <= not w13107 and w13110;
w13112 <= not pi0181 and not w13111;
w13113 <= pi0189 and not w12615;
w13114 <= not pi0189 and w12613;
w13115 <= pi0178 and not w13114;
w13116 <= not w13113 and w13115;
w13117 <= w13112 and not w13116;
w13118 <= pi0189 and w12605;
w13119 <= not pi0189 and not w12596;
w13120 <= not w12006 and w13119;
w13121 <= not w13118 and not w13120;
w13122 <= not pi0178 and not w13121;
w13123 <= not pi0189 and w12634;
w13124 <= w12629 and not w12940;
w13125 <= pi0178 and not w13123;
w13126 <= not w13124 and w13125;
w13127 <= pi0181 and not w13122;
w13128 <= not w13126 and w13127;
w13129 <= w9396 and not w13117;
w13130 <= not w13128 and w13129;
w13131 <= w12647 and w13109;
w13132 <= not pi0189 and not w12621;
w13133 <= pi0189 and w12619;
w13134 <= pi0178 and not w13132;
w13135 <= not w13133 and w13134;
w13136 <= w13112 and not w13131;
w13137 <= not w13135 and w13136;
w13138 <= pi0189 and w12627;
w13139 <= not w13123 and not w13138;
w13140 <= pi0178 and not w13139;
w13141 <= pi0189 and not w12602;
w13142 <= not pi0178 and not w13119;
w13143 <= not w13141 and w13142;
w13144 <= not w13140 and not w13143;
w13145 <= pi0181 and not w13144;
w13146 <= w9328 and not w13137;
w13147 <= not w13145 and w13146;
w13148 <= not w13106 and not w13130;
w13149 <= not w13089 and w13148;
w13150 <= not w13147 and w13149;
w13151 <= pi0232 and not w13150;
w13152 <= w12502 and not w13151;
w13153 <= w12895 and not w13072;
w13154 <= not w13152 and w13153;
w13155 <= w171 and not w13027;
w13156 <= not w13154 and w13155;
w13157 <= w98 and not w12897;
w13158 <= not w12891 and w13157;
w13159 <= not w13156 and w13158;
w13160 <= w12018 and not w12890;
w13161 <= not pi0150 and pi0299;
w13162 <= not pi0185 and not pi0299;
w13163 <= not w13161 and not w13162;
w13164 <= w5036 and w13163;
w13165 <= pi0087 and not w13164;
w13166 <= not w13160 and not w13165;
w13167 <= w12003 and not w12895;
w13168 <= not w13166 and not w13167;
w13169 <= w4989 and not w13168;
w13170 <= not w13159 and w13169;
w13171 <= pi0232 and not w12882;
w13172 <= w12895 and not w13171;
w13173 <= not pi0232 and not w12002;
w13174 <= not w12886 and not w13173;
w13175 <= not w13172 and w13174;
w13176 <= not pi0087 and not w13175;
w13177 <= pi0087 and not w11248;
w13178 <= not w4989 and not w13177;
w13179 <= not w13176 and w13178;
w13180 <= not w13170 and not w13179;
w13181 <= w100 and w6450;
w13182 <= w92 and w13181;
w13183 <= not w891 and not w13182;
w13184 <= not w92 and not w13181;
w13185 <= pi0129 and w4864;
w13186 <= w3886 and w13185;
w13187 <= pi0074 and not w13186;
w13188 <= pi0054 and w174;
w13189 <= w6450 and w13188;
w13190 <= pi0092 and not pi0129;
w13191 <= pi0075 and w13185;
w13192 <= not w188 and not w6528;
w13193 <= w6450 and not w13192;
w13194 <= not w131 and not w13193;
w13195 <= pi0129 and w3698;
w13196 <= pi0038 and not w13195;
w13197 <= pi0039 and w6450;
w13198 <= not w292 and not w669;
w13199 <= w351 and not w422;
w13200 <= w25 and not w13199;
w13201 <= w436 and not w13200;
w13202 <= w348 and not w13201;
w13203 <= w440 and not w13202;
w13204 <= w282 and not w13203;
w13205 <= not w285 and not w13204;
w13206 <= not pi0086 and not w13205;
w13207 <= w346 and not w13206;
w13208 <= not pi0097 and not w13207;
w13209 <= not w339 and not w13208;
w13210 <= not pi0108 and not w13209;
w13211 <= w338 and not w13210;
w13212 <= w452 and not w13211;
w13213 <= not w329 and not w13212;
w13214 <= w328 and not w13213;
w13215 <= w327 and not w13214;
w13216 <= w3841 and w13215;
w13217 <= pi0250 and not w5037;
w13218 <= w7640 and w13217;
w13219 <= w344 and not w13207;
w13220 <= not w339 and not w13219;
w13221 <= not pi0108 and not w13220;
w13222 <= w338 and not w13221;
w13223 <= w452 and not w13222;
w13224 <= not w329 and not w13223;
w13225 <= w328 and not w13224;
w13226 <= w327 and not w13225;
w13227 <= not w3841 and w13226;
w13228 <= not w13216 and w13218;
w13229 <= not w13227 and w13228;
w13230 <= not pi0127 and w13215;
w13231 <= pi0127 and w13226;
w13232 <= not w13218 and not w13230;
w13233 <= not w13231 and w13232;
w13234 <= not w13229 and not w13233;
w13235 <= w320 and not w13234;
w13236 <= w671 and not w13235;
w13237 <= w67 and not w13236;
w13238 <= w13198 and not w13237;
w13239 <= not pi0070 and not w13238;
w13240 <= not w662 and not w13239;
w13241 <= not pi0051 and not w13240;
w13242 <= w311 and not w13241;
w13243 <= w731 and not w13242;
w13244 <= not w308 and not w13243;
w13245 <= w73 and not w13244;
w13246 <= w976 and not w13245;
w13247 <= not pi0095 and not w13246;
w13248 <= not pi0039 and pi0129;
w13249 <= not w304 and w13248;
w13250 <= not w13247 and w13249;
w13251 <= not pi0038 and not w13197;
w13252 <= not w13250 and w13251;
w13253 <= not w13196 and not w13252;
w13254 <= w131 and not w13253;
w13255 <= not pi0075 and not w13194;
w13256 <= not w13254 and w13255;
w13257 <= not pi0092 and not w13191;
w13258 <= not w13256 and w13257;
w13259 <= w11217 and not w13190;
w13260 <= not w13258 and w13259;
w13261 <= not pi0074 and not w13189;
w13262 <= not w13260 and w13261;
w13263 <= not pi0055 and not w13187;
w13264 <= not w13262 and w13263;
w13265 <= pi0055 and w133;
w13266 <= w13185 and w13265;
w13267 <= not w13264 and not w13266;
w13268 <= not pi0056 and not w13267;
w13269 <= not w8873 and not w8881;
w13270 <= not w13268 and w13269;
w13271 <= not w13184 and not w13270;
w13272 <= w891 and not w13271;
w13273 <= not w3683 and not w13183;
w13274 <= not w13272 and w13273;
w13275 <= not w3693 and not w4910;
w13276 <= w6451 and w7954;
w13277 <= w3841 and w13276;
w13278 <= not pi0129 and not w13276;
w13279 <= w6530 and not w13277;
w13280 <= not w13278 and w13279;
w13281 <= w84 and w13280;
w13282 <= not pi0038 and not w981;
w13283 <= w3700 and not w13282;
w13284 <= not w3843 and w3849;
w13285 <= not pi0087 and not w13284;
w13286 <= not w13283 and w13285;
w13287 <= w3696 and not w13286;
w13288 <= w3697 and not w13281;
w13289 <= not w13287 and w13288;
w13290 <= not w4868 and not w4904;
w13291 <= not w13289 and w13290;
w13292 <= w6442 and not w13291;
w13293 <= w13275 and not w13292;
w13294 <= not pi0056 and not w13293;
w13295 <= not w3690 and not w13294;
w13296 <= not pi0062 and not w13295;
w13297 <= not w3862 and not w13296;
w13298 <= w891 and not w13297;
w13299 <= w3686 and not w13298;
w13300 <= pi0087 and not w7310;
w13301 <= w5036 and not w6585;
w13302 <= w12159 and not w13301;
w13303 <= not w12882 and not w13302;
w13304 <= w12018 and not w13303;
w13305 <= not w13300 and not w13304;
w13306 <= not w12003 and not w13305;
w13307 <= not pi0132 and w12892;
w13308 <= pi0130 and not w13307;
w13309 <= not pi0130 and w13307;
w13310 <= not w13308 and not w13309;
w13311 <= not w11992 and not w13310;
w13312 <= pi0100 and w13303;
w13313 <= w98 and not w13312;
w13314 <= not w8545 and w13302;
w13315 <= not pi0051 and not w12860;
w13316 <= not pi0232 and not w13315;
w13317 <= w8545 and not w13316;
w13318 <= not pi0191 and not pi0299;
w13319 <= not pi0051 and not w12819;
w13320 <= pi0140 and w12845;
w13321 <= w13319 and not w13320;
w13322 <= w13318 and not w13321;
w13323 <= not pi0051 and w12826;
w13324 <= pi0140 and w12220;
w13325 <= w13323 and not w13324;
w13326 <= w6583 and not w13325;
w13327 <= pi0169 and w3760;
w13328 <= not w6599 and w12159;
w13329 <= not w13327 and w13328;
w13330 <= pi0162 and w6599;
w13331 <= not pi0051 and not w12241;
w13332 <= not w12220 and w13331;
w13333 <= pi0169 and not w13332;
w13334 <= not pi0169 and not w12844;
w13335 <= w13330 and not w13334;
w13336 <= not w13333 and w13335;
w13337 <= not w84 and w13327;
w13338 <= not w12218 and not w13327;
w13339 <= not pi0162 and w6599;
w13340 <= not w13338 and w13339;
w13341 <= not w13337 and w13340;
w13342 <= pi0299 and not w13329;
w13343 <= not w13341 and w13342;
w13344 <= not w13336 and w13343;
w13345 <= not w13322 and not w13326;
w13346 <= not w13344 and w13345;
w13347 <= pi0232 and not w13346;
w13348 <= w13317 and not w13347;
w13349 <= not pi0100 and not w13314;
w13350 <= not w13348 and w13349;
w13351 <= not w12030 and w13313;
w13352 <= not w13350 and w13351;
w13353 <= not w13306 and not w13311;
w13354 <= not w13352 and w13353;
w13355 <= not w12239 and not w13327;
w13356 <= pi0169 and w12511;
w13357 <= not w13355 and not w13356;
w13358 <= not pi0216 and not w13357;
w13359 <= not w12229 and w12525;
w13360 <= pi0169 and w13359;
w13361 <= not pi0051 and not w12527;
w13362 <= not pi0169 and w13361;
w13363 <= pi0162 and pi0216;
w13364 <= not w13360 and w13363;
w13365 <= not w13362 and w13364;
w13366 <= not w13358 and not w13365;
w13367 <= w3942 and not w13366;
w13368 <= pi0169 and w12160;
w13369 <= not pi0051 and not w13368;
w13370 <= not w5133 and not w13330;
w13371 <= not w13369 and w13370;
w13372 <= not w13367 and not w13371;
w13373 <= pi0299 and not w13372;
w13374 <= w5114 and w12238;
w13375 <= not pi0051 and not w13374;
w13376 <= not pi0140 and w13375;
w13377 <= w12238 and w12559;
w13378 <= not pi0051 and not w13377;
w13379 <= pi0140 and w13378;
w13380 <= w13318 and not w13376;
w13381 <= not w13379 and w13380;
w13382 <= not w3760 and not w12239;
w13383 <= not w12511 and not w13382;
w13384 <= w5114 and not w13383;
w13385 <= not w5114 and not w12882;
w13386 <= not w13384 and not w13385;
w13387 <= not pi0140 and w13386;
w13388 <= pi0224 and not w13359;
w13389 <= not pi0224 and not w13383;
w13390 <= not w13388 and not w13389;
w13391 <= w3968 and not w13390;
w13392 <= not w3968 and not w12882;
w13393 <= not w13391 and not w13392;
w13394 <= pi0140 and w13393;
w13395 <= w6583 and not w13387;
w13396 <= not w13394 and w13395;
w13397 <= not w13373 and not w13381;
w13398 <= not w13396 and w13397;
w13399 <= pi0232 and not w13398;
w13400 <= w12238 and w12505;
w13401 <= not pi0051 and not w13400;
w13402 <= not pi0232 and not w13401;
w13403 <= pi0039 and not w13402;
w13404 <= not w13399 and w13403;
w13405 <= not pi0232 and not w12141;
w13406 <= not pi0039 and not w13405;
w13407 <= not w3760 and w12141;
w13408 <= not w12633 and not w13407;
w13409 <= not w6585 and not w13408;
w13410 <= w6585 and w12141;
w13411 <= pi0232 and not w13410;
w13412 <= not w13409 and w13411;
w13413 <= w13406 and not w13412;
w13414 <= not w13404 and not w13413;
w13415 <= not pi0038 and not w13414;
w13416 <= pi0038 and not w13303;
w13417 <= not pi0100 and not w13416;
w13418 <= not w13415 and w13417;
w13419 <= w13313 and not w13418;
w13420 <= w13305 and w13311;
w13421 <= not w13419 and w13420;
w13422 <= not w13354 and not w13421;
w13423 <= w4989 and not w13422;
w13424 <= pi0087 and not w7268;
w13425 <= pi0169 and w5036;
w13426 <= not pi0087 and w12159;
w13427 <= not w13425 and w13426;
w13428 <= not pi0051 and not pi0087;
w13429 <= not w13368 and w13428;
w13430 <= w13311 and w13429;
w13431 <= not w4989 and not w13424;
w13432 <= not w13427 and w13431;
w13433 <= not w13430 and w13432;
w13434 <= not w13423 and not w13433;
w13435 <= not pi0100 and not w11572;
w13436 <= not pi0087 and not w4897;
w13437 <= not w13435 and w13436;
w13438 <= not pi0075 and not w13437;
w13439 <= not w4865 and not w13438;
w13440 <= not pi0092 and not w13439;
w13441 <= w6443 and w11217;
w13442 <= not w13440 and w13441;
w13443 <= pi0164 and w12483;
w13444 <= pi0051 and not pi0151;
w13445 <= not w11315 and not w12006;
w13446 <= not w13444 and not w13445;
w13447 <= w12009 and w13446;
w13448 <= pi0232 and w13447;
w13449 <= pi0132 and not w12892;
w13450 <= not w13307 and not w13449;
w13451 <= not w11993 and not w13450;
w13452 <= w12002 and not w13451;
w13453 <= not w13448 and not w13452;
w13454 <= not pi0087 and not w13453;
w13455 <= not w4989 and not w13443;
w13456 <= not w13454 and w13455;
w13457 <= pi0173 and w12006;
w13458 <= pi0190 and w12160;
w13459 <= not pi0299 and not w13457;
w13460 <= not w13458 and w13459;
w13461 <= pi0299 and not w13447;
w13462 <= pi0232 and not w13460;
w13463 <= not w13461 and w13462;
w13464 <= w12018 and not w13463;
w13465 <= pi0087 and not w6593;
w13466 <= not w171 and w13463;
w13467 <= not w11315 and w12171;
w13468 <= pi0168 and w12155;
w13469 <= not pi0151 and not w13468;
w13470 <= not w13467 and w13469;
w13471 <= not w3760 and not w12171;
w13472 <= pi0168 and not w12612;
w13473 <= not w13471 and w13472;
w13474 <= not w3760 and w12171;
w13475 <= w12176 and not w13474;
w13476 <= not pi0168 and not w13475;
w13477 <= pi0151 and not w13473;
w13478 <= not w13476 and w13477;
w13479 <= not pi0160 and not w13470;
w13480 <= not w13478 and w13479;
w13481 <= pi0151 and w12141;
w13482 <= not pi0151 and not w12147;
w13483 <= not pi0168 and not w13481;
w13484 <= not w13482 and w13483;
w13485 <= pi0168 and not w13444;
w13486 <= not w12069 and w13485;
w13487 <= w3760 and not w13486;
w13488 <= not w13484 and w13487;
w13489 <= pi0160 and not w13471;
w13490 <= not w13488 and w13489;
w13491 <= pi0299 and not w13480;
w13492 <= not w13490 and w13491;
w13493 <= pi0190 and not pi0299;
w13494 <= pi0051 and not pi0173;
w13495 <= pi0182 and w12049;
w13496 <= w12068 and not w13495;
w13497 <= w3760 and not w13494;
w13498 <= not w13496 and w13497;
w13499 <= w13493 and not w13498;
w13500 <= not w13474 and w13499;
w13501 <= not pi0190 and not pi0299;
w13502 <= not pi0182 and w12171;
w13503 <= pi0182 and not w13471;
w13504 <= not w12148 and w13503;
w13505 <= not pi0173 and not w13502;
w13506 <= not w13504 and w13505;
w13507 <= not pi0182 and not w13475;
w13508 <= not w12142 and not w13474;
w13509 <= pi0182 and not w13508;
w13510 <= pi0173 and not w13507;
w13511 <= not w13509 and w13510;
w13512 <= not w13506 and not w13511;
w13513 <= w13501 and not w13512;
w13514 <= pi0232 and not w13500;
w13515 <= not w13492 and w13514;
w13516 <= not w13513 and w13515;
w13517 <= not pi0232 and w12171;
w13518 <= not w13516 and not w13517;
w13519 <= not pi0039 and not w13518;
w13520 <= not pi0183 and w12542;
w13521 <= pi0183 and not w12573;
w13522 <= not pi0183 and not w12544;
w13523 <= not pi0173 and not w13522;
w13524 <= not w13521 and w13523;
w13525 <= not pi0183 and not w12552;
w13526 <= pi0173 and not w12556;
w13527 <= not w13525 and w13526;
w13528 <= not w13520 and not w13527;
w13529 <= not w13524 and w13528;
w13530 <= w13493 and not w13529;
w13531 <= not pi0183 and not w5114;
w13532 <= not pi0173 and not w13531;
w13533 <= w12567 and w13532;
w13534 <= pi0183 and w12562;
w13535 <= not pi0183 and not w12006;
w13536 <= not w12547 and w13535;
w13537 <= pi0173 and not w13536;
w13538 <= not w13534 and w13537;
w13539 <= w13501 and not w13533;
w13540 <= not w13538 and w13539;
w13541 <= not pi0149 and pi0216;
w13542 <= w3942 and not w13541;
w13543 <= w13447 and not w13542;
w13544 <= not pi0168 and w12339;
w13545 <= pi0168 and w12222;
w13546 <= not pi0151 and not w13545;
w13547 <= not w13544 and w13546;
w13548 <= not pi0168 and not w12528;
w13549 <= pi0168 and not w12525;
w13550 <= pi0151 and not w13549;
w13551 <= not w13548 and w13550;
w13552 <= pi0149 and not w13547;
w13553 <= not w13551 and w13552;
w13554 <= pi0216 and not w13553;
w13555 <= pi0168 and not w12512;
w13556 <= not pi0168 and not w12514;
w13557 <= not w13555 and not w13556;
w13558 <= not w13444 and not w13557;
w13559 <= not pi0216 and not w13558;
w13560 <= w3942 and not w13554;
w13561 <= not w13559 and w13560;
w13562 <= pi0299 and not w13543;
w13563 <= not w13561 and w13562;
w13564 <= not w13530 and not w13540;
w13565 <= not w13563 and w13564;
w13566 <= pi0232 and not w13565;
w13567 <= w12508 and not w13566;
w13568 <= not w13519 and not w13567;
w13569 <= w171 and not w13568;
w13570 <= w98 and not w13466;
w13571 <= not w13569 and w13570;
w13572 <= w13451 and not w13465;
w13573 <= not w13464 and w13572;
w13574 <= not w13571 and w13573;
w13575 <= w12019 and not w13463;
w13576 <= not w12002 and w13461;
w13577 <= not w10693 and not w13576;
w13578 <= not pi0168 and not w12230;
w13579 <= pi0168 and not w12236;
w13580 <= pi0151 and not w13578;
w13581 <= not w13579 and w13580;
w13582 <= pi0168 and w12240;
w13583 <= not w11315 and not w12217;
w13584 <= not pi0151 and not w13583;
w13585 <= not w13582 and w13584;
w13586 <= not pi0149 and not w13585;
w13587 <= not w13581 and w13586;
w13588 <= not w12277 and not w13446;
w13589 <= not pi0168 and not w13588;
w13590 <= not w12528 and not w13444;
w13591 <= not w12241 and not w13590;
w13592 <= pi0168 and not w13591;
w13593 <= pi0149 and not w13589;
w13594 <= not w13592 and w13593;
w13595 <= w6599 and not w13587;
w13596 <= not w13594 and w13595;
w13597 <= not w13577 and not w13596;
w13598 <= not pi0183 and not w12834;
w13599 <= pi0183 and not w12842;
w13600 <= pi0173 and not w13599;
w13601 <= not w13598 and w13600;
w13602 <= pi0183 and w12246;
w13603 <= not pi0173 and not w13602;
w13604 <= w12826 and w13603;
w13605 <= not w13601 and not w13604;
w13606 <= w13493 and not w13605;
w13607 <= pi0183 and w12277;
w13608 <= not w13457 and w13501;
w13609 <= not w12819 and w13608;
w13610 <= not w13607 and w13609;
w13611 <= not w13597 and not w13610;
w13612 <= not w13606 and w13611;
w13613 <= pi0232 and not w13612;
w13614 <= not w12861 and not w13613;
w13615 <= pi0039 and not w13614;
w13616 <= not pi0232 and w12076;
w13617 <= pi0182 and w12710;
w13618 <= not w12076 and w13608;
w13619 <= not w13617 and w13618;
w13620 <= not pi0182 and w12100;
w13621 <= not w12709 and not w13494;
w13622 <= not w13620 and w13621;
w13623 <= w13493 and not w13622;
w13624 <= not pi0168 and w12160;
w13625 <= not w12709 and not w13624;
w13626 <= pi0151 and not w13625;
w13627 <= not pi0151 and not w13447;
w13628 <= not w12710 and w13627;
w13629 <= pi0160 and not w13626;
w13630 <= not w13628 and w13629;
w13631 <= not pi0151 and not w12076;
w13632 <= pi0151 and w12313;
w13633 <= not pi0168 and not w13631;
w13634 <= not w13632 and w13633;
w13635 <= not pi0151 and w12006;
w13636 <= pi0168 and not w13635;
w13637 <= not w12100 and w13636;
w13638 <= not w13634 and not w13637;
w13639 <= not pi0160 and not w12709;
w13640 <= not w13638 and w13639;
w13641 <= pi0299 and not w13630;
w13642 <= not w13640 and w13641;
w13643 <= pi0232 and not w13619;
w13644 <= not w13623 and w13643;
w13645 <= not w13642 and w13644;
w13646 <= not pi0039 and not w13616;
w13647 <= not w13645 and w13646;
w13648 <= w171 and not w13647;
w13649 <= not w13615 and w13648;
w13650 <= w98 and not w12896;
w13651 <= not w13466 and w13650;
w13652 <= not w13649 and w13651;
w13653 <= not w13451 and not w13465;
w13654 <= not w13575 and w13653;
w13655 <= not w13652 and w13654;
w13656 <= w4989 and not w13655;
w13657 <= not w13574 and w13656;
w13658 <= not w13456 and not w13657;
w13659 <= not pi0133 and not w12472;
w13660 <= pi0145 and w12277;
w13661 <= w12856 and not w13660;
w13662 <= pi0197 and w12220;
w13663 <= w12857 and not w13662;
w13664 <= w12002 and not w13663;
w13665 <= pi0299 and not w13664;
w13666 <= not w13661 and not w13665;
w13667 <= pi0232 and not w13666;
w13668 <= w12862 and not w13667;
w13669 <= not w6775 and w12066;
w13670 <= not pi0039 and w12002;
w13671 <= not w13669 and w13670;
w13672 <= not pi0038 and not w13671;
w13673 <= not w13668 and w13672;
w13674 <= w12036 and not w13673;
w13675 <= w12031 and not w13674;
w13676 <= not w12019 and not w13675;
w13677 <= not w13659 and not w13676;
w13678 <= not pi0183 and not pi0299;
w13679 <= not pi0149 and pi0299;
w13680 <= not w13678 and not w13679;
w13681 <= w5036 and w13680;
w13682 <= pi0087 and not w13681;
w13683 <= not w6772 and w12095;
w13684 <= not w3760 and not w12095;
w13685 <= not w12148 and not w13684;
w13686 <= w6772 and w13685;
w13687 <= not pi0039 and pi0176;
w13688 <= not w13683 and w13687;
w13689 <= not w13686 and w13688;
w13690 <= not w3340 and not w13662;
w13691 <= w4203 and not w13690;
w13692 <= not pi0145 and not w5114;
w13693 <= not pi0299 and not w13692;
w13694 <= not w12566 and w13693;
w13695 <= not w13691 and not w13694;
w13696 <= w84 and not w13695;
w13697 <= pi0232 and not w13696;
w13698 <= not w12507 and not w13697;
w13699 <= pi0039 and not w13698;
w13700 <= pi0154 and pi0232;
w13701 <= pi0299 and w13700;
w13702 <= w12095 and not w13701;
w13703 <= w13685 and w13701;
w13704 <= not pi0039 and not pi0176;
w13705 <= not w13702 and w13704;
w13706 <= not w13703 and w13705;
w13707 <= w8937 and not w13699;
w13708 <= not w13689 and w13707;
w13709 <= not w13706 and w13708;
w13710 <= not pi0087 and w13659;
w13711 <= not w13709 and w13710;
w13712 <= not w13677 and not w13682;
w13713 <= not w13711 and w13712;
w13714 <= w4989 and not w13713;
w13715 <= pi0149 and w12483;
w13716 <= w12003 and not w13659;
w13717 <= not w4989 and not w13715;
w13718 <= not w13716 and w13717;
w13719 <= not w13714 and not w13718;
w13720 <= not w4989 and w13428;
w13721 <= not pi0136 and w13309;
w13722 <= not pi0135 and w13721;
w13723 <= pi0134 and not w13722;
w13724 <= w12001 and not w13723;
w13725 <= pi0171 and w3760;
w13726 <= not w12001 and w13725;
w13727 <= pi0232 and w13726;
w13728 <= w13720 and not w13727;
w13729 <= not w13724 and w13728;
w13730 <= pi0192 and not pi0299;
w13731 <= pi0171 and pi0299;
w13732 <= not w13730 and not w13731;
w13733 <= w5036 and not w13732;
w13734 <= w12159 and not w13733;
w13735 <= not w12882 and not w13734;
w13736 <= w12018 and not w13735;
w13737 <= not w171 and w13735;
w13738 <= w98 and not w13737;
w13739 <= not pi0051 and not w13726;
w13740 <= not pi0164 and pi0216;
w13741 <= w3942 and not w13740;
w13742 <= not w13739 and not w13741;
w13743 <= not w12239 and not w13725;
w13744 <= pi0171 and w12511;
w13745 <= not w13743 and not w13744;
w13746 <= not pi0216 and not w13745;
w13747 <= pi0171 and w13359;
w13748 <= not pi0171 and w13361;
w13749 <= pi0164 and pi0216;
w13750 <= not w13747 and w13749;
w13751 <= not w13748 and w13750;
w13752 <= not w13746 and not w13751;
w13753 <= w3942 and not w13752;
w13754 <= not w13742 and not w13753;
w13755 <= pi0299 and not w13754;
w13756 <= not pi0192 and not pi0299;
w13757 <= not w13375 and w13756;
w13758 <= pi0039 and pi0186;
w13759 <= not w13386 and w13730;
w13760 <= not w13757 and not w13758;
w13761 <= not w13759 and w13760;
w13762 <= not w13378 and w13756;
w13763 <= not w13393 and w13730;
w13764 <= pi0186 and not w13762;
w13765 <= not w13763 and w13764;
w13766 <= not w13761 and not w13765;
w13767 <= not w13755 and not w13766;
w13768 <= pi0232 and not w13767;
w13769 <= w13403 and not w13768;
w13770 <= pi0232 and not w13732;
w13771 <= not w12141 and not w13770;
w13772 <= w13408 and w13770;
w13773 <= not pi0039 and not w13771;
w13774 <= not w13772 and w13773;
w13775 <= w171 and not w13769;
w13776 <= not w13774 and w13775;
w13777 <= w13738 and not w13776;
w13778 <= w13723 and not w13736;
w13779 <= not w13777 and w13778;
w13780 <= w12018 and w13734;
w13781 <= pi0039 and not pi0186;
w13782 <= not w13323 and w13730;
w13783 <= not w13319 and w13756;
w13784 <= not w13782 and not w13783;
w13785 <= w13328 and not w13725;
w13786 <= pi0299 and not w13785;
w13787 <= not w12218 and not w13725;
w13788 <= w1755 and w3760;
w13789 <= w6599 and not w13787;
w13790 <= not w13788 and w13789;
w13791 <= w13786 and not w13790;
w13792 <= w13784 and not w13791;
w13793 <= pi0232 and not w13792;
w13794 <= not w13316 and not w13793;
w13795 <= w13781 and not w13794;
w13796 <= not pi0039 and not w13734;
w13797 <= not w12220 and w13323;
w13798 <= w13730 and not w13797;
w13799 <= not w12845 and w13319;
w13800 <= w13756 and not w13799;
w13801 <= not w13798 and not w13800;
w13802 <= not w13791 and w13801;
w13803 <= pi0232 and not w13802;
w13804 <= not w13316 and not w13803;
w13805 <= w13758 and not w13804;
w13806 <= not pi0164 and not w13796;
w13807 <= not w13795 and w13806;
w13808 <= not w13805 and w13807;
w13809 <= not pi0171 and not w12844;
w13810 <= pi0171 and not w13332;
w13811 <= w6599 and not w13809;
w13812 <= not w13810 and w13811;
w13813 <= w13786 and not w13812;
w13814 <= w13784 and not w13813;
w13815 <= pi0232 and not w13814;
w13816 <= not w13316 and not w13815;
w13817 <= w13781 and not w13816;
w13818 <= w13801 and not w13813;
w13819 <= pi0232 and not w13818;
w13820 <= not w13316 and not w13819;
w13821 <= w13758 and not w13820;
w13822 <= pi0164 and not w13796;
w13823 <= not w13817 and w13822;
w13824 <= not w13821 and w13823;
w13825 <= w171 and not w13808;
w13826 <= not w13824 and w13825;
w13827 <= not w12896 and w13738;
w13828 <= not w13826 and w13827;
w13829 <= not w13723 and not w13780;
w13830 <= not w13828 and w13829;
w13831 <= w4989 and not w13779;
w13832 <= not w13830 and w13831;
w13833 <= not w13729 and not w13832;
w13834 <= pi0135 and not w13721;
w13835 <= pi0134 and w13722;
w13836 <= not w13834 and not w13835;
w13837 <= pi0170 and w3760;
w13838 <= w8161 and w13837;
w13839 <= w12159 and not w13838;
w13840 <= pi0194 and w6756;
w13841 <= w13839 and not w13840;
w13842 <= w12018 and w13841;
w13843 <= pi0185 and w12845;
w13844 <= w13319 and not w13843;
w13845 <= not w8545 and w13839;
w13846 <= not pi0194 and not w13845;
w13847 <= not w13844 and w13846;
w13848 <= not pi0185 and w13323;
w13849 <= pi0170 and w5036;
w13850 <= not w6756 and not w13849;
w13851 <= w12159 and w13850;
w13852 <= not w8545 and w13851;
w13853 <= pi0194 and not w13852;
w13854 <= not w13797 and w13853;
w13855 <= not w13848 and w13854;
w13856 <= not w13847 and not w13855;
w13857 <= not pi0299 and not w13856;
w13858 <= w13328 and not w13837;
w13859 <= pi0150 and pi0299;
w13860 <= not pi0170 and not w12844;
w13861 <= pi0170 and not w13332;
w13862 <= w6599 and not w13860;
w13863 <= not w13861 and w13862;
w13864 <= w13859 and not w13863;
w13865 <= not w12218 and not w13837;
w13866 <= w1978 and w3760;
w13867 <= w6599 and not w13865;
w13868 <= not w13866 and w13867;
w13869 <= w13161 and not w13868;
w13870 <= not w13864 and not w13869;
w13871 <= not w13846 and not w13853;
w13872 <= not w13858 and not w13871;
w13873 <= not w13870 and w13872;
w13874 <= not w13857 and not w13873;
w13875 <= pi0232 and not w13874;
w13876 <= not w13317 and not w13871;
w13877 <= not w13875 and not w13876;
w13878 <= not pi0100 and not w13877;
w13879 <= not w12882 and not w13841;
w13880 <= pi0100 and w13879;
w13881 <= w98 and not w13880;
w13882 <= not w12030 and w13881;
w13883 <= not w13878 and w13882;
w13884 <= w13836 and not w13842;
w13885 <= not w13883 and w13884;
w13886 <= not w12882 and not w13839;
w13887 <= pi0038 and not w13886;
w13888 <= not w12001 and w13837;
w13889 <= not pi0051 and not w13888;
w13890 <= not w3942 and w13889;
w13891 <= pi0170 and w12511;
w13892 <= not w12239 and not w13837;
w13893 <= w5133 and not w13891;
w13894 <= not w13892 and w13893;
w13895 <= not w6599 and not w13894;
w13896 <= not pi0170 and w13361;
w13897 <= pi0170 and w13359;
w13898 <= pi0216 and not w13897;
w13899 <= not w13896 and w13898;
w13900 <= not w13895 and not w13899;
w13901 <= w13859 and not w13890;
w13902 <= not w13900 and w13901;
w13903 <= not w5133 and w13889;
w13904 <= w13161 and not w13903;
w13905 <= not w13894 and w13904;
w13906 <= not w13902 and not w13905;
w13907 <= not pi0185 and w13375;
w13908 <= pi0185 and w13378;
w13909 <= not pi0299 and not w13907;
w13910 <= not w13908 and w13909;
w13911 <= w13906 and not w13910;
w13912 <= pi0232 and not w13911;
w13913 <= w13403 and not w13912;
w13914 <= not pi0299 and not w12141;
w13915 <= pi0170 and not w13408;
w13916 <= not pi0170 and w12141;
w13917 <= w8161 and not w13916;
w13918 <= not w13915 and w13917;
w13919 <= w13406 and not w13918;
w13920 <= not w13914 and w13919;
w13921 <= not w13913 and not w13920;
w13922 <= not pi0038 and not w13921;
w13923 <= not pi0194 and not w13887;
w13924 <= not w13922 and w13923;
w13925 <= not w12882 and not w13851;
w13926 <= pi0038 and not w13925;
w13927 <= not pi0185 and w13386;
w13928 <= pi0185 and w13393;
w13929 <= not pi0299 and not w13927;
w13930 <= not w13928 and w13929;
w13931 <= w13906 and not w13930;
w13932 <= pi0232 and not w13931;
w13933 <= w13403 and not w13932;
w13934 <= w8165 and w13408;
w13935 <= w13919 and not w13934;
w13936 <= not w13933 and not w13935;
w13937 <= not pi0038 and not w13936;
w13938 <= pi0194 and not w13926;
w13939 <= not w13937 and w13938;
w13940 <= not w13924 and not w13939;
w13941 <= not pi0100 and not w13940;
w13942 <= w13881 and not w13941;
w13943 <= w12018 and not w13879;
w13944 <= not w13836 and not w13943;
w13945 <= not w13942 and w13944;
w13946 <= w4989 and not w13885;
w13947 <= not w13945 and w13946;
w13948 <= w12001 and w13836;
w13949 <= not w12001 and w13849;
w13950 <= w13720 and not w13949;
w13951 <= not w13948 and w13950;
w13952 <= not w13947 and not w13951;
w13953 <= pi0136 and not w13309;
w13954 <= not w13721 and not w13953;
w13955 <= not w11991 and not w13954;
w13956 <= not w12159 and w13955;
w13957 <= pi0148 and w5036;
w13958 <= not w12001 and not w13957;
w13959 <= not w13956 and not w13958;
w13960 <= w13720 and not w13959;
w13961 <= w7302 and not w12001;
w13962 <= not pi0051 and not w13961;
w13963 <= w12018 and w13962;
w13964 <= not w171 and not w13962;
w13965 <= not w7301 and not w13408;
w13966 <= w7301 and w12141;
w13967 <= pi0232 and not w13966;
w13968 <= not w13965 and w13967;
w13969 <= w13406 and not w13968;
w13970 <= not pi0184 and w13386;
w13971 <= pi0184 and w13393;
w13972 <= w7299 and not w13970;
w13973 <= not w13971 and w13972;
w13974 <= not pi0141 and not pi0299;
w13975 <= not pi0184 and w13375;
w13976 <= pi0184 and w13378;
w13977 <= w13974 and not w13975;
w13978 <= not w13976 and w13977;
w13979 <= not pi0287 and w11228;
w13980 <= pi0216 and not w13979;
w13981 <= w3942 and not w13980;
w13982 <= w12238 and w13981;
w13983 <= not pi0051 and not pi0148;
w13984 <= not w13982 and w13983;
w13985 <= not w3942 and w12882;
w13986 <= not w5133 and not w12882;
w13987 <= not pi0163 and not w13986;
w13988 <= pi0163 and w3942;
w13989 <= w13359 and w13988;
w13990 <= not w13985 and not w13987;
w13991 <= not w13989 and w13990;
w13992 <= w5133 and not w13383;
w13993 <= pi0148 and not w13991;
w13994 <= not w13992 and w13993;
w13995 <= pi0299 and not w13984;
w13996 <= not w13994 and w13995;
w13997 <= not w13978 and not w13996;
w13998 <= not w13973 and w13997;
w13999 <= pi0232 and not w13998;
w14000 <= w13403 and not w13999;
w14001 <= w171 and not w14000;
w14002 <= not w13969 and w14001;
w14003 <= w98 and not w13964;
w14004 <= not w14002 and w14003;
w14005 <= w13955 and not w13963;
w14006 <= not w14004 and w14005;
w14007 <= not w12001 and w13963;
w14008 <= not w8774 and not w12001;
w14009 <= w13962 and w14008;
w14010 <= pi0184 and w12845;
w14011 <= w13319 and not w14010;
w14012 <= w13974 and not w14011;
w14013 <= pi0184 and w12220;
w14014 <= w13323 and not w14013;
w14015 <= w7299 and not w14014;
w14016 <= not w3760 and w13328;
w14017 <= w6599 and w13331;
w14018 <= pi0148 and not w14016;
w14019 <= not w14017 and w14018;
w14020 <= not pi0051 and w12857;
w14021 <= not pi0148 and not w14020;
w14022 <= not w13979 and not w14021;
w14023 <= not pi0148 and w12159;
w14024 <= not w14022 and not w14023;
w14025 <= not w14019 and not w14024;
w14026 <= pi0299 and not w14025;
w14027 <= not w14012 and not w14015;
w14028 <= not w14026 and w14027;
w14029 <= pi0232 and not w14028;
w14030 <= not pi0100 and w13317;
w14031 <= not w14029 and w14030;
w14032 <= not w14009 and not w14031;
w14033 <= w98 and not w14032;
w14034 <= not w13955 and not w14007;
w14035 <= not w14033 and w14034;
w14036 <= w4989 and not w14035;
w14037 <= not w14006 and w14036;
w14038 <= not w13960 and not w14037;
w14039 <= not pi0039 and pi0137;
w14040 <= w7931 and w12436;
w14041 <= w3731 and w9131;
w14042 <= not pi0299 and w4989;
w14043 <= not pi0198 and w9142;
w14044 <= w14042 and w14043;
w14045 <= not w14041 and not w14044;
w14046 <= not w14040 and not w14045;
w14047 <= not pi0210 and w9131;
w14048 <= not w4989 and w14047;
w14049 <= not w14046 and not w14048;
w14050 <= w8041 and not w14049;
w14051 <= not w14039 and not w14050;
w14052 <= not w7302 and w11473;
w14053 <= not pi0039 and not w14052;
w14054 <= not pi0232 and not w9044;
w14055 <= w3761 and w3959;
w14056 <= w6614 and w14055;
w14057 <= w7299 and not w14056;
w14058 <= not w3761 and w7300;
w14059 <= not w7299 and not w9044;
w14060 <= not w14057 and not w14058;
w14061 <= not w14059 and w14060;
w14062 <= pi0232 and not w14061;
w14063 <= not w14054 and not w14062;
w14064 <= pi0039 and not w14063;
w14065 <= w7763 and not w14053;
w14066 <= not w14064 and w14065;
w14067 <= not pi0138 and w14066;
w14068 <= w6813 and not w6845;
w14069 <= pi0092 and not w14068;
w14070 <= w95 and not w14069;
w14071 <= not pi0075 and not w6851;
w14072 <= not w6889 and not w9455;
w14073 <= w6900 and not w14072;
w14074 <= w11378 and not w14073;
w14075 <= not w3805 and not w6889;
w14076 <= w6599 and not w14072;
w14077 <= not w14075 and w14076;
w14078 <= w6854 and not w14077;
w14079 <= not w14074 and not w14078;
w14080 <= not pi0232 and not w14079;
w14081 <= not pi0141 and w14074;
w14082 <= not w6868 and w14073;
w14083 <= w11378 and not w14082;
w14084 <= pi0141 and w14083;
w14085 <= not w6863 and not w14072;
w14086 <= not w6853 and not w14085;
w14087 <= pi0148 and not w14086;
w14088 <= not w7300 and not w14078;
w14089 <= not w14087 and not w14088;
w14090 <= not w14081 and not w14084;
w14091 <= not w14089 and w14090;
w14092 <= pi0232 and not w14091;
w14093 <= not w14080 and not w14092;
w14094 <= pi0039 and not w14093;
w14095 <= pi0299 and not w7168;
w14096 <= not pi0299 and not w7512;
w14097 <= not pi0232 and not w14095;
w14098 <= not w14096 and w14097;
w14099 <= not pi0039 and not w14098;
w14100 <= not w3760 and not w7512;
w14101 <= not w11335 and not w14100;
w14102 <= not pi0299 and not w14101;
w14103 <= pi0141 and w14102;
w14104 <= pi0148 and w3760;
w14105 <= not w7168 and not w14104;
w14106 <= pi0148 and w11300;
w14107 <= not w14105 and not w14106;
w14108 <= pi0299 and not w14107;
w14109 <= not pi0141 and w14096;
w14110 <= pi0232 and not w14109;
w14111 <= not w14103 and w14110;
w14112 <= not w14108 and w14111;
w14113 <= w14099 and not w14112;
w14114 <= w171 and not w14094;
w14115 <= not w14113 and w14114;
w14116 <= not pi0087 and not w14115;
w14117 <= w14071 and not w14116;
w14118 <= not pi0092 and not w14117;
w14119 <= w14070 and not w14118;
w14120 <= not pi0055 and not w14119;
w14121 <= w6814 and not w11249;
w14122 <= pi0055 and not w14121;
w14123 <= not w14120 and not w14122;
w14124 <= w92 and not w14123;
w14125 <= w7446 and not w14124;
w14126 <= pi0138 and w14125;
w14127 <= not pi0118 and w11227;
w14128 <= not pi0139 and w14127;
w14129 <= not w14067 and not w14128;
w14130 <= not w14126 and w14129;
w14131 <= not pi0138 and not w6537;
w14132 <= w14066 and not w14131;
w14133 <= w14125 and w14131;
w14134 <= w14128 and not w14132;
w14135 <= not w14133 and w14134;
w14136 <= not w14130 and not w14135;
w14137 <= w11473 and not w13301;
w14138 <= not pi0039 and not w14137;
w14139 <= not w9040 and w13318;
w14140 <= not w3761 and w6584;
w14141 <= w6583 and not w14056;
w14142 <= not w9043 and not w14140;
w14143 <= not w14139 and not w14141;
w14144 <= w14142 and w14143;
w14145 <= pi0232 and not w14144;
w14146 <= not w14054 and not w14145;
w14147 <= pi0039 and not w14146;
w14148 <= w7763 and not w14138;
w14149 <= not w14147 and w14148;
w14150 <= not pi0139 and w14149;
w14151 <= not pi0169 and w6889;
w14152 <= not w14085 and not w14151;
w14153 <= w6599 and not w14152;
w14154 <= w6854 and not w14153;
w14155 <= not pi0191 and w14074;
w14156 <= pi0191 and w14083;
w14157 <= not w14154 and not w14155;
w14158 <= not w14156 and w14157;
w14159 <= pi0232 and not w14158;
w14160 <= not w14080 and not w14159;
w14161 <= pi0039 and not w14160;
w14162 <= pi0191 and w14102;
w14163 <= not w7168 and not w13327;
w14164 <= pi0169 and w11300;
w14165 <= not w14163 and not w14164;
w14166 <= pi0299 and not w14165;
w14167 <= not pi0191 and w14096;
w14168 <= pi0232 and not w14167;
w14169 <= not w14162 and w14168;
w14170 <= not w14166 and w14169;
w14171 <= w14099 and not w14170;
w14172 <= w171 and not w14161;
w14173 <= not w14171 and w14172;
w14174 <= not pi0087 and not w14173;
w14175 <= w14071 and not w14174;
w14176 <= not pi0092 and not w14175;
w14177 <= w14070 and not w14176;
w14178 <= not pi0055 and not w14177;
w14179 <= not w14122 and not w14178;
w14180 <= w92 and not w14179;
w14181 <= w7446 and not w14180;
w14182 <= pi0139 and w14181;
w14183 <= not w14127 and not w14150;
w14184 <= not w14182 and w14183;
w14185 <= not pi0139 and not w6538;
w14186 <= w14149 and not w14185;
w14187 <= w14181 and w14185;
w14188 <= w14127 and not w14186;
w14189 <= not w14187 and w14188;
w14190 <= not w14184 and not w14189;
w14191 <= not pi0641 and pi1158;
w14192 <= pi0641 and not pi1158;
w14193 <= not w14191 and not w14192;
w14194 <= pi0788 and not w14193;
w14195 <= not pi0648 and pi1159;
w14196 <= pi0648 and not pi1159;
w14197 <= not w14195 and not w14196;
w14198 <= pi0789 and not w14197;
w14199 <= pi0627 and pi1154;
w14200 <= not pi0627 and not pi1154;
w14201 <= pi0781 and not w14199;
w14202 <= not w14200 and w14201;
w14203 <= pi0140 and not w134;
w14204 <= w489 and w3847;
w14205 <= not pi0140 and not w14204;
w14206 <= pi0665 and pi1091;
w14207 <= pi0680 and not w14206;
w14208 <= w489 and w14207;
w14209 <= w3847 and w14208;
w14210 <= pi0038 and not w14209;
w14211 <= not w14205 and w14210;
w14212 <= not w3747 and w3943;
w14213 <= not pi0120 and not w14212;
w14214 <= pi0120 and not w84;
w14215 <= not w14213 and not w14214;
w14216 <= w489 and w14215;
w14217 <= w166 and w14216;
w14218 <= w14207 and w14217;
w14219 <= not pi0661 and not pi0681;
w14220 <= not pi0662 and w14219;
w14221 <= not w14206 and w14216;
w14222 <= not w3755 and w14221;
w14223 <= not pi0824 and not w14212;
w14224 <= w3943 and not w7767;
w14225 <= pi1092 and w14224;
w14226 <= not w8594 and not w14225;
w14227 <= not w14223 and not w14226;
w14228 <= pi1093 and w14227;
w14229 <= not pi0120 and not w14228;
w14230 <= w84 and w489;
w14231 <= pi0120 and not w14230;
w14232 <= not pi1091 and not w14231;
w14233 <= not w14229 and w14232;
w14234 <= w489 and w14212;
w14235 <= w486 and w14234;
w14236 <= pi0829 and not w14225;
w14237 <= not pi0829 and not w14227;
w14238 <= w5080 and not w14236;
w14239 <= not w14237 and w14238;
w14240 <= not w14235 and not w14239;
w14241 <= pi1091 and not w14240;
w14242 <= not pi0120 and not w14241;
w14243 <= not w14231 and not w14242;
w14244 <= not w14233 and not w14243;
w14245 <= not w3760 and w14244;
w14246 <= w3760 and not w14216;
w14247 <= not w14245 and not w14246;
w14248 <= pi0665 and not w14233;
w14249 <= not w14244 and not w14248;
w14250 <= not w14221 and not w14249;
w14251 <= w14247 and not w14250;
w14252 <= w3755 and w14251;
w14253 <= not w14222 and not w14252;
w14254 <= not w14220 and w14253;
w14255 <= w14220 and not w14251;
w14256 <= pi0680 and not w14255;
w14257 <= not w14254 and w14256;
w14258 <= w3768 and not w14257;
w14259 <= w3758 and w14249;
w14260 <= w3760 and not w14244;
w14261 <= not w3760 and w14216;
w14262 <= not w14260 and not w14261;
w14263 <= not w3755 and w14262;
w14264 <= w3755 and w14244;
w14265 <= not w14263 and not w14264;
w14266 <= w14207 and w14265;
w14267 <= not w14220 and w14266;
w14268 <= not w14259 and not w14267;
w14269 <= not w3768 and w14268;
w14270 <= not w166 and not w14258;
w14271 <= not w14269 and w14270;
w14272 <= not w14218 and not w14271;
w14273 <= not pi0223 and not w14272;
w14274 <= w3750 and w11768;
w14275 <= w14230 and not w14274;
w14276 <= pi0120 and not w14275;
w14277 <= not pi0120 and not w14234;
w14278 <= pi1091 and not w14276;
w14279 <= not w14277 and w14278;
w14280 <= pi0120 and pi0824;
w14281 <= w3750 and w14280;
w14282 <= w14232 and not w14281;
w14283 <= not w14277 and w14282;
w14284 <= not w14279 and not w14283;
w14285 <= w3760 and not w14284;
w14286 <= not w14261 and not w14285;
w14287 <= not w3768 and w14286;
w14288 <= not w3760 and w14284;
w14289 <= w14221 and not w14288;
w14290 <= not w14222 and not w14289;
w14291 <= pi0680 and not w14290;
w14292 <= not w14287 and w14291;
w14293 <= w14220 and not w14289;
w14294 <= pi0223 and not w14293;
w14295 <= w14292 and w14294;
w14296 <= not w14273 and not w14295;
w14297 <= not pi0299 and not w14296;
w14298 <= not w3805 and w14268;
w14299 <= w3805 and not w14257;
w14300 <= not w1011 and not w14298;
w14301 <= not w14299 and w14300;
w14302 <= w14207 and w14216;
w14303 <= w1011 and w14302;
w14304 <= not w14301 and not w14303;
w14305 <= not pi0215 and not w14304;
w14306 <= not w3805 and w14286;
w14307 <= w14291 and not w14306;
w14308 <= pi0215 and not w14293;
w14309 <= w14307 and w14308;
w14310 <= not w14305 and not w14309;
w14311 <= pi0299 and not w14310;
w14312 <= not w14297 and not w14311;
w14313 <= pi0140 and not w14312;
w14314 <= pi0039 and pi0140;
w14315 <= not w14207 and w14217;
w14316 <= not pi0680 and not w14265;
w14317 <= w14206 and w14243;
w14318 <= not w3789 and w14317;
w14319 <= w14206 and w14261;
w14320 <= not w3755 and w14319;
w14321 <= not w14318 and not w14320;
w14322 <= not w14220 and not w14321;
w14323 <= w14220 and w14317;
w14324 <= pi0680 and not w14323;
w14325 <= not w14322 and w14324;
w14326 <= not w14316 and not w14325;
w14327 <= not w3768 and not w14326;
w14328 <= pi0616 and not w14216;
w14329 <= pi0614 and not w14216;
w14330 <= not pi0603 and not w14216;
w14331 <= pi0603 and not w14247;
w14332 <= not w14330 and not w14331;
w14333 <= not pi0642 and not w14332;
w14334 <= not w3753 and not w14216;
w14335 <= not w14333 and not w14334;
w14336 <= not pi0614 and not w14335;
w14337 <= not w14329 and not w14336;
w14338 <= not pi0616 and not w14337;
w14339 <= not w14328 and not w14338;
w14340 <= not pi0680 and not w14339;
w14341 <= w14206 and w14216;
w14342 <= w3760 and not w14341;
w14343 <= not w3760 and not w14317;
w14344 <= not w14342 and not w14343;
w14345 <= w3755 and w14344;
w14346 <= not w3755 and w14341;
w14347 <= pi0680 and not w14346;
w14348 <= not w14345 and w14347;
w14349 <= not w14340 and not w14348;
w14350 <= not w14220 and w14349;
w14351 <= pi0680 and not w14344;
w14352 <= w14220 and not w14351;
w14353 <= not w14340 and w14352;
w14354 <= not w14350 and not w14353;
w14355 <= w3768 and w14354;
w14356 <= not w166 and not w14327;
w14357 <= not w14355 and w14356;
w14358 <= not pi0223 and not w14315;
w14359 <= not w14357 and w14358;
w14360 <= not w14246 and not w14288;
w14361 <= w3753 and not w14360;
w14362 <= not w14334 and not w14361;
w14363 <= not pi0614 and not w14362;
w14364 <= not w14329 and not w14363;
w14365 <= not pi0616 and not w14364;
w14366 <= not w14328 and not w14365;
w14367 <= not pi0680 and not w14366;
w14368 <= pi0665 and w14279;
w14369 <= not w3760 and not w14368;
w14370 <= not w14342 and not w14369;
w14371 <= w3758 and not w14370;
w14372 <= w14347 and not w14370;
w14373 <= not w14371 and not w14372;
w14374 <= not w14367 and w14373;
w14375 <= w3768 and w14374;
w14376 <= not pi0616 and w14363;
w14377 <= not w14286 and not w14376;
w14378 <= not pi0680 and not w14377;
w14379 <= pi0680 and not w14368;
w14380 <= not w14320 and w14379;
w14381 <= not w14378 and not w14380;
w14382 <= w14373 and w14381;
w14383 <= not w3768 and w14382;
w14384 <= pi0223 and not w14375;
w14385 <= not w14383 and w14384;
w14386 <= not w14359 and not w14385;
w14387 <= not pi0299 and not w14386;
w14388 <= w1011 and w14215;
w14389 <= w489 and not w14207;
w14390 <= w14388 and w14389;
w14391 <= not w3805 and not w14326;
w14392 <= w3805 and w14354;
w14393 <= not w1011 and not w14391;
w14394 <= not w14392 and w14393;
w14395 <= not pi0215 and not w14390;
w14396 <= not w14394 and w14395;
w14397 <= w3805 and w14374;
w14398 <= not w3805 and w14382;
w14399 <= pi0215 and not w14397;
w14400 <= not w14398 and w14399;
w14401 <= not w14396 and not w14400;
w14402 <= pi0299 and not w14401;
w14403 <= not w14387 and not w14402;
w14404 <= pi0039 and w14403;
w14405 <= not w14314 and not w14404;
w14406 <= not w14313 and not w14405;
w14407 <= not pi0102 and not w8862;
w14408 <= not pi0098 and not w350;
w14409 <= not w14407 and w14408;
w14410 <= w5001 and w9938;
w14411 <= w14409 and w14410;
w14412 <= w6460 and w6704;
w14413 <= w14411 and w14412;
w14414 <= not pi0040 and not w14413;
w14415 <= w7852 and not w14414;
w14416 <= not pi0252 and not w14415;
w14417 <= w326 and w501;
w14418 <= w6459 and w14411;
w14419 <= not pi0047 and not w14418;
w14420 <= pi0314 and w7804;
w14421 <= w14419 and not w14420;
w14422 <= w14417 and not w14421;
w14423 <= not pi0035 and not w14422;
w14424 <= not pi0040 and w7837;
w14425 <= not w14423 and w14424;
w14426 <= pi0252 and not w306;
w14427 <= not w14425 and w14426;
w14428 <= not w14416 and not w14427;
w14429 <= w81 and w14428;
w14430 <= pi1092 and not w9936;
w14431 <= w14429 and w14430;
w14432 <= not pi0088 and not w14409;
w14433 <= w8583 and not w14432;
w14434 <= not pi0252 and w7063;
w14435 <= w14433 and w14434;
w14436 <= w63 and w14433;
w14437 <= not pi0047 and not w14420;
w14438 <= not w14436 and w14437;
w14439 <= w14417 and not w14438;
w14440 <= not pi0035 and not w14439;
w14441 <= pi0252 and w7837;
w14442 <= not w14440 and w14441;
w14443 <= not pi0040 and not w14435;
w14444 <= not w14442 and w14443;
w14445 <= w4980 and w7852;
w14446 <= not w14444 and w14445;
w14447 <= not w14431 and not w14446;
w14448 <= pi1093 and not w14447;
w14449 <= not w486 and not w14448;
w14450 <= pi1092 and w493;
w14451 <= w486 and w14450;
w14452 <= w14429 and w14451;
w14453 <= not w487 and not w14452;
w14454 <= not w14449 and not w14453;
w14455 <= not pi1091 and w14448;
w14456 <= not w14454 and not w14455;
w14457 <= pi0665 and not w14455;
w14458 <= not w14456 and not w14457;
w14459 <= not pi0198 and not w14458;
w14460 <= not w974 and not w14444;
w14461 <= not pi0032 and not w14460;
w14462 <= pi0032 and not w4048;
w14463 <= not pi0095 and w495;
w14464 <= not w14462 and w14463;
w14465 <= not w14461 and w14464;
w14466 <= pi0824 and w14465;
w14467 <= not w14431 and not w14466;
w14468 <= w5189 and not w14467;
w14469 <= not pi0032 and not w14428;
w14470 <= w14464 and not w14469;
w14471 <= not pi0824 and pi0829;
w14472 <= w14470 and w14471;
w14473 <= w14467 and not w14472;
w14474 <= pi1093 and not w14473;
w14475 <= not w486 and not w14474;
w14476 <= not w14453 and not w14475;
w14477 <= not w14468 and not w14476;
w14478 <= pi0665 and not w14468;
w14479 <= not w14477 and not w14478;
w14480 <= pi0198 and not w14479;
w14481 <= not w14459 and not w14480;
w14482 <= pi0680 and w14481;
w14483 <= not pi0299 and not w14482;
w14484 <= pi0210 and not w14479;
w14485 <= not pi0210 and not w14458;
w14486 <= not w14484 and not w14485;
w14487 <= pi0680 and w14486;
w14488 <= pi0299 and not w14487;
w14489 <= not w14483 and not w14488;
w14490 <= pi0140 and w14489;
w14491 <= not pi0198 and w14456;
w14492 <= pi0198 and w14477;
w14493 <= not w14491 and not w14492;
w14494 <= pi0665 and w14476;
w14495 <= pi0198 and not w14494;
w14496 <= pi0665 and w14454;
w14497 <= not pi0198 and not w14496;
w14498 <= not w14495 and not w14497;
w14499 <= pi0680 and not w14498;
w14500 <= w14493 and not w14499;
w14501 <= not pi0299 and not w14500;
w14502 <= not pi0210 and w14456;
w14503 <= pi0210 and w14477;
w14504 <= not w14502 and not w14503;
w14505 <= not pi0210 and not w14496;
w14506 <= pi0210 and not w14494;
w14507 <= not w14505 and not w14506;
w14508 <= pi0680 and not w14507;
w14509 <= w14504 and not w14508;
w14510 <= pi0299 and not w14509;
w14511 <= not w14501 and not w14510;
w14512 <= not pi0140 and not w14511;
w14513 <= not pi0039 and not w14490;
w14514 <= not w14512 and w14513;
w14515 <= not w14406 and not w14514;
w14516 <= not pi0038 and not w14515;
w14517 <= not pi0738 and not w14211;
w14518 <= not w14516 and w14517;
w14519 <= pi0299 and not w14504;
w14520 <= not pi0299 and not w14493;
w14521 <= not w14519 and not w14520;
w14522 <= not pi0039 and not w14521;
w14523 <= pi0681 and not w14377;
w14524 <= pi0661 and w14377;
w14525 <= not w3756 and not w14366;
w14526 <= w3756 and w14284;
w14527 <= not w3760 and not w14526;
w14528 <= not w14525 and w14527;
w14529 <= not w14285 and not w14528;
w14530 <= not pi0661 and not w14529;
w14531 <= not pi0681 and not w14524;
w14532 <= not w14530 and w14531;
w14533 <= not w14523 and not w14532;
w14534 <= not w3768 and not w14533;
w14535 <= pi0681 and not w14366;
w14536 <= pi0680 and not w14360;
w14537 <= not pi0680 and not w14216;
w14538 <= pi0616 and w14220;
w14539 <= not w14537 and w14538;
w14540 <= not w14536 and w14539;
w14541 <= pi0616 and w14216;
w14542 <= not w14220 and w14541;
w14543 <= not w14540 and not w14542;
w14544 <= not pi0616 and not w14220;
w14545 <= w14364 and w14544;
w14546 <= not pi0680 and w14365;
w14547 <= not pi0616 and w14220;
w14548 <= not w14536 and w14547;
w14549 <= not w14546 and w14548;
w14550 <= not w14545 and not w14549;
w14551 <= not pi0681 and w14543;
w14552 <= w14550 and w14551;
w14553 <= not w14535 and not w14552;
w14554 <= w3768 and not w14553;
w14555 <= not w14534 and not w14554;
w14556 <= pi0223 and not w14555;
w14557 <= pi0681 and not w14339;
w14558 <= pi0680 and not w14247;
w14559 <= pi0614 and w14220;
w14560 <= not w14537 and w14559;
w14561 <= not w14558 and w14560;
w14562 <= pi0614 and w14216;
w14563 <= not w14220 and w14562;
w14564 <= not w14561 and not w14563;
w14565 <= not pi0614 and not w3758;
w14566 <= not pi0616 and not w14335;
w14567 <= not w14328 and w14565;
w14568 <= not w14566 and w14567;
w14569 <= not pi0614 and w3758;
w14570 <= w14247 and w14569;
w14571 <= not w14568 and not w14570;
w14572 <= not pi0681 and w14564;
w14573 <= w14571 and w14572;
w14574 <= not w14557 and not w14573;
w14575 <= w3768 and not w14574;
w14576 <= pi0681 and not w14265;
w14577 <= w3757 and not w14244;
w14578 <= not w3757 and w14265;
w14579 <= not pi0681 and not w14577;
w14580 <= not w14578 and w14579;
w14581 <= not w14576 and not w14580;
w14582 <= not w3768 and not w14581;
w14583 <= not w14575 and not w14582;
w14584 <= not w166 and w14583;
w14585 <= not pi0223 and not w14217;
w14586 <= not w14584 and w14585;
w14587 <= not w14556 and not w14586;
w14588 <= not pi0299 and not w14587;
w14589 <= w1011 and w14216;
w14590 <= w3804 and not w14574;
w14591 <= not w3804 and not w14581;
w14592 <= w3799 and not w14591;
w14593 <= not w14590 and w14592;
w14594 <= not w1011 and w14593;
w14595 <= not w3799 and w14581;
w14596 <= not w1011 and w14595;
w14597 <= not pi0215 and not w14589;
w14598 <= not w14596 and w14597;
w14599 <= not w14594 and w14598;
w14600 <= not w3799 and w14533;
w14601 <= not w3804 and not w14533;
w14602 <= w3804 and not w14553;
w14603 <= w3799 and not w14602;
w14604 <= not w14601 and w14603;
w14605 <= not w14600 and not w14604;
w14606 <= pi0215 and w14605;
w14607 <= not w14599 and not w14606;
w14608 <= pi0299 and not w14607;
w14609 <= not w14588 and not w14608;
w14610 <= pi0039 and not w14609;
w14611 <= not w14522 and not w14610;
w14612 <= not pi0038 and not w14611;
w14613 <= w489 and w3698;
w14614 <= pi0038 and not w14613;
w14615 <= not w14612 and not w14614;
w14616 <= not pi0140 and pi0738;
w14617 <= not w14615 and w14616;
w14618 <= w134 and not w14617;
w14619 <= not w14518 and w14618;
w14620 <= not w14203 and not w14619;
w14621 <= not pi0778 and not w14620;
w14622 <= w134 and w14615;
w14623 <= not pi0140 and not w14622;
w14624 <= not pi0625 and w14623;
w14625 <= pi0625 and w14620;
w14626 <= pi1153 and not w14624;
w14627 <= not w14625 and w14626;
w14628 <= not pi0625 and w14620;
w14629 <= pi0625 and w14623;
w14630 <= not pi1153 and not w14629;
w14631 <= not w14628 and w14630;
w14632 <= not w14627 and not w14631;
w14633 <= pi0778 and not w14632;
w14634 <= not w14621 and not w14633;
w14635 <= pi0660 and pi1155;
w14636 <= not pi0660 and not pi1155;
w14637 <= pi0785 and not w14635;
w14638 <= not w14636 and w14637;
w14639 <= not w14634 and not w14638;
w14640 <= not w14623 and w14638;
w14641 <= not w14639 and not w14640;
w14642 <= not w14202 and w14641;
w14643 <= w14202 and w14623;
w14644 <= not w14642 and not w14643;
w14645 <= not w14198 and w14644;
w14646 <= w14198 and not w14623;
w14647 <= not w14645 and not w14646;
w14648 <= not w14194 and w14647;
w14649 <= w14194 and w14623;
w14650 <= not w14648 and not w14649;
w14651 <= not pi0792 and w14650;
w14652 <= not pi0628 and w14623;
w14653 <= pi0628 and not w14650;
w14654 <= pi1156 and not w14652;
w14655 <= not w14653 and w14654;
w14656 <= pi0628 and w14623;
w14657 <= not pi0628 and not w14650;
w14658 <= not pi1156 and not w14656;
w14659 <= not w14657 and w14658;
w14660 <= not w14655 and not w14659;
w14661 <= pi0792 and not w14660;
w14662 <= not w14651 and not w14661;
w14663 <= not pi0787 and not w14662;
w14664 <= not pi0647 and w14623;
w14665 <= pi0647 and w14662;
w14666 <= pi1157 and not w14664;
w14667 <= not w14665 and w14666;
w14668 <= not pi0647 and w14662;
w14669 <= pi0647 and w14623;
w14670 <= not pi1157 and not w14669;
w14671 <= not w14668 and w14670;
w14672 <= not w14667 and not w14671;
w14673 <= pi0787 and not w14672;
w14674 <= not w14663 and not w14673;
w14675 <= not pi0644 and w14674;
w14676 <= not pi0619 and w14623;
w14677 <= not pi0608 and pi1153;
w14678 <= pi0608 and not pi1153;
w14679 <= not w14677 and not w14678;
w14680 <= pi0778 and not w14679;
w14681 <= pi0621 and w14454;
w14682 <= not pi0210 and not w14681;
w14683 <= pi0621 and w14476;
w14684 <= pi0210 and not w14683;
w14685 <= not w14682 and not w14684;
w14686 <= pi0603 and not w14685;
w14687 <= w14504 and not w14686;
w14688 <= pi0299 and not w14687;
w14689 <= not pi0198 and not w14681;
w14690 <= pi0198 and not w14683;
w14691 <= not w14689 and not w14690;
w14692 <= pi0621 and not w14455;
w14693 <= not w14456 and not w14692;
w14694 <= not pi0198 and w14693;
w14695 <= pi0621 and not w14468;
w14696 <= not w14477 and not w14695;
w14697 <= pi0198 and w14696;
w14698 <= not w14694 and not w14697;
w14699 <= not pi0603 and not w14698;
w14700 <= not w14691 and not w14699;
w14701 <= not pi0299 and w14700;
w14702 <= not w14688 and not w14701;
w14703 <= not pi0039 and not w14702;
w14704 <= not w3758 and not w14265;
w14705 <= w3758 and w14244;
w14706 <= not w14704 and not w14705;
w14707 <= pi0621 and pi1091;
w14708 <= w14243 and w14707;
w14709 <= pi0621 and not w14233;
w14710 <= not w14244 and not w14709;
w14711 <= not pi0603 and w14710;
w14712 <= not pi0603 and w14262;
w14713 <= w3760 and w14708;
w14714 <= w14261 and w14707;
w14715 <= pi0603 and not w14714;
w14716 <= not w14713 and w14715;
w14717 <= not w14712 and not w14716;
w14718 <= not w14708 and not w14711;
w14719 <= not w14717 and w14718;
w14720 <= w14706 and not w14719;
w14721 <= not w3805 and not w14720;
w14722 <= w14216 and w14707;
w14723 <= w3760 and not w14722;
w14724 <= not w3760 and not w14708;
w14725 <= not w14723 and not w14724;
w14726 <= pi0603 and not w14725;
w14727 <= w14247 and not w14726;
w14728 <= w3758 and not w14727;
w14729 <= not pi0614 and not pi0642;
w14730 <= not pi0616 and w14729;
w14731 <= pi0603 and not w14707;
w14732 <= w14216 and not w14731;
w14733 <= not w14730 and w14732;
w14734 <= not w14330 and w14730;
w14735 <= not w14726 and w14734;
w14736 <= not w14733 and not w14735;
w14737 <= not w3758 and w14736;
w14738 <= not w14728 and not w14737;
w14739 <= w3805 and not w14738;
w14740 <= not w1011 and not w14721;
w14741 <= not w14739 and w14740;
w14742 <= w1011 and w14732;
w14743 <= not w14741 and not w14742;
w14744 <= not pi0215 and not w14743;
w14745 <= w489 and not w14731;
w14746 <= not w14286 and w14745;
w14747 <= w3755 and not w14279;
w14748 <= w14746 and not w14747;
w14749 <= not w3758 and not w14748;
w14750 <= not w14284 and w14745;
w14751 <= w3758 and not w14750;
w14752 <= not w14749 and not w14751;
w14753 <= not w3805 and not w14752;
w14754 <= pi0621 and w14279;
w14755 <= not w3760 and not w14754;
w14756 <= not w14723 and not w14755;
w14757 <= pi0603 and not w14756;
w14758 <= w14734 and not w14757;
w14759 <= not w14733 and not w14758;
w14760 <= not w3758 and not w14759;
w14761 <= w3758 and w14360;
w14762 <= not w14757 and w14761;
w14763 <= not w14760 and not w14762;
w14764 <= w3805 and w14763;
w14765 <= pi0215 and not w14753;
w14766 <= not w14764 and w14765;
w14767 <= not w14744 and not w14766;
w14768 <= pi0299 and not w14767;
w14769 <= not w3768 and not w14720;
w14770 <= w3768 and not w14738;
w14771 <= not w166 and not w14769;
w14772 <= not w14770 and w14771;
w14773 <= w166 and w14732;
w14774 <= not w14772 and not w14773;
w14775 <= not pi0223 and not w14774;
w14776 <= not w3768 and not w14752;
w14777 <= w3768 and w14763;
w14778 <= pi0223 and not w14776;
w14779 <= not w14777 and w14778;
w14780 <= not w14775 and not w14779;
w14781 <= not pi0299 and not w14780;
w14782 <= not w14768 and not w14781;
w14783 <= pi0039 and w14782;
w14784 <= not w14703 and not w14783;
w14785 <= not pi0761 and w14784;
w14786 <= pi0761 and w14611;
w14787 <= not pi0140 and not w14785;
w14788 <= not w14786 and w14787;
w14789 <= pi0603 and not w14698;
w14790 <= not pi0299 and not w14789;
w14791 <= not pi0210 and not w14693;
w14792 <= pi0210 and not w14696;
w14793 <= not w14791 and not w14792;
w14794 <= pi0603 and w14793;
w14795 <= pi0299 and not w14794;
w14796 <= not w14790 and not w14795;
w14797 <= not pi0039 and not w14796;
w14798 <= w14216 and w14731;
w14799 <= not w14288 and w14798;
w14800 <= not w14286 and w14798;
w14801 <= w14288 and w14730;
w14802 <= w14800 and not w14801;
w14803 <= not w3758 and w14802;
w14804 <= not w14799 and not w14803;
w14805 <= not w14306 and not w14804;
w14806 <= pi0215 and not w14805;
w14807 <= w489 and w14731;
w14808 <= w14388 and w14807;
w14809 <= w14247 and w14731;
w14810 <= w3758 and w14809;
w14811 <= not w14730 and w14798;
w14812 <= w14730 and w14809;
w14813 <= not w14811 and not w14812;
w14814 <= not w3758 and not w14813;
w14815 <= not w14810 and not w14814;
w14816 <= w3805 and w14815;
w14817 <= w14706 and w14731;
w14818 <= not w3805 and not w14817;
w14819 <= not w1011 and not w14816;
w14820 <= not w14818 and w14819;
w14821 <= not pi0215 and not w14808;
w14822 <= not w14820 and w14821;
w14823 <= pi0299 and not w14806;
w14824 <= not w14822 and w14823;
w14825 <= not w14287 and not w14804;
w14826 <= pi0223 and not w14825;
w14827 <= w3768 and w14815;
w14828 <= not w3768 and not w14817;
w14829 <= not w166 and not w14827;
w14830 <= not w14828 and w14829;
w14831 <= w14217 and w14731;
w14832 <= not pi0223 and not w14831;
w14833 <= not w14830 and w14832;
w14834 <= not pi0299 and not w14826;
w14835 <= not w14833 and w14834;
w14836 <= not w14824 and not w14835;
w14837 <= pi0039 and w14836;
w14838 <= not w14797 and not w14837;
w14839 <= pi0140 and not pi0761;
w14840 <= w14838 and w14839;
w14841 <= not w14788 and not w14840;
w14842 <= not pi0038 and not w14841;
w14843 <= w3847 and w14807;
w14844 <= not pi0761 and w14843;
w14845 <= not w14205 and not w14844;
w14846 <= pi0038 and not w14845;
w14847 <= not w14842 and not w14846;
w14848 <= w134 and w14847;
w14849 <= not w14203 and not w14848;
w14850 <= not w14680 and not w14849;
w14851 <= not w14623 and w14680;
w14852 <= not w14850 and not w14851;
w14853 <= not pi0785 and not w14852;
w14854 <= pi0609 and not w14680;
w14855 <= not w14623 and not w14854;
w14856 <= pi0609 and w14850;
w14857 <= not w14855 and not w14856;
w14858 <= pi1155 and not w14857;
w14859 <= not pi0609 and not w14680;
w14860 <= not w14623 and not w14859;
w14861 <= not pi0609 and w14850;
w14862 <= not w14860 and not w14861;
w14863 <= not pi1155 and not w14862;
w14864 <= not w14858 and not w14863;
w14865 <= pi0785 and not w14864;
w14866 <= not w14853 and not w14865;
w14867 <= not pi0781 and not w14866;
w14868 <= not pi0618 and w14623;
w14869 <= pi0618 and w14866;
w14870 <= pi1154 and not w14868;
w14871 <= not w14869 and w14870;
w14872 <= not pi0618 and w14866;
w14873 <= pi0618 and w14623;
w14874 <= not pi1154 and not w14873;
w14875 <= not w14872 and w14874;
w14876 <= not w14871 and not w14875;
w14877 <= pi0781 and not w14876;
w14878 <= not w14867 and not w14877;
w14879 <= pi0619 and w14878;
w14880 <= pi1159 and not w14676;
w14881 <= not w14879 and w14880;
w14882 <= pi0738 and not w14847;
w14883 <= not w14284 and w14798;
w14884 <= not w14368 and not w14883;
w14885 <= w3758 and w14884;
w14886 <= pi0680 and not w14220;
w14887 <= not w14319 and not w14368;
w14888 <= not w14800 and w14887;
w14889 <= not w14730 and w14888;
w14890 <= not pi0603 and w14319;
w14891 <= w14884 and not w14890;
w14892 <= w14730 and w14891;
w14893 <= not w14889 and not w14892;
w14894 <= w14886 and not w14893;
w14895 <= not w14885 and not w14894;
w14896 <= not w14378 and w14895;
w14897 <= not w3768 and not w14896;
w14898 <= w14371 and not w14799;
w14899 <= not w14206 and not w14731;
w14900 <= w14216 and not w14899;
w14901 <= pi0616 and not w14900;
w14902 <= pi0614 and not w14900;
w14903 <= pi0642 and not w14900;
w14904 <= not pi0642 and not w14370;
w14905 <= not w14799 and w14904;
w14906 <= w14891 and w14905;
w14907 <= not w14903 and not w14906;
w14908 <= not pi0614 and not w14907;
w14909 <= not w14902 and not w14908;
w14910 <= not pi0616 and not w14909;
w14911 <= not w14901 and not w14910;
w14912 <= w14886 and not w14911;
w14913 <= not w14367 and not w14898;
w14914 <= not w14912 and w14913;
w14915 <= w3768 and not w14914;
w14916 <= pi0223 and not w14897;
w14917 <= not w14915 and w14916;
w14918 <= pi0680 and w14899;
w14919 <= w14216 and not w14918;
w14920 <= w166 and not w14919;
w14921 <= w14332 and not w14899;
w14922 <= not pi0642 and not w14921;
w14923 <= not w14903 and not w14922;
w14924 <= not pi0614 and not w14923;
w14925 <= not w14902 and not w14924;
w14926 <= not pi0616 and not w14925;
w14927 <= not w14901 and not w14926;
w14928 <= w14886 and not w14927;
w14929 <= not pi0603 and not w14344;
w14930 <= pi0603 and not pi0665;
w14931 <= w14707 and w14930;
w14932 <= not w14331 and not w14931;
w14933 <= not w14929 and w14932;
w14934 <= w3758 and not w14933;
w14935 <= not w14340 and not w14934;
w14936 <= not w14928 and w14935;
w14937 <= w3768 and w14936;
w14938 <= pi0603 and w14710;
w14939 <= pi0603 and not pi0621;
w14940 <= w14317 and not w14939;
w14941 <= w3758 and not w14940;
w14942 <= not w14938 and w14941;
w14943 <= w14265 and not w14899;
w14944 <= w14886 and not w14943;
w14945 <= not w14316 and not w14942;
w14946 <= not w14944 and w14945;
w14947 <= not w3768 and w14946;
w14948 <= not w166 and not w14947;
w14949 <= not w14937 and w14948;
w14950 <= not pi0223 and not w14920;
w14951 <= not w14949 and w14950;
w14952 <= not w14917 and not w14951;
w14953 <= not pi0299 and not w14952;
w14954 <= w1011 and not w14919;
w14955 <= not w3805 and not w14946;
w14956 <= w3805 and not w14936;
w14957 <= not w14955 and not w14956;
w14958 <= not w1011 and not w14957;
w14959 <= not pi0215 and not w14954;
w14960 <= not w14958 and w14959;
w14961 <= w3805 and not w14914;
w14962 <= not w3805 and not w14896;
w14963 <= pi0215 and not w14962;
w14964 <= not w14961 and w14963;
w14965 <= not w14960 and not w14964;
w14966 <= pi0299 and not w14965;
w14967 <= not w14953 and not w14966;
w14968 <= not pi0140 and w14967;
w14969 <= w14589 and w14918;
w14970 <= not w14206 and w14732;
w14971 <= pi0616 and not w14970;
w14972 <= w14886 and not w14971;
w14973 <= not w14729 and w14970;
w14974 <= pi0603 and pi0665;
w14975 <= not pi0603 and not w14221;
w14976 <= not w14974 and not w14975;
w14977 <= not w14726 and w14976;
w14978 <= w14729 and w14977;
w14979 <= not pi0616 and not w14973;
w14980 <= not w14978 and w14979;
w14981 <= w14972 and not w14980;
w14982 <= w14247 and w14934;
w14983 <= not w14981 and not w14982;
w14984 <= w3805 and w14983;
w14985 <= not w14250 and w14717;
w14986 <= pi0616 and not w14985;
w14987 <= not pi0665 and w14708;
w14988 <= pi0603 and not w14987;
w14989 <= not w14250 and not w14262;
w14990 <= not pi0603 and not w14989;
w14991 <= not w14988 and not w14990;
w14992 <= w14729 and w14991;
w14993 <= w14730 and not w14991;
w14994 <= w14985 and not w14993;
w14995 <= not pi0616 and not w14992;
w14996 <= not w14994 and w14995;
w14997 <= not w14986 and not w14996;
w14998 <= not w14220 and not w14997;
w14999 <= w14259 and not w14988;
w15000 <= not w14886 and not w14999;
w15001 <= not w14998 and not w15000;
w15002 <= not w3805 and not w15001;
w15003 <= not w1011 and not w14984;
w15004 <= not w15002 and w15003;
w15005 <= not pi0215 and not w14969;
w15006 <= not w15004 and w15005;
w15007 <= not w14206 and not w14759;
w15008 <= not pi0616 and not w15007;
w15009 <= w14972 and not w15008;
w15010 <= w14762 and w14976;
w15011 <= not w15009 and not w15010;
w15012 <= w3805 and not w15011;
w15013 <= w14746 and w14976;
w15014 <= pi0616 and not w15013;
w15015 <= pi0614 and not pi0616;
w15016 <= not w15013 and w15015;
w15017 <= not w14757 and w14976;
w15018 <= not pi0642 and not w15017;
w15019 <= w15013 and not w15018;
w15020 <= w3754 and not w15019;
w15021 <= not w15016 and not w15020;
w15022 <= not w15014 and w15021;
w15023 <= not w14220 and not w15022;
w15024 <= not w14284 and w14918;
w15025 <= not w14886 and not w15024;
w15026 <= not w15023 and not w15025;
w15027 <= not w3805 and w15026;
w15028 <= pi0215 and not w15012;
w15029 <= not w15027 and w15028;
w15030 <= not w15006 and not w15029;
w15031 <= pi0299 and not w15030;
w15032 <= w14208 and not w14731;
w15033 <= not w14807 and not w15032;
w15034 <= w14216 and not w15033;
w15035 <= w166 and not w15034;
w15036 <= not w3768 and w15001;
w15037 <= w3768 and not w14983;
w15038 <= not w166 and not w15037;
w15039 <= not w15036 and w15038;
w15040 <= w14832 and not w15035;
w15041 <= not w15039 and w15040;
w15042 <= w3768 and w15011;
w15043 <= not w3768 and not w15026;
w15044 <= pi0223 and not w15042;
w15045 <= not w15043 and w15044;
w15046 <= not pi0299 and not w15045;
w15047 <= not w15041 and w15046;
w15048 <= not w15031 and not w15047;
w15049 <= pi0140 and w15048;
w15050 <= pi0761 and not w15049;
w15051 <= not w14968 and w15050;
w15052 <= not w14207 and not w14731;
w15053 <= w14230 and w15052;
w15054 <= not w14213 and w15053;
w15055 <= w166 and w15054;
w15056 <= w14206 and not w14939;
w15057 <= not w14321 and w15056;
w15058 <= w14886 and not w15057;
w15059 <= w14265 and not w14731;
w15060 <= not pi0680 and not w15059;
w15061 <= not w14941 and not w15058;
w15062 <= not w15060 and w15061;
w15063 <= not w3768 and w15062;
w15064 <= not pi0680 and w14736;
w15065 <= w14344 and w15056;
w15066 <= w3758 and not w15065;
w15067 <= w14341 and not w14939;
w15068 <= not w14730 and w15067;
w15069 <= w14206 and w14735;
w15070 <= w14886 and not w15068;
w15071 <= not w15069 and w15070;
w15072 <= not w15064 and not w15066;
w15073 <= not w15071 and w15072;
w15074 <= w3768 and w15073;
w15075 <= not w15063 and not w15074;
w15076 <= not w166 and not w15075;
w15077 <= not pi0223 and not w15055;
w15078 <= not w15076 and w15077;
w15079 <= not w14207 and w14760;
w15080 <= w3758 and not w14939;
w15081 <= w14370 and w15080;
w15082 <= not w15079 and not w15081;
w15083 <= w3768 and not w15082;
w15084 <= not pi0680 and not w14748;
w15085 <= not w14379 and not w14939;
w15086 <= w3758 and not w15085;
w15087 <= not w14759 and not w14887;
w15088 <= w14886 and not w15087;
w15089 <= not w15084 and not w15086;
w15090 <= not w15088 and w15089;
w15091 <= not w3768 and w15090;
w15092 <= pi0223 and not w15083;
w15093 <= not w15091 and w15092;
w15094 <= not w15078 and not w15093;
w15095 <= not pi0299 and not w15094;
w15096 <= w1011 and w15054;
w15097 <= not w3805 and w15062;
w15098 <= w3805 and w15073;
w15099 <= not w15097 and not w15098;
w15100 <= not w1011 and not w15099;
w15101 <= not pi0215 and not w15096;
w15102 <= not w15100 and w15101;
w15103 <= w3805 and not w15082;
w15104 <= not w3805 and w15090;
w15105 <= pi0215 and not w15103;
w15106 <= not w15104 and w15105;
w15107 <= not w15102 and not w15106;
w15108 <= pi0299 and not w15107;
w15109 <= not w15095 and not w15108;
w15110 <= not pi0140 and not w15109;
w15111 <= w14216 and not w15056;
w15112 <= not w14730 and w15111;
w15113 <= w14886 and not w15112;
w15114 <= w14290 and not w14799;
w15115 <= w14730 and not w15114;
w15116 <= w15113 and not w15115;
w15117 <= pi0680 and not w14293;
w15118 <= w14804 and not w15117;
w15119 <= not w15116 and not w15118;
w15120 <= w3768 and not w15119;
w15121 <= not w14803 and not w14883;
w15122 <= w14221 and not w14286;
w15123 <= not w14290 and w15117;
w15124 <= w15122 and w15123;
w15125 <= w15121 and not w15124;
w15126 <= not w3768 and w15125;
w15127 <= pi0223 and not w15126;
w15128 <= not w15120 and w15127;
w15129 <= not pi0680 and w14813;
w15130 <= not w14809 and not w14977;
w15131 <= w14730 and not w15130;
w15132 <= w15113 and not w15131;
w15133 <= w3758 and not w14251;
w15134 <= not w14809 and w15133;
w15135 <= not w15129 and not w15134;
w15136 <= not w15132 and w15135;
w15137 <= w3768 and w15136;
w15138 <= not w14938 and not w14991;
w15139 <= w14730 and not w15138;
w15140 <= not w14262 and w14731;
w15141 <= not w14989 and not w15140;
w15142 <= not w14730 and not w15141;
w15143 <= w14886 and not w15142;
w15144 <= not w15139 and w15143;
w15145 <= not w14259 and not w14886;
w15146 <= not w14817 and w15145;
w15147 <= not w15144 and not w15146;
w15148 <= not w3768 and w15147;
w15149 <= not w166 and not w15137;
w15150 <= not w15148 and w15149;
w15151 <= not pi0223 and not w15035;
w15152 <= not w15150 and w15151;
w15153 <= not pi0299 and not w15128;
w15154 <= not w15152 and w15153;
w15155 <= w1011 and w15034;
w15156 <= not w3805 and w15147;
w15157 <= w3805 and w15136;
w15158 <= not w15156 and not w15157;
w15159 <= not w1011 and not w15158;
w15160 <= not pi0215 and not w15155;
w15161 <= not w15159 and w15160;
w15162 <= not w3805 and not w15125;
w15163 <= w3805 and w15119;
w15164 <= pi0215 and not w15162;
w15165 <= not w15163 and w15164;
w15166 <= not w15161 and not w15165;
w15167 <= pi0299 and not w15166;
w15168 <= not w15154 and not w15167;
w15169 <= pi0140 and w15168;
w15170 <= not pi0761 and not w15110;
w15171 <= not w15169 and w15170;
w15172 <= not w15051 and not w15171;
w15173 <= pi0039 and not w15172;
w15174 <= pi0680 and w14796;
w15175 <= not w14511 and not w15174;
w15176 <= not pi0140 and not w15175;
w15177 <= pi0603 and not w14691;
w15178 <= not pi0603 and not w14481;
w15179 <= not w14974 and not w15177;
w15180 <= not w15178 and w15179;
w15181 <= pi0680 and w15180;
w15182 <= not pi0299 and not w15181;
w15183 <= not pi0603 and not w14486;
w15184 <= not w14686 and not w14974;
w15185 <= not w15183 and w15184;
w15186 <= pi0680 and w15185;
w15187 <= pi0299 and not w15186;
w15188 <= not w15182 and not w15187;
w15189 <= pi0140 and not w15188;
w15190 <= pi0761 and not w15176;
w15191 <= not w15189 and w15190;
w15192 <= w14511 and w14702;
w15193 <= not pi0140 and w15192;
w15194 <= not w14489 and not w14796;
w15195 <= pi0140 and w15194;
w15196 <= not pi0761 and not w15195;
w15197 <= not w15193 and w15196;
w15198 <= not pi0039 and not w15197;
w15199 <= not w15191 and w15198;
w15200 <= not pi0038 and not w15199;
w15201 <= not w15173 and w15200;
w15202 <= pi0140 and not w15033;
w15203 <= w84 and w15202;
w15204 <= not pi0140 and not w15053;
w15205 <= not pi0761 and not w15203;
w15206 <= not w15204 and w15205;
w15207 <= not pi0140 and not w14230;
w15208 <= w14230 and w14918;
w15209 <= pi0761 and not w15207;
w15210 <= not w15208 and w15209;
w15211 <= not w15206 and not w15210;
w15212 <= not pi0039 and not w15211;
w15213 <= pi0038 and not w14314;
w15214 <= not w15212 and w15213;
w15215 <= not w15201 and not w15214;
w15216 <= not pi0738 and not w15215;
w15217 <= w134 and not w14882;
w15218 <= not w15216 and w15217;
w15219 <= not w14203 and not w15218;
w15220 <= not pi0625 and w15219;
w15221 <= pi0625 and w14849;
w15222 <= not pi1153 and not w15221;
w15223 <= not w15220 and w15222;
w15224 <= not pi0608 and not w14627;
w15225 <= not w15223 and w15224;
w15226 <= not pi0625 and w14849;
w15227 <= pi0625 and w15219;
w15228 <= pi1153 and not w15226;
w15229 <= not w15227 and w15228;
w15230 <= pi0608 and not w14631;
w15231 <= not w15229 and w15230;
w15232 <= not w15225 and not w15231;
w15233 <= pi0778 and not w15232;
w15234 <= not pi0778 and w15219;
w15235 <= not w15233 and not w15234;
w15236 <= not pi0609 and not w15235;
w15237 <= pi0609 and w14634;
w15238 <= not pi1155 and not w15237;
w15239 <= not w15236 and w15238;
w15240 <= not pi0660 and not w14858;
w15241 <= not w15239 and w15240;
w15242 <= not pi0609 and w14634;
w15243 <= pi0609 and not w15235;
w15244 <= pi1155 and not w15242;
w15245 <= not w15243 and w15244;
w15246 <= pi0660 and not w14863;
w15247 <= not w15245 and w15246;
w15248 <= not w15241 and not w15247;
w15249 <= pi0785 and not w15248;
w15250 <= not pi0785 and not w15235;
w15251 <= not w15249 and not w15250;
w15252 <= not pi0618 and not w15251;
w15253 <= pi0618 and w14641;
w15254 <= not pi1154 and not w15253;
w15255 <= not w15252 and w15254;
w15256 <= not pi0627 and not w14871;
w15257 <= not w15255 and w15256;
w15258 <= not pi0618 and w14641;
w15259 <= pi0618 and not w15251;
w15260 <= pi1154 and not w15258;
w15261 <= not w15259 and w15260;
w15262 <= pi0627 and not w14875;
w15263 <= not w15261 and w15262;
w15264 <= not w15257 and not w15263;
w15265 <= pi0781 and not w15264;
w15266 <= not pi0781 and not w15251;
w15267 <= not w15265 and not w15266;
w15268 <= not pi0619 and not w15267;
w15269 <= pi0619 and not w14644;
w15270 <= not pi1159 and not w15269;
w15271 <= not w15268 and w15270;
w15272 <= not pi0648 and not w14881;
w15273 <= not w15271 and w15272;
w15274 <= not pi0619 and w14878;
w15275 <= pi0619 and w14623;
w15276 <= not pi1159 and not w15275;
w15277 <= not w15274 and w15276;
w15278 <= pi0619 and not w15267;
w15279 <= not pi0619 and not w14644;
w15280 <= pi1159 and not w15279;
w15281 <= not w15278 and w15280;
w15282 <= pi0648 and not w15277;
w15283 <= not w15281 and w15282;
w15284 <= not w15273 and not w15283;
w15285 <= pi0789 and not w15284;
w15286 <= not pi0789 and not w15267;
w15287 <= not w15285 and not w15286;
w15288 <= not pi0788 and w15287;
w15289 <= not pi0626 and w15287;
w15290 <= pi0626 and not w14647;
w15291 <= not pi0641 and not w15290;
w15292 <= not w15289 and w15291;
w15293 <= not pi0641 and not pi1158;
w15294 <= not pi0789 and not w14878;
w15295 <= not w14881 and not w15277;
w15296 <= pi0789 and not w15295;
w15297 <= not w15294 and not w15296;
w15298 <= not pi0626 and w15297;
w15299 <= pi0626 and w14623;
w15300 <= not pi1158 and not w15299;
w15301 <= not w15298 and w15300;
w15302 <= not w15293 and not w15301;
w15303 <= not w15292 and not w15302;
w15304 <= pi0626 and w15287;
w15305 <= not pi0626 and not w14647;
w15306 <= pi0641 and not w15305;
w15307 <= not w15304 and w15306;
w15308 <= pi0641 and pi1158;
w15309 <= not pi0626 and w14623;
w15310 <= pi0626 and w15297;
w15311 <= pi1158 and not w15309;
w15312 <= not w15310 and w15311;
w15313 <= not w15308 and not w15312;
w15314 <= not w15307 and not w15313;
w15315 <= not w15303 and not w15314;
w15316 <= pi0788 and not w15315;
w15317 <= not w15288 and not w15316;
w15318 <= not pi0628 and w15317;
w15319 <= not w15301 and not w15312;
w15320 <= pi0788 and not w15319;
w15321 <= not pi0788 and not w15297;
w15322 <= not w15320 and not w15321;
w15323 <= pi0628 and w15322;
w15324 <= not pi1156 and not w15323;
w15325 <= not w15318 and w15324;
w15326 <= not pi0629 and not w14655;
w15327 <= not w15325 and w15326;
w15328 <= pi0628 and w15317;
w15329 <= not pi0628 and w15322;
w15330 <= pi1156 and not w15329;
w15331 <= not w15328 and w15330;
w15332 <= pi0629 and not w14659;
w15333 <= not w15331 and w15332;
w15334 <= not w15327 and not w15333;
w15335 <= pi0792 and not w15334;
w15336 <= not pi0792 and w15317;
w15337 <= not w15335 and not w15336;
w15338 <= not pi0647 and not w15337;
w15339 <= not pi0629 and pi1156;
w15340 <= pi0629 and not pi1156;
w15341 <= not w15339 and not w15340;
w15342 <= pi0792 and not w15341;
w15343 <= w15322 and not w15342;
w15344 <= w14623 and w15342;
w15345 <= not w15343 and not w15344;
w15346 <= pi0647 and not w15345;
w15347 <= not pi1157 and not w15346;
w15348 <= not w15338 and w15347;
w15349 <= not pi0630 and not w14667;
w15350 <= not w15348 and w15349;
w15351 <= pi0647 and not w15337;
w15352 <= not pi0647 and not w15345;
w15353 <= pi1157 and not w15352;
w15354 <= not w15351 and w15353;
w15355 <= pi0630 and not w14671;
w15356 <= not w15354 and w15355;
w15357 <= not w15350 and not w15356;
w15358 <= pi0787 and not w15357;
w15359 <= not pi0787 and not w15337;
w15360 <= not w15358 and not w15359;
w15361 <= pi0644 and not w15360;
w15362 <= pi0715 and not w14675;
w15363 <= not w15361 and w15362;
w15364 <= not pi0630 and pi1157;
w15365 <= pi0630 and not pi1157;
w15366 <= not w15364 and not w15365;
w15367 <= pi0787 and not w15366;
w15368 <= w15345 and not w15367;
w15369 <= not w14623 and w15367;
w15370 <= not w15368 and not w15369;
w15371 <= pi0644 and w15370;
w15372 <= not pi0644 and w14623;
w15373 <= not pi0715 and not w15372;
w15374 <= not w15371 and w15373;
w15375 <= pi1160 and not w15374;
w15376 <= not w15363 and w15375;
w15377 <= not pi0644 and not w15360;
w15378 <= pi0644 and w14674;
w15379 <= not pi0715 and not w15378;
w15380 <= not w15377 and w15379;
w15381 <= not pi0644 and w15370;
w15382 <= pi0644 and w14623;
w15383 <= pi0715 and not w15382;
w15384 <= not w15381 and w15383;
w15385 <= not pi1160 and not w15384;
w15386 <= not w15380 and w15385;
w15387 <= pi0790 and not w15376;
w15388 <= not w15386 and w15387;
w15389 <= not pi0790 and w15360;
w15390 <= w4989 and not w15389;
w15391 <= not w15388 and w15390;
w15392 <= not pi0140 and not w4989;
w15393 <= not pi0832 and not w15392;
w15394 <= not w15391 and w15393;
w15395 <= not pi0140 and not w489;
w15396 <= not pi0647 and w15395;
w15397 <= not pi0738 and w14208;
w15398 <= not w15395 and not w15397;
w15399 <= not pi0778 and w15398;
w15400 <= not pi0625 and w15397;
w15401 <= not w15398 and not w15400;
w15402 <= pi1153 and not w15401;
w15403 <= not pi1153 and not w15395;
w15404 <= not w15400 and w15403;
w15405 <= not w15402 and not w15404;
w15406 <= pi0778 and not w15405;
w15407 <= not w15399 and not w15406;
w15408 <= w489 and w14638;
w15409 <= w15407 and not w15408;
w15410 <= w489 and w14202;
w15411 <= w15409 and not w15410;
w15412 <= w489 and w14198;
w15413 <= w15411 and not w15412;
w15414 <= w489 and w14194;
w15415 <= w15413 and not w15414;
w15416 <= not pi0628 and pi1156;
w15417 <= pi0628 and not pi1156;
w15418 <= not w15416 and not w15417;
w15419 <= pi0792 and not w15418;
w15420 <= w489 and w15419;
w15421 <= w15415 and not w15420;
w15422 <= pi0647 and w15421;
w15423 <= pi1157 and not w15396;
w15424 <= not w15422 and w15423;
w15425 <= not pi0628 and w489;
w15426 <= w15415 and not w15425;
w15427 <= pi1156 and not w15426;
w15428 <= not pi0626 and pi1158;
w15429 <= pi0626 and not pi1158;
w15430 <= not w15428 and not w15429;
w15431 <= not pi0626 and pi0641;
w15432 <= pi0626 and not pi0641;
w15433 <= not w15431 and not w15432;
w15434 <= not w15430 and not w15433;
w15435 <= w15413 and w15434;
w15436 <= not pi0626 and w15395;
w15437 <= w489 and w14680;
w15438 <= not pi0761 and w14807;
w15439 <= not w15395 and not w15438;
w15440 <= not w15437 and not w15439;
w15441 <= not pi0785 and not w15440;
w15442 <= w489 and not w14854;
w15443 <= not w15439 and not w15442;
w15444 <= pi1155 and not w15443;
w15445 <= pi0609 and w489;
w15446 <= w15440 and not w15445;
w15447 <= not pi1155 and not w15446;
w15448 <= not w15444 and not w15447;
w15449 <= pi0785 and not w15448;
w15450 <= not w15441 and not w15449;
w15451 <= not pi0781 and not w15450;
w15452 <= not pi0618 and w489;
w15453 <= w15450 and not w15452;
w15454 <= pi1154 and not w15453;
w15455 <= pi0618 and w489;
w15456 <= w15450 and not w15455;
w15457 <= not pi1154 and not w15456;
w15458 <= not w15454 and not w15457;
w15459 <= pi0781 and not w15458;
w15460 <= not w15451 and not w15459;
w15461 <= not pi0789 and not w15460;
w15462 <= not pi0619 and w15395;
w15463 <= pi0619 and w15460;
w15464 <= pi1159 and not w15462;
w15465 <= not w15463 and w15464;
w15466 <= not pi0619 and w15460;
w15467 <= pi0619 and w15395;
w15468 <= not pi1159 and not w15467;
w15469 <= not w15466 and w15468;
w15470 <= not w15465 and not w15469;
w15471 <= pi0789 and not w15470;
w15472 <= not w15461 and not w15471;
w15473 <= pi0626 and w15472;
w15474 <= pi1158 and not w15436;
w15475 <= not w15473 and w15474;
w15476 <= not pi0626 and w15472;
w15477 <= pi0626 and w15395;
w15478 <= not pi1158 and not w15477;
w15479 <= not w15476 and w15478;
w15480 <= not w15475 and not w15479;
w15481 <= not w14193 and w15480;
w15482 <= not w15435 and not w15481;
w15483 <= pi0788 and not w15482;
w15484 <= pi0618 and w15409;
w15485 <= pi0609 and w15407;
w15486 <= not w14731 and not w15398;
w15487 <= pi0625 and w15486;
w15488 <= w15439 and not w15486;
w15489 <= not w15487 and not w15488;
w15490 <= w15403 and not w15489;
w15491 <= not pi0608 and not w15402;
w15492 <= not w15490 and w15491;
w15493 <= pi1153 and w15439;
w15494 <= not w15487 and w15493;
w15495 <= pi0608 and not w15404;
w15496 <= not w15494 and w15495;
w15497 <= not w15492 and not w15496;
w15498 <= pi0778 and not w15497;
w15499 <= not pi0778 and not w15488;
w15500 <= not w15498 and not w15499;
w15501 <= not pi0609 and not w15500;
w15502 <= not pi1155 and not w15485;
w15503 <= not w15501 and w15502;
w15504 <= not pi0660 and not w15444;
w15505 <= not w15503 and w15504;
w15506 <= not pi0609 and w15407;
w15507 <= pi0609 and not w15500;
w15508 <= pi1155 and not w15506;
w15509 <= not w15507 and w15508;
w15510 <= pi0660 and not w15447;
w15511 <= not w15509 and w15510;
w15512 <= not w15505 and not w15511;
w15513 <= pi0785 and not w15512;
w15514 <= not pi0785 and not w15500;
w15515 <= not w15513 and not w15514;
w15516 <= not pi0618 and not w15515;
w15517 <= not pi1154 and not w15484;
w15518 <= not w15516 and w15517;
w15519 <= not pi0627 and not w15454;
w15520 <= not w15518 and w15519;
w15521 <= not pi0618 and w15409;
w15522 <= pi0618 and not w15515;
w15523 <= pi1154 and not w15521;
w15524 <= not w15522 and w15523;
w15525 <= pi0627 and not w15457;
w15526 <= not w15524 and w15525;
w15527 <= not w15520 and not w15526;
w15528 <= pi0781 and not w15527;
w15529 <= not pi0781 and not w15515;
w15530 <= not w15528 and not w15529;
w15531 <= not pi0789 and w15530;
w15532 <= pi0788 and not w15430;
w15533 <= not w14194 and not w15532;
w15534 <= not pi0619 and not w15530;
w15535 <= pi0619 and w15411;
w15536 <= not pi1159 and not w15535;
w15537 <= not w15534 and w15536;
w15538 <= not pi0648 and not w15465;
w15539 <= not w15537 and w15538;
w15540 <= not pi0619 and w15411;
w15541 <= pi0619 and not w15530;
w15542 <= pi1159 and not w15540;
w15543 <= not w15541 and w15542;
w15544 <= pi0648 and not w15469;
w15545 <= not w15543 and w15544;
w15546 <= pi0789 and not w15539;
w15547 <= not w15545 and w15546;
w15548 <= not w15531 and w15533;
w15549 <= not w15547 and w15548;
w15550 <= not w15483 and not w15549;
w15551 <= not pi0628 and not w15550;
w15552 <= not pi0788 and not w15472;
w15553 <= pi0788 and not w15480;
w15554 <= not w15552 and not w15553;
w15555 <= pi0628 and w15554;
w15556 <= not pi1156 and not w15555;
w15557 <= not w15551 and w15556;
w15558 <= not pi0629 and not w15427;
w15559 <= not w15557 and w15558;
w15560 <= pi0628 and w489;
w15561 <= w15415 and not w15560;
w15562 <= not pi1156 and not w15561;
w15563 <= not pi0628 and w15554;
w15564 <= pi0628 and not w15550;
w15565 <= pi1156 and not w15563;
w15566 <= not w15564 and w15565;
w15567 <= pi0629 and not w15562;
w15568 <= not w15566 and w15567;
w15569 <= not w15559 and not w15568;
w15570 <= pi0792 and not w15569;
w15571 <= not pi0792 and not w15550;
w15572 <= not w15570 and not w15571;
w15573 <= not pi0647 and not w15572;
w15574 <= not w15342 and w15554;
w15575 <= w15342 and w15395;
w15576 <= not w15574 and not w15575;
w15577 <= pi0647 and not w15576;
w15578 <= not pi1157 and not w15577;
w15579 <= not w15573 and w15578;
w15580 <= not pi0630 and not w15424;
w15581 <= not w15579 and w15580;
w15582 <= not pi0647 and w15421;
w15583 <= pi0647 and w15395;
w15584 <= not pi1157 and not w15583;
w15585 <= not w15582 and w15584;
w15586 <= pi0647 and not w15572;
w15587 <= not pi0647 and not w15576;
w15588 <= pi1157 and not w15587;
w15589 <= not w15586 and w15588;
w15590 <= pi0630 and not w15585;
w15591 <= not w15589 and w15590;
w15592 <= not w15581 and not w15591;
w15593 <= pi0787 and not w15592;
w15594 <= not pi0787 and not w15572;
w15595 <= not w15593 and not w15594;
w15596 <= not pi0790 and not w15595;
w15597 <= not pi0787 and not w15421;
w15598 <= not w15424 and not w15585;
w15599 <= pi0787 and not w15598;
w15600 <= not w15597 and not w15599;
w15601 <= not pi0644 and w15600;
w15602 <= pi0644 and not w15595;
w15603 <= pi0715 and not w15601;
w15604 <= not w15602 and w15603;
w15605 <= w15367 and not w15395;
w15606 <= not w15367 and w15576;
w15607 <= not w15605 and not w15606;
w15608 <= pi0644 and w15607;
w15609 <= not pi0644 and w15395;
w15610 <= not pi0715 and not w15609;
w15611 <= not w15608 and w15610;
w15612 <= pi1160 and not w15611;
w15613 <= not w15604 and w15612;
w15614 <= not pi0644 and w15607;
w15615 <= pi0644 and w15395;
w15616 <= pi0715 and not w15615;
w15617 <= not w15614 and w15616;
w15618 <= pi0644 and w15600;
w15619 <= not pi0644 and not w15595;
w15620 <= not pi0715 and not w15618;
w15621 <= not w15619 and w15620;
w15622 <= not pi1160 and not w15617;
w15623 <= not w15621 and w15622;
w15624 <= not w15613 and not w15623;
w15625 <= pi0790 and not w15624;
w15626 <= pi0832 and not w15596;
w15627 <= not w15625 and w15626;
w15628 <= not w15394 and not w15627;
w15629 <= not pi0141 and not w14622;
w15630 <= w14198 and not w15629;
w15631 <= pi0141 and not w134;
w15632 <= not pi0141 and not w14204;
w15633 <= w14210 and not w15632;
w15634 <= not pi0039 and w14511;
w15635 <= not w14404 and not w15634;
w15636 <= not pi0141 and w15635;
w15637 <= pi0039 and not w14312;
w15638 <= not pi0039 and w14489;
w15639 <= not w15637 and not w15638;
w15640 <= pi0141 and not w15639;
w15641 <= not pi0038 and not w15640;
w15642 <= not w15636 and w15641;
w15643 <= pi0706 and not w15633;
w15644 <= not w15642 and w15643;
w15645 <= not pi0141 and not pi0706;
w15646 <= not w14615 and w15645;
w15647 <= w134 and not w15646;
w15648 <= not w15644 and w15647;
w15649 <= not w15631 and not w15648;
w15650 <= not pi0778 and not w15649;
w15651 <= not pi0625 and w15629;
w15652 <= pi0625 and w15649;
w15653 <= pi1153 and not w15651;
w15654 <= not w15652 and w15653;
w15655 <= not pi0625 and w15649;
w15656 <= pi0625 and w15629;
w15657 <= not pi1153 and not w15656;
w15658 <= not w15655 and w15657;
w15659 <= not w15654 and not w15658;
w15660 <= pi0778 and not w15659;
w15661 <= not w15650 and not w15660;
w15662 <= not w14638 and not w15661;
w15663 <= w14638 and not w15629;
w15664 <= not w15662 and not w15663;
w15665 <= not w14202 and w15664;
w15666 <= w14202 and w15629;
w15667 <= not w15665 and not w15666;
w15668 <= not w14198 and w15667;
w15669 <= not w15630 and not w15668;
w15670 <= not w14194 and w15669;
w15671 <= w14194 and w15629;
w15672 <= not w15670 and not w15671;
w15673 <= not pi0792 and w15672;
w15674 <= not pi0628 and w15629;
w15675 <= pi0628 and not w15672;
w15676 <= pi1156 and not w15674;
w15677 <= not w15675 and w15676;
w15678 <= pi0628 and w15629;
w15679 <= not pi0628 and not w15672;
w15680 <= not pi1156 and not w15678;
w15681 <= not w15679 and w15680;
w15682 <= not w15677 and not w15681;
w15683 <= pi0792 and not w15682;
w15684 <= not w15673 and not w15683;
w15685 <= not pi0787 and not w15684;
w15686 <= not pi0647 and w15629;
w15687 <= pi0647 and w15684;
w15688 <= pi1157 and not w15686;
w15689 <= not w15687 and w15688;
w15690 <= not pi0647 and w15684;
w15691 <= pi0647 and w15629;
w15692 <= not pi1157 and not w15691;
w15693 <= not w15690 and w15692;
w15694 <= not w15689 and not w15693;
w15695 <= pi0787 and not w15694;
w15696 <= not w15685 and not w15695;
w15697 <= not pi0644 and w15696;
w15698 <= not pi0618 and w15629;
w15699 <= pi0749 and w14843;
w15700 <= not w15632 and not w15699;
w15701 <= pi0038 and not w15700;
w15702 <= not pi0749 and w14609;
w15703 <= pi0141 and w14836;
w15704 <= not w15702 and not w15703;
w15705 <= pi0039 and not w15704;
w15706 <= not pi0141 and w14784;
w15707 <= pi0141 and w14797;
w15708 <= pi0749 and not w15707;
w15709 <= not w15706 and w15708;
w15710 <= not pi0039 and w14521;
w15711 <= not pi0141 and not pi0749;
w15712 <= not w15710 and w15711;
w15713 <= not w15709 and not w15712;
w15714 <= not pi0038 and not w15713;
w15715 <= not w15705 and w15714;
w15716 <= not w15701 and not w15715;
w15717 <= w134 and w15716;
w15718 <= not w15631 and not w15717;
w15719 <= not w14680 and not w15718;
w15720 <= w14680 and not w15629;
w15721 <= not w15719 and not w15720;
w15722 <= not pi0785 and not w15721;
w15723 <= not w14854 and not w15629;
w15724 <= pi0609 and w15719;
w15725 <= not w15723 and not w15724;
w15726 <= pi1155 and not w15725;
w15727 <= not w14859 and not w15629;
w15728 <= not pi0609 and w15719;
w15729 <= not w15727 and not w15728;
w15730 <= not pi1155 and not w15729;
w15731 <= not w15726 and not w15730;
w15732 <= pi0785 and not w15731;
w15733 <= not w15722 and not w15732;
w15734 <= pi0618 and w15733;
w15735 <= pi1154 and not w15698;
w15736 <= not w15734 and w15735;
w15737 <= not pi0706 and not w15716;
w15738 <= not pi0039 and w15208;
w15739 <= pi0038 and not w15738;
w15740 <= w15700 and w15739;
w15741 <= not pi0141 and not w15192;
w15742 <= pi0141 and not w15194;
w15743 <= pi0749 and not w15742;
w15744 <= not w15741 and w15743;
w15745 <= not pi0141 and w15175;
w15746 <= pi0141 and w15188;
w15747 <= not pi0749 and not w15745;
w15748 <= not w15746 and w15747;
w15749 <= not pi0039 and not w15744;
w15750 <= not w15748 and w15749;
w15751 <= pi0141 and w15168;
w15752 <= not pi0141 and not w15109;
w15753 <= pi0749 and not w15752;
w15754 <= not w15751 and w15753;
w15755 <= not pi0141 and w14967;
w15756 <= pi0141 and w15048;
w15757 <= not pi0749 and not w15756;
w15758 <= not w15755 and w15757;
w15759 <= pi0039 and not w15754;
w15760 <= not w15758 and w15759;
w15761 <= not pi0038 and not w15750;
w15762 <= not w15760 and w15761;
w15763 <= pi0706 and not w15740;
w15764 <= not w15762 and w15763;
w15765 <= w134 and not w15737;
w15766 <= not w15764 and w15765;
w15767 <= not w15631 and not w15766;
w15768 <= not pi0625 and w15767;
w15769 <= pi0625 and w15718;
w15770 <= not pi1153 and not w15769;
w15771 <= not w15768 and w15770;
w15772 <= not pi0608 and not w15654;
w15773 <= not w15771 and w15772;
w15774 <= not pi0625 and w15718;
w15775 <= pi0625 and w15767;
w15776 <= pi1153 and not w15774;
w15777 <= not w15775 and w15776;
w15778 <= pi0608 and not w15658;
w15779 <= not w15777 and w15778;
w15780 <= not w15773 and not w15779;
w15781 <= pi0778 and not w15780;
w15782 <= not pi0778 and w15767;
w15783 <= not w15781 and not w15782;
w15784 <= not pi0609 and not w15783;
w15785 <= pi0609 and w15661;
w15786 <= not pi1155 and not w15785;
w15787 <= not w15784 and w15786;
w15788 <= not pi0660 and not w15726;
w15789 <= not w15787 and w15788;
w15790 <= not pi0609 and w15661;
w15791 <= pi0609 and not w15783;
w15792 <= pi1155 and not w15790;
w15793 <= not w15791 and w15792;
w15794 <= pi0660 and not w15730;
w15795 <= not w15793 and w15794;
w15796 <= not w15789 and not w15795;
w15797 <= pi0785 and not w15796;
w15798 <= not pi0785 and not w15783;
w15799 <= not w15797 and not w15798;
w15800 <= not pi0618 and not w15799;
w15801 <= pi0618 and w15664;
w15802 <= not pi1154 and not w15801;
w15803 <= not w15800 and w15802;
w15804 <= not pi0627 and not w15736;
w15805 <= not w15803 and w15804;
w15806 <= not pi0618 and w15733;
w15807 <= pi0618 and w15629;
w15808 <= not pi1154 and not w15807;
w15809 <= not w15806 and w15808;
w15810 <= not pi0618 and w15664;
w15811 <= pi0618 and not w15799;
w15812 <= pi1154 and not w15810;
w15813 <= not w15811 and w15812;
w15814 <= pi0627 and not w15809;
w15815 <= not w15813 and w15814;
w15816 <= not w15805 and not w15815;
w15817 <= pi0781 and not w15816;
w15818 <= not pi0781 and not w15799;
w15819 <= not w15817 and not w15818;
w15820 <= not pi0619 and not w15819;
w15821 <= pi0619 and not w15667;
w15822 <= not pi1159 and not w15821;
w15823 <= not w15820 and w15822;
w15824 <= not pi0619 and w15629;
w15825 <= not pi0781 and not w15733;
w15826 <= not w15736 and not w15809;
w15827 <= pi0781 and not w15826;
w15828 <= not w15825 and not w15827;
w15829 <= pi0619 and w15828;
w15830 <= pi1159 and not w15824;
w15831 <= not w15829 and w15830;
w15832 <= not pi0648 and not w15831;
w15833 <= not w15823 and w15832;
w15834 <= pi0619 and not w15819;
w15835 <= not pi0619 and not w15667;
w15836 <= pi1159 and not w15835;
w15837 <= not w15834 and w15836;
w15838 <= not pi0619 and w15828;
w15839 <= pi0619 and w15629;
w15840 <= not pi1159 and not w15839;
w15841 <= not w15838 and w15840;
w15842 <= pi0648 and not w15841;
w15843 <= not w15837 and w15842;
w15844 <= not w15833 and not w15843;
w15845 <= pi0789 and not w15844;
w15846 <= not pi0789 and not w15819;
w15847 <= not w15845 and not w15846;
w15848 <= not pi0788 and w15847;
w15849 <= not pi0626 and w15847;
w15850 <= pi0626 and not w15669;
w15851 <= not pi0641 and not w15850;
w15852 <= not w15849 and w15851;
w15853 <= not pi0789 and not w15828;
w15854 <= not w15831 and not w15841;
w15855 <= pi0789 and not w15854;
w15856 <= not w15853 and not w15855;
w15857 <= not pi0626 and w15856;
w15858 <= pi0626 and w15629;
w15859 <= not pi1158 and not w15858;
w15860 <= not w15857 and w15859;
w15861 <= not w15293 and not w15860;
w15862 <= not w15852 and not w15861;
w15863 <= pi0626 and w15847;
w15864 <= not pi0626 and not w15669;
w15865 <= pi0641 and not w15864;
w15866 <= not w15863 and w15865;
w15867 <= not pi0626 and w15629;
w15868 <= pi0626 and w15856;
w15869 <= pi1158 and not w15867;
w15870 <= not w15868 and w15869;
w15871 <= not w15308 and not w15870;
w15872 <= not w15866 and not w15871;
w15873 <= not w15862 and not w15872;
w15874 <= pi0788 and not w15873;
w15875 <= not w15848 and not w15874;
w15876 <= not pi0628 and w15875;
w15877 <= not w15860 and not w15870;
w15878 <= pi0788 and not w15877;
w15879 <= not pi0788 and not w15856;
w15880 <= not w15878 and not w15879;
w15881 <= pi0628 and w15880;
w15882 <= not pi1156 and not w15881;
w15883 <= not w15876 and w15882;
w15884 <= not pi0629 and not w15677;
w15885 <= not w15883 and w15884;
w15886 <= pi0628 and w15875;
w15887 <= not pi0628 and w15880;
w15888 <= pi1156 and not w15887;
w15889 <= not w15886 and w15888;
w15890 <= pi0629 and not w15681;
w15891 <= not w15889 and w15890;
w15892 <= not w15885 and not w15891;
w15893 <= pi0792 and not w15892;
w15894 <= not pi0792 and w15875;
w15895 <= not w15893 and not w15894;
w15896 <= not pi0647 and not w15895;
w15897 <= not w15342 and w15880;
w15898 <= w15342 and w15629;
w15899 <= not w15897 and not w15898;
w15900 <= pi0647 and not w15899;
w15901 <= not pi1157 and not w15900;
w15902 <= not w15896 and w15901;
w15903 <= not pi0630 and not w15689;
w15904 <= not w15902 and w15903;
w15905 <= pi0647 and not w15895;
w15906 <= not pi0647 and not w15899;
w15907 <= pi1157 and not w15906;
w15908 <= not w15905 and w15907;
w15909 <= pi0630 and not w15693;
w15910 <= not w15908 and w15909;
w15911 <= not w15904 and not w15910;
w15912 <= pi0787 and not w15911;
w15913 <= not pi0787 and not w15895;
w15914 <= not w15912 and not w15913;
w15915 <= pi0644 and not w15914;
w15916 <= pi0715 and not w15697;
w15917 <= not w15915 and w15916;
w15918 <= w15367 and not w15629;
w15919 <= not w15367 and w15899;
w15920 <= not w15918 and not w15919;
w15921 <= pi0644 and w15920;
w15922 <= not pi0644 and w15629;
w15923 <= not pi0715 and not w15922;
w15924 <= not w15921 and w15923;
w15925 <= pi1160 and not w15924;
w15926 <= not w15917 and w15925;
w15927 <= not pi0644 and not w15914;
w15928 <= pi0644 and w15696;
w15929 <= not pi0715 and not w15928;
w15930 <= not w15927 and w15929;
w15931 <= not pi0644 and w15920;
w15932 <= pi0644 and w15629;
w15933 <= pi0715 and not w15932;
w15934 <= not w15931 and w15933;
w15935 <= not pi1160 and not w15934;
w15936 <= not w15930 and w15935;
w15937 <= pi0790 and not w15926;
w15938 <= not w15936 and w15937;
w15939 <= not pi0790 and w15914;
w15940 <= w4989 and not w15939;
w15941 <= not w15938 and w15940;
w15942 <= not pi0141 and not w4989;
w15943 <= not pi0832 and not w15942;
w15944 <= not w15941 and w15943;
w15945 <= not pi0141 and not w489;
w15946 <= not pi0647 and w15945;
w15947 <= pi0706 and w14208;
w15948 <= not w15945 and not w15947;
w15949 <= not pi0778 and w15948;
w15950 <= not pi0625 and w15947;
w15951 <= not w15948 and not w15950;
w15952 <= pi1153 and not w15951;
w15953 <= not pi1153 and not w15945;
w15954 <= not w15950 and w15953;
w15955 <= not w15952 and not w15954;
w15956 <= pi0778 and not w15955;
w15957 <= not w15949 and not w15956;
w15958 <= not w15408 and w15957;
w15959 <= not w15410 and w15958;
w15960 <= not w15412 and w15959;
w15961 <= not w15414 and w15960;
w15962 <= not w15420 and w15961;
w15963 <= pi0647 and w15962;
w15964 <= pi1157 and not w15946;
w15965 <= not w15963 and w15964;
w15966 <= not w15425 and w15961;
w15967 <= pi1156 and not w15966;
w15968 <= w15434 and w15960;
w15969 <= not pi0626 and w15945;
w15970 <= pi0749 and w14807;
w15971 <= not w15945 and not w15970;
w15972 <= not w15437 and not w15971;
w15973 <= not pi0785 and not w15972;
w15974 <= not w15442 and not w15971;
w15975 <= pi1155 and not w15974;
w15976 <= not w15445 and w15972;
w15977 <= not pi1155 and not w15976;
w15978 <= not w15975 and not w15977;
w15979 <= pi0785 and not w15978;
w15980 <= not w15973 and not w15979;
w15981 <= not pi0781 and not w15980;
w15982 <= not w15452 and w15980;
w15983 <= pi1154 and not w15982;
w15984 <= not w15455 and w15980;
w15985 <= not pi1154 and not w15984;
w15986 <= not w15983 and not w15985;
w15987 <= pi0781 and not w15986;
w15988 <= not w15981 and not w15987;
w15989 <= not pi0789 and not w15988;
w15990 <= not pi0619 and w15945;
w15991 <= pi0619 and w15988;
w15992 <= pi1159 and not w15990;
w15993 <= not w15991 and w15992;
w15994 <= not pi0619 and w15988;
w15995 <= pi0619 and w15945;
w15996 <= not pi1159 and not w15995;
w15997 <= not w15994 and w15996;
w15998 <= not w15993 and not w15997;
w15999 <= pi0789 and not w15998;
w16000 <= not w15989 and not w15999;
w16001 <= pi0626 and w16000;
w16002 <= pi1158 and not w15969;
w16003 <= not w16001 and w16002;
w16004 <= not pi0626 and w16000;
w16005 <= pi0626 and w15945;
w16006 <= not pi1158 and not w16005;
w16007 <= not w16004 and w16006;
w16008 <= not w16003 and not w16007;
w16009 <= not w14193 and w16008;
w16010 <= not w15968 and not w16009;
w16011 <= pi0788 and not w16010;
w16012 <= pi0618 and w15958;
w16013 <= pi0609 and w15957;
w16014 <= not w14731 and not w15948;
w16015 <= pi0625 and w16014;
w16016 <= w15971 and not w16014;
w16017 <= not w16015 and not w16016;
w16018 <= w15953 and not w16017;
w16019 <= not pi0608 and not w15952;
w16020 <= not w16018 and w16019;
w16021 <= pi1153 and w15971;
w16022 <= not w16015 and w16021;
w16023 <= pi0608 and not w15954;
w16024 <= not w16022 and w16023;
w16025 <= not w16020 and not w16024;
w16026 <= pi0778 and not w16025;
w16027 <= not pi0778 and not w16016;
w16028 <= not w16026 and not w16027;
w16029 <= not pi0609 and not w16028;
w16030 <= not pi1155 and not w16013;
w16031 <= not w16029 and w16030;
w16032 <= not pi0660 and not w15975;
w16033 <= not w16031 and w16032;
w16034 <= not pi0609 and w15957;
w16035 <= pi0609 and not w16028;
w16036 <= pi1155 and not w16034;
w16037 <= not w16035 and w16036;
w16038 <= pi0660 and not w15977;
w16039 <= not w16037 and w16038;
w16040 <= not w16033 and not w16039;
w16041 <= pi0785 and not w16040;
w16042 <= not pi0785 and not w16028;
w16043 <= not w16041 and not w16042;
w16044 <= not pi0618 and not w16043;
w16045 <= not pi1154 and not w16012;
w16046 <= not w16044 and w16045;
w16047 <= not pi0627 and not w15983;
w16048 <= not w16046 and w16047;
w16049 <= not pi0618 and w15958;
w16050 <= pi0618 and not w16043;
w16051 <= pi1154 and not w16049;
w16052 <= not w16050 and w16051;
w16053 <= pi0627 and not w15985;
w16054 <= not w16052 and w16053;
w16055 <= not w16048 and not w16054;
w16056 <= pi0781 and not w16055;
w16057 <= not pi0781 and not w16043;
w16058 <= not w16056 and not w16057;
w16059 <= not pi0789 and w16058;
w16060 <= not pi0619 and not w16058;
w16061 <= pi0619 and w15959;
w16062 <= not pi1159 and not w16061;
w16063 <= not w16060 and w16062;
w16064 <= not pi0648 and not w15993;
w16065 <= not w16063 and w16064;
w16066 <= not pi0619 and w15959;
w16067 <= pi0619 and not w16058;
w16068 <= pi1159 and not w16066;
w16069 <= not w16067 and w16068;
w16070 <= pi0648 and not w15997;
w16071 <= not w16069 and w16070;
w16072 <= pi0789 and not w16065;
w16073 <= not w16071 and w16072;
w16074 <= w15533 and not w16059;
w16075 <= not w16073 and w16074;
w16076 <= not w16011 and not w16075;
w16077 <= not pi0628 and not w16076;
w16078 <= not pi0788 and not w16000;
w16079 <= pi0788 and not w16008;
w16080 <= not w16078 and not w16079;
w16081 <= pi0628 and w16080;
w16082 <= not pi1156 and not w16081;
w16083 <= not w16077 and w16082;
w16084 <= not pi0629 and not w15967;
w16085 <= not w16083 and w16084;
w16086 <= not w15560 and w15961;
w16087 <= not pi1156 and not w16086;
w16088 <= not pi0628 and w16080;
w16089 <= pi0628 and not w16076;
w16090 <= pi1156 and not w16088;
w16091 <= not w16089 and w16090;
w16092 <= pi0629 and not w16087;
w16093 <= not w16091 and w16092;
w16094 <= not w16085 and not w16093;
w16095 <= pi0792 and not w16094;
w16096 <= not pi0792 and not w16076;
w16097 <= not w16095 and not w16096;
w16098 <= not pi0647 and not w16097;
w16099 <= not w15342 and w16080;
w16100 <= w15342 and w15945;
w16101 <= not w16099 and not w16100;
w16102 <= pi0647 and not w16101;
w16103 <= not pi1157 and not w16102;
w16104 <= not w16098 and w16103;
w16105 <= not pi0630 and not w15965;
w16106 <= not w16104 and w16105;
w16107 <= not pi0647 and w15962;
w16108 <= pi0647 and w15945;
w16109 <= not pi1157 and not w16108;
w16110 <= not w16107 and w16109;
w16111 <= pi0647 and not w16097;
w16112 <= not pi0647 and not w16101;
w16113 <= pi1157 and not w16112;
w16114 <= not w16111 and w16113;
w16115 <= pi0630 and not w16110;
w16116 <= not w16114 and w16115;
w16117 <= not w16106 and not w16116;
w16118 <= pi0787 and not w16117;
w16119 <= not pi0787 and not w16097;
w16120 <= not w16118 and not w16119;
w16121 <= not pi0790 and not w16120;
w16122 <= not pi0787 and not w15962;
w16123 <= not w15965 and not w16110;
w16124 <= pi0787 and not w16123;
w16125 <= not w16122 and not w16124;
w16126 <= not pi0644 and w16125;
w16127 <= pi0644 and not w16120;
w16128 <= pi0715 and not w16126;
w16129 <= not w16127 and w16128;
w16130 <= w15367 and not w15945;
w16131 <= not w15367 and w16101;
w16132 <= not w16130 and not w16131;
w16133 <= pi0644 and w16132;
w16134 <= not pi0644 and w15945;
w16135 <= not pi0715 and not w16134;
w16136 <= not w16133 and w16135;
w16137 <= pi1160 and not w16136;
w16138 <= not w16129 and w16137;
w16139 <= not pi0644 and w16132;
w16140 <= pi0644 and w15945;
w16141 <= pi0715 and not w16140;
w16142 <= not w16139 and w16141;
w16143 <= pi0644 and w16125;
w16144 <= not pi0644 and not w16120;
w16145 <= not pi0715 and not w16143;
w16146 <= not w16144 and w16145;
w16147 <= not pi1160 and not w16142;
w16148 <= not w16146 and w16147;
w16149 <= not w16138 and not w16148;
w16150 <= pi0790 and not w16149;
w16151 <= pi0832 and not w16121;
w16152 <= not w16150 and w16151;
w16153 <= not w15944 and not w16152;
w16154 <= w134 and not w14614;
w16155 <= pi0142 and not w16154;
w16156 <= pi0039 and not w14588;
w16157 <= pi0142 and not w15710;
w16158 <= not w16156 and w16157;
w16159 <= pi0142 and not w14533;
w16160 <= not w3805 and not w16159;
w16161 <= pi0142 and not w14553;
w16162 <= w3805 and not w16161;
w16163 <= pi0215 and not w16162;
w16164 <= not w16160 and w16163;
w16165 <= pi0142 and not w14216;
w16166 <= w1011 and not w16165;
w16167 <= pi0142 and not w14581;
w16168 <= not w3805 and not w16167;
w16169 <= pi0142 and not w14574;
w16170 <= w3805 and not w16169;
w16171 <= not w16168 and not w16170;
w16172 <= not w1011 and not w16171;
w16173 <= not pi0215 and not w16166;
w16174 <= not w16172 and w16173;
w16175 <= not w16164 and not w16174;
w16176 <= pi0039 and pi0299;
w16177 <= not w16175 and w16176;
w16178 <= not w16158 and not w16177;
w16179 <= w12436 and not w16178;
w16180 <= not w16155 and not w16179;
w16181 <= w14202 and not w16180;
w16182 <= pi0142 and not w134;
w16183 <= pi0039 and pi0142;
w16184 <= pi0038 and not w16183;
w16185 <= pi0142 and not w14230;
w16186 <= pi0735 and w14208;
w16187 <= w84 and w16186;
w16188 <= not w16185 and not w16187;
w16189 <= not pi0039 and not w16188;
w16190 <= w16184 and not w16189;
w16191 <= not pi0142 and not w14489;
w16192 <= pi0142 and w14511;
w16193 <= pi0735 and not w16191;
w16194 <= not w16192 and w16193;
w16195 <= pi0142 and not pi0735;
w16196 <= not w14521 and w16195;
w16197 <= not w16194 and not w16196;
w16198 <= not pi0039 and not w16197;
w16199 <= w14215 and w16186;
w16200 <= not w16165 and not w16199;
w16201 <= w1011 and w16200;
w16202 <= not pi0142 and not w14257;
w16203 <= pi0142 and not w14354;
w16204 <= not w16202 and not w16203;
w16205 <= pi0735 and not w16204;
w16206 <= not pi0735 and not w16169;
w16207 <= not w16205 and not w16206;
w16208 <= w3805 and w16207;
w16209 <= not pi0142 and w14268;
w16210 <= pi0142 and w14326;
w16211 <= not w16209 and not w16210;
w16212 <= pi0735 and not w16211;
w16213 <= not pi0735 and not w16167;
w16214 <= not w16212 and not w16213;
w16215 <= not w3805 and w16214;
w16216 <= not w1011 and not w16215;
w16217 <= not w16208 and w16216;
w16218 <= not pi0215 and not w16201;
w16219 <= not w16217 and w16218;
w16220 <= not pi0735 and not w16161;
w16221 <= not pi0142 and w15123;
w16222 <= pi0142 and not w14374;
w16223 <= pi0735 and not w16221;
w16224 <= not w16222 and w16223;
w16225 <= not w16220 and not w16224;
w16226 <= w3805 and not w16225;
w16227 <= not pi0735 and not w16159;
w16228 <= pi0142 and not w14382;
w16229 <= w15122 and w16221;
w16230 <= pi0735 and not w16229;
w16231 <= not w16228 and w16230;
w16232 <= not w16227 and not w16231;
w16233 <= not w3805 and not w16232;
w16234 <= pi0215 and not w16226;
w16235 <= not w16233 and w16234;
w16236 <= pi0299 and not w16235;
w16237 <= not w16219 and w16236;
w16238 <= w3768 and not w16225;
w16239 <= not w3768 and not w16232;
w16240 <= pi0223 and not w16238;
w16241 <= not w16239 and w16240;
w16242 <= w166 and w16200;
w16243 <= w3768 and w16207;
w16244 <= not w3768 and w16214;
w16245 <= not w166 and not w16244;
w16246 <= not w16243 and w16245;
w16247 <= not pi0223 and not w16242;
w16248 <= not w16246 and w16247;
w16249 <= not pi0299 and not w16241;
w16250 <= not w16248 and w16249;
w16251 <= pi0039 and not w16237;
w16252 <= not w16250 and w16251;
w16253 <= not pi0038 and not w16198;
w16254 <= not w16252 and w16253;
w16255 <= w134 and not w16190;
w16256 <= not w16254 and w16255;
w16257 <= not w16182 and not w16256;
w16258 <= not pi0778 and not w16257;
w16259 <= not pi0625 and w16257;
w16260 <= pi0625 and w16180;
w16261 <= not pi1153 and not w16260;
w16262 <= not w16259 and w16261;
w16263 <= not pi0625 and w16180;
w16264 <= pi0625 and w16257;
w16265 <= pi1153 and not w16263;
w16266 <= not w16264 and w16265;
w16267 <= not w16262 and not w16266;
w16268 <= pi0778 and not w16267;
w16269 <= not w16258 and not w16268;
w16270 <= not w14638 and w16269;
w16271 <= w14638 and w16180;
w16272 <= not w16270 and not w16271;
w16273 <= not w14202 and w16272;
w16274 <= not w16181 and not w16273;
w16275 <= not w14198 and w16274;
w16276 <= w14198 and w16180;
w16277 <= not w16275 and not w16276;
w16278 <= not w14194 and not w16277;
w16279 <= w14194 and w16180;
w16280 <= not w16278 and not w16279;
w16281 <= not pi0792 and w16280;
w16282 <= not pi0628 and w16180;
w16283 <= pi0628 and not w16280;
w16284 <= pi1156 and not w16282;
w16285 <= not w16283 and w16284;
w16286 <= pi0628 and w16180;
w16287 <= not pi0628 and not w16280;
w16288 <= not pi1156 and not w16286;
w16289 <= not w16287 and w16288;
w16290 <= not w16285 and not w16289;
w16291 <= pi0792 and not w16290;
w16292 <= not w16281 and not w16291;
w16293 <= not pi0787 and not w16292;
w16294 <= not pi0647 and w16180;
w16295 <= pi0647 and w16292;
w16296 <= pi1157 and not w16294;
w16297 <= not w16295 and w16296;
w16298 <= not pi0647 and w16292;
w16299 <= pi0647 and w16180;
w16300 <= not pi1157 and not w16299;
w16301 <= not w16298 and w16300;
w16302 <= not w16297 and not w16301;
w16303 <= pi0787 and not w16302;
w16304 <= not w16293 and not w16303;
w16305 <= not pi0644 and w16304;
w16306 <= not pi0618 and w16180;
w16307 <= pi0743 and w14807;
w16308 <= w84 and w16307;
w16309 <= not w16185 and not w16308;
w16310 <= not pi0039 and not w16309;
w16311 <= w16184 and not w16310;
w16312 <= pi0142 and not pi0743;
w16313 <= not w14493 and w16312;
w16314 <= not pi0142 and not w14789;
w16315 <= pi0142 and not w14700;
w16316 <= pi0743 and not w16314;
w16317 <= not w16315 and w16316;
w16318 <= not pi0299 and not w16313;
w16319 <= not w16317 and w16318;
w16320 <= not pi0142 and not w14794;
w16321 <= pi0142 and not w14504;
w16322 <= not pi0743 and not w16321;
w16323 <= pi0142 and w14687;
w16324 <= not w16320 and not w16322;
w16325 <= not w16323 and w16324;
w16326 <= pi0299 and not w16325;
w16327 <= not w16319 and not w16326;
w16328 <= not pi0039 and w16327;
w16329 <= not pi0743 and not w16159;
w16330 <= pi0142 and not w14752;
w16331 <= pi0743 and w15121;
w16332 <= not w16330 and w16331;
w16333 <= not w16329 and not w16332;
w16334 <= not w3768 and not w16333;
w16335 <= not pi0743 and not w16161;
w16336 <= pi0142 and w14763;
w16337 <= pi0743 and w14804;
w16338 <= not w16336 and w16337;
w16339 <= not w16335 and not w16338;
w16340 <= w3768 and not w16339;
w16341 <= pi0223 and not w16340;
w16342 <= not w16334 and w16341;
w16343 <= not pi0743 and not w16167;
w16344 <= pi0142 and not w14720;
w16345 <= pi0743 and not w14817;
w16346 <= not w16344 and w16345;
w16347 <= not w16343 and not w16346;
w16348 <= not w3768 and w16347;
w16349 <= not pi0142 and w14815;
w16350 <= pi0142 and w14738;
w16351 <= not w16349 and not w16350;
w16352 <= pi0743 and not w16351;
w16353 <= not pi0743 and not w16169;
w16354 <= not w16352 and not w16353;
w16355 <= w3768 and w16354;
w16356 <= not w166 and not w16348;
w16357 <= not w16355 and w16356;
w16358 <= pi0743 and w14798;
w16359 <= not w16165 and not w16358;
w16360 <= w166 and w16359;
w16361 <= not pi0223 and not w16360;
w16362 <= not w16357 and w16361;
w16363 <= not pi0299 and not w16342;
w16364 <= not w16362 and w16363;
w16365 <= w1011 and not w16359;
w16366 <= not w3805 and w16347;
w16367 <= w3805 and w16354;
w16368 <= not w16366 and not w16367;
w16369 <= not w1011 and not w16368;
w16370 <= not pi0215 and not w16365;
w16371 <= not w16369 and w16370;
w16372 <= not w3805 and w16333;
w16373 <= w3805 and w16339;
w16374 <= pi0215 and not w16373;
w16375 <= not w16372 and w16374;
w16376 <= not w16371 and not w16375;
w16377 <= pi0299 and not w16376;
w16378 <= pi0039 and not w16364;
w16379 <= not w16377 and w16378;
w16380 <= not pi0038 and not w16328;
w16381 <= not w16379 and w16380;
w16382 <= w134 and not w16311;
w16383 <= not w16381 and w16382;
w16384 <= not w16182 and not w16383;
w16385 <= not w14680 and not w16384;
w16386 <= w14680 and not w16180;
w16387 <= not w16385 and not w16386;
w16388 <= not pi0785 and not w16387;
w16389 <= not w14854 and not w16180;
w16390 <= pi0609 and w16385;
w16391 <= not w16389 and not w16390;
w16392 <= pi1155 and not w16391;
w16393 <= not w14859 and not w16180;
w16394 <= not pi0609 and w16385;
w16395 <= not w16393 and not w16394;
w16396 <= not pi1155 and not w16395;
w16397 <= not w16392 and not w16396;
w16398 <= pi0785 and not w16397;
w16399 <= not w16388 and not w16398;
w16400 <= pi0618 and w16399;
w16401 <= pi1154 and not w16306;
w16402 <= not w16400 and w16401;
w16403 <= pi0609 and w16269;
w16404 <= not pi0625 and w16384;
w16405 <= not pi0735 and w16327;
w16406 <= w14500 and w16315;
w16407 <= not w14482 and w16314;
w16408 <= not w16406 and not w16407;
w16409 <= pi0743 and not w16408;
w16410 <= pi0142 and not w14500;
w16411 <= not w14789 and w16410;
w16412 <= not pi0142 and w15181;
w16413 <= not pi0743 and not w16411;
w16414 <= not w16412 and w16413;
w16415 <= not pi0299 and not w16414;
w16416 <= not w16409 and w16415;
w16417 <= not w14487 and w16320;
w16418 <= not w14508 and w16323;
w16419 <= not w16417 and not w16418;
w16420 <= pi0743 and not w16419;
w16421 <= not pi0142 and w15186;
w16422 <= pi0142 and not w14509;
w16423 <= not w14794 and w16422;
w16424 <= not pi0743 and not w16423;
w16425 <= not w16421 and w16424;
w16426 <= pi0299 and not w16420;
w16427 <= not w16425 and w16426;
w16428 <= not w16416 and not w16427;
w16429 <= pi0735 and not w16428;
w16430 <= not pi0039 and not w16405;
w16431 <= not w16429 and w16430;
w16432 <= not pi0142 and not w15119;
w16433 <= pi0142 and not w15082;
w16434 <= pi0743 and not w16432;
w16435 <= not w16433 and w16434;
w16436 <= not pi0142 and w15011;
w16437 <= pi0142 and w14914;
w16438 <= not pi0743 and not w16436;
w16439 <= not w16437 and w16438;
w16440 <= not w16435 and not w16439;
w16441 <= pi0735 and not w16440;
w16442 <= not pi0735 and w16339;
w16443 <= not w16441 and not w16442;
w16444 <= w3768 and w16443;
w16445 <= not pi0142 and w15125;
w16446 <= pi0142 and w15090;
w16447 <= pi0743 and not w16445;
w16448 <= not w16446 and w16447;
w16449 <= not pi0142 and not w15026;
w16450 <= pi0142 and w14896;
w16451 <= not pi0743 and not w16450;
w16452 <= not w16449 and w16451;
w16453 <= not w16448 and not w16452;
w16454 <= pi0735 and not w16453;
w16455 <= not pi0735 and w16333;
w16456 <= not w16454 and not w16455;
w16457 <= not w3768 and w16456;
w16458 <= pi0223 and not w16444;
w16459 <= not w16457 and w16458;
w16460 <= not pi0735 and w16359;
w16461 <= not w15208 and w16309;
w16462 <= not w14213 and not w16461;
w16463 <= pi0735 and not w16462;
w16464 <= not w16165 and w16463;
w16465 <= not w16460 and not w16464;
w16466 <= w166 and not w16465;
w16467 <= pi0142 and w15073;
w16468 <= not pi0142 and not w15136;
w16469 <= pi0743 and not w16467;
w16470 <= not w16468 and w16469;
w16471 <= not pi0142 and w14983;
w16472 <= pi0142 and w14936;
w16473 <= not pi0743 and not w16471;
w16474 <= not w16472 and w16473;
w16475 <= not w16470 and not w16474;
w16476 <= pi0735 and not w16475;
w16477 <= not pi0735 and w16354;
w16478 <= not w16476 and not w16477;
w16479 <= w3768 and not w16478;
w16480 <= not pi0142 and not w15147;
w16481 <= pi0142 and w15062;
w16482 <= pi0743 and not w16481;
w16483 <= not w16480 and w16482;
w16484 <= not pi0142 and not w15001;
w16485 <= pi0142 and w14946;
w16486 <= not pi0743 and not w16485;
w16487 <= not w16484 and w16486;
w16488 <= not w16483 and not w16487;
w16489 <= pi0735 and not w16488;
w16490 <= not pi0735 and w16347;
w16491 <= not w16489 and not w16490;
w16492 <= not w3768 and not w16491;
w16493 <= not w166 and not w16492;
w16494 <= not w16479 and w16493;
w16495 <= not pi0223 and not w16466;
w16496 <= not w16494 and w16495;
w16497 <= not w16459 and not w16496;
w16498 <= not pi0299 and not w16497;
w16499 <= w3805 and w16443;
w16500 <= not w3805 and w16456;
w16501 <= pi0215 and not w16499;
w16502 <= not w16500 and w16501;
w16503 <= w1011 and not w16465;
w16504 <= not w3805 and not w16491;
w16505 <= w3805 and not w16478;
w16506 <= not w1011 and not w16504;
w16507 <= not w16505 and w16506;
w16508 <= not pi0215 and not w16503;
w16509 <= not w16507 and w16508;
w16510 <= not w16502 and not w16509;
w16511 <= pi0299 and not w16510;
w16512 <= pi0039 and not w16498;
w16513 <= not w16511 and w16512;
w16514 <= not w16431 and not w16513;
w16515 <= not pi0038 and not w16514;
w16516 <= pi0735 and w15208;
w16517 <= w16309 and not w16516;
w16518 <= not pi0039 and not w16517;
w16519 <= w16184 and not w16518;
w16520 <= w134 and not w16519;
w16521 <= not w16515 and w16520;
w16522 <= not w16182 and not w16521;
w16523 <= pi0625 and w16522;
w16524 <= pi1153 and not w16404;
w16525 <= not w16523 and w16524;
w16526 <= pi0608 and not w16262;
w16527 <= not w16525 and w16526;
w16528 <= not pi0625 and w16522;
w16529 <= pi0625 and w16384;
w16530 <= not pi1153 and not w16529;
w16531 <= not w16528 and w16530;
w16532 <= not pi0608 and not w16266;
w16533 <= not w16531 and w16532;
w16534 <= not w16527 and not w16533;
w16535 <= pi0778 and not w16534;
w16536 <= not pi0778 and w16522;
w16537 <= not w16535 and not w16536;
w16538 <= not pi0609 and not w16537;
w16539 <= not pi1155 and not w16403;
w16540 <= not w16538 and w16539;
w16541 <= not pi0660 and not w16392;
w16542 <= not w16540 and w16541;
w16543 <= not pi0609 and w16269;
w16544 <= pi0609 and not w16537;
w16545 <= pi1155 and not w16543;
w16546 <= not w16544 and w16545;
w16547 <= pi0660 and not w16396;
w16548 <= not w16546 and w16547;
w16549 <= not w16542 and not w16548;
w16550 <= pi0785 and not w16549;
w16551 <= not pi0785 and not w16537;
w16552 <= not w16550 and not w16551;
w16553 <= not pi0618 and not w16552;
w16554 <= pi0618 and not w16272;
w16555 <= not pi1154 and not w16554;
w16556 <= not w16553 and w16555;
w16557 <= not pi0627 and not w16402;
w16558 <= not w16556 and w16557;
w16559 <= not pi0618 and w16399;
w16560 <= pi0618 and w16180;
w16561 <= not pi1154 and not w16560;
w16562 <= not w16559 and w16561;
w16563 <= pi0618 and not w16552;
w16564 <= not pi0618 and not w16272;
w16565 <= pi1154 and not w16564;
w16566 <= not w16563 and w16565;
w16567 <= pi0627 and not w16562;
w16568 <= not w16566 and w16567;
w16569 <= not w16558 and not w16568;
w16570 <= pi0781 and not w16569;
w16571 <= not pi0781 and not w16552;
w16572 <= not w16570 and not w16571;
w16573 <= not pi0619 and not w16572;
w16574 <= pi0619 and w16274;
w16575 <= not pi1159 and not w16574;
w16576 <= not w16573 and w16575;
w16577 <= not pi0619 and w16180;
w16578 <= not pi0781 and not w16399;
w16579 <= not w16402 and not w16562;
w16580 <= pi0781 and not w16579;
w16581 <= not w16578 and not w16580;
w16582 <= pi0619 and w16581;
w16583 <= pi1159 and not w16577;
w16584 <= not w16582 and w16583;
w16585 <= not pi0648 and not w16584;
w16586 <= not w16576 and w16585;
w16587 <= pi0619 and not w16572;
w16588 <= not pi0619 and w16274;
w16589 <= pi1159 and not w16588;
w16590 <= not w16587 and w16589;
w16591 <= not pi0619 and w16581;
w16592 <= pi0619 and w16180;
w16593 <= not pi1159 and not w16592;
w16594 <= not w16591 and w16593;
w16595 <= pi0648 and not w16594;
w16596 <= not w16590 and w16595;
w16597 <= not w16586 and not w16596;
w16598 <= pi0789 and not w16597;
w16599 <= not pi0789 and not w16572;
w16600 <= not w16598 and not w16599;
w16601 <= not pi0788 and w16600;
w16602 <= not pi0626 and w16600;
w16603 <= pi0626 and w16277;
w16604 <= not pi0641 and not w16603;
w16605 <= not w16602 and w16604;
w16606 <= not pi0789 and not w16581;
w16607 <= not w16584 and not w16594;
w16608 <= pi0789 and not w16607;
w16609 <= not w16606 and not w16608;
w16610 <= not pi0626 and w16609;
w16611 <= pi0626 and w16180;
w16612 <= not pi1158 and not w16611;
w16613 <= not w16610 and w16612;
w16614 <= not w15293 and not w16613;
w16615 <= not w16605 and not w16614;
w16616 <= pi0626 and w16600;
w16617 <= not pi0626 and w16277;
w16618 <= pi0641 and not w16617;
w16619 <= not w16616 and w16618;
w16620 <= not pi0626 and w16180;
w16621 <= pi0626 and w16609;
w16622 <= pi1158 and not w16620;
w16623 <= not w16621 and w16622;
w16624 <= not w15308 and not w16623;
w16625 <= not w16619 and not w16624;
w16626 <= not w16615 and not w16625;
w16627 <= pi0788 and not w16626;
w16628 <= not w16601 and not w16627;
w16629 <= not pi0628 and w16628;
w16630 <= not w16613 and not w16623;
w16631 <= pi0788 and not w16630;
w16632 <= not pi0788 and not w16609;
w16633 <= not w16631 and not w16632;
w16634 <= pi0628 and w16633;
w16635 <= not pi1156 and not w16634;
w16636 <= not w16629 and w16635;
w16637 <= not pi0629 and not w16285;
w16638 <= not w16636 and w16637;
w16639 <= pi0628 and w16628;
w16640 <= not pi0628 and w16633;
w16641 <= pi1156 and not w16640;
w16642 <= not w16639 and w16641;
w16643 <= pi0629 and not w16289;
w16644 <= not w16642 and w16643;
w16645 <= not w16638 and not w16644;
w16646 <= pi0792 and not w16645;
w16647 <= not pi0792 and w16628;
w16648 <= not w16646 and not w16647;
w16649 <= not pi0647 and not w16648;
w16650 <= not w15342 and w16633;
w16651 <= w15342 and w16180;
w16652 <= not w16650 and not w16651;
w16653 <= pi0647 and not w16652;
w16654 <= not pi1157 and not w16653;
w16655 <= not w16649 and w16654;
w16656 <= not pi0630 and not w16297;
w16657 <= not w16655 and w16656;
w16658 <= pi0647 and not w16648;
w16659 <= not pi0647 and not w16652;
w16660 <= pi1157 and not w16659;
w16661 <= not w16658 and w16660;
w16662 <= pi0630 and not w16301;
w16663 <= not w16661 and w16662;
w16664 <= not w16657 and not w16663;
w16665 <= pi0787 and not w16664;
w16666 <= not pi0787 and not w16648;
w16667 <= not w16665 and not w16666;
w16668 <= pi0644 and not w16667;
w16669 <= pi0715 and not w16305;
w16670 <= not w16668 and w16669;
w16671 <= w15367 and not w16180;
w16672 <= not w15367 and w16652;
w16673 <= not w16671 and not w16672;
w16674 <= pi0644 and w16673;
w16675 <= not pi0644 and w16180;
w16676 <= not pi0715 and not w16675;
w16677 <= not w16674 and w16676;
w16678 <= pi1160 and not w16677;
w16679 <= not w16670 and w16678;
w16680 <= not pi0644 and not w16667;
w16681 <= pi0644 and w16304;
w16682 <= not pi0715 and not w16681;
w16683 <= not w16680 and w16682;
w16684 <= not pi0644 and w16673;
w16685 <= pi0644 and w16180;
w16686 <= pi0715 and not w16685;
w16687 <= not w16684 and w16686;
w16688 <= not pi1160 and not w16687;
w16689 <= not w16683 and w16688;
w16690 <= pi0790 and not w16679;
w16691 <= not w16689 and w16690;
w16692 <= not pi0790 and w16667;
w16693 <= w3868 and not w16692;
w16694 <= not w16691 and w16693;
w16695 <= not pi0142 and not w3868;
w16696 <= not pi0057 and not w16695;
w16697 <= not w16694 and w16696;
w16698 <= pi0057 and pi0142;
w16699 <= not pi0832 and not w16698;
w16700 <= not w16697 and w16699;
w16701 <= pi0142 and not w489;
w16702 <= pi0628 and pi1156;
w16703 <= not pi0628 and not pi1156;
w16704 <= pi0792 and not w16702;
w16705 <= not w16703 and w16704;
w16706 <= not pi0625 and pi1153;
w16707 <= pi0625 and not pi1153;
w16708 <= not w16706 and not w16707;
w16709 <= pi0778 and not w16708;
w16710 <= w16186 and not w16709;
w16711 <= not w16701 and not w16710;
w16712 <= not w14194 and not w14198;
w16713 <= not w14202 and not w14638;
w16714 <= w16712 and w16713;
w16715 <= not w16711 and w16714;
w16716 <= not w16705 and w16715;
w16717 <= pi0647 and w16716;
w16718 <= pi1157 and not w16701;
w16719 <= not w16717 and w16718;
w16720 <= pi0628 and w16715;
w16721 <= not w16701 and not w16720;
w16722 <= pi1156 and not w16721;
w16723 <= not pi0626 and w16701;
w16724 <= not w14680 and w16307;
w16725 <= pi0609 and w16724;
w16726 <= pi1155 and not w16701;
w16727 <= not w16725 and w16726;
w16728 <= not pi0609 and w16724;
w16729 <= not pi1155 and not w16701;
w16730 <= not w16728 and w16729;
w16731 <= not w16727 and not w16730;
w16732 <= pi0785 and not w16731;
w16733 <= not pi0785 and not w16701;
w16734 <= not w16724 and w16733;
w16735 <= not w16732 and not w16734;
w16736 <= not pi0781 and not w16735;
w16737 <= not pi0618 and w16701;
w16738 <= pi0618 and w16735;
w16739 <= pi1154 and not w16737;
w16740 <= not w16738 and w16739;
w16741 <= not pi0618 and w16735;
w16742 <= pi0618 and w16701;
w16743 <= not pi1154 and not w16742;
w16744 <= not w16741 and w16743;
w16745 <= not w16740 and not w16744;
w16746 <= pi0781 and not w16745;
w16747 <= not w16736 and not w16746;
w16748 <= not pi0789 and not w16747;
w16749 <= not pi0619 and w16701;
w16750 <= pi0619 and w16747;
w16751 <= pi1159 and not w16749;
w16752 <= not w16750 and w16751;
w16753 <= not pi0619 and w16747;
w16754 <= pi0619 and w16701;
w16755 <= not pi1159 and not w16754;
w16756 <= not w16753 and w16755;
w16757 <= not w16752 and not w16756;
w16758 <= pi0789 and not w16757;
w16759 <= not w16748 and not w16758;
w16760 <= pi0626 and w16759;
w16761 <= pi1158 and not w16723;
w16762 <= not w16760 and w16761;
w16763 <= not pi0626 and w16759;
w16764 <= pi0626 and w16701;
w16765 <= not pi1158 and not w16764;
w16766 <= not w16763 and w16765;
w16767 <= not w16762 and not w16766;
w16768 <= not w14193 and w16767;
w16769 <= w14198 and not w16701;
w16770 <= not w14638 and not w16711;
w16771 <= not w14202 and w16770;
w16772 <= not w16701 and not w16771;
w16773 <= w15434 and not w16769;
w16774 <= not w16772 and w16773;
w16775 <= not w16768 and not w16774;
w16776 <= pi0788 and not w16775;
w16777 <= not w16701 and not w16770;
w16778 <= pi0618 and not w16777;
w16779 <= pi0625 and w16186;
w16780 <= pi1153 and not w16701;
w16781 <= not w16779 and w16780;
w16782 <= pi0735 and w15032;
w16783 <= pi0625 and w16782;
w16784 <= not w16307 and not w16701;
w16785 <= not w16782 and w16784;
w16786 <= not w16783 and not w16785;
w16787 <= not pi1153 and not w16786;
w16788 <= not pi0608 and not w16781;
w16789 <= not w16787 and w16788;
w16790 <= not w16307 and not w16783;
w16791 <= pi1153 and not w16790;
w16792 <= not pi0625 and not pi1153;
w16793 <= w16186 and w16792;
w16794 <= not w16701 and not w16793;
w16795 <= not w16791 and w16794;
w16796 <= pi0608 and not w16795;
w16797 <= not w16789 and not w16796;
w16798 <= pi0778 and not w16797;
w16799 <= not pi0778 and not w16785;
w16800 <= not w16798 and not w16799;
w16801 <= not pi0609 and not w16800;
w16802 <= pi0609 and not w16711;
w16803 <= not pi1155 and not w16802;
w16804 <= not w16801 and w16803;
w16805 <= not pi0660 and not w16727;
w16806 <= not w16804 and w16805;
w16807 <= pi0609 and not w16800;
w16808 <= not pi0609 and not w16711;
w16809 <= pi1155 and not w16808;
w16810 <= not w16807 and w16809;
w16811 <= pi0660 and not w16730;
w16812 <= not w16810 and w16811;
w16813 <= not w16806 and not w16812;
w16814 <= pi0785 and not w16813;
w16815 <= not pi0785 and not w16800;
w16816 <= not w16814 and not w16815;
w16817 <= not pi0618 and not w16816;
w16818 <= not pi1154 and not w16778;
w16819 <= not w16817 and w16818;
w16820 <= not pi0627 and not w16740;
w16821 <= not w16819 and w16820;
w16822 <= not pi0618 and not w16777;
w16823 <= pi0618 and not w16816;
w16824 <= pi1154 and not w16822;
w16825 <= not w16823 and w16824;
w16826 <= pi0627 and not w16744;
w16827 <= not w16825 and w16826;
w16828 <= not w16821 and not w16827;
w16829 <= pi0781 and not w16828;
w16830 <= not pi0781 and not w16816;
w16831 <= not w16829 and not w16830;
w16832 <= not pi0789 and w16831;
w16833 <= not pi0619 and not w16831;
w16834 <= pi0619 and not w16772;
w16835 <= not pi1159 and not w16834;
w16836 <= not w16833 and w16835;
w16837 <= not pi0648 and not w16752;
w16838 <= not w16836 and w16837;
w16839 <= pi0619 and not w16831;
w16840 <= not pi0619 and not w16772;
w16841 <= pi1159 and not w16840;
w16842 <= not w16839 and w16841;
w16843 <= pi0648 and not w16756;
w16844 <= not w16842 and w16843;
w16845 <= pi0789 and not w16838;
w16846 <= not w16844 and w16845;
w16847 <= w15533 and not w16832;
w16848 <= not w16846 and w16847;
w16849 <= not w16776 and not w16848;
w16850 <= not pi0628 and w16849;
w16851 <= not pi0788 and not w16759;
w16852 <= pi0788 and not w16767;
w16853 <= not w16851 and not w16852;
w16854 <= pi0628 and not w16853;
w16855 <= not pi1156 and not w16854;
w16856 <= not w16850 and w16855;
w16857 <= not pi0629 and not w16722;
w16858 <= not w16856 and w16857;
w16859 <= not pi0628 and w16715;
w16860 <= not w16701 and not w16859;
w16861 <= not pi1156 and not w16860;
w16862 <= pi0628 and w16849;
w16863 <= not pi0628 and not w16853;
w16864 <= pi1156 and not w16863;
w16865 <= not w16862 and w16864;
w16866 <= pi0629 and not w16861;
w16867 <= not w16865 and w16866;
w16868 <= not w16858 and not w16867;
w16869 <= pi0792 and not w16868;
w16870 <= not pi0792 and w16849;
w16871 <= not w16869 and not w16870;
w16872 <= not pi0647 and w16871;
w16873 <= not w15342 and w16853;
w16874 <= w15342 and w16701;
w16875 <= not w16873 and not w16874;
w16876 <= pi0647 and not w16875;
w16877 <= not pi1157 and not w16876;
w16878 <= not w16872 and w16877;
w16879 <= not pi0630 and not w16719;
w16880 <= not w16878 and w16879;
w16881 <= not pi0647 and w16716;
w16882 <= not pi1157 and not w16701;
w16883 <= not w16881 and w16882;
w16884 <= not pi0647 and not w16875;
w16885 <= pi0647 and w16871;
w16886 <= pi1157 and not w16884;
w16887 <= not w16885 and w16886;
w16888 <= pi0630 and not w16883;
w16889 <= not w16887 and w16888;
w16890 <= not w16880 and not w16889;
w16891 <= pi0787 and not w16890;
w16892 <= not pi0787 and w16871;
w16893 <= not w16891 and not w16892;
w16894 <= not pi0790 and not w16893;
w16895 <= w15367 and not w16701;
w16896 <= not w15367 and w16875;
w16897 <= not w16895 and not w16896;
w16898 <= pi0644 and w16897;
w16899 <= not pi0644 and w16701;
w16900 <= not pi0715 and not w16899;
w16901 <= not w16898 and w16900;
w16902 <= not pi0647 and pi1157;
w16903 <= pi0647 and not pi1157;
w16904 <= not w16902 and not w16903;
w16905 <= pi0787 and not w16904;
w16906 <= w16716 and not w16905;
w16907 <= not w16701 and not w16906;
w16908 <= not pi0644 and not w16907;
w16909 <= pi0644 and not w16893;
w16910 <= pi0715 and not w16908;
w16911 <= not w16909 and w16910;
w16912 <= pi1160 and not w16901;
w16913 <= not w16911 and w16912;
w16914 <= not pi0644 and w16897;
w16915 <= pi0644 and w16701;
w16916 <= pi0715 and not w16915;
w16917 <= not w16914 and w16916;
w16918 <= pi0644 and not w16907;
w16919 <= not pi0644 and not w16893;
w16920 <= not pi0715 and not w16918;
w16921 <= not w16919 and w16920;
w16922 <= not pi1160 and not w16917;
w16923 <= not w16921 and w16922;
w16924 <= not w16913 and not w16923;
w16925 <= pi0790 and not w16924;
w16926 <= pi0832 and not w16894;
w16927 <= not w16925 and w16926;
w16928 <= not w16700 and not w16927;
w16929 <= not pi0143 and not w14622;
w16930 <= w14198 and not w16929;
w16931 <= pi0143 and not w134;
w16932 <= not pi0143 and not w14615;
w16933 <= not pi0687 and w16932;
w16934 <= not pi0143 and not w14204;
w16935 <= w14210 and not w16934;
w16936 <= not pi0143 and w15635;
w16937 <= pi0143 and not w15639;
w16938 <= not pi0038 and not w16937;
w16939 <= not w16936 and w16938;
w16940 <= pi0687 and not w16935;
w16941 <= not w16939 and w16940;
w16942 <= w134 and not w16933;
w16943 <= not w16941 and w16942;
w16944 <= not w16931 and not w16943;
w16945 <= not pi0778 and not w16944;
w16946 <= not pi0625 and w16929;
w16947 <= pi0625 and w16944;
w16948 <= pi1153 and not w16946;
w16949 <= not w16947 and w16948;
w16950 <= not pi0625 and w16944;
w16951 <= pi0625 and w16929;
w16952 <= not pi1153 and not w16951;
w16953 <= not w16950 and w16952;
w16954 <= not w16949 and not w16953;
w16955 <= pi0778 and not w16954;
w16956 <= not w16945 and not w16955;
w16957 <= not w14638 and not w16956;
w16958 <= w14638 and not w16929;
w16959 <= not w16957 and not w16958;
w16960 <= not w14202 and w16959;
w16961 <= w14202 and w16929;
w16962 <= not w16960 and not w16961;
w16963 <= not w14198 and w16962;
w16964 <= not w16930 and not w16963;
w16965 <= not w14194 and w16964;
w16966 <= w14194 and w16929;
w16967 <= not w16965 and not w16966;
w16968 <= not pi0792 and w16967;
w16969 <= not pi0628 and w16929;
w16970 <= pi0628 and not w16967;
w16971 <= pi1156 and not w16969;
w16972 <= not w16970 and w16971;
w16973 <= pi0628 and w16929;
w16974 <= not pi0628 and not w16967;
w16975 <= not pi1156 and not w16973;
w16976 <= not w16974 and w16975;
w16977 <= not w16972 and not w16976;
w16978 <= pi0792 and not w16977;
w16979 <= not w16968 and not w16978;
w16980 <= not pi0787 and not w16979;
w16981 <= not pi0647 and w16929;
w16982 <= pi0647 and w16979;
w16983 <= pi1157 and not w16981;
w16984 <= not w16982 and w16983;
w16985 <= not pi0647 and w16979;
w16986 <= pi0647 and w16929;
w16987 <= not pi1157 and not w16986;
w16988 <= not w16985 and w16987;
w16989 <= not w16984 and not w16988;
w16990 <= pi0787 and not w16989;
w16991 <= not w16980 and not w16990;
w16992 <= not pi0644 and w16991;
w16993 <= not pi0618 and w16929;
w16994 <= pi0774 and not w16932;
w16995 <= w3698 and w14807;
w16996 <= pi0038 and w16995;
w16997 <= not pi0038 and w14838;
w16998 <= pi0143 and not w16997;
w16999 <= not pi0038 and not w14784;
w17000 <= w3847 and w14745;
w17001 <= pi0038 and not w17000;
w17002 <= not w16999 and not w17001;
w17003 <= not pi0143 and not pi0774;
w17004 <= w17002 and w17003;
w17005 <= not w16998 and not w17004;
w17006 <= not w16996 and not w17005;
w17007 <= not w16994 and not w17006;
w17008 <= w134 and not w17007;
w17009 <= not w16931 and not w17008;
w17010 <= not w14680 and not w17009;
w17011 <= w14680 and not w16929;
w17012 <= not w17010 and not w17011;
w17013 <= not pi0785 and not w17012;
w17014 <= not w14854 and not w16929;
w17015 <= pi0609 and w17010;
w17016 <= not w17014 and not w17015;
w17017 <= pi1155 and not w17016;
w17018 <= not w14859 and not w16929;
w17019 <= not pi0609 and w17010;
w17020 <= not w17018 and not w17019;
w17021 <= not pi1155 and not w17020;
w17022 <= not w17017 and not w17021;
w17023 <= pi0785 and not w17022;
w17024 <= not w17013 and not w17023;
w17025 <= pi0618 and w17024;
w17026 <= pi1154 and not w16993;
w17027 <= not w17025 and w17026;
w17028 <= not pi0039 and not w15188;
w17029 <= pi0039 and not w15048;
w17030 <= not w17028 and not w17029;
w17031 <= not pi0038 and w17030;
w17032 <= pi0143 and w17031;
w17033 <= pi0038 and w15738;
w17034 <= w14204 and not w14918;
w17035 <= pi0038 and w17034;
w17036 <= pi0039 and not w14967;
w17037 <= not pi0039 and not w15175;
w17038 <= not w17036 and not w17037;
w17039 <= not pi0038 and not w17038;
w17040 <= not w17035 and not w17039;
w17041 <= not pi0143 and w17040;
w17042 <= pi0774 and not w17033;
w17043 <= not w17032 and w17042;
w17044 <= not w17041 and w17043;
w17045 <= not pi0039 and not w15192;
w17046 <= not pi0038 and w17045;
w17047 <= pi0039 and not w15109;
w17048 <= not pi0039 and w15053;
w17049 <= pi0038 and not w17048;
w17050 <= not w17046 and not w17049;
w17051 <= not w17047 and w17050;
w17052 <= not pi0143 and not w17051;
w17053 <= w3847 and not w15033;
w17054 <= pi0038 and not w17053;
w17055 <= pi0039 and not w15168;
w17056 <= not w14489 and w14797;
w17057 <= not w17055 and not w17056;
w17058 <= not pi0038 and not w17057;
w17059 <= not w17054 and not w17058;
w17060 <= pi0143 and w17059;
w17061 <= not pi0774 and not w17052;
w17062 <= not w17060 and w17061;
w17063 <= pi0687 and not w17062;
w17064 <= not w17044 and w17063;
w17065 <= not pi0687 and w17007;
w17066 <= w134 and not w17064;
w17067 <= not w17065 and w17066;
w17068 <= not w16931 and not w17067;
w17069 <= not pi0625 and w17068;
w17070 <= pi0625 and w17009;
w17071 <= not pi1153 and not w17070;
w17072 <= not w17069 and w17071;
w17073 <= not pi0608 and not w16949;
w17074 <= not w17072 and w17073;
w17075 <= not pi0625 and w17009;
w17076 <= pi0625 and w17068;
w17077 <= pi1153 and not w17075;
w17078 <= not w17076 and w17077;
w17079 <= pi0608 and not w16953;
w17080 <= not w17078 and w17079;
w17081 <= not w17074 and not w17080;
w17082 <= pi0778 and not w17081;
w17083 <= not pi0778 and w17068;
w17084 <= not w17082 and not w17083;
w17085 <= not pi0609 and not w17084;
w17086 <= pi0609 and w16956;
w17087 <= not pi1155 and not w17086;
w17088 <= not w17085 and w17087;
w17089 <= not pi0660 and not w17017;
w17090 <= not w17088 and w17089;
w17091 <= not pi0609 and w16956;
w17092 <= pi0609 and not w17084;
w17093 <= pi1155 and not w17091;
w17094 <= not w17092 and w17093;
w17095 <= pi0660 and not w17021;
w17096 <= not w17094 and w17095;
w17097 <= not w17090 and not w17096;
w17098 <= pi0785 and not w17097;
w17099 <= not pi0785 and not w17084;
w17100 <= not w17098 and not w17099;
w17101 <= not pi0618 and not w17100;
w17102 <= pi0618 and w16959;
w17103 <= not pi1154 and not w17102;
w17104 <= not w17101 and w17103;
w17105 <= not pi0627 and not w17027;
w17106 <= not w17104 and w17105;
w17107 <= not pi0618 and w17024;
w17108 <= pi0618 and w16929;
w17109 <= not pi1154 and not w17108;
w17110 <= not w17107 and w17109;
w17111 <= not pi0618 and w16959;
w17112 <= pi0618 and not w17100;
w17113 <= pi1154 and not w17111;
w17114 <= not w17112 and w17113;
w17115 <= pi0627 and not w17110;
w17116 <= not w17114 and w17115;
w17117 <= not w17106 and not w17116;
w17118 <= pi0781 and not w17117;
w17119 <= not pi0781 and not w17100;
w17120 <= not w17118 and not w17119;
w17121 <= not pi0619 and not w17120;
w17122 <= pi0619 and not w16962;
w17123 <= not pi1159 and not w17122;
w17124 <= not w17121 and w17123;
w17125 <= not pi0619 and w16929;
w17126 <= not pi0781 and not w17024;
w17127 <= not w17027 and not w17110;
w17128 <= pi0781 and not w17127;
w17129 <= not w17126 and not w17128;
w17130 <= pi0619 and w17129;
w17131 <= pi1159 and not w17125;
w17132 <= not w17130 and w17131;
w17133 <= not pi0648 and not w17132;
w17134 <= not w17124 and w17133;
w17135 <= pi0619 and not w17120;
w17136 <= not pi0619 and not w16962;
w17137 <= pi1159 and not w17136;
w17138 <= not w17135 and w17137;
w17139 <= not pi0619 and w17129;
w17140 <= pi0619 and w16929;
w17141 <= not pi1159 and not w17140;
w17142 <= not w17139 and w17141;
w17143 <= pi0648 and not w17142;
w17144 <= not w17138 and w17143;
w17145 <= not w17134 and not w17144;
w17146 <= pi0789 and not w17145;
w17147 <= not pi0789 and not w17120;
w17148 <= not w17146 and not w17147;
w17149 <= not pi0788 and w17148;
w17150 <= not pi0626 and w17148;
w17151 <= pi0626 and not w16964;
w17152 <= not pi0641 and not w17151;
w17153 <= not w17150 and w17152;
w17154 <= not pi0789 and not w17129;
w17155 <= not w17132 and not w17142;
w17156 <= pi0789 and not w17155;
w17157 <= not w17154 and not w17156;
w17158 <= not pi0626 and w17157;
w17159 <= pi0626 and w16929;
w17160 <= not pi1158 and not w17159;
w17161 <= not w17158 and w17160;
w17162 <= not w15293 and not w17161;
w17163 <= not w17153 and not w17162;
w17164 <= pi0626 and w17148;
w17165 <= not pi0626 and not w16964;
w17166 <= pi0641 and not w17165;
w17167 <= not w17164 and w17166;
w17168 <= not pi0626 and w16929;
w17169 <= pi0626 and w17157;
w17170 <= pi1158 and not w17168;
w17171 <= not w17169 and w17170;
w17172 <= not w15308 and not w17171;
w17173 <= not w17167 and not w17172;
w17174 <= not w17163 and not w17173;
w17175 <= pi0788 and not w17174;
w17176 <= not w17149 and not w17175;
w17177 <= not pi0628 and w17176;
w17178 <= not w17161 and not w17171;
w17179 <= pi0788 and not w17178;
w17180 <= not pi0788 and not w17157;
w17181 <= not w17179 and not w17180;
w17182 <= pi0628 and w17181;
w17183 <= not pi1156 and not w17182;
w17184 <= not w17177 and w17183;
w17185 <= not pi0629 and not w16972;
w17186 <= not w17184 and w17185;
w17187 <= pi0628 and w17176;
w17188 <= not pi0628 and w17181;
w17189 <= pi1156 and not w17188;
w17190 <= not w17187 and w17189;
w17191 <= pi0629 and not w16976;
w17192 <= not w17190 and w17191;
w17193 <= not w17186 and not w17192;
w17194 <= pi0792 and not w17193;
w17195 <= not pi0792 and w17176;
w17196 <= not w17194 and not w17195;
w17197 <= not pi0647 and not w17196;
w17198 <= not w15342 and w17181;
w17199 <= w15342 and w16929;
w17200 <= not w17198 and not w17199;
w17201 <= pi0647 and not w17200;
w17202 <= not pi1157 and not w17201;
w17203 <= not w17197 and w17202;
w17204 <= not pi0630 and not w16984;
w17205 <= not w17203 and w17204;
w17206 <= pi0647 and not w17196;
w17207 <= not pi0647 and not w17200;
w17208 <= pi1157 and not w17207;
w17209 <= not w17206 and w17208;
w17210 <= pi0630 and not w16988;
w17211 <= not w17209 and w17210;
w17212 <= not w17205 and not w17211;
w17213 <= pi0787 and not w17212;
w17214 <= not pi0787 and not w17196;
w17215 <= not w17213 and not w17214;
w17216 <= pi0644 and not w17215;
w17217 <= pi0715 and not w16992;
w17218 <= not w17216 and w17217;
w17219 <= w15367 and not w16929;
w17220 <= not w15367 and w17200;
w17221 <= not w17219 and not w17220;
w17222 <= pi0644 and w17221;
w17223 <= not pi0644 and w16929;
w17224 <= not pi0715 and not w17223;
w17225 <= not w17222 and w17224;
w17226 <= pi1160 and not w17225;
w17227 <= not w17218 and w17226;
w17228 <= not pi0644 and not w17215;
w17229 <= pi0644 and w16991;
w17230 <= not pi0715 and not w17229;
w17231 <= not w17228 and w17230;
w17232 <= not pi0644 and w17221;
w17233 <= pi0644 and w16929;
w17234 <= pi0715 and not w17233;
w17235 <= not w17232 and w17234;
w17236 <= not pi1160 and not w17235;
w17237 <= not w17231 and w17236;
w17238 <= pi0790 and not w17227;
w17239 <= not w17237 and w17238;
w17240 <= not pi0790 and w17215;
w17241 <= w4989 and not w17240;
w17242 <= not w17239 and w17241;
w17243 <= not pi0143 and not w4989;
w17244 <= not pi0832 and not w17243;
w17245 <= not w17242 and w17244;
w17246 <= not pi0143 and not w489;
w17247 <= not pi0647 and w17246;
w17248 <= pi0687 and w14208;
w17249 <= not w17246 and not w17248;
w17250 <= not pi0778 and w17249;
w17251 <= not pi0625 and w17248;
w17252 <= not w17249 and not w17251;
w17253 <= pi1153 and not w17252;
w17254 <= not pi1153 and not w17246;
w17255 <= not w17251 and w17254;
w17256 <= not w17253 and not w17255;
w17257 <= pi0778 and not w17256;
w17258 <= not w17250 and not w17257;
w17259 <= not w15408 and w17258;
w17260 <= not w15410 and w17259;
w17261 <= not w15412 and w17260;
w17262 <= not w15414 and w17261;
w17263 <= not w15420 and w17262;
w17264 <= pi0647 and w17263;
w17265 <= pi1157 and not w17247;
w17266 <= not w17264 and w17265;
w17267 <= not w15425 and w17262;
w17268 <= pi1156 and not w17267;
w17269 <= w15434 and w17261;
w17270 <= not pi0626 and w17246;
w17271 <= not pi0774 and w14807;
w17272 <= not w17246 and not w17271;
w17273 <= not w15437 and not w17272;
w17274 <= not pi0785 and not w17273;
w17275 <= not w15442 and not w17272;
w17276 <= pi1155 and not w17275;
w17277 <= not w15445 and w17273;
w17278 <= not pi1155 and not w17277;
w17279 <= not w17276 and not w17278;
w17280 <= pi0785 and not w17279;
w17281 <= not w17274 and not w17280;
w17282 <= not pi0781 and not w17281;
w17283 <= not w15452 and w17281;
w17284 <= pi1154 and not w17283;
w17285 <= not w15455 and w17281;
w17286 <= not pi1154 and not w17285;
w17287 <= not w17284 and not w17286;
w17288 <= pi0781 and not w17287;
w17289 <= not w17282 and not w17288;
w17290 <= not pi0789 and not w17289;
w17291 <= not pi0619 and w17246;
w17292 <= pi0619 and w17289;
w17293 <= pi1159 and not w17291;
w17294 <= not w17292 and w17293;
w17295 <= not pi0619 and w17289;
w17296 <= pi0619 and w17246;
w17297 <= not pi1159 and not w17296;
w17298 <= not w17295 and w17297;
w17299 <= not w17294 and not w17298;
w17300 <= pi0789 and not w17299;
w17301 <= not w17290 and not w17300;
w17302 <= pi0626 and w17301;
w17303 <= pi1158 and not w17270;
w17304 <= not w17302 and w17303;
w17305 <= not pi0626 and w17301;
w17306 <= pi0626 and w17246;
w17307 <= not pi1158 and not w17306;
w17308 <= not w17305 and w17307;
w17309 <= not w17304 and not w17308;
w17310 <= not w14193 and w17309;
w17311 <= not w17269 and not w17310;
w17312 <= pi0788 and not w17311;
w17313 <= pi0618 and w17259;
w17314 <= pi0609 and w17258;
w17315 <= not w14731 and not w17249;
w17316 <= pi0625 and w17315;
w17317 <= w17272 and not w17315;
w17318 <= not w17316 and not w17317;
w17319 <= w17254 and not w17318;
w17320 <= not pi0608 and not w17253;
w17321 <= not w17319 and w17320;
w17322 <= pi1153 and w17272;
w17323 <= not w17316 and w17322;
w17324 <= pi0608 and not w17255;
w17325 <= not w17323 and w17324;
w17326 <= not w17321 and not w17325;
w17327 <= pi0778 and not w17326;
w17328 <= not pi0778 and not w17317;
w17329 <= not w17327 and not w17328;
w17330 <= not pi0609 and not w17329;
w17331 <= not pi1155 and not w17314;
w17332 <= not w17330 and w17331;
w17333 <= not pi0660 and not w17276;
w17334 <= not w17332 and w17333;
w17335 <= not pi0609 and w17258;
w17336 <= pi0609 and not w17329;
w17337 <= pi1155 and not w17335;
w17338 <= not w17336 and w17337;
w17339 <= pi0660 and not w17278;
w17340 <= not w17338 and w17339;
w17341 <= not w17334 and not w17340;
w17342 <= pi0785 and not w17341;
w17343 <= not pi0785 and not w17329;
w17344 <= not w17342 and not w17343;
w17345 <= not pi0618 and not w17344;
w17346 <= not pi1154 and not w17313;
w17347 <= not w17345 and w17346;
w17348 <= not pi0627 and not w17284;
w17349 <= not w17347 and w17348;
w17350 <= not pi0618 and w17259;
w17351 <= pi0618 and not w17344;
w17352 <= pi1154 and not w17350;
w17353 <= not w17351 and w17352;
w17354 <= pi0627 and not w17286;
w17355 <= not w17353 and w17354;
w17356 <= not w17349 and not w17355;
w17357 <= pi0781 and not w17356;
w17358 <= not pi0781 and not w17344;
w17359 <= not w17357 and not w17358;
w17360 <= not pi0789 and w17359;
w17361 <= not pi0619 and not w17359;
w17362 <= pi0619 and w17260;
w17363 <= not pi1159 and not w17362;
w17364 <= not w17361 and w17363;
w17365 <= not pi0648 and not w17294;
w17366 <= not w17364 and w17365;
w17367 <= not pi0619 and w17260;
w17368 <= pi0619 and not w17359;
w17369 <= pi1159 and not w17367;
w17370 <= not w17368 and w17369;
w17371 <= pi0648 and not w17298;
w17372 <= not w17370 and w17371;
w17373 <= pi0789 and not w17366;
w17374 <= not w17372 and w17373;
w17375 <= w15533 and not w17360;
w17376 <= not w17374 and w17375;
w17377 <= not w17312 and not w17376;
w17378 <= not pi0628 and not w17377;
w17379 <= not pi0788 and not w17301;
w17380 <= pi0788 and not w17309;
w17381 <= not w17379 and not w17380;
w17382 <= pi0628 and w17381;
w17383 <= not pi1156 and not w17382;
w17384 <= not w17378 and w17383;
w17385 <= not pi0629 and not w17268;
w17386 <= not w17384 and w17385;
w17387 <= not w15560 and w17262;
w17388 <= not pi1156 and not w17387;
w17389 <= not pi0628 and w17381;
w17390 <= pi0628 and not w17377;
w17391 <= pi1156 and not w17389;
w17392 <= not w17390 and w17391;
w17393 <= pi0629 and not w17388;
w17394 <= not w17392 and w17393;
w17395 <= not w17386 and not w17394;
w17396 <= pi0792 and not w17395;
w17397 <= not pi0792 and not w17377;
w17398 <= not w17396 and not w17397;
w17399 <= not pi0647 and not w17398;
w17400 <= not w15342 and w17381;
w17401 <= w15342 and w17246;
w17402 <= not w17400 and not w17401;
w17403 <= pi0647 and not w17402;
w17404 <= not pi1157 and not w17403;
w17405 <= not w17399 and w17404;
w17406 <= not pi0630 and not w17266;
w17407 <= not w17405 and w17406;
w17408 <= not pi0647 and w17263;
w17409 <= pi0647 and w17246;
w17410 <= not pi1157 and not w17409;
w17411 <= not w17408 and w17410;
w17412 <= pi0647 and not w17398;
w17413 <= not pi0647 and not w17402;
w17414 <= pi1157 and not w17413;
w17415 <= not w17412 and w17414;
w17416 <= pi0630 and not w17411;
w17417 <= not w17415 and w17416;
w17418 <= not w17407 and not w17417;
w17419 <= pi0787 and not w17418;
w17420 <= not pi0787 and not w17398;
w17421 <= not w17419 and not w17420;
w17422 <= not pi0790 and not w17421;
w17423 <= not pi0787 and not w17263;
w17424 <= not w17266 and not w17411;
w17425 <= pi0787 and not w17424;
w17426 <= not w17423 and not w17425;
w17427 <= not pi0644 and w17426;
w17428 <= pi0644 and not w17421;
w17429 <= pi0715 and not w17427;
w17430 <= not w17428 and w17429;
w17431 <= w15367 and not w17246;
w17432 <= not w15367 and w17402;
w17433 <= not w17431 and not w17432;
w17434 <= pi0644 and w17433;
w17435 <= not pi0644 and w17246;
w17436 <= not pi0715 and not w17435;
w17437 <= not w17434 and w17436;
w17438 <= pi1160 and not w17437;
w17439 <= not w17430 and w17438;
w17440 <= not pi0644 and w17433;
w17441 <= pi0644 and w17246;
w17442 <= pi0715 and not w17441;
w17443 <= not w17440 and w17442;
w17444 <= pi0644 and w17426;
w17445 <= not pi0644 and not w17421;
w17446 <= not pi0715 and not w17444;
w17447 <= not w17445 and w17446;
w17448 <= not pi1160 and not w17443;
w17449 <= not w17447 and w17448;
w17450 <= not w17439 and not w17449;
w17451 <= pi0790 and not w17450;
w17452 <= pi0832 and not w17422;
w17453 <= not w17451 and w17452;
w17454 <= not w17245 and not w17453;
w17455 <= pi0144 and not w14622;
w17456 <= w14198 and not w17455;
w17457 <= w14638 and not w17455;
w17458 <= pi0736 and w134;
w17459 <= not w17455 and not w17458;
w17460 <= not pi0144 and not w14204;
w17461 <= w14204 and not w14207;
w17462 <= pi0038 and not w17461;
w17463 <= not w17460 and w17462;
w17464 <= not pi0144 and w15639;
w17465 <= pi0144 and not w15635;
w17466 <= not pi0038 and not w17464;
w17467 <= not w17465 and w17466;
w17468 <= w17458 and not w17463;
w17469 <= not w17467 and w17468;
w17470 <= not w17459 and not w17469;
w17471 <= not pi0778 and w17470;
w17472 <= not pi0625 and not w17455;
w17473 <= pi0625 and not w17470;
w17474 <= pi1153 and not w17472;
w17475 <= not w17473 and w17474;
w17476 <= not pi0625 and not w17470;
w17477 <= pi0625 and not w17455;
w17478 <= not pi1153 and not w17477;
w17479 <= not w17476 and w17478;
w17480 <= not w17475 and not w17479;
w17481 <= pi0778 and not w17480;
w17482 <= not w17471 and not w17481;
w17483 <= not w14638 and w17482;
w17484 <= not w17457 and not w17483;
w17485 <= not w14202 and w17484;
w17486 <= w14202 and w17455;
w17487 <= not w17485 and not w17486;
w17488 <= not w14198 and w17487;
w17489 <= not w17456 and not w17488;
w17490 <= not w14194 and w17489;
w17491 <= w14194 and w17455;
w17492 <= not w17490 and not w17491;
w17493 <= not pi0792 and not w17492;
w17494 <= not pi0628 and not w17455;
w17495 <= pi0628 and w17492;
w17496 <= pi1156 and not w17494;
w17497 <= not w17495 and w17496;
w17498 <= pi0628 and not w17455;
w17499 <= not pi0628 and w17492;
w17500 <= not pi1156 and not w17498;
w17501 <= not w17499 and w17500;
w17502 <= not w17497 and not w17501;
w17503 <= pi0792 and not w17502;
w17504 <= not w17493 and not w17503;
w17505 <= not pi0787 and not w17504;
w17506 <= not pi0647 and not w17455;
w17507 <= pi0647 and w17504;
w17508 <= pi1157 and not w17506;
w17509 <= not w17507 and w17508;
w17510 <= pi0647 and not w17455;
w17511 <= not pi0647 and w17504;
w17512 <= not pi1157 and not w17510;
w17513 <= not w17511 and w17512;
w17514 <= not w17509 and not w17513;
w17515 <= pi0787 and not w17514;
w17516 <= not w17505 and not w17515;
w17517 <= not pi0644 and w17516;
w17518 <= not pi0619 and not w17455;
w17519 <= w14680 and not w17455;
w17520 <= pi0144 and not w134;
w17521 <= not pi0758 and not w14609;
w17522 <= pi0758 and w14782;
w17523 <= not w17521 and not w17522;
w17524 <= pi0039 and not w17523;
w17525 <= not pi0758 and w14521;
w17526 <= pi0758 and w14702;
w17527 <= not pi0039 and not w17525;
w17528 <= not w17526 and w17527;
w17529 <= not w17524 and not w17528;
w17530 <= pi0144 and not w17529;
w17531 <= not pi0144 and pi0758;
w17532 <= w14838 and w17531;
w17533 <= not w17530 and not w17532;
w17534 <= not pi0038 and not w17533;
w17535 <= pi0758 and w14731;
w17536 <= w14204 and not w17535;
w17537 <= pi0038 and not w17460;
w17538 <= not w17536 and w17537;
w17539 <= not w17534 and not w17538;
w17540 <= w134 and not w17539;
w17541 <= not w17520 and not w17540;
w17542 <= not w14680 and w17541;
w17543 <= not w17519 and not w17542;
w17544 <= not pi0785 and w17543;
w17545 <= not pi0609 and not w17455;
w17546 <= pi0609 and not w17543;
w17547 <= pi1155 and not w17545;
w17548 <= not w17546 and w17547;
w17549 <= not pi0609 and not w17543;
w17550 <= pi0609 and not w17455;
w17551 <= not pi1155 and not w17550;
w17552 <= not w17549 and w17551;
w17553 <= not w17548 and not w17552;
w17554 <= pi0785 and not w17553;
w17555 <= not w17544 and not w17554;
w17556 <= not pi0781 and not w17555;
w17557 <= not pi0618 and not w17455;
w17558 <= pi0618 and w17555;
w17559 <= pi1154 and not w17557;
w17560 <= not w17558 and w17559;
w17561 <= pi0618 and not w17455;
w17562 <= not pi0618 and w17555;
w17563 <= not pi1154 and not w17561;
w17564 <= not w17562 and w17563;
w17565 <= not w17560 and not w17564;
w17566 <= pi0781 and not w17565;
w17567 <= not w17556 and not w17566;
w17568 <= pi0619 and w17567;
w17569 <= pi1159 and not w17518;
w17570 <= not w17568 and w17569;
w17571 <= not pi0736 and w17539;
w17572 <= not pi0144 and not w15168;
w17573 <= pi0144 and w15109;
w17574 <= pi0758 and not w17573;
w17575 <= not w17572 and w17574;
w17576 <= pi0144 and not w14967;
w17577 <= not pi0144 and not w15048;
w17578 <= not pi0758 and not w17577;
w17579 <= not w17576 and w17578;
w17580 <= pi0039 and not w17575;
w17581 <= not w17579 and w17580;
w17582 <= not pi0144 and w15194;
w17583 <= pi0144 and w15192;
w17584 <= pi0758 and not w17582;
w17585 <= not w17583 and w17584;
w17586 <= not pi0144 and not w15188;
w17587 <= pi0144 and not w15175;
w17588 <= not pi0758 and not w17586;
w17589 <= not w17587 and w17588;
w17590 <= not pi0039 and not w17585;
w17591 <= not w17589 and w17590;
w17592 <= not pi0038 and not w17591;
w17593 <= not w17581 and w17592;
w17594 <= pi0736 and not w17033;
w17595 <= not w17538 and w17594;
w17596 <= not w17593 and w17595;
w17597 <= w134 and not w17596;
w17598 <= not w17571 and w17597;
w17599 <= not w17520 and not w17598;
w17600 <= not pi0625 and w17599;
w17601 <= pi0625 and w17541;
w17602 <= not pi1153 and not w17601;
w17603 <= not w17600 and w17602;
w17604 <= not pi0608 and not w17475;
w17605 <= not w17603 and w17604;
w17606 <= not pi0625 and w17541;
w17607 <= pi0625 and w17599;
w17608 <= pi1153 and not w17606;
w17609 <= not w17607 and w17608;
w17610 <= pi0608 and not w17479;
w17611 <= not w17609 and w17610;
w17612 <= not w17605 and not w17611;
w17613 <= pi0778 and not w17612;
w17614 <= not pi0778 and w17599;
w17615 <= not w17613 and not w17614;
w17616 <= not pi0609 and not w17615;
w17617 <= pi0609 and w17482;
w17618 <= not pi1155 and not w17617;
w17619 <= not w17616 and w17618;
w17620 <= not pi0660 and not w17548;
w17621 <= not w17619 and w17620;
w17622 <= not pi0609 and w17482;
w17623 <= pi0609 and not w17615;
w17624 <= pi1155 and not w17622;
w17625 <= not w17623 and w17624;
w17626 <= pi0660 and not w17552;
w17627 <= not w17625 and w17626;
w17628 <= not w17621 and not w17627;
w17629 <= pi0785 and not w17628;
w17630 <= not pi0785 and not w17615;
w17631 <= not w17629 and not w17630;
w17632 <= not pi0618 and not w17631;
w17633 <= pi0618 and not w17484;
w17634 <= not pi1154 and not w17633;
w17635 <= not w17632 and w17634;
w17636 <= not pi0627 and not w17560;
w17637 <= not w17635 and w17636;
w17638 <= pi0618 and not w17631;
w17639 <= not pi0618 and not w17484;
w17640 <= pi1154 and not w17639;
w17641 <= not w17638 and w17640;
w17642 <= pi0627 and not w17564;
w17643 <= not w17641 and w17642;
w17644 <= not w17637 and not w17643;
w17645 <= pi0781 and not w17644;
w17646 <= not pi0781 and not w17631;
w17647 <= not w17645 and not w17646;
w17648 <= not pi0619 and not w17647;
w17649 <= pi0619 and w17487;
w17650 <= not pi1159 and not w17649;
w17651 <= not w17648 and w17650;
w17652 <= not pi0648 and not w17570;
w17653 <= not w17651 and w17652;
w17654 <= pi0619 and not w17455;
w17655 <= not pi0619 and w17567;
w17656 <= not pi1159 and not w17654;
w17657 <= not w17655 and w17656;
w17658 <= not pi0619 and w17487;
w17659 <= pi0619 and not w17647;
w17660 <= pi1159 and not w17658;
w17661 <= not w17659 and w17660;
w17662 <= pi0648 and not w17657;
w17663 <= not w17661 and w17662;
w17664 <= not w17653 and not w17663;
w17665 <= pi0789 and not w17664;
w17666 <= not pi0789 and not w17647;
w17667 <= not w17665 and not w17666;
w17668 <= not pi0788 and w17667;
w17669 <= not pi0626 and w17667;
w17670 <= pi0626 and w17489;
w17671 <= not pi0641 and not w17670;
w17672 <= not w17669 and w17671;
w17673 <= not pi0789 and not w17567;
w17674 <= not w17570 and not w17657;
w17675 <= pi0789 and not w17674;
w17676 <= not w17673 and not w17675;
w17677 <= not pi0626 and w17676;
w17678 <= pi0626 and not w17455;
w17679 <= not pi1158 and not w17678;
w17680 <= not w17677 and w17679;
w17681 <= not w15293 and not w17680;
w17682 <= not w17672 and not w17681;
w17683 <= pi0626 and w17667;
w17684 <= not pi0626 and w17489;
w17685 <= pi0641 and not w17684;
w17686 <= not w17683 and w17685;
w17687 <= pi0626 and w17676;
w17688 <= not pi0626 and not w17455;
w17689 <= pi1158 and not w17688;
w17690 <= not w17687 and w17689;
w17691 <= not w15308 and not w17690;
w17692 <= not w17686 and not w17691;
w17693 <= not w17682 and not w17692;
w17694 <= pi0788 and not w17693;
w17695 <= not w17668 and not w17694;
w17696 <= not pi0628 and w17695;
w17697 <= not w17680 and not w17690;
w17698 <= pi0788 and not w17697;
w17699 <= not pi0788 and not w17676;
w17700 <= not w17698 and not w17699;
w17701 <= pi0628 and w17700;
w17702 <= not pi1156 and not w17701;
w17703 <= not w17696 and w17702;
w17704 <= not pi0629 and not w17497;
w17705 <= not w17703 and w17704;
w17706 <= pi0628 and w17695;
w17707 <= not pi0628 and w17700;
w17708 <= pi1156 and not w17707;
w17709 <= not w17706 and w17708;
w17710 <= pi0629 and not w17501;
w17711 <= not w17709 and w17710;
w17712 <= not w17705 and not w17711;
w17713 <= pi0792 and not w17712;
w17714 <= not pi0792 and w17695;
w17715 <= not w17713 and not w17714;
w17716 <= not pi0647 and not w17715;
w17717 <= not w15342 and not w17700;
w17718 <= w15342 and w17455;
w17719 <= not w17717 and not w17718;
w17720 <= pi0647 and w17719;
w17721 <= not pi1157 and not w17720;
w17722 <= not w17716 and w17721;
w17723 <= not pi0630 and not w17509;
w17724 <= not w17722 and w17723;
w17725 <= pi0647 and not w17715;
w17726 <= not pi0647 and w17719;
w17727 <= pi1157 and not w17726;
w17728 <= not w17725 and w17727;
w17729 <= pi0630 and not w17513;
w17730 <= not w17728 and w17729;
w17731 <= not w17724 and not w17730;
w17732 <= pi0787 and not w17731;
w17733 <= not pi0787 and not w17715;
w17734 <= not w17732 and not w17733;
w17735 <= pi0644 and not w17734;
w17736 <= pi0715 and not w17517;
w17737 <= not w17735 and w17736;
w17738 <= w15367 and not w17455;
w17739 <= not w15367 and w17719;
w17740 <= not w17738 and not w17739;
w17741 <= pi0644 and not w17740;
w17742 <= not pi0644 and not w17455;
w17743 <= not pi0715 and not w17742;
w17744 <= not w17741 and w17743;
w17745 <= pi1160 and not w17744;
w17746 <= not w17737 and w17745;
w17747 <= not pi0644 and not w17734;
w17748 <= pi0644 and w17516;
w17749 <= not pi0715 and not w17748;
w17750 <= not w17747 and w17749;
w17751 <= not pi0644 and not w17740;
w17752 <= pi0644 and not w17455;
w17753 <= pi0715 and not w17752;
w17754 <= not w17751 and w17753;
w17755 <= not pi1160 and not w17754;
w17756 <= not w17750 and w17755;
w17757 <= pi0790 and not w17746;
w17758 <= not w17756 and w17757;
w17759 <= not pi0790 and w17734;
w17760 <= w3868 and not w17759;
w17761 <= not w17758 and w17760;
w17762 <= not pi0144 and not w3868;
w17763 <= not pi0057 and not w17762;
w17764 <= not w17761 and w17763;
w17765 <= pi0057 and pi0144;
w17766 <= not pi0832 and not w17765;
w17767 <= not w17764 and w17766;
w17768 <= w15366 and w16904;
w17769 <= pi0787 and not w17768;
w17770 <= pi0144 and not w489;
w17771 <= pi0736 and w14208;
w17772 <= not w17770 and not w17771;
w17773 <= not pi0778 and w17772;
w17774 <= pi0625 and w17771;
w17775 <= not w17772 and not w17774;
w17776 <= not pi1153 and not w17775;
w17777 <= pi1153 and not w17770;
w17778 <= not w17774 and w17777;
w17779 <= not w17776 and not w17778;
w17780 <= pi0778 and not w17779;
w17781 <= not w17773 and not w17780;
w17782 <= w16714 and w17781;
w17783 <= not pi0628 and w17782;
w17784 <= pi0629 and not w17783;
w17785 <= not pi0609 and not pi1155;
w17786 <= pi0609 and pi1155;
w17787 <= pi0785 and not w17785;
w17788 <= not w17786 and w17787;
w17789 <= pi0758 and w14807;
w17790 <= not w17788 and w17789;
w17791 <= not pi0619 and pi1159;
w17792 <= pi0619 and not pi1159;
w17793 <= not w17791 and not w17792;
w17794 <= pi0789 and not w17793;
w17795 <= not pi0618 and not pi1154;
w17796 <= pi0618 and pi1154;
w17797 <= pi0781 and not w17795;
w17798 <= not w17796 and w17797;
w17799 <= not w14680 and not w17794;
w17800 <= not w17798 and w17799;
w17801 <= w17790 and w17800;
w17802 <= not w15532 and w17801;
w17803 <= pi0628 and not w17802;
w17804 <= not w17784 and not w17803;
w17805 <= not pi1156 and not w17804;
w17806 <= pi0628 and w17782;
w17807 <= not pi0628 and not w17802;
w17808 <= pi0629 and not w17807;
w17809 <= pi1156 and not w17808;
w17810 <= not w17806 and w17809;
w17811 <= not w17805 and not w17810;
w17812 <= not w17770 and not w17811;
w17813 <= pi0792 and w17812;
w17814 <= w14198 and not w17770;
w17815 <= not w14638 and w17781;
w17816 <= not w14202 and w17815;
w17817 <= not w17770 and not w17816;
w17818 <= not w17814 and not w17817;
w17819 <= w15428 and w17818;
w17820 <= not pi0626 and w17801;
w17821 <= not w17770 and not w17820;
w17822 <= not pi1158 and not w17821;
w17823 <= pi0641 and not w17822;
w17824 <= not w17819 and w17823;
w17825 <= pi0626 and w17801;
w17826 <= not w17770 and not w17825;
w17827 <= pi1158 and not w17826;
w17828 <= w15429 and w17818;
w17829 <= not pi0641 and not w17827;
w17830 <= not w17828 and w17829;
w17831 <= pi0788 and not w17824;
w17832 <= not w17830 and w17831;
w17833 <= pi0618 and not w14680;
w17834 <= w17790 and w17833;
w17835 <= pi1154 and not w17770;
w17836 <= not w17834 and w17835;
w17837 <= not w17770 and not w17815;
w17838 <= pi0618 and not w17837;
w17839 <= w14854 and w17789;
w17840 <= pi1155 and not w17770;
w17841 <= not w17839 and w17840;
w17842 <= pi0609 and w17781;
w17843 <= not w17770 and not w17789;
w17844 <= pi0736 and w15032;
w17845 <= w17843 and not w17844;
w17846 <= pi0625 and w17844;
w17847 <= not w17845 and not w17846;
w17848 <= not pi1153 and not w17847;
w17849 <= not pi0608 and not w17778;
w17850 <= not w17848 and w17849;
w17851 <= pi1153 and w17843;
w17852 <= not w17846 and w17851;
w17853 <= pi0608 and not w17776;
w17854 <= not w17852 and w17853;
w17855 <= not w17850 and not w17854;
w17856 <= pi0778 and not w17855;
w17857 <= not pi0778 and not w17845;
w17858 <= not w17856 and not w17857;
w17859 <= not pi0609 and not w17858;
w17860 <= not pi1155 and not w17842;
w17861 <= not w17859 and w17860;
w17862 <= not pi0660 and not w17841;
w17863 <= not w17861 and w17862;
w17864 <= w14859 and w17789;
w17865 <= not pi1155 and not w17770;
w17866 <= not w17864 and w17865;
w17867 <= not pi0609 and w17781;
w17868 <= pi0609 and not w17858;
w17869 <= pi1155 and not w17867;
w17870 <= not w17868 and w17869;
w17871 <= pi0660 and not w17866;
w17872 <= not w17870 and w17871;
w17873 <= not w17863 and not w17872;
w17874 <= pi0785 and not w17873;
w17875 <= not pi0785 and not w17858;
w17876 <= not w17874 and not w17875;
w17877 <= not pi0618 and not w17876;
w17878 <= not pi1154 and not w17838;
w17879 <= not w17877 and w17878;
w17880 <= not pi0627 and not w17836;
w17881 <= not w17879 and w17880;
w17882 <= not pi0618 and not w14680;
w17883 <= w17790 and w17882;
w17884 <= not pi1154 and not w17770;
w17885 <= not w17883 and w17884;
w17886 <= not pi0618 and not w17837;
w17887 <= pi0618 and not w17876;
w17888 <= pi1154 and not w17886;
w17889 <= not w17887 and w17888;
w17890 <= pi0627 and not w17885;
w17891 <= not w17889 and w17890;
w17892 <= not w17881 and not w17891;
w17893 <= pi0781 and not w17892;
w17894 <= not pi0781 and not w17876;
w17895 <= not w17893 and not w17894;
w17896 <= not pi0789 and w17895;
w17897 <= w17790 and not w17798;
w17898 <= pi0619 and not w14680;
w17899 <= w17897 and w17898;
w17900 <= pi1159 and not w17770;
w17901 <= not w17899 and w17900;
w17902 <= pi0619 and not w17817;
w17903 <= not pi0619 and not w17895;
w17904 <= not pi1159 and not w17902;
w17905 <= not w17903 and w17904;
w17906 <= not pi0648 and not w17901;
w17907 <= not w17905 and w17906;
w17908 <= not pi0619 and not w14680;
w17909 <= w17897 and w17908;
w17910 <= not pi1159 and not w17770;
w17911 <= not w17909 and w17910;
w17912 <= not pi0619 and not w17817;
w17913 <= pi0619 and not w17895;
w17914 <= pi1159 and not w17912;
w17915 <= not w17913 and w17914;
w17916 <= pi0648 and not w17911;
w17917 <= not w17915 and w17916;
w17918 <= pi0789 and not w17907;
w17919 <= not w17917 and w17918;
w17920 <= w15533 and not w17896;
w17921 <= not w17919 and w17920;
w17922 <= not w17832 and not w17921;
w17923 <= not w17813 and not w17922;
w17924 <= pi0629 and w16702;
w17925 <= not pi0629 and w16703;
w17926 <= pi0792 and not w17924;
w17927 <= not w17925 and w17926;
w17928 <= not w17812 and w17927;
w17929 <= not w17769 and not w17928;
w17930 <= not w17923 and w17929;
w17931 <= not w15342 and w17802;
w17932 <= not pi0630 and w17931;
w17933 <= pi0647 and not w17932;
w17934 <= not w16705 and w17782;
w17935 <= pi0630 and not w17934;
w17936 <= not w17933 and not w17935;
w17937 <= not pi1157 and not w17936;
w17938 <= pi0630 and w17931;
w17939 <= not pi0630 and not w17934;
w17940 <= pi0647 and not w17939;
w17941 <= pi1157 and not w17938;
w17942 <= not w17940 and w17941;
w17943 <= not w17937 and not w17942;
w17944 <= pi0787 and not w17770;
w17945 <= not w17943 and w17944;
w17946 <= not w17930 and not w17945;
w17947 <= not pi0790 and w17946;
w17948 <= not w15367 and w17931;
w17949 <= pi0644 and w17948;
w17950 <= not pi0715 and not w17770;
w17951 <= not w17949 and w17950;
w17952 <= not w16905 and w17934;
w17953 <= not w17770 and not w17952;
w17954 <= not pi0644 and not w17953;
w17955 <= pi0644 and w17946;
w17956 <= pi0715 and not w17954;
w17957 <= not w17955 and w17956;
w17958 <= pi1160 and not w17951;
w17959 <= not w17957 and w17958;
w17960 <= not pi0644 and w17948;
w17961 <= pi0715 and not w17770;
w17962 <= not w17960 and w17961;
w17963 <= not pi0644 and w17946;
w17964 <= pi0644 and not w17953;
w17965 <= not pi0715 and not w17964;
w17966 <= not w17963 and w17965;
w17967 <= not pi1160 and not w17962;
w17968 <= not w17966 and w17967;
w17969 <= not w17959 and not w17968;
w17970 <= pi0790 and not w17969;
w17971 <= pi0832 and not w17947;
w17972 <= not w17970 and w17971;
w17973 <= not w17767 and not w17972;
w17974 <= not pi0145 and not w4989;
w17975 <= not pi0145 and not w14622;
w17976 <= w14198 and not w17975;
w17977 <= not pi0698 and w134;
w17978 <= w17975 and not w17977;
w17979 <= not pi0145 and not w14204;
w17980 <= w14210 and not w17979;
w17981 <= pi0145 and not w15639;
w17982 <= not pi0038 and not w17981;
w17983 <= w134 and not w17982;
w17984 <= not pi0145 and w15635;
w17985 <= not w17983 and not w17984;
w17986 <= not pi0698 and not w17980;
w17987 <= not w17985 and w17986;
w17988 <= not w17978 and not w17987;
w17989 <= not pi0778 and w17988;
w17990 <= not pi0625 and w17975;
w17991 <= pi0625 and not w17988;
w17992 <= pi1153 and not w17990;
w17993 <= not w17991 and w17992;
w17994 <= pi0625 and w17975;
w17995 <= not pi0625 and not w17988;
w17996 <= not pi1153 and not w17994;
w17997 <= not w17995 and w17996;
w17998 <= not w17993 and not w17997;
w17999 <= pi0778 and not w17998;
w18000 <= not w17989 and not w17999;
w18001 <= not w14638 and not w18000;
w18002 <= w14638 and not w17975;
w18003 <= not w18001 and not w18002;
w18004 <= not w14202 and w18003;
w18005 <= w14202 and w17975;
w18006 <= not w18004 and not w18005;
w18007 <= not w14198 and w18006;
w18008 <= not w17976 and not w18007;
w18009 <= not w14194 and w18008;
w18010 <= w14194 and w17975;
w18011 <= not w18009 and not w18010;
w18012 <= not pi0792 and w18011;
w18013 <= pi0628 and not w18011;
w18014 <= not pi0628 and w17975;
w18015 <= pi1156 and not w18014;
w18016 <= not w18013 and w18015;
w18017 <= pi0628 and w17975;
w18018 <= not pi0628 and not w18011;
w18019 <= not pi1156 and not w18017;
w18020 <= not w18018 and w18019;
w18021 <= not w18016 and not w18020;
w18022 <= pi0792 and not w18021;
w18023 <= not w18012 and not w18022;
w18024 <= not pi0647 and not w18023;
w18025 <= pi0647 and not w17975;
w18026 <= not w18024 and not w18025;
w18027 <= not pi1157 and w18026;
w18028 <= pi0647 and not w18023;
w18029 <= not pi0647 and not w17975;
w18030 <= not w18028 and not w18029;
w18031 <= pi1157 and w18030;
w18032 <= not w18027 and not w18031;
w18033 <= pi0787 and not w18032;
w18034 <= not pi0787 and w18023;
w18035 <= not w18033 and not w18034;
w18036 <= not pi0644 and not w18035;
w18037 <= pi0715 and not w18036;
w18038 <= pi0145 and not w134;
w18039 <= pi0145 and not w14838;
w18040 <= not pi0145 and not w14611;
w18041 <= pi0767 and not w18040;
w18042 <= not pi0145 and not pi0767;
w18043 <= w14784 and w18042;
w18044 <= not w18039 and not w18043;
w18045 <= not w18041 and w18044;
w18046 <= not pi0038 and not w18045;
w18047 <= not pi0767 and w14843;
w18048 <= pi0038 and not w17979;
w18049 <= not w18047 and w18048;
w18050 <= not w18046 and not w18049;
w18051 <= w134 and not w18050;
w18052 <= not w18038 and not w18051;
w18053 <= not w14680 and not w18052;
w18054 <= w14680 and not w17975;
w18055 <= not w18053 and not w18054;
w18056 <= not pi0785 and not w18055;
w18057 <= not w14854 and not w17975;
w18058 <= pi0609 and w18053;
w18059 <= not w18057 and not w18058;
w18060 <= pi1155 and not w18059;
w18061 <= not w14859 and not w17975;
w18062 <= not pi0609 and w18053;
w18063 <= not w18061 and not w18062;
w18064 <= not pi1155 and not w18063;
w18065 <= not w18060 and not w18064;
w18066 <= pi0785 and not w18065;
w18067 <= not w18056 and not w18066;
w18068 <= not pi0781 and not w18067;
w18069 <= not pi0618 and w17975;
w18070 <= pi0618 and w18067;
w18071 <= pi1154 and not w18069;
w18072 <= not w18070 and w18071;
w18073 <= not pi0618 and w18067;
w18074 <= pi0618 and w17975;
w18075 <= not pi1154 and not w18074;
w18076 <= not w18073 and w18075;
w18077 <= not w18072 and not w18076;
w18078 <= pi0781 and not w18077;
w18079 <= not w18068 and not w18078;
w18080 <= not pi0789 and not w18079;
w18081 <= not pi0619 and w17975;
w18082 <= pi0619 and w18079;
w18083 <= pi1159 and not w18081;
w18084 <= not w18082 and w18083;
w18085 <= not pi0619 and w18079;
w18086 <= pi0619 and w17975;
w18087 <= not pi1159 and not w18086;
w18088 <= not w18085 and w18087;
w18089 <= not w18084 and not w18088;
w18090 <= pi0789 and not w18089;
w18091 <= not w18080 and not w18090;
w18092 <= not pi0788 and not w18091;
w18093 <= not pi0626 and w17975;
w18094 <= pi0626 and w18091;
w18095 <= pi1158 and not w18093;
w18096 <= not w18094 and w18095;
w18097 <= not pi0626 and w18091;
w18098 <= pi0626 and w17975;
w18099 <= not pi1158 and not w18098;
w18100 <= not w18097 and w18099;
w18101 <= not w18096 and not w18100;
w18102 <= pi0788 and not w18101;
w18103 <= not w18092 and not w18102;
w18104 <= not w15342 and w18103;
w18105 <= w15342 and w17975;
w18106 <= not w18104 and not w18105;
w18107 <= not w15367 and not w18106;
w18108 <= w15367 and w17975;
w18109 <= not w18107 and not w18108;
w18110 <= pi0644 and not w18109;
w18111 <= not pi0644 and w17975;
w18112 <= not pi0715 and not w18111;
w18113 <= not w18110 and w18112;
w18114 <= pi1160 and not w18113;
w18115 <= not w18037 and w18114;
w18116 <= pi0644 and not w18035;
w18117 <= w15365 and not w18026;
w18118 <= pi0630 and not pi0647;
w18119 <= pi1157 and w18118;
w18120 <= not pi0630 and pi0647;
w18121 <= not pi1157 and w18120;
w18122 <= not w18119 and not w18121;
w18123 <= w18106 and not w18122;
w18124 <= w15364 and not w18030;
w18125 <= not w18117 and not w18124;
w18126 <= not w18123 and w18125;
w18127 <= pi0787 and not w18126;
w18128 <= not pi0629 and w18016;
w18129 <= not pi0628 and pi0629;
w18130 <= pi1156 and w18129;
w18131 <= pi0628 and not pi0629;
w18132 <= not pi1156 and w18131;
w18133 <= not w18130 and not w18132;
w18134 <= not w18103 and not w18133;
w18135 <= pi0629 and w18020;
w18136 <= not w18128 and not w18135;
w18137 <= not w18134 and w18136;
w18138 <= pi0792 and not w18137;
w18139 <= pi0609 and w18000;
w18140 <= pi0145 and not w15188;
w18141 <= not pi0145 and not w15175;
w18142 <= pi0767 and not w18140;
w18143 <= not w18141 and w18142;
w18144 <= not pi0145 and w15192;
w18145 <= pi0145 and w15194;
w18146 <= not pi0767 and not w18145;
w18147 <= not w18144 and w18146;
w18148 <= not w18143 and not w18147;
w18149 <= not pi0039 and not w18148;
w18150 <= pi0145 and w15168;
w18151 <= not pi0145 and not w15109;
w18152 <= not pi0767 and not w18151;
w18153 <= not w18150 and w18152;
w18154 <= not pi0145 and w14967;
w18155 <= pi0145 and w15048;
w18156 <= pi0767 and not w18155;
w18157 <= not w18154 and w18156;
w18158 <= pi0039 and not w18153;
w18159 <= not w18157 and w18158;
w18160 <= not pi0038 and not w18149;
w18161 <= not w18159 and w18160;
w18162 <= not pi0767 and not w15053;
w18163 <= w17034 and not w18162;
w18164 <= not pi0145 and not w18163;
w18165 <= not pi0767 and w14807;
w18166 <= not w15032 and not w18165;
w18167 <= pi0145 and not w18166;
w18168 <= w3847 and w18167;
w18169 <= pi0038 and not w18168;
w18170 <= not w18164 and w18169;
w18171 <= not pi0698 and not w18170;
w18172 <= not w18161 and w18171;
w18173 <= pi0698 and w18050;
w18174 <= w134 and not w18172;
w18175 <= not w18173 and w18174;
w18176 <= not w18038 and not w18175;
w18177 <= not pi0625 and w18176;
w18178 <= pi0625 and w18052;
w18179 <= not pi1153 and not w18178;
w18180 <= not w18177 and w18179;
w18181 <= not pi0608 and not w17993;
w18182 <= not w18180 and w18181;
w18183 <= not pi0625 and w18052;
w18184 <= pi0625 and w18176;
w18185 <= pi1153 and not w18183;
w18186 <= not w18184 and w18185;
w18187 <= pi0608 and not w17997;
w18188 <= not w18186 and w18187;
w18189 <= not w18182 and not w18188;
w18190 <= pi0778 and not w18189;
w18191 <= not pi0778 and w18176;
w18192 <= not w18190 and not w18191;
w18193 <= not pi0609 and not w18192;
w18194 <= not pi1155 and not w18139;
w18195 <= not w18193 and w18194;
w18196 <= not pi0660 and not w18060;
w18197 <= not w18195 and w18196;
w18198 <= not pi0609 and w18000;
w18199 <= pi0609 and not w18192;
w18200 <= pi1155 and not w18198;
w18201 <= not w18199 and w18200;
w18202 <= pi0660 and not w18064;
w18203 <= not w18201 and w18202;
w18204 <= not w18197 and not w18203;
w18205 <= pi0785 and not w18204;
w18206 <= not pi0785 and not w18192;
w18207 <= not w18205 and not w18206;
w18208 <= not pi0618 and not w18207;
w18209 <= pi0618 and w18003;
w18210 <= not pi1154 and not w18209;
w18211 <= not w18208 and w18210;
w18212 <= not pi0627 and not w18072;
w18213 <= not w18211 and w18212;
w18214 <= not pi0618 and w18003;
w18215 <= pi0618 and not w18207;
w18216 <= pi1154 and not w18214;
w18217 <= not w18215 and w18216;
w18218 <= pi0627 and not w18076;
w18219 <= not w18217 and w18218;
w18220 <= not w18213 and not w18219;
w18221 <= pi0781 and not w18220;
w18222 <= not pi0781 and not w18207;
w18223 <= not w18221 and not w18222;
w18224 <= not pi0789 and w18223;
w18225 <= pi0619 and not w18006;
w18226 <= not pi0619 and not w18223;
w18227 <= not pi1159 and not w18225;
w18228 <= not w18226 and w18227;
w18229 <= not pi0648 and not w18084;
w18230 <= not w18228 and w18229;
w18231 <= pi0619 and not w18223;
w18232 <= not pi0619 and not w18006;
w18233 <= pi1159 and not w18232;
w18234 <= not w18231 and w18233;
w18235 <= pi0648 and not w18088;
w18236 <= not w18234 and w18235;
w18237 <= pi0789 and not w18230;
w18238 <= not w18236 and w18237;
w18239 <= w15533 and not w18224;
w18240 <= not w18238 and w18239;
w18241 <= w15434 and w18008;
w18242 <= not w14193 and w18101;
w18243 <= not w18241 and not w18242;
w18244 <= pi0788 and not w18243;
w18245 <= not w17927 and not w18244;
w18246 <= not w18240 and w18245;
w18247 <= not w18138 and not w18246;
w18248 <= not w17769 and not w18247;
w18249 <= not w18127 and not w18248;
w18250 <= not pi0644 and w18249;
w18251 <= not pi0715 and not w18116;
w18252 <= not w18250 and w18251;
w18253 <= pi0644 and w17975;
w18254 <= not pi0644 and not w18109;
w18255 <= pi0715 and not w18253;
w18256 <= not w18254 and w18255;
w18257 <= not pi1160 and not w18256;
w18258 <= not w18252 and w18257;
w18259 <= not w18115 and not w18258;
w18260 <= pi0790 and not w18259;
w18261 <= pi0644 and w18114;
w18262 <= pi0790 and not w18261;
w18263 <= w18249 and not w18262;
w18264 <= not w18260 and not w18263;
w18265 <= w4989 and not w18264;
w18266 <= not pi0832 and not w17974;
w18267 <= not w18265 and w18266;
w18268 <= not pi0145 and not w489;
w18269 <= not pi0698 and w14208;
w18270 <= not w18268 and not w18269;
w18271 <= not pi0778 and w18270;
w18272 <= not pi0625 and w18269;
w18273 <= not w18270 and not w18272;
w18274 <= pi1153 and not w18273;
w18275 <= not pi1153 and not w18268;
w18276 <= not w18272 and w18275;
w18277 <= not w18274 and not w18276;
w18278 <= pi0778 and not w18277;
w18279 <= not w18271 and not w18278;
w18280 <= not w15408 and w18279;
w18281 <= not w15410 and w18280;
w18282 <= not w15412 and w18281;
w18283 <= not w15414 and w18282;
w18284 <= not w15420 and w18283;
w18285 <= not pi0647 and w18284;
w18286 <= pi0647 and w18268;
w18287 <= not pi1157 and not w18286;
w18288 <= not w18285 and w18287;
w18289 <= pi0630 and w18288;
w18290 <= not w18165 and not w18268;
w18291 <= not w15437 and not w18290;
w18292 <= not pi0785 and not w18291;
w18293 <= not w15442 and not w18290;
w18294 <= pi1155 and not w18293;
w18295 <= not w15445 and w18291;
w18296 <= not pi1155 and not w18295;
w18297 <= not w18294 and not w18296;
w18298 <= pi0785 and not w18297;
w18299 <= not w18292 and not w18298;
w18300 <= not pi0781 and not w18299;
w18301 <= not w15452 and w18299;
w18302 <= pi1154 and not w18301;
w18303 <= not w15455 and w18299;
w18304 <= not pi1154 and not w18303;
w18305 <= not w18302 and not w18304;
w18306 <= pi0781 and not w18305;
w18307 <= not w18300 and not w18306;
w18308 <= not pi0789 and not w18307;
w18309 <= not pi0619 and w18268;
w18310 <= pi0619 and w18307;
w18311 <= pi1159 and not w18309;
w18312 <= not w18310 and w18311;
w18313 <= not pi0619 and w18307;
w18314 <= pi0619 and w18268;
w18315 <= not pi1159 and not w18314;
w18316 <= not w18313 and w18315;
w18317 <= not w18312 and not w18316;
w18318 <= pi0789 and not w18317;
w18319 <= not w18308 and not w18318;
w18320 <= not pi0788 and not w18319;
w18321 <= not pi0626 and w18268;
w18322 <= pi0626 and w18319;
w18323 <= pi1158 and not w18321;
w18324 <= not w18322 and w18323;
w18325 <= not pi0626 and w18319;
w18326 <= pi0626 and w18268;
w18327 <= not pi1158 and not w18326;
w18328 <= not w18325 and w18327;
w18329 <= not w18324 and not w18328;
w18330 <= pi0788 and not w18329;
w18331 <= not w18320 and not w18330;
w18332 <= not w15342 and w18331;
w18333 <= w15342 and w18268;
w18334 <= not w18332 and not w18333;
w18335 <= not w18122 and w18334;
w18336 <= pi0647 and not w18284;
w18337 <= not pi0647 and not w18268;
w18338 <= not w18336 and not w18337;
w18339 <= w15364 and not w18338;
w18340 <= not w18289 and not w18339;
w18341 <= not w18335 and w18340;
w18342 <= pi0787 and not w18341;
w18343 <= w15434 and w18282;
w18344 <= not w14193 and w18329;
w18345 <= not w18343 and not w18344;
w18346 <= pi0788 and not w18345;
w18347 <= pi0618 and w18280;
w18348 <= pi0609 and w18279;
w18349 <= not w14731 and not w18270;
w18350 <= pi0625 and w18349;
w18351 <= w18290 and not w18349;
w18352 <= not w18350 and not w18351;
w18353 <= w18275 and not w18352;
w18354 <= not pi0608 and not w18274;
w18355 <= not w18353 and w18354;
w18356 <= pi1153 and w18290;
w18357 <= not w18350 and w18356;
w18358 <= pi0608 and not w18276;
w18359 <= not w18357 and w18358;
w18360 <= not w18355 and not w18359;
w18361 <= pi0778 and not w18360;
w18362 <= not pi0778 and not w18351;
w18363 <= not w18361 and not w18362;
w18364 <= not pi0609 and not w18363;
w18365 <= not pi1155 and not w18348;
w18366 <= not w18364 and w18365;
w18367 <= not pi0660 and not w18294;
w18368 <= not w18366 and w18367;
w18369 <= not pi0609 and w18279;
w18370 <= pi0609 and not w18363;
w18371 <= pi1155 and not w18369;
w18372 <= not w18370 and w18371;
w18373 <= pi0660 and not w18296;
w18374 <= not w18372 and w18373;
w18375 <= not w18368 and not w18374;
w18376 <= pi0785 and not w18375;
w18377 <= not pi0785 and not w18363;
w18378 <= not w18376 and not w18377;
w18379 <= not pi0618 and not w18378;
w18380 <= not pi1154 and not w18347;
w18381 <= not w18379 and w18380;
w18382 <= not pi0627 and not w18302;
w18383 <= not w18381 and w18382;
w18384 <= not pi0618 and w18280;
w18385 <= pi0618 and not w18378;
w18386 <= pi1154 and not w18384;
w18387 <= not w18385 and w18386;
w18388 <= pi0627 and not w18304;
w18389 <= not w18387 and w18388;
w18390 <= not w18383 and not w18389;
w18391 <= pi0781 and not w18390;
w18392 <= not pi0781 and not w18378;
w18393 <= not w18391 and not w18392;
w18394 <= not pi0789 and w18393;
w18395 <= not pi0619 and not w18393;
w18396 <= pi0619 and w18281;
w18397 <= not pi1159 and not w18396;
w18398 <= not w18395 and w18397;
w18399 <= not pi0648 and not w18312;
w18400 <= not w18398 and w18399;
w18401 <= not pi0619 and w18281;
w18402 <= pi0619 and not w18393;
w18403 <= pi1159 and not w18401;
w18404 <= not w18402 and w18403;
w18405 <= pi0648 and not w18316;
w18406 <= not w18404 and w18405;
w18407 <= pi0789 and not w18400;
w18408 <= not w18406 and w18407;
w18409 <= w15533 and not w18394;
w18410 <= not w18408 and w18409;
w18411 <= not w18346 and not w18410;
w18412 <= not w17927 and not w18411;
w18413 <= w15417 and w18331;
w18414 <= pi1156 and not w15425;
w18415 <= w18283 and w18414;
w18416 <= not w18413 and not w18415;
w18417 <= not pi0629 and not w18416;
w18418 <= not pi1156 and not w15560;
w18419 <= w18283 and w18418;
w18420 <= w15416 and w18331;
w18421 <= not w18419 and not w18420;
w18422 <= pi0629 and not w18421;
w18423 <= not w18417 and not w18422;
w18424 <= pi0792 and not w18423;
w18425 <= not w17769 and not w18424;
w18426 <= not w18412 and w18425;
w18427 <= not w18342 and not w18426;
w18428 <= not pi0790 and w18427;
w18429 <= not pi0787 and not w18284;
w18430 <= pi1157 and not w18338;
w18431 <= not w18288 and not w18430;
w18432 <= pi0787 and not w18431;
w18433 <= not w18429 and not w18432;
w18434 <= not pi0644 and w18433;
w18435 <= pi0644 and w18427;
w18436 <= pi0715 and not w18434;
w18437 <= not w18435 and w18436;
w18438 <= not w15367 and not w18334;
w18439 <= w15367 and w18268;
w18440 <= not w18438 and not w18439;
w18441 <= pi0644 and not w18440;
w18442 <= not pi0644 and w18268;
w18443 <= not pi0715 and not w18442;
w18444 <= not w18441 and w18443;
w18445 <= pi1160 and not w18444;
w18446 <= not w18437 and w18445;
w18447 <= not pi0644 and not w18440;
w18448 <= pi0644 and w18268;
w18449 <= pi0715 and not w18448;
w18450 <= not w18447 and w18449;
w18451 <= pi0644 and w18433;
w18452 <= not pi0644 and w18427;
w18453 <= not pi0715 and not w18451;
w18454 <= not w18452 and w18453;
w18455 <= not pi1160 and not w18450;
w18456 <= not w18454 and w18455;
w18457 <= not w18446 and not w18456;
w18458 <= pi0790 and not w18457;
w18459 <= pi0832 and not w18428;
w18460 <= not w18458 and w18459;
w18461 <= not w18267 and not w18460;
w18462 <= not pi0146 and not w7760;
w18463 <= not pi0146 and not w14204;
w18464 <= pi0743 and pi0947;
w18465 <= pi0907 and not pi0947;
w18466 <= pi0735 and w18465;
w18467 <= not w18464 and not w18466;
w18468 <= w489 and w18467;
w18469 <= w3847 and w18468;
w18470 <= pi0038 and not w18469;
w18471 <= not w18463 and w18470;
w18472 <= not pi0146 and not w14504;
w18473 <= w14504 and w18467;
w18474 <= pi0299 and not w18472;
w18475 <= not w18473 and w18474;
w18476 <= not pi0146 and not w14493;
w18477 <= w14493 and w18467;
w18478 <= not pi0299 and not w18476;
w18479 <= not w18477 and w18478;
w18480 <= not pi0039 and not w18475;
w18481 <= not w18479 and w18480;
w18482 <= w14216 and not w18467;
w18483 <= pi0146 and not w14216;
w18484 <= not w18482 and not w18483;
w18485 <= w1011 and not w18484;
w18486 <= not pi0907 and w3804;
w18487 <= pi0146 and not w14581;
w18488 <= not w18486 and w18487;
w18489 <= pi0735 and pi0907;
w18490 <= w14581 and w18489;
w18491 <= pi0146 and not w14574;
w18492 <= w18486 and w18491;
w18493 <= not pi0947 and not w18490;
w18494 <= not w18492 and w18493;
w18495 <= pi0743 and w14581;
w18496 <= pi0947 and not w18487;
w18497 <= not w18495 and w18496;
w18498 <= not w18494 and not w18497;
w18499 <= not w18488 and not w18498;
w18500 <= not w1011 and not w18499;
w18501 <= not pi0215 and not w18485;
w18502 <= not w18500 and w18501;
w18503 <= w14533 and not w18467;
w18504 <= pi0146 and w14605;
w18505 <= pi0215 and not w18503;
w18506 <= not w18504 and w18505;
w18507 <= not w18502 and not w18506;
w18508 <= pi0299 and not w18507;
w18509 <= pi0146 and not w14533;
w18510 <= not w18503 and not w18509;
w18511 <= not w3768 and not w18510;
w18512 <= not pi0146 and not w14553;
w18513 <= w14553 and w18467;
w18514 <= w3768 and not w18512;
w18515 <= not w18513 and w18514;
w18516 <= not w18511 and not w18515;
w18517 <= pi0223 and not w18516;
w18518 <= w166 and w18484;
w18519 <= w14581 and not w18467;
w18520 <= not w3768 and not w18487;
w18521 <= not w18519 and w18520;
w18522 <= w14574 and not w18467;
w18523 <= w3768 and not w18491;
w18524 <= not w18522 and w18523;
w18525 <= not w18521 and not w18524;
w18526 <= not w166 and not w18525;
w18527 <= not pi0223 and not w18518;
w18528 <= not w18526 and w18527;
w18529 <= not pi0299 and not w18517;
w18530 <= not w18528 and w18529;
w18531 <= not w18508 and not w18530;
w18532 <= pi0039 and not w18531;
w18533 <= not pi0038 and not w18481;
w18534 <= not w18532 and w18533;
w18535 <= w7760 and not w18471;
w18536 <= not w18534 and w18535;
w18537 <= not pi0832 and not w18462;
w18538 <= not w18536 and w18537;
w18539 <= not pi0146 and not w489;
w18540 <= pi0832 and not w18539;
w18541 <= not w18468 and w18540;
w18542 <= not w18538 and not w18541;
w18543 <= not pi0147 and not w489;
w18544 <= not pi0770 and pi0947;
w18545 <= pi0726 and w18465;
w18546 <= not w18544 and not w18545;
w18547 <= w489 and not w18546;
w18548 <= pi0832 and not w18543;
w18549 <= not w18547 and w18548;
w18550 <= not pi0147 and not w7760;
w18551 <= not pi0947 and w14521;
w18552 <= not pi0039 and not w18551;
w18553 <= not pi0299 and w14587;
w18554 <= pi0947 and w18553;
w18555 <= not pi0947 and w14589;
w18556 <= w14581 and w18465;
w18557 <= not w14593 and not w18556;
w18558 <= not w1011 and not w18557;
w18559 <= not pi0215 and not w18558;
w18560 <= not w18555 and w18559;
w18561 <= pi0215 and not w14604;
w18562 <= w14533 and w18465;
w18563 <= w18561 and not w18562;
w18564 <= not w18560 and not w18563;
w18565 <= pi0299 and not w18564;
w18566 <= not w14588 and not w18565;
w18567 <= not w18554 and w18566;
w18568 <= pi0039 and not w18567;
w18569 <= not w18552 and not w18568;
w18570 <= not pi0038 and w18569;
w18571 <= pi0038 and not pi0947;
w18572 <= w14613 and w18571;
w18573 <= not w18570 and not w18572;
w18574 <= not pi0770 and w18573;
w18575 <= pi0770 and not w14615;
w18576 <= not w18574 and not w18575;
w18577 <= not pi0147 and not w18576;
w18578 <= not w14614 and not w18572;
w18579 <= pi0947 and w14521;
w18580 <= not pi0039 and not w18579;
w18581 <= pi0947 and w14587;
w18582 <= not pi0299 and not w18581;
w18583 <= pi0215 and pi0947;
w18584 <= w14533 and w18583;
w18585 <= pi0299 and not w18584;
w18586 <= pi0947 and w14581;
w18587 <= not w1011 and not w18586;
w18588 <= pi0947 and w14216;
w18589 <= w1011 and not w18588;
w18590 <= not pi0215 and not w18589;
w18591 <= not w18587 and w18590;
w18592 <= w18585 and not w18591;
w18593 <= not w18582 and not w18592;
w18594 <= pi0039 and not w18593;
w18595 <= not w18580 and not w18594;
w18596 <= not pi0038 and not w18595;
w18597 <= w18578 and not w18596;
w18598 <= pi0147 and not pi0770;
w18599 <= w18597 and w18598;
w18600 <= not pi0726 and not w18599;
w18601 <= not w18577 and w18600;
w18602 <= w3799 and w14613;
w18603 <= not pi0147 and not w18602;
w18604 <= not w3799 and w14204;
w18605 <= pi0038 and not w18604;
w18606 <= not w18603 and w18605;
w18607 <= pi0299 and pi0947;
w18608 <= w14589 and not w18465;
w18609 <= not w14593 and not w18586;
w18610 <= not w1011 and not w18609;
w18611 <= not pi0215 and not w18610;
w18612 <= not w18608 and w18611;
w18613 <= not w18561 and not w18612;
w18614 <= pi0299 and not w18613;
w18615 <= not pi0947 and w14555;
w18616 <= pi0223 and not w18615;
w18617 <= w14555 and not w18465;
w18618 <= pi0223 and not w18617;
w18619 <= w84 and w14217;
w18620 <= not w14584 and not w18619;
w18621 <= w3799 and not w18620;
w18622 <= not pi0223 and not w18621;
w18623 <= not w18616 and not w18618;
w18624 <= not w18622 and w18623;
w18625 <= not pi0299 and not w18624;
w18626 <= not w18607 and not w18614;
w18627 <= not w18625 and w18626;
w18628 <= pi0039 and w18627;
w18629 <= not w3799 and w14521;
w18630 <= not pi0039 and not w18629;
w18631 <= w14521 and w18630;
w18632 <= not w18628 and not w18631;
w18633 <= not pi0147 and w18632;
w18634 <= not w3799 and w14587;
w18635 <= not pi0299 and w18634;
w18636 <= pi0215 and not w14600;
w18637 <= not w3799 and w14216;
w18638 <= w1011 and w18637;
w18639 <= not pi0215 and not w18638;
w18640 <= not w14596 and w18639;
w18641 <= pi0299 and not w18636;
w18642 <= not w18640 and w18641;
w18643 <= not w18635 and not w18642;
w18644 <= pi0039 and w18643;
w18645 <= not w18630 and not w18644;
w18646 <= pi0147 and w18645;
w18647 <= not pi0038 and not w18646;
w18648 <= not w18633 and w18647;
w18649 <= not pi0770 and not w18606;
w18650 <= not w18648 and w18649;
w18651 <= not pi0147 and not w14204;
w18652 <= w14204 and w18465;
w18653 <= pi0038 and not w18652;
w18654 <= not w18651 and w18653;
w18655 <= not w18584 and not w18613;
w18656 <= pi0299 and not w18655;
w18657 <= not w18465 and w18553;
w18658 <= not w18656 and not w18657;
w18659 <= pi0039 and not w18658;
w18660 <= w14521 and not w18465;
w18661 <= not pi0039 and w18660;
w18662 <= not w18659 and not w18661;
w18663 <= not pi0147 and w18662;
w18664 <= pi0215 and not w18562;
w18665 <= not w1011 and not w18556;
w18666 <= pi0907 and w14216;
w18667 <= not pi0947 and w18666;
w18668 <= w1011 and not w18667;
w18669 <= not w18665 and not w18668;
w18670 <= not pi0215 and not w18669;
w18671 <= not w18664 and not w18670;
w18672 <= pi0299 and not w18671;
w18673 <= w14587 and w18465;
w18674 <= not pi0299 and not w18673;
w18675 <= not w18672 and not w18674;
w18676 <= pi0039 and not w18675;
w18677 <= w14521 and w18465;
w18678 <= not pi0039 and not w18677;
w18679 <= not w18676 and not w18678;
w18680 <= pi0147 and w18679;
w18681 <= not pi0038 and not w18680;
w18682 <= not w18663 and w18681;
w18683 <= pi0770 and not w18654;
w18684 <= not w18682 and w18683;
w18685 <= pi0726 and not w18650;
w18686 <= not w18684 and w18685;
w18687 <= w7760 and not w18686;
w18688 <= not w18601 and w18687;
w18689 <= not pi0832 and not w18550;
w18690 <= not w18688 and w18689;
w18691 <= not w18549 and not w18690;
w18692 <= pi0057 and pi0148;
w18693 <= w134 and w3868;
w18694 <= not pi0148 and not w18693;
w18695 <= not pi0749 and pi0947;
w18696 <= w18604 and not w18695;
w18697 <= not pi0148 and not w14204;
w18698 <= not w18696 and not w18697;
w18699 <= pi0038 and not w18698;
w18700 <= not w14588 and not w18672;
w18701 <= pi0148 and not w18700;
w18702 <= not w7300 and not w18658;
w18703 <= not pi0749 and not w18701;
w18704 <= not w18702 and w18703;
w18705 <= not pi0148 and w18627;
w18706 <= pi0148 and w18643;
w18707 <= pi0749 and not w18706;
w18708 <= not w18705 and w18707;
w18709 <= pi0039 and not w18704;
w18710 <= not w18708 and w18709;
w18711 <= not pi0148 and not w14521;
w18712 <= not pi0039 and not w18711;
w18713 <= w18629 and not w18695;
w18714 <= w18712 and not w18713;
w18715 <= not pi0038 and not w18714;
w18716 <= not w18710 and w18715;
w18717 <= pi0706 and not w18699;
w18718 <= not w18716 and w18717;
w18719 <= pi0749 and pi0947;
w18720 <= w14521 and w18719;
w18721 <= w18712 and not w18720;
w18722 <= not pi0148 and not pi0749;
w18723 <= not w14609 and w18722;
w18724 <= not pi0148 and not w18564;
w18725 <= not w18584 and not w18591;
w18726 <= pi0148 and not w18725;
w18727 <= pi0299 and not w18726;
w18728 <= not w18724 and w18727;
w18729 <= not pi0148 and not w14587;
w18730 <= w18582 and not w18729;
w18731 <= pi0749 and not w18730;
w18732 <= not w18728 and w18731;
w18733 <= pi0039 and not w18723;
w18734 <= not w18732 and w18733;
w18735 <= not pi0038 and not w18721;
w18736 <= not w18734 and w18735;
w18737 <= w14204 and not w18719;
w18738 <= pi0148 and not w14613;
w18739 <= pi0038 and not w18737;
w18740 <= not w18738 and w18739;
w18741 <= not pi0706 and not w18740;
w18742 <= not w18736 and w18741;
w18743 <= w18693 and not w18742;
w18744 <= not w18718 and w18743;
w18745 <= not pi0057 and not w18694;
w18746 <= not w18744 and w18745;
w18747 <= not pi0832 and not w18692;
w18748 <= not w18746 and w18747;
w18749 <= pi0706 and w18465;
w18750 <= w489 and not w18719;
w18751 <= not w18749 and w18750;
w18752 <= pi0148 and not w489;
w18753 <= pi0832 and not w18752;
w18754 <= not w18751 and w18753;
w18755 <= not w18748 and not w18754;
w18756 <= not pi0149 and not w489;
w18757 <= not pi0755 and pi0947;
w18758 <= not pi0725 and w18465;
w18759 <= not w18757 and not w18758;
w18760 <= w489 and not w18759;
w18761 <= pi0832 and not w18756;
w18762 <= not w18760 and w18761;
w18763 <= not pi0149 and not w7760;
w18764 <= w14204 and not w18757;
w18765 <= pi0149 and not w14613;
w18766 <= pi0038 and not w18764;
w18767 <= not w18765 and w18766;
w18768 <= not pi0149 and not w14521;
w18769 <= w14521 and w18757;
w18770 <= not pi0039 and not w18768;
w18771 <= not w18769 and w18770;
w18772 <= not pi0149 and not w14587;
w18773 <= w18582 and not w18772;
w18774 <= not pi0149 and not w18564;
w18775 <= not w13679 and not w18592;
w18776 <= not w18774 and not w18775;
w18777 <= not pi0755 and not w18773;
w18778 <= not w18776 and w18777;
w18779 <= not pi0149 and pi0755;
w18780 <= not w14609 and w18779;
w18781 <= pi0039 and not w18780;
w18782 <= not w18778 and w18781;
w18783 <= not pi0038 and not w18771;
w18784 <= not w18782 and w18783;
w18785 <= not w18767 and not w18784;
w18786 <= pi0725 and not w18785;
w18787 <= not w18677 and w18771;
w18788 <= not pi0149 and w18627;
w18789 <= pi0149 and w18643;
w18790 <= not pi0755 and not w18789;
w18791 <= not w18788 and w18790;
w18792 <= not pi0149 and w18656;
w18793 <= pi0149 and not w18700;
w18794 <= pi0755 and not w18657;
w18795 <= not w18793 and w18794;
w18796 <= not w18792 and w18795;
w18797 <= pi0039 and not w18796;
w18798 <= not w18791 and w18797;
w18799 <= not w18787 and not w18798;
w18800 <= not pi0038 and not w18799;
w18801 <= not pi0149 and not w14204;
w18802 <= not w3799 and w14230;
w18803 <= pi0755 and pi0947;
w18804 <= not pi0039 and not w18803;
w18805 <= w18802 and w18804;
w18806 <= pi0038 and not w18801;
w18807 <= not w18805 and w18806;
w18808 <= not pi0725 and not w18807;
w18809 <= not w18800 and w18808;
w18810 <= not w18786 and not w18809;
w18811 <= w7760 and not w18810;
w18812 <= not pi0832 and not w18763;
w18813 <= not w18811 and w18812;
w18814 <= not w18762 and not w18813;
w18815 <= not pi0150 and not w7760;
w18816 <= pi0150 and not w14613;
w18817 <= not pi0751 and pi0947;
w18818 <= w14204 and not w18817;
w18819 <= not w18816 and not w18818;
w18820 <= pi0038 and not w18819;
w18821 <= pi0150 and not w14521;
w18822 <= pi0751 and w14521;
w18823 <= not w18821 and not w18822;
w18824 <= w18552 and w18823;
w18825 <= not pi0150 and w18567;
w18826 <= pi0150 and not w18593;
w18827 <= not pi0751 and not w18826;
w18828 <= not w18825 and w18827;
w18829 <= not pi0150 and pi0751;
w18830 <= not w14609 and w18829;
w18831 <= not w18828 and not w18830;
w18832 <= pi0039 and not w18831;
w18833 <= not pi0038 and not w18824;
w18834 <= not w18832 and w18833;
w18835 <= pi0701 and not w18820;
w18836 <= not w18834 and w18835;
w18837 <= not pi0150 and not w14204;
w18838 <= pi0751 and pi0947;
w18839 <= not pi0039 and not w18838;
w18840 <= w18802 and w18839;
w18841 <= pi0038 and not w18837;
w18842 <= not w18840 and w18841;
w18843 <= w18660 and not w18817;
w18844 <= not pi0039 and not w18821;
w18845 <= not w18843 and w18844;
w18846 <= not pi0150 and not w18658;
w18847 <= pi0150 and not w18675;
w18848 <= pi0751 and not w18847;
w18849 <= not w18846 and w18848;
w18850 <= not pi0150 and w18627;
w18851 <= pi0150 and w18643;
w18852 <= not pi0751 and not w18851;
w18853 <= not w18850 and w18852;
w18854 <= not w18849 and not w18853;
w18855 <= pi0039 and not w18854;
w18856 <= not pi0038 and not w18845;
w18857 <= not w18855 and w18856;
w18858 <= not pi0701 and not w18842;
w18859 <= not w18857 and w18858;
w18860 <= not w18836 and not w18859;
w18861 <= w7760 and not w18860;
w18862 <= not pi0832 and not w18815;
w18863 <= not w18861 and w18862;
w18864 <= not pi0150 and not w489;
w18865 <= not pi0701 and w18465;
w18866 <= not w18817 and not w18865;
w18867 <= w489 and not w18866;
w18868 <= pi0832 and not w18864;
w18869 <= not w18867 and w18868;
w18870 <= not w18863 and not w18869;
w18871 <= not pi0151 and not w489;
w18872 <= not pi0745 and pi0947;
w18873 <= not pi0723 and w18465;
w18874 <= not w18872 and not w18873;
w18875 <= w489 and not w18874;
w18876 <= pi0832 and not w18871;
w18877 <= not w18875 and w18876;
w18878 <= not pi0151 and not w7760;
w18879 <= not pi0151 and not w14204;
w18880 <= pi0745 and pi0947;
w18881 <= not pi0039 and not w18880;
w18882 <= w18802 and w18881;
w18883 <= pi0038 and not w18879;
w18884 <= not w18882 and w18883;
w18885 <= not pi0151 and not w14521;
w18886 <= not pi0745 and w18579;
w18887 <= not w18885 and not w18886;
w18888 <= w18678 and w18887;
w18889 <= not w14604 and not w18562;
w18890 <= not pi0151 and w18889;
w18891 <= not w14600 and not w18890;
w18892 <= pi0215 and not w18891;
w18893 <= pi0151 and not w1011;
w18894 <= not w14595 and w18893;
w18895 <= not w14594 and not w18894;
w18896 <= not pi0151 and not w14216;
w18897 <= w18668 and not w18896;
w18898 <= not w18637 and w18897;
w18899 <= not pi0215 and not w18898;
w18900 <= w18895 and w18899;
w18901 <= not w18892 and not w18900;
w18902 <= pi0299 and not w18901;
w18903 <= pi0151 and not w18634;
w18904 <= w18625 and not w18903;
w18905 <= not w18902 and not w18904;
w18906 <= not pi0745 and not w18905;
w18907 <= w18895 and not w18897;
w18908 <= w18611 and w18907;
w18909 <= not w18892 and not w18908;
w18910 <= not w18584 and not w18909;
w18911 <= pi0299 and not w18910;
w18912 <= not pi0151 and not w14587;
w18913 <= w18674 and not w18912;
w18914 <= pi0745 and not w18913;
w18915 <= not w18911 and w18914;
w18916 <= pi0039 and not w18915;
w18917 <= not w18906 and w18916;
w18918 <= not w18888 and not w18917;
w18919 <= not pi0038 and not w18918;
w18920 <= not pi0723 and not w18884;
w18921 <= not w18919 and w18920;
w18922 <= pi0151 and not w14613;
w18923 <= w14204 and not w18872;
w18924 <= not w18922 and not w18923;
w18925 <= pi0038 and not w18924;
w18926 <= not pi0039 and not w18887;
w18927 <= not pi0745 and not w14588;
w18928 <= not pi0151 and not w14609;
w18929 <= not w18927 and w18928;
w18930 <= w18589 and not w18896;
w18931 <= w18895 and not w18930;
w18932 <= w18559 and w18931;
w18933 <= w18664 and not w18891;
w18934 <= pi0299 and not w18933;
w18935 <= not w18932 and w18934;
w18936 <= not pi0745 and not w18582;
w18937 <= not w18935 and w18936;
w18938 <= not w18929 and not w18937;
w18939 <= pi0039 and not w18938;
w18940 <= not pi0038 and not w18926;
w18941 <= not w18939 and w18940;
w18942 <= pi0723 and not w18925;
w18943 <= not w18941 and w18942;
w18944 <= not w18921 and not w18943;
w18945 <= w7760 and not w18944;
w18946 <= not pi0832 and not w18878;
w18947 <= not w18945 and w18946;
w18948 <= not w18877 and not w18947;
w18949 <= not pi0152 and not w7760;
w18950 <= not pi0152 and not w14204;
w18951 <= pi0759 and pi0947;
w18952 <= not pi0039 and not w18951;
w18953 <= w14230 and not w18465;
w18954 <= w18952 and w18953;
w18955 <= pi0038 and not w18950;
w18956 <= not w18954 and w18955;
w18957 <= pi0152 and not w14521;
w18958 <= not w14522 and not w18952;
w18959 <= not w18957 and not w18958;
w18960 <= not w18677 and w18959;
w18961 <= not pi0152 and not w14600;
w18962 <= w18561 and not w18961;
w18963 <= not w18465 and not w18636;
w18964 <= w18962 and not w18963;
w18965 <= pi0152 and w18609;
w18966 <= w18665 and not w18965;
w18967 <= pi0152 and not w14216;
w18968 <= not w18637 and not w18967;
w18969 <= w1011 and w18968;
w18970 <= not pi0215 and not w18969;
w18971 <= not w18608 and w18970;
w18972 <= not w18966 and w18971;
w18973 <= pi0299 and not w18964;
w18974 <= not w18972 and w18973;
w18975 <= not w18667 and not w18967;
w18976 <= w166 and not w18975;
w18977 <= not pi0152 and not w14583;
w18978 <= w14583 and not w18465;
w18979 <= not w166 and not w18978;
w18980 <= not w18977 and w18979;
w18981 <= not w18976 and not w18980;
w18982 <= not pi0223 and not w18981;
w18983 <= not pi0152 and not w14555;
w18984 <= w18618 and not w18983;
w18985 <= not pi0299 and not w18984;
w18986 <= not w18982 and w18985;
w18987 <= not pi0759 and not w18974;
w18988 <= not w18986 and w18987;
w18989 <= not w14595 and w18966;
w18990 <= w18970 and not w18989;
w18991 <= pi0299 and not w18962;
w18992 <= not w18990 and w18991;
w18993 <= w166 and w18968;
w18994 <= not pi0947 and w14583;
w18995 <= not w166 and not w18994;
w18996 <= not w18977 and w18995;
w18997 <= not w3799 and w14583;
w18998 <= not w166 and not w18997;
w18999 <= not w18996 and w18998;
w19000 <= not pi0223 and not w18993;
w19001 <= not w18999 and w19000;
w19002 <= w18616 and not w18983;
w19003 <= not pi0299 and not w19002;
w19004 <= not w18984 and w19003;
w19005 <= not w19001 and w19004;
w19006 <= pi0759 and not w18992;
w19007 <= not w19005 and w19006;
w19008 <= pi0039 and not w18988;
w19009 <= not w19007 and w19008;
w19010 <= not pi0038 and not w18960;
w19011 <= not w19009 and w19010;
w19012 <= pi0696 and not w18956;
w19013 <= not w19011 and w19012;
w19014 <= not pi0152 and not w14613;
w19015 <= w14204 and not w18951;
w19016 <= pi0038 and not w19015;
w19017 <= not w19014 and w19016;
w19018 <= not w18588 and not w18967;
w19019 <= w166 and not w19018;
w19020 <= not w18996 and not w19019;
w19021 <= not pi0223 and not w19020;
w19022 <= w19003 and not w19021;
w19023 <= pi0152 and w18563;
w19024 <= w1011 and w19018;
w19025 <= not w18558 and not w18966;
w19026 <= not w18586 and not w19025;
w19027 <= not pi0215 and not w19024;
w19028 <= not w19026 and w19027;
w19029 <= w18585 and not w19023;
w19030 <= not w19028 and w19029;
w19031 <= pi0759 and not w19022;
w19032 <= not w19030 and w19031;
w19033 <= not pi0759 and not w14609;
w19034 <= pi0152 and w19033;
w19035 <= pi0039 and not w19034;
w19036 <= not w19032 and w19035;
w19037 <= not pi0038 and not w18959;
w19038 <= not w19036 and w19037;
w19039 <= not pi0696 and not w19017;
w19040 <= not w19038 and w19039;
w19041 <= not w19013 and not w19040;
w19042 <= w7760 and not w19041;
w19043 <= not pi0832 and not w18949;
w19044 <= not w19042 and w19043;
w19045 <= not pi0152 and not w489;
w19046 <= pi0696 and w18465;
w19047 <= w489 and not w18951;
w19048 <= not w19046 and w19047;
w19049 <= pi0832 and not w19045;
w19050 <= not w19048 and w19049;
w19051 <= not w19044 and not w19050;
w19052 <= pi0153 and not w489;
w19053 <= pi0766 and pi0947;
w19054 <= w489 and not w19053;
w19055 <= pi0700 and w18465;
w19056 <= w19054 and not w19055;
w19057 <= pi0832 and not w19052;
w19058 <= not w19056 and w19057;
w19059 <= pi0057 and pi0153;
w19060 <= not pi0153 and not w18693;
w19061 <= not pi0153 and not w14521;
w19062 <= not pi0766 and w15710;
w19063 <= not w18580 and not w19062;
w19064 <= not w19061 and not w19063;
w19065 <= not w18677 and w19064;
w19066 <= not pi0153 and not w14587;
w19067 <= w18674 and not w19066;
w19068 <= pi0153 and not w14600;
w19069 <= w18561 and not w19068;
w19070 <= w18636 and not w19069;
w19071 <= pi0153 and not w1011;
w19072 <= not w14595 and w19071;
w19073 <= not w14594 and not w19072;
w19074 <= not pi0153 and not w14216;
w19075 <= w18668 and not w19074;
w19076 <= not w18610 and not w19075;
w19077 <= w19073 and w19076;
w19078 <= not pi0215 and not w19077;
w19079 <= not w18584 and not w19070;
w19080 <= not w19078 and w19079;
w19081 <= pi0299 and not w19080;
w19082 <= not pi0766 and not w19067;
w19083 <= not w19081 and w19082;
w19084 <= w18589 and not w19074;
w19085 <= not w18666 and w19084;
w19086 <= not pi0215 and not w19085;
w19087 <= w19073 and w19086;
w19088 <= not w19069 and not w19087;
w19089 <= pi0299 and not w19088;
w19090 <= pi0153 and not w18634;
w19091 <= w18625 and not w19090;
w19092 <= not w19089 and not w19091;
w19093 <= pi0766 and not w19092;
w19094 <= pi0039 and not w19083;
w19095 <= not w19093 and w19094;
w19096 <= not w19065 and not w19095;
w19097 <= not pi0038 and not w19096;
w19098 <= not pi0153 and not w14204;
w19099 <= not pi0766 and pi0947;
w19100 <= not pi0039 and not w19099;
w19101 <= w18802 and w19100;
w19102 <= pi0038 and not w19098;
w19103 <= not w19101 and w19102;
w19104 <= not w19097 and not w19103;
w19105 <= pi0700 and not w19104;
w19106 <= w3847 and w19054;
w19107 <= pi0153 and not w14613;
w19108 <= pi0038 and not w19106;
w19109 <= not w19107 and w19108;
w19110 <= w18582 and not w19066;
w19111 <= w18563 and not w19068;
w19112 <= w19073 and not w19084;
w19113 <= w18559 and w19112;
w19114 <= pi0299 and not w19111;
w19115 <= not w19113 and w19114;
w19116 <= pi0766 and not w19115;
w19117 <= not w19110 and w19116;
w19118 <= not pi0153 and not pi0766;
w19119 <= not w14609 and w19118;
w19120 <= pi0039 and not w19119;
w19121 <= not w19117 and w19120;
w19122 <= not pi0038 and not w19064;
w19123 <= not w19121 and w19122;
w19124 <= not pi0700 and not w19109;
w19125 <= not w19123 and w19124;
w19126 <= w18693 and not w19125;
w19127 <= not w19105 and w19126;
w19128 <= not pi0057 and not w19060;
w19129 <= not w19127 and w19128;
w19130 <= not pi0832 and not w19059;
w19131 <= not w19129 and w19130;
w19132 <= not w19058 and not w19131;
w19133 <= not pi0154 and not w489;
w19134 <= not pi0742 and pi0947;
w19135 <= not pi0704 and w18465;
w19136 <= not w19134 and not w19135;
w19137 <= w489 and not w19136;
w19138 <= pi0832 and not w19133;
w19139 <= not w19137 and w19138;
w19140 <= not pi0154 and not w7760;
w19141 <= not pi0154 and not w14204;
w19142 <= w18653 and not w19141;
w19143 <= not pi0154 and not w14521;
w19144 <= w18678 and not w19143;
w19145 <= not pi0154 and w18658;
w19146 <= pi0154 and w18675;
w19147 <= pi0039 and not w19146;
w19148 <= not w19145 and w19147;
w19149 <= not w19144 and not w19148;
w19150 <= not pi0038 and not w19149;
w19151 <= pi0742 and not w19142;
w19152 <= not w19150 and w19151;
w19153 <= w18605 and not w19141;
w19154 <= not w18629 and w19144;
w19155 <= not pi0154 and not w18627;
w19156 <= pi0154 and not w18643;
w19157 <= pi0039 and not w19156;
w19158 <= not w19155 and w19157;
w19159 <= not w19154 and not w19158;
w19160 <= not pi0038 and not w19159;
w19161 <= not pi0742 and not w19153;
w19162 <= not w19160 and w19161;
w19163 <= not pi0704 and not w19152;
w19164 <= not w19162 and w19163;
w19165 <= not pi0154 and not w14613;
w19166 <= not w18578 and not w19165;
w19167 <= w18580 and not w19143;
w19168 <= pi0154 and w18593;
w19169 <= not pi0154 and not w18567;
w19170 <= pi0039 and not w19168;
w19171 <= not w19169 and w19170;
w19172 <= not w19167 and not w19171;
w19173 <= not pi0038 and not w19172;
w19174 <= not pi0742 and not w19166;
w19175 <= not w19173 and w19174;
w19176 <= not pi0154 and pi0742;
w19177 <= not w14615 and w19176;
w19178 <= pi0704 and not w19177;
w19179 <= not w19175 and w19178;
w19180 <= w7760 and not w19179;
w19181 <= not w19164 and w19180;
w19182 <= not pi0832 and not w19140;
w19183 <= not w19181 and w19182;
w19184 <= not w19139 and not w19183;
w19185 <= not pi0757 and w18597;
w19186 <= pi0686 and not w19185;
w19187 <= not pi0038 and not w18645;
w19188 <= not w18605 and not w19187;
w19189 <= not pi0757 and w19188;
w19190 <= not pi0038 and not w18679;
w19191 <= not w18653 and not w19190;
w19192 <= pi0757 and w19191;
w19193 <= not pi0686 and not w19189;
w19194 <= not w19192 and w19193;
w19195 <= w7760 and not w19186;
w19196 <= not w19194 and w19195;
w19197 <= pi0155 and not w19196;
w19198 <= not pi0038 and not w18632;
w19199 <= pi0038 and w18602;
w19200 <= not w19198 and not w19199;
w19201 <= not pi0757 and w19200;
w19202 <= not pi0038 and not w18662;
w19203 <= w14204 and w18653;
w19204 <= not w19202 and not w19203;
w19205 <= pi0757 and w19204;
w19206 <= not pi0686 and not w19201;
w19207 <= not w19205 and w19206;
w19208 <= not pi0757 and w18573;
w19209 <= pi0757 and not w14615;
w19210 <= pi0686 and not w19209;
w19211 <= not w19208 and w19210;
w19212 <= not w19207 and not w19211;
w19213 <= not pi0155 and w7760;
w19214 <= not w19212 and w19213;
w19215 <= not w19197 and not w19214;
w19216 <= not pi0832 and not w19215;
w19217 <= not pi0155 and not w489;
w19218 <= not pi0757 and pi0947;
w19219 <= not pi0686 and w18465;
w19220 <= not w19218 and not w19219;
w19221 <= w489 and not w19220;
w19222 <= pi0832 and not w19217;
w19223 <= not w19221 and w19222;
w19224 <= not w19216 and not w19223;
w19225 <= not pi0156 and not w489;
w19226 <= not pi0741 and pi0947;
w19227 <= not pi0724 and w18465;
w19228 <= not w19226 and not w19227;
w19229 <= w489 and not w19228;
w19230 <= pi0832 and not w19225;
w19231 <= not w19229 and w19230;
w19232 <= not pi0741 and not w19200;
w19233 <= pi0741 and not w19204;
w19234 <= not pi0724 and not w19232;
w19235 <= not w19233 and w19234;
w19236 <= not pi0741 and not w18573;
w19237 <= pi0741 and w14615;
w19238 <= pi0724 and not w19237;
w19239 <= not w19236 and w19238;
w19240 <= w7760 and not w19239;
w19241 <= not w19235 and w19240;
w19242 <= not pi0156 and not w19241;
w19243 <= not pi0741 and not w19188;
w19244 <= pi0741 and not w19191;
w19245 <= not pi0724 and not w19243;
w19246 <= not w19244 and w19245;
w19247 <= pi0724 and not pi0741;
w19248 <= w18597 and w19247;
w19249 <= not w19246 and not w19248;
w19250 <= pi0156 and w7760;
w19251 <= not w19249 and w19250;
w19252 <= not pi0832 and not w19251;
w19253 <= not w19242 and w19252;
w19254 <= not w19231 and not w19253;
w19255 <= not pi0157 and not w489;
w19256 <= not pi0760 and pi0947;
w19257 <= not pi0688 and w18465;
w19258 <= not w19256 and not w19257;
w19259 <= w489 and not w19258;
w19260 <= pi0832 and not w19255;
w19261 <= not w19259 and w19260;
w19262 <= not pi0157 and not w7760;
w19263 <= w14204 and not w19256;
w19264 <= pi0157 and not w14613;
w19265 <= pi0038 and not w19263;
w19266 <= not w19264 and w19265;
w19267 <= not pi0157 and pi0760;
w19268 <= not w14609 and w19267;
w19269 <= not pi0157 and not w14587;
w19270 <= w18582 and not w19269;
w19271 <= not pi0157 and not w18564;
w19272 <= not w11280 and not w18592;
w19273 <= not w19271 and not w19272;
w19274 <= not pi0760 and not w19270;
w19275 <= not w19273 and w19274;
w19276 <= pi0039 and not w19268;
w19277 <= not w19275 and w19276;
w19278 <= not pi0157 and not w14521;
w19279 <= w14521 and w19256;
w19280 <= not pi0039 and not w19278;
w19281 <= not w19279 and w19280;
w19282 <= not pi0038 and not w19281;
w19283 <= not w19277 and w19282;
w19284 <= not w19266 and not w19283;
w19285 <= pi0688 and not w19284;
w19286 <= not w18677 and w19281;
w19287 <= not pi0760 and w18643;
w19288 <= pi0760 and not w18675;
w19289 <= pi0157 and not w19287;
w19290 <= not w19288 and w19289;
w19291 <= pi0760 and not w18658;
w19292 <= not pi0760 and w18627;
w19293 <= not pi0157 and not w19291;
w19294 <= not w19292 and w19293;
w19295 <= pi0039 and not w19290;
w19296 <= not w19294 and w19295;
w19297 <= not w19286 and not w19296;
w19298 <= not pi0038 and not w19297;
w19299 <= not pi0157 and not w14204;
w19300 <= pi0760 and pi0947;
w19301 <= not pi0039 and not w19300;
w19302 <= w18802 and w19301;
w19303 <= pi0038 and not w19299;
w19304 <= not w19302 and w19303;
w19305 <= not pi0688 and not w19304;
w19306 <= not w19298 and w19305;
w19307 <= not w19285 and not w19306;
w19308 <= w7760 and not w19307;
w19309 <= not pi0832 and not w19262;
w19310 <= not w19308 and w19309;
w19311 <= not w19261 and not w19310;
w19312 <= not pi0158 and not w7760;
w19313 <= pi0158 and not w14613;
w19314 <= not pi0753 and pi0947;
w19315 <= w14204 and not w19314;
w19316 <= not w19313 and not w19315;
w19317 <= pi0038 and not w19316;
w19318 <= pi0158 and not w14521;
w19319 <= pi0753 and w14521;
w19320 <= not w19318 and not w19319;
w19321 <= w18552 and w19320;
w19322 <= not pi0158 and w18567;
w19323 <= pi0158 and not w18593;
w19324 <= not pi0753 and not w19323;
w19325 <= not w19322 and w19324;
w19326 <= not pi0158 and pi0753;
w19327 <= not w14609 and w19326;
w19328 <= not w19325 and not w19327;
w19329 <= pi0039 and not w19328;
w19330 <= not pi0038 and not w19321;
w19331 <= not w19329 and w19330;
w19332 <= pi0702 and not w19317;
w19333 <= not w19331 and w19332;
w19334 <= not pi0158 and not w14204;
w19335 <= pi0753 and pi0947;
w19336 <= not pi0039 and not w19335;
w19337 <= w18802 and w19336;
w19338 <= pi0038 and not w19334;
w19339 <= not w19337 and w19338;
w19340 <= w18660 and not w19314;
w19341 <= not pi0039 and not w19318;
w19342 <= not w19340 and w19341;
w19343 <= not pi0158 and not w18658;
w19344 <= pi0158 and not w18675;
w19345 <= pi0753 and not w19344;
w19346 <= not w19343 and w19345;
w19347 <= not pi0158 and w18627;
w19348 <= pi0158 and w18643;
w19349 <= not pi0753 and not w19348;
w19350 <= not w19347 and w19349;
w19351 <= not w19346 and not w19350;
w19352 <= pi0039 and not w19351;
w19353 <= not pi0038 and not w19342;
w19354 <= not w19352 and w19353;
w19355 <= not pi0702 and not w19339;
w19356 <= not w19354 and w19355;
w19357 <= not w19333 and not w19356;
w19358 <= w7760 and not w19357;
w19359 <= not pi0832 and not w19312;
w19360 <= not w19358 and w19359;
w19361 <= not pi0158 and not w489;
w19362 <= not pi0702 and w18465;
w19363 <= not w19314 and not w19362;
w19364 <= w489 and not w19363;
w19365 <= pi0832 and not w19361;
w19366 <= not w19364 and w19365;
w19367 <= not w19360 and not w19366;
w19368 <= not pi0159 and not w7760;
w19369 <= pi0159 and not w14613;
w19370 <= not pi0754 and pi0947;
w19371 <= w14204 and not w19370;
w19372 <= not w19369 and not w19371;
w19373 <= pi0038 and not w19372;
w19374 <= pi0159 and not w14521;
w19375 <= pi0754 and w14521;
w19376 <= not w19374 and not w19375;
w19377 <= w18552 and w19376;
w19378 <= not pi0159 and w18567;
w19379 <= pi0159 and not w18593;
w19380 <= not pi0754 and not w19379;
w19381 <= not w19378 and w19380;
w19382 <= not pi0159 and pi0754;
w19383 <= not w14609 and w19382;
w19384 <= not w19381 and not w19383;
w19385 <= pi0039 and not w19384;
w19386 <= not pi0038 and not w19377;
w19387 <= not w19385 and w19386;
w19388 <= pi0709 and not w19373;
w19389 <= not w19387 and w19388;
w19390 <= not pi0159 and not w14204;
w19391 <= pi0754 and pi0947;
w19392 <= not pi0039 and not w19391;
w19393 <= w18802 and w19392;
w19394 <= pi0038 and not w19390;
w19395 <= not w19393 and w19394;
w19396 <= w18660 and not w19370;
w19397 <= not pi0039 and not w19374;
w19398 <= not w19396 and w19397;
w19399 <= not pi0159 and not w18658;
w19400 <= pi0159 and not w18675;
w19401 <= pi0754 and not w19400;
w19402 <= not w19399 and w19401;
w19403 <= not pi0159 and w18627;
w19404 <= pi0159 and w18643;
w19405 <= not pi0754 and not w19404;
w19406 <= not w19403 and w19405;
w19407 <= not w19402 and not w19406;
w19408 <= pi0039 and not w19407;
w19409 <= not pi0038 and not w19398;
w19410 <= not w19408 and w19409;
w19411 <= not pi0709 and not w19395;
w19412 <= not w19410 and w19411;
w19413 <= not w19389 and not w19412;
w19414 <= w7760 and not w19413;
w19415 <= not pi0832 and not w19368;
w19416 <= not w19414 and w19415;
w19417 <= not pi0159 and not w489;
w19418 <= not pi0709 and w18465;
w19419 <= not w19370 and not w19418;
w19420 <= w489 and not w19419;
w19421 <= pi0832 and not w19417;
w19422 <= not w19420 and w19421;
w19423 <= not w19416 and not w19422;
w19424 <= not pi0160 and not w489;
w19425 <= not pi0756 and pi0947;
w19426 <= not pi0734 and w18465;
w19427 <= not w19425 and not w19426;
w19428 <= w489 and not w19427;
w19429 <= pi0832 and not w19424;
w19430 <= not w19428 and w19429;
w19431 <= not pi0160 and not w7760;
w19432 <= w14204 and not w19425;
w19433 <= pi0160 and not w14613;
w19434 <= pi0038 and not w19432;
w19435 <= not w19433 and w19434;
w19436 <= not pi0160 and not w14521;
w19437 <= w14521 and w19425;
w19438 <= not pi0039 and not w19436;
w19439 <= not w19437 and w19438;
w19440 <= not pi0160 and not w18564;
w19441 <= pi0160 and not w18725;
w19442 <= pi0299 and not w19441;
w19443 <= not w19440 and w19442;
w19444 <= not pi0160 and not w14587;
w19445 <= w18582 and not w19444;
w19446 <= not pi0756 and not w19445;
w19447 <= not w19443 and w19446;
w19448 <= not pi0160 and pi0756;
w19449 <= not w14609 and w19448;
w19450 <= pi0039 and not w19449;
w19451 <= not w19447 and w19450;
w19452 <= not pi0038 and not w19439;
w19453 <= not w19451 and w19452;
w19454 <= not w19435 and not w19453;
w19455 <= pi0734 and not w19454;
w19456 <= not w18677 and w19439;
w19457 <= not pi0160 and w18627;
w19458 <= pi0160 and w18643;
w19459 <= not pi0756 and not w19458;
w19460 <= not w19457 and w19459;
w19461 <= pi0160 and not w18700;
w19462 <= not pi0160 and w18656;
w19463 <= pi0756 and not w18657;
w19464 <= not w19461 and w19463;
w19465 <= not w19462 and w19464;
w19466 <= pi0039 and not w19465;
w19467 <= not w19460 and w19466;
w19468 <= not w19456 and not w19467;
w19469 <= not pi0038 and not w19468;
w19470 <= not pi0160 and not w14204;
w19471 <= pi0756 and pi0947;
w19472 <= not pi0039 and not w19471;
w19473 <= w18802 and w19472;
w19474 <= pi0038 and not w19470;
w19475 <= not w19473 and w19474;
w19476 <= not pi0734 and not w19475;
w19477 <= not w19469 and w19476;
w19478 <= not w19455 and not w19477;
w19479 <= w7760 and not w19478;
w19480 <= not pi0832 and not w19431;
w19481 <= not w19479 and w19480;
w19482 <= not w19430 and not w19481;
w19483 <= not pi0161 and not w7760;
w19484 <= not pi0161 and not w14204;
w19485 <= pi0758 and pi0947;
w19486 <= not pi0039 and not w19485;
w19487 <= w18953 and w19486;
w19488 <= pi0038 and not w19484;
w19489 <= not w19487 and w19488;
w19490 <= w14521 and w19485;
w19491 <= pi0161 and not w14521;
w19492 <= not pi0039 and not w19490;
w19493 <= not w19491 and w19492;
w19494 <= not w18677 and w19493;
w19495 <= not pi0161 and not w14600;
w19496 <= w18561 and not w19495;
w19497 <= not w18963 and w19496;
w19498 <= pi0161 and w18609;
w19499 <= w18665 and not w19498;
w19500 <= pi0161 and not w14216;
w19501 <= not w18637 and not w19500;
w19502 <= w1011 and w19501;
w19503 <= not pi0215 and not w19502;
w19504 <= not w18608 and w19503;
w19505 <= not w19499 and w19504;
w19506 <= pi0299 and not w19497;
w19507 <= not w19505 and w19506;
w19508 <= not w18667 and not w19500;
w19509 <= w166 and not w19508;
w19510 <= not pi0161 and not w14583;
w19511 <= w18979 and not w19510;
w19512 <= not w19509 and not w19511;
w19513 <= not pi0223 and not w19512;
w19514 <= not pi0161 and not w14555;
w19515 <= w18618 and not w19514;
w19516 <= not pi0299 and not w19515;
w19517 <= not w19513 and w19516;
w19518 <= not pi0758 and not w19507;
w19519 <= not w19517 and w19518;
w19520 <= not w14595 and w19499;
w19521 <= w19503 and not w19520;
w19522 <= pi0299 and not w19496;
w19523 <= not w19521 and w19522;
w19524 <= w166 and w19501;
w19525 <= w18995 and not w19510;
w19526 <= w18998 and not w19525;
w19527 <= not pi0223 and not w19524;
w19528 <= not w19526 and w19527;
w19529 <= w18616 and not w19514;
w19530 <= not pi0299 and not w19529;
w19531 <= not w19515 and w19530;
w19532 <= not w19528 and w19531;
w19533 <= pi0758 and not w19523;
w19534 <= not w19532 and w19533;
w19535 <= pi0039 and not w19519;
w19536 <= not w19534 and w19535;
w19537 <= not pi0038 and not w19494;
w19538 <= not w19536 and w19537;
w19539 <= pi0736 and not w19489;
w19540 <= not w19538 and w19539;
w19541 <= not pi0161 and not w14613;
w19542 <= w14204 and not w19485;
w19543 <= pi0038 and not w19542;
w19544 <= not w19541 and w19543;
w19545 <= not w18588 and not w19500;
w19546 <= w166 and not w19545;
w19547 <= not w19525 and not w19546;
w19548 <= not pi0223 and not w19547;
w19549 <= w19530 and not w19548;
w19550 <= pi0161 and w18563;
w19551 <= w1011 and w19545;
w19552 <= not w18558 and not w19499;
w19553 <= not w18586 and not w19552;
w19554 <= not pi0215 and not w19551;
w19555 <= not w19553 and w19554;
w19556 <= w18585 and not w19550;
w19557 <= not w19555 and w19556;
w19558 <= pi0758 and not w19549;
w19559 <= not w19557 and w19558;
w19560 <= pi0161 and w17521;
w19561 <= pi0039 and not w19560;
w19562 <= not w19559 and w19561;
w19563 <= not pi0038 and not w19493;
w19564 <= not w19562 and w19563;
w19565 <= not pi0736 and not w19544;
w19566 <= not w19564 and w19565;
w19567 <= not w19540 and not w19566;
w19568 <= w7760 and not w19567;
w19569 <= not pi0832 and not w19483;
w19570 <= not w19568 and w19569;
w19571 <= not pi0161 and not w489;
w19572 <= pi0736 and w18465;
w19573 <= w489 and not w19485;
w19574 <= not w19572 and w19573;
w19575 <= pi0832 and not w19571;
w19576 <= not w19574 and w19575;
w19577 <= not w19570 and not w19576;
w19578 <= not pi0162 and not w7760;
w19579 <= not pi0761 and pi0947;
w19580 <= w14204 and not w19579;
w19581 <= pi0162 and not w14613;
w19582 <= pi0038 and not w19580;
w19583 <= not w19581 and w19582;
w19584 <= not pi0162 and not w14521;
w19585 <= w14521 and w19579;
w19586 <= not pi0039 and not w19584;
w19587 <= not w19585 and w19586;
w19588 <= w12496 and not w18725;
w19589 <= not w18554 and not w19588;
w19590 <= not pi0761 and not w19589;
w19591 <= not pi0761 and w18566;
w19592 <= pi0761 and w14609;
w19593 <= not pi0162 and not w19592;
w19594 <= not w19591 and w19593;
w19595 <= pi0039 and not w19590;
w19596 <= not w19594 and w19595;
w19597 <= not pi0038 and not w19587;
w19598 <= not w19596 and w19597;
w19599 <= not w19583 and not w19598;
w19600 <= pi0738 and not w19599;
w19601 <= not w18677 and w19587;
w19602 <= pi0162 and not w18700;
w19603 <= not w12496 and not w18658;
w19604 <= pi0761 and not w19602;
w19605 <= not w19603 and w19604;
w19606 <= not pi0162 and w18627;
w19607 <= pi0162 and w18643;
w19608 <= not pi0761 and not w19607;
w19609 <= not w19606 and w19608;
w19610 <= pi0039 and not w19605;
w19611 <= not w19609 and w19610;
w19612 <= not w19601 and not w19611;
w19613 <= not pi0038 and not w19612;
w19614 <= not pi0162 and not w14204;
w19615 <= pi0761 and pi0947;
w19616 <= not pi0039 and not w19615;
w19617 <= w18802 and w19616;
w19618 <= pi0038 and not w19614;
w19619 <= not w19617 and w19618;
w19620 <= not pi0738 and not w19619;
w19621 <= not w19613 and w19620;
w19622 <= not w19600 and not w19621;
w19623 <= w7760 and not w19622;
w19624 <= not pi0832 and not w19578;
w19625 <= not w19623 and w19624;
w19626 <= not pi0162 and not w489;
w19627 <= not pi0738 and w18465;
w19628 <= not w19579 and not w19627;
w19629 <= w489 and not w19628;
w19630 <= pi0832 and not w19626;
w19631 <= not w19629 and w19630;
w19632 <= not w19625 and not w19631;
w19633 <= not pi0163 and not w489;
w19634 <= not pi0777 and pi0947;
w19635 <= not pi0737 and w18465;
w19636 <= not w19634 and not w19635;
w19637 <= w489 and not w19636;
w19638 <= pi0832 and not w19633;
w19639 <= not w19637 and w19638;
w19640 <= not pi0163 and not w7760;
w19641 <= w14204 and not w19634;
w19642 <= pi0163 and not w14613;
w19643 <= pi0038 and not w19641;
w19644 <= not w19642 and w19643;
w19645 <= not pi0163 and not w14521;
w19646 <= w14521 and w19634;
w19647 <= not pi0039 and not w19645;
w19648 <= not w19646 and w19647;
w19649 <= not pi0163 and not w14587;
w19650 <= w18582 and not w19649;
w19651 <= not pi0163 and not w18564;
w19652 <= not w12298 and not w18592;
w19653 <= not w19651 and not w19652;
w19654 <= not pi0777 and not w19650;
w19655 <= not w19653 and w19654;
w19656 <= not pi0163 and pi0777;
w19657 <= not w14609 and w19656;
w19658 <= pi0039 and not w19657;
w19659 <= not w19655 and w19658;
w19660 <= not pi0038 and not w19648;
w19661 <= not w19659 and w19660;
w19662 <= not w19644 and not w19661;
w19663 <= pi0737 and not w19662;
w19664 <= not w18677 and w19648;
w19665 <= not pi0163 and w18627;
w19666 <= pi0163 and w18643;
w19667 <= not pi0777 and not w19666;
w19668 <= not w19665 and w19667;
w19669 <= not pi0163 and w18656;
w19670 <= pi0163 and not w18700;
w19671 <= pi0777 and not w18657;
w19672 <= not w19670 and w19671;
w19673 <= not w19669 and w19672;
w19674 <= pi0039 and not w19673;
w19675 <= not w19668 and w19674;
w19676 <= not w19664 and not w19675;
w19677 <= not pi0038 and not w19676;
w19678 <= not pi0163 and not w14204;
w19679 <= pi0777 and pi0947;
w19680 <= not pi0039 and not w19679;
w19681 <= w18802 and w19680;
w19682 <= pi0038 and not w19678;
w19683 <= not w19681 and w19682;
w19684 <= not pi0737 and not w19683;
w19685 <= not w19677 and w19684;
w19686 <= not w19663 and not w19685;
w19687 <= w7760 and not w19686;
w19688 <= not pi0832 and not w19640;
w19689 <= not w19687 and w19688;
w19690 <= not w19639 and not w19689;
w19691 <= not pi0164 and not w489;
w19692 <= not pi0752 and pi0947;
w19693 <= pi0703 and w18465;
w19694 <= not w19692 and not w19693;
w19695 <= w489 and not w19694;
w19696 <= pi0832 and not w19691;
w19697 <= not w19695 and w19696;
w19698 <= not pi0164 and not w7760;
w19699 <= not pi0164 and not w18602;
w19700 <= w18605 and not w19699;
w19701 <= not pi0164 and w18632;
w19702 <= pi0164 and w18645;
w19703 <= not pi0038 and not w19702;
w19704 <= not w19701 and w19703;
w19705 <= not pi0752 and not w19700;
w19706 <= not w19704 and w19705;
w19707 <= not pi0164 and not w14204;
w19708 <= w18653 and not w19707;
w19709 <= not pi0164 and w18662;
w19710 <= pi0164 and w18679;
w19711 <= not pi0038 and not w19710;
w19712 <= not w19709 and w19711;
w19713 <= pi0752 and not w19708;
w19714 <= not w19712 and w19713;
w19715 <= not w19706 and not w19714;
w19716 <= pi0703 and not w19715;
w19717 <= pi0752 and w14615;
w19718 <= not pi0752 and w18597;
w19719 <= pi0164 and not w19718;
w19720 <= pi0164 and not w18572;
w19721 <= not pi0752 and not w19720;
w19722 <= not w18573 and w19721;
w19723 <= not pi0703 and not w19717;
w19724 <= not w19719 and w19723;
w19725 <= not w19722 and w19724;
w19726 <= not w19716 and not w19725;
w19727 <= w7760 and not w19726;
w19728 <= not pi0832 and not w19698;
w19729 <= not w19727 and w19728;
w19730 <= not w19697 and not w19729;
w19731 <= not pi0165 and not w489;
w19732 <= not pi0774 and pi0947;
w19733 <= pi0687 and w18465;
w19734 <= not w19732 and not w19733;
w19735 <= w489 and not w19734;
w19736 <= pi0832 and not w19731;
w19737 <= not w19735 and w19736;
w19738 <= not pi0165 and not w7760;
w19739 <= not pi0165 and not w18602;
w19740 <= w18605 and not w19739;
w19741 <= not pi0165 and w18632;
w19742 <= pi0165 and w18645;
w19743 <= not pi0038 and not w19742;
w19744 <= not w19741 and w19743;
w19745 <= not pi0774 and not w19740;
w19746 <= not w19744 and w19745;
w19747 <= not pi0165 and not w14204;
w19748 <= w18653 and not w19747;
w19749 <= not pi0165 and w18662;
w19750 <= pi0165 and w18679;
w19751 <= not pi0038 and not w19750;
w19752 <= not w19749 and w19751;
w19753 <= pi0774 and not w19748;
w19754 <= not w19752 and w19753;
w19755 <= not w19746 and not w19754;
w19756 <= pi0687 and not w19755;
w19757 <= pi0774 and w14615;
w19758 <= not pi0774 and w18597;
w19759 <= pi0165 and not w19758;
w19760 <= pi0165 and not w18572;
w19761 <= not pi0774 and not w19760;
w19762 <= not w18573 and w19761;
w19763 <= not pi0687 and not w19757;
w19764 <= not w19759 and w19763;
w19765 <= not w19762 and w19764;
w19766 <= not w19756 and not w19765;
w19767 <= w7760 and not w19766;
w19768 <= not pi0832 and not w19738;
w19769 <= not w19767 and w19768;
w19770 <= not w19737 and not w19769;
w19771 <= not pi0166 and not w7760;
w19772 <= not pi0166 and not w14613;
w19773 <= pi0772 and pi0947;
w19774 <= w14204 and not w19773;
w19775 <= pi0038 and not w19774;
w19776 <= not w19772 and w19775;
w19777 <= pi0166 and not w14521;
w19778 <= not pi0039 and not w19773;
w19779 <= not w14522 and not w19778;
w19780 <= not w19777 and not w19779;
w19781 <= not pi0166 and not w14555;
w19782 <= w18616 and not w19781;
w19783 <= not pi0299 and not w19782;
w19784 <= pi0166 and not w14216;
w19785 <= not w18588 and not w19784;
w19786 <= w166 and not w19785;
w19787 <= not pi0166 and not w14583;
w19788 <= w18995 and not w19787;
w19789 <= not w19786 and not w19788;
w19790 <= not pi0223 and not w19789;
w19791 <= w19783 and not w19790;
w19792 <= pi0166 and w18563;
w19793 <= w1011 and w19785;
w19794 <= pi0166 and w18609;
w19795 <= w18665 and not w19794;
w19796 <= not w18558 and not w19795;
w19797 <= not w18586 and not w19796;
w19798 <= not pi0215 and not w19793;
w19799 <= not w19797 and w19798;
w19800 <= w18585 and not w19792;
w19801 <= not w19799 and w19800;
w19802 <= pi0772 and not w19791;
w19803 <= not w19801 and w19802;
w19804 <= not pi0772 and not w14609;
w19805 <= pi0166 and w19804;
w19806 <= pi0039 and not w19805;
w19807 <= not w19803 and w19806;
w19808 <= not pi0038 and not w19780;
w19809 <= not w19807 and w19808;
w19810 <= not pi0727 and not w19776;
w19811 <= not w19809 and w19810;
w19812 <= w18953 and w19778;
w19813 <= not pi0166 and not w14204;
w19814 <= pi0038 and not w19812;
w19815 <= not w19813 and w19814;
w19816 <= not w18677 and w19780;
w19817 <= not w3799 and w14555;
w19818 <= not pi0166 and not w19817;
w19819 <= w18618 and not w19818;
w19820 <= not w18637 and not w19784;
w19821 <= w166 and w19820;
w19822 <= not pi0223 and not w19821;
w19823 <= not w18978 and not w19787;
w19824 <= w18998 and not w19823;
w19825 <= w19822 and not w19824;
w19826 <= w19783 and not w19819;
w19827 <= not w19825 and w19826;
w19828 <= not pi0166 and not w14600;
w19829 <= w18561 and not w19828;
w19830 <= w1011 and w19820;
w19831 <= not pi0215 and not w19830;
w19832 <= not w14595 and w19795;
w19833 <= w19831 and not w19832;
w19834 <= pi0299 and not w19829;
w19835 <= not w19833 and w19834;
w19836 <= pi0772 and not w19827;
w19837 <= not w19835 and w19836;
w19838 <= not w166 and not w19823;
w19839 <= w166 and w18588;
w19840 <= w19822 and not w19839;
w19841 <= not w19838 and w19840;
w19842 <= not pi0299 and not w19819;
w19843 <= not w19841 and w19842;
w19844 <= not w18608 and w19831;
w19845 <= not w19795 and w19844;
w19846 <= not w18963 and w19829;
w19847 <= pi0299 and not w19846;
w19848 <= not w19845 and w19847;
w19849 <= not pi0772 and not w19843;
w19850 <= not w19848 and w19849;
w19851 <= pi0039 and not w19837;
w19852 <= not w19850 and w19851;
w19853 <= not pi0038 and not w19816;
w19854 <= not w19852 and w19853;
w19855 <= pi0727 and not w19815;
w19856 <= not w19854 and w19855;
w19857 <= not w19811 and not w19856;
w19858 <= w7760 and not w19857;
w19859 <= not pi0832 and not w19771;
w19860 <= not w19858 and w19859;
w19861 <= not pi0166 and not w489;
w19862 <= pi0727 and w18465;
w19863 <= w489 and not w19773;
w19864 <= not w19862 and w19863;
w19865 <= pi0832 and not w19861;
w19866 <= not w19864 and w19865;
w19867 <= not w19860 and not w19866;
w19868 <= not pi0167 and not w489;
w19869 <= not pi0768 and pi0947;
w19870 <= pi0705 and w18465;
w19871 <= not w19869 and not w19870;
w19872 <= w489 and not w19871;
w19873 <= pi0832 and not w19868;
w19874 <= not w19872 and w19873;
w19875 <= not pi0167 and not w7760;
w19876 <= pi0768 and not w14615;
w19877 <= not pi0167 and w19876;
w19878 <= not pi0167 and not w14613;
w19879 <= not w18578 and not w19878;
w19880 <= pi0167 and w18595;
w19881 <= not pi0167 and not w18569;
w19882 <= not pi0038 and not w19880;
w19883 <= not w19881 and w19882;
w19884 <= not pi0768 and not w19879;
w19885 <= not w19883 and w19884;
w19886 <= not pi0705 and not w19877;
w19887 <= not w19885 and w19886;
w19888 <= not pi0167 and not w14204;
w19889 <= w18653 and not w19888;
w19890 <= not pi0167 and w18662;
w19891 <= pi0167 and w18679;
w19892 <= not pi0038 and not w19891;
w19893 <= not w19890 and w19892;
w19894 <= pi0768 and not w19889;
w19895 <= not w19893 and w19894;
w19896 <= not pi0167 and not w18602;
w19897 <= w18605 and not w19896;
w19898 <= not pi0167 and w18632;
w19899 <= pi0167 and w18645;
w19900 <= not pi0038 and not w19899;
w19901 <= not w19898 and w19900;
w19902 <= not pi0768 and not w19897;
w19903 <= not w19901 and w19902;
w19904 <= pi0705 and not w19895;
w19905 <= not w19903 and w19904;
w19906 <= w7760 and not w19887;
w19907 <= not w19905 and w19906;
w19908 <= not pi0832 and not w19875;
w19909 <= not w19907 and w19908;
w19910 <= not w19874 and not w19909;
w19911 <= pi0168 and not w489;
w19912 <= pi0763 and pi0947;
w19913 <= w489 and not w19912;
w19914 <= pi0699 and w18465;
w19915 <= w19913 and not w19914;
w19916 <= pi0832 and not w19911;
w19917 <= not w19915 and w19916;
w19918 <= pi0057 and pi0168;
w19919 <= not pi0168 and not w18693;
w19920 <= not pi0168 and not w14521;
w19921 <= not pi0763 and w15710;
w19922 <= not w18580 and not w19921;
w19923 <= not w19920 and not w19922;
w19924 <= not w18677 and w19923;
w19925 <= not pi0168 and not w14587;
w19926 <= w18674 and not w19925;
w19927 <= pi0168 and not w14600;
w19928 <= w18561 and not w19927;
w19929 <= w18636 and not w19928;
w19930 <= pi0168 and not w1011;
w19931 <= not w14595 and w19930;
w19932 <= not w14594 and not w19931;
w19933 <= not pi0168 and not w14216;
w19934 <= w18668 and not w19933;
w19935 <= not w18610 and not w19934;
w19936 <= w19932 and w19935;
w19937 <= not pi0215 and not w19936;
w19938 <= not w18584 and not w19929;
w19939 <= not w19937 and w19938;
w19940 <= pi0299 and not w19939;
w19941 <= not pi0763 and not w19926;
w19942 <= not w19940 and w19941;
w19943 <= w18589 and not w19933;
w19944 <= not w18666 and w19943;
w19945 <= not pi0215 and not w19944;
w19946 <= w19932 and w19945;
w19947 <= not w19928 and not w19946;
w19948 <= pi0299 and not w19947;
w19949 <= pi0168 and not w18634;
w19950 <= w18625 and not w19949;
w19951 <= not w19948 and not w19950;
w19952 <= pi0763 and not w19951;
w19953 <= pi0039 and not w19942;
w19954 <= not w19952 and w19953;
w19955 <= not w19924 and not w19954;
w19956 <= not pi0038 and not w19955;
w19957 <= not pi0168 and not w14204;
w19958 <= not pi0763 and pi0947;
w19959 <= not pi0039 and not w19958;
w19960 <= w18802 and w19959;
w19961 <= pi0038 and not w19957;
w19962 <= not w19960 and w19961;
w19963 <= not w19956 and not w19962;
w19964 <= pi0699 and not w19963;
w19965 <= w3847 and w19913;
w19966 <= pi0168 and not w14613;
w19967 <= pi0038 and not w19965;
w19968 <= not w19966 and w19967;
w19969 <= w18582 and not w19925;
w19970 <= w18563 and not w19927;
w19971 <= w19932 and not w19943;
w19972 <= w18559 and w19971;
w19973 <= pi0299 and not w19970;
w19974 <= not w19972 and w19973;
w19975 <= pi0763 and not w19974;
w19976 <= not w19969 and w19975;
w19977 <= not pi0168 and not pi0763;
w19978 <= not w14609 and w19977;
w19979 <= pi0039 and not w19978;
w19980 <= not w19976 and w19979;
w19981 <= not pi0038 and not w19923;
w19982 <= not w19980 and w19981;
w19983 <= not pi0699 and not w19968;
w19984 <= not w19982 and w19983;
w19985 <= w18693 and not w19984;
w19986 <= not w19964 and w19985;
w19987 <= not pi0057 and not w19919;
w19988 <= not w19986 and w19987;
w19989 <= not pi0832 and not w19918;
w19990 <= not w19988 and w19989;
w19991 <= not w19917 and not w19990;
w19992 <= pi0169 and not w489;
w19993 <= pi0746 and pi0947;
w19994 <= w489 and not w19993;
w19995 <= pi0729 and w18465;
w19996 <= w19994 and not w19995;
w19997 <= pi0832 and not w19992;
w19998 <= not w19996 and w19997;
w19999 <= pi0057 and pi0169;
w20000 <= not pi0169 and not w18693;
w20001 <= not pi0169 and not w14521;
w20002 <= not pi0746 and w15710;
w20003 <= not w18580 and not w20002;
w20004 <= not w20001 and not w20003;
w20005 <= not w18677 and w20004;
w20006 <= not pi0169 and not w14587;
w20007 <= w18674 and not w20006;
w20008 <= pi0169 and not w14600;
w20009 <= w18561 and not w20008;
w20010 <= w18636 and not w20009;
w20011 <= pi0169 and not w1011;
w20012 <= not w14595 and w20011;
w20013 <= not w14594 and not w20012;
w20014 <= not pi0169 and not w14216;
w20015 <= w18668 and not w20014;
w20016 <= not w18610 and not w20015;
w20017 <= w20013 and w20016;
w20018 <= not pi0215 and not w20017;
w20019 <= not w18584 and not w20010;
w20020 <= not w20018 and w20019;
w20021 <= pi0299 and not w20020;
w20022 <= not pi0746 and not w20007;
w20023 <= not w20021 and w20022;
w20024 <= w18589 and not w20014;
w20025 <= not w18666 and w20024;
w20026 <= not pi0215 and not w20025;
w20027 <= w20013 and w20026;
w20028 <= not w20009 and not w20027;
w20029 <= pi0299 and not w20028;
w20030 <= pi0169 and not w18634;
w20031 <= w18625 and not w20030;
w20032 <= not w20029 and not w20031;
w20033 <= pi0746 and not w20032;
w20034 <= pi0039 and not w20023;
w20035 <= not w20033 and w20034;
w20036 <= not w20005 and not w20035;
w20037 <= not pi0038 and not w20036;
w20038 <= not pi0169 and not w14204;
w20039 <= not pi0746 and pi0947;
w20040 <= not pi0039 and not w20039;
w20041 <= w18802 and w20040;
w20042 <= pi0038 and not w20038;
w20043 <= not w20041 and w20042;
w20044 <= not w20037 and not w20043;
w20045 <= pi0729 and not w20044;
w20046 <= w3847 and w19994;
w20047 <= pi0169 and not w14613;
w20048 <= pi0038 and not w20046;
w20049 <= not w20047 and w20048;
w20050 <= w18582 and not w20006;
w20051 <= w18563 and not w20008;
w20052 <= w20013 and not w20024;
w20053 <= w18559 and w20052;
w20054 <= pi0299 and not w20051;
w20055 <= not w20053 and w20054;
w20056 <= pi0746 and not w20055;
w20057 <= not w20050 and w20056;
w20058 <= not pi0169 and not pi0746;
w20059 <= not w14609 and w20058;
w20060 <= pi0039 and not w20059;
w20061 <= not w20057 and w20060;
w20062 <= not pi0038 and not w20004;
w20063 <= not w20061 and w20062;
w20064 <= not pi0729 and not w20049;
w20065 <= not w20063 and w20064;
w20066 <= w18693 and not w20065;
w20067 <= not w20045 and w20066;
w20068 <= not pi0057 and not w20000;
w20069 <= not w20067 and w20068;
w20070 <= not pi0832 and not w19999;
w20071 <= not w20069 and w20070;
w20072 <= not w19998 and not w20071;
w20073 <= pi0730 and w18465;
w20074 <= pi0748 and pi0947;
w20075 <= w489 and not w20074;
w20076 <= not w20073 and w20075;
w20077 <= pi0170 and not w489;
w20078 <= pi0832 and not w20077;
w20079 <= not w20076 and w20078;
w20080 <= pi0057 and pi0170;
w20081 <= not pi0170 and not w18693;
w20082 <= not pi0170 and not w14204;
w20083 <= w18653 and not w20082;
w20084 <= pi0170 and not w14600;
w20085 <= w18561 and not w20084;
w20086 <= w18636 and not w20085;
w20087 <= pi0170 and not w1011;
w20088 <= not w14595 and w20087;
w20089 <= not w14594 and not w20088;
w20090 <= not pi0170 and not w14216;
w20091 <= w18668 and not w20090;
w20092 <= not w18610 and not w20091;
w20093 <= w20089 and w20092;
w20094 <= not pi0215 and not w20093;
w20095 <= not w18584 and not w20086;
w20096 <= not w20094 and w20095;
w20097 <= pi0299 and not w20096;
w20098 <= not pi0170 and not w14587;
w20099 <= not pi0299 and not w20098;
w20100 <= not w18673 and w20099;
w20101 <= not w20097 and not w20100;
w20102 <= pi0039 and not w20101;
w20103 <= not pi0170 and not w14521;
w20104 <= w18678 and not w20103;
w20105 <= not w20102 and not w20104;
w20106 <= not pi0038 and not w20105;
w20107 <= not pi0748 and not w20083;
w20108 <= not w20106 and w20107;
w20109 <= w18605 and not w20082;
w20110 <= w18630 and not w20103;
w20111 <= w18589 and not w20090;
w20112 <= not w18666 and w20111;
w20113 <= not pi0215 and not w20112;
w20114 <= w20089 and w20113;
w20115 <= not w20085 and not w20114;
w20116 <= pi0299 and not w20115;
w20117 <= pi0170 and not w18634;
w20118 <= w18625 and not w20117;
w20119 <= pi0039 and not w20116;
w20120 <= not w20118 and w20119;
w20121 <= not w20110 and not w20120;
w20122 <= not pi0038 and not w20121;
w20123 <= pi0748 and not w20109;
w20124 <= not w20122 and w20123;
w20125 <= pi0730 and not w20124;
w20126 <= not w20108 and w20125;
w20127 <= not pi0170 and not w14613;
w20128 <= not w18578 and not w20127;
w20129 <= w18580 and not w20103;
w20130 <= w18563 and not w20084;
w20131 <= w20089 and not w20111;
w20132 <= w18559 and w20131;
w20133 <= pi0299 and not w20130;
w20134 <= not w20132 and w20133;
w20135 <= not w18581 and w20099;
w20136 <= not w20134 and not w20135;
w20137 <= pi0039 and not w20136;
w20138 <= not w20129 and not w20137;
w20139 <= not pi0038 and not w20138;
w20140 <= pi0748 and not w20128;
w20141 <= not w20139 and w20140;
w20142 <= not pi0170 and not pi0748;
w20143 <= not w14615 and w20142;
w20144 <= not pi0730 and not w20143;
w20145 <= not w20141 and w20144;
w20146 <= w18693 and not w20145;
w20147 <= not w20126 and w20146;
w20148 <= not pi0057 and not w20081;
w20149 <= not w20147 and w20148;
w20150 <= not pi0832 and not w20080;
w20151 <= not w20149 and w20150;
w20152 <= not w20079 and not w20151;
w20153 <= pi0171 and not w489;
w20154 <= pi0764 and pi0947;
w20155 <= w489 and not w20154;
w20156 <= pi0691 and w18465;
w20157 <= w20155 and not w20156;
w20158 <= pi0832 and not w20153;
w20159 <= not w20157 and w20158;
w20160 <= pi0057 and pi0171;
w20161 <= not pi0171 and not w18693;
w20162 <= not pi0171 and not w14521;
w20163 <= not pi0764 and w15710;
w20164 <= not w18580 and not w20163;
w20165 <= not w20162 and not w20164;
w20166 <= not w18677 and w20165;
w20167 <= not pi0171 and not w14587;
w20168 <= w18674 and not w20167;
w20169 <= pi0171 and not w14600;
w20170 <= w18561 and not w20169;
w20171 <= w18636 and not w20170;
w20172 <= pi0171 and not w1011;
w20173 <= not w14595 and w20172;
w20174 <= not w14594 and not w20173;
w20175 <= not pi0171 and not w14216;
w20176 <= w18668 and not w20175;
w20177 <= not w18610 and not w20176;
w20178 <= w20174 and w20177;
w20179 <= not pi0215 and not w20178;
w20180 <= not w18584 and not w20171;
w20181 <= not w20179 and w20180;
w20182 <= pi0299 and not w20181;
w20183 <= not pi0764 and not w20168;
w20184 <= not w20182 and w20183;
w20185 <= w18589 and not w20175;
w20186 <= not w18666 and w20185;
w20187 <= not pi0215 and not w20186;
w20188 <= w20174 and w20187;
w20189 <= not w20170 and not w20188;
w20190 <= pi0299 and not w20189;
w20191 <= pi0171 and not w18634;
w20192 <= w18625 and not w20191;
w20193 <= not w20190 and not w20192;
w20194 <= pi0764 and not w20193;
w20195 <= pi0039 and not w20184;
w20196 <= not w20194 and w20195;
w20197 <= not w20166 and not w20196;
w20198 <= not pi0038 and not w20197;
w20199 <= not pi0171 and not w14204;
w20200 <= not pi0764 and pi0947;
w20201 <= not pi0039 and not w20200;
w20202 <= w18802 and w20201;
w20203 <= pi0038 and not w20199;
w20204 <= not w20202 and w20203;
w20205 <= not w20198 and not w20204;
w20206 <= pi0691 and not w20205;
w20207 <= w3847 and w20155;
w20208 <= pi0171 and not w14613;
w20209 <= pi0038 and not w20207;
w20210 <= not w20208 and w20209;
w20211 <= w18582 and not w20167;
w20212 <= w18563 and not w20169;
w20213 <= w20174 and not w20185;
w20214 <= w18559 and w20213;
w20215 <= pi0299 and not w20212;
w20216 <= not w20214 and w20215;
w20217 <= pi0764 and not w20216;
w20218 <= not w20211 and w20217;
w20219 <= not pi0171 and not pi0764;
w20220 <= not w14609 and w20219;
w20221 <= pi0039 and not w20220;
w20222 <= not w20218 and w20221;
w20223 <= not pi0038 and not w20165;
w20224 <= not w20222 and w20223;
w20225 <= not pi0691 and not w20210;
w20226 <= not w20224 and w20225;
w20227 <= w18693 and not w20226;
w20228 <= not w20206 and w20227;
w20229 <= not pi0057 and not w20161;
w20230 <= not w20228 and w20229;
w20231 <= not pi0832 and not w20160;
w20232 <= not w20230 and w20231;
w20233 <= not w20159 and not w20232;
w20234 <= pi0172 and not w489;
w20235 <= pi0739 and pi0947;
w20236 <= w489 and not w20235;
w20237 <= pi0690 and w18465;
w20238 <= w20236 and not w20237;
w20239 <= pi0832 and not w20234;
w20240 <= not w20238 and w20239;
w20241 <= pi0057 and pi0172;
w20242 <= not pi0172 and not w18693;
w20243 <= not pi0172 and not w14521;
w20244 <= w14521 and w20235;
w20245 <= not pi0039 and not w20243;
w20246 <= not w20244 and w20245;
w20247 <= not w18677 and w20246;
w20248 <= not pi0172 and not w14587;
w20249 <= w18674 and not w20248;
w20250 <= pi0172 and not w14600;
w20251 <= w18561 and not w20250;
w20252 <= w18636 and not w20251;
w20253 <= pi0172 and not w1011;
w20254 <= not w14595 and w20253;
w20255 <= not w14594 and not w20254;
w20256 <= not pi0172 and not w14216;
w20257 <= w18668 and not w20256;
w20258 <= not w18610 and not w20257;
w20259 <= w20255 and w20258;
w20260 <= not pi0215 and not w20259;
w20261 <= not w18584 and not w20252;
w20262 <= not w20260 and w20261;
w20263 <= pi0299 and not w20262;
w20264 <= not pi0739 and not w20249;
w20265 <= not w20263 and w20264;
w20266 <= w18589 and not w20256;
w20267 <= not w18666 and w20266;
w20268 <= not pi0215 and not w20267;
w20269 <= w20255 and w20268;
w20270 <= not w20251 and not w20269;
w20271 <= pi0299 and not w20270;
w20272 <= pi0172 and not w18634;
w20273 <= w18625 and not w20272;
w20274 <= not w20271 and not w20273;
w20275 <= pi0739 and not w20274;
w20276 <= pi0039 and not w20265;
w20277 <= not w20275 and w20276;
w20278 <= not w20247 and not w20277;
w20279 <= not pi0038 and not w20278;
w20280 <= not pi0172 and not w14204;
w20281 <= not pi0739 and pi0947;
w20282 <= not pi0039 and not w20281;
w20283 <= w18802 and w20282;
w20284 <= pi0038 and not w20280;
w20285 <= not w20283 and w20284;
w20286 <= not w20279 and not w20285;
w20287 <= pi0690 and not w20286;
w20288 <= w3847 and w20236;
w20289 <= pi0172 and not w14613;
w20290 <= pi0038 and not w20288;
w20291 <= not w20289 and w20290;
w20292 <= w18582 and not w20248;
w20293 <= w18563 and not w20250;
w20294 <= w20255 and not w20266;
w20295 <= w18559 and w20294;
w20296 <= pi0299 and not w20293;
w20297 <= not w20295 and w20296;
w20298 <= pi0739 and not w20297;
w20299 <= not w20292 and w20298;
w20300 <= not pi0172 and not pi0739;
w20301 <= not w14609 and w20300;
w20302 <= pi0039 and not w20301;
w20303 <= not w20299 and w20302;
w20304 <= not pi0038 and not w20246;
w20305 <= not w20303 and w20304;
w20306 <= not pi0690 and not w20291;
w20307 <= not w20305 and w20306;
w20308 <= w18693 and not w20307;
w20309 <= not w20287 and w20308;
w20310 <= not pi0057 and not w20242;
w20311 <= not w20309 and w20310;
w20312 <= not pi0832 and not w20241;
w20313 <= not w20311 and w20312;
w20314 <= not w20240 and not w20313;
w20315 <= not pi0173 and not w4989;
w20316 <= not pi0173 and not w14622;
w20317 <= w14198 and not w20316;
w20318 <= not pi0723 and w134;
w20319 <= w20316 and not w20318;
w20320 <= not pi0173 and not w14204;
w20321 <= w14210 and not w20320;
w20322 <= pi0173 and not w15639;
w20323 <= not pi0038 and not w20322;
w20324 <= w134 and not w20323;
w20325 <= not pi0173 and w15635;
w20326 <= not w20324 and not w20325;
w20327 <= not pi0723 and not w20321;
w20328 <= not w20326 and w20327;
w20329 <= not w20319 and not w20328;
w20330 <= not pi0778 and w20329;
w20331 <= not pi0625 and w20316;
w20332 <= pi0625 and not w20329;
w20333 <= pi1153 and not w20331;
w20334 <= not w20332 and w20333;
w20335 <= pi0625 and w20316;
w20336 <= not pi0625 and not w20329;
w20337 <= not pi1153 and not w20335;
w20338 <= not w20336 and w20337;
w20339 <= not w20334 and not w20338;
w20340 <= pi0778 and not w20339;
w20341 <= not w20330 and not w20340;
w20342 <= not w14638 and not w20341;
w20343 <= w14638 and not w20316;
w20344 <= not w20342 and not w20343;
w20345 <= not w14202 and w20344;
w20346 <= w14202 and w20316;
w20347 <= not w20345 and not w20346;
w20348 <= not w14198 and w20347;
w20349 <= not w20317 and not w20348;
w20350 <= not w14194 and w20349;
w20351 <= w14194 and w20316;
w20352 <= not w20350 and not w20351;
w20353 <= not pi0792 and w20352;
w20354 <= pi0628 and not w20352;
w20355 <= not pi0628 and w20316;
w20356 <= pi1156 and not w20355;
w20357 <= not w20354 and w20356;
w20358 <= pi0628 and w20316;
w20359 <= not pi0628 and not w20352;
w20360 <= not pi1156 and not w20358;
w20361 <= not w20359 and w20360;
w20362 <= not w20357 and not w20361;
w20363 <= pi0792 and not w20362;
w20364 <= not w20353 and not w20363;
w20365 <= not pi0647 and not w20364;
w20366 <= pi0647 and not w20316;
w20367 <= not w20365 and not w20366;
w20368 <= not pi1157 and w20367;
w20369 <= pi0647 and not w20364;
w20370 <= not pi0647 and not w20316;
w20371 <= not w20369 and not w20370;
w20372 <= pi1157 and w20371;
w20373 <= not w20368 and not w20372;
w20374 <= pi0787 and not w20373;
w20375 <= not pi0787 and w20364;
w20376 <= not w20374 and not w20375;
w20377 <= not pi0644 and not w20376;
w20378 <= pi0715 and not w20377;
w20379 <= pi0173 and not w134;
w20380 <= pi0173 and not w14838;
w20381 <= not pi0173 and not w14611;
w20382 <= pi0745 and not w20381;
w20383 <= not pi0173 and not pi0745;
w20384 <= w14784 and w20383;
w20385 <= not w20380 and not w20384;
w20386 <= not w20382 and w20385;
w20387 <= not pi0038 and not w20386;
w20388 <= not pi0745 and w14843;
w20389 <= pi0038 and not w20320;
w20390 <= not w20388 and w20389;
w20391 <= not w20387 and not w20390;
w20392 <= w134 and not w20391;
w20393 <= not w20379 and not w20392;
w20394 <= not w14680 and not w20393;
w20395 <= w14680 and not w20316;
w20396 <= not w20394 and not w20395;
w20397 <= not pi0785 and not w20396;
w20398 <= not w14854 and not w20316;
w20399 <= pi0609 and w20394;
w20400 <= not w20398 and not w20399;
w20401 <= pi1155 and not w20400;
w20402 <= not w14859 and not w20316;
w20403 <= not pi0609 and w20394;
w20404 <= not w20402 and not w20403;
w20405 <= not pi1155 and not w20404;
w20406 <= not w20401 and not w20405;
w20407 <= pi0785 and not w20406;
w20408 <= not w20397 and not w20407;
w20409 <= not pi0781 and not w20408;
w20410 <= not pi0618 and w20316;
w20411 <= pi0618 and w20408;
w20412 <= pi1154 and not w20410;
w20413 <= not w20411 and w20412;
w20414 <= not pi0618 and w20408;
w20415 <= pi0618 and w20316;
w20416 <= not pi1154 and not w20415;
w20417 <= not w20414 and w20416;
w20418 <= not w20413 and not w20417;
w20419 <= pi0781 and not w20418;
w20420 <= not w20409 and not w20419;
w20421 <= not pi0789 and not w20420;
w20422 <= not pi0619 and w20316;
w20423 <= pi0619 and w20420;
w20424 <= pi1159 and not w20422;
w20425 <= not w20423 and w20424;
w20426 <= not pi0619 and w20420;
w20427 <= pi0619 and w20316;
w20428 <= not pi1159 and not w20427;
w20429 <= not w20426 and w20428;
w20430 <= not w20425 and not w20429;
w20431 <= pi0789 and not w20430;
w20432 <= not w20421 and not w20431;
w20433 <= not pi0788 and not w20432;
w20434 <= not pi0626 and w20316;
w20435 <= pi0626 and w20432;
w20436 <= pi1158 and not w20434;
w20437 <= not w20435 and w20436;
w20438 <= not pi0626 and w20432;
w20439 <= pi0626 and w20316;
w20440 <= not pi1158 and not w20439;
w20441 <= not w20438 and w20440;
w20442 <= not w20437 and not w20441;
w20443 <= pi0788 and not w20442;
w20444 <= not w20433 and not w20443;
w20445 <= not w15342 and w20444;
w20446 <= w15342 and w20316;
w20447 <= not w20445 and not w20446;
w20448 <= not w15367 and not w20447;
w20449 <= w15367 and w20316;
w20450 <= not w20448 and not w20449;
w20451 <= pi0644 and not w20450;
w20452 <= not pi0644 and w20316;
w20453 <= not pi0715 and not w20452;
w20454 <= not w20451 and w20453;
w20455 <= pi1160 and not w20454;
w20456 <= not w20378 and w20455;
w20457 <= pi0644 and not w20376;
w20458 <= w15365 and not w20367;
w20459 <= not w18122 and w20447;
w20460 <= w15364 and not w20371;
w20461 <= not w20458 and not w20460;
w20462 <= not w20459 and w20461;
w20463 <= pi0787 and not w20462;
w20464 <= not pi0629 and w20357;
w20465 <= not w18133 and not w20444;
w20466 <= pi0629 and w20361;
w20467 <= not w20464 and not w20466;
w20468 <= not w20465 and w20467;
w20469 <= pi0792 and not w20468;
w20470 <= pi0609 and w20341;
w20471 <= pi0173 and not w15188;
w20472 <= not pi0173 and not w15175;
w20473 <= pi0745 and not w20471;
w20474 <= not w20472 and w20473;
w20475 <= not pi0173 and w15192;
w20476 <= pi0173 and w15194;
w20477 <= not pi0745 and not w20476;
w20478 <= not w20475 and w20477;
w20479 <= not w20474 and not w20478;
w20480 <= not pi0039 and not w20479;
w20481 <= pi0173 and w15168;
w20482 <= not pi0173 and not w15109;
w20483 <= not pi0745 and not w20482;
w20484 <= not w20481 and w20483;
w20485 <= not pi0173 and w14967;
w20486 <= pi0173 and w15048;
w20487 <= pi0745 and not w20486;
w20488 <= not w20485 and w20487;
w20489 <= pi0039 and not w20484;
w20490 <= not w20488 and w20489;
w20491 <= not pi0038 and not w20480;
w20492 <= not w20490 and w20491;
w20493 <= not pi0745 and not w15053;
w20494 <= w17034 and not w20493;
w20495 <= not pi0173 and not w20494;
w20496 <= not pi0745 and w14807;
w20497 <= not w15032 and not w20496;
w20498 <= pi0173 and not w20497;
w20499 <= w3847 and w20498;
w20500 <= pi0038 and not w20499;
w20501 <= not w20495 and w20500;
w20502 <= not pi0723 and not w20501;
w20503 <= not w20492 and w20502;
w20504 <= pi0723 and w20391;
w20505 <= w134 and not w20503;
w20506 <= not w20504 and w20505;
w20507 <= not w20379 and not w20506;
w20508 <= not pi0625 and w20507;
w20509 <= pi0625 and w20393;
w20510 <= not pi1153 and not w20509;
w20511 <= not w20508 and w20510;
w20512 <= not pi0608 and not w20334;
w20513 <= not w20511 and w20512;
w20514 <= not pi0625 and w20393;
w20515 <= pi0625 and w20507;
w20516 <= pi1153 and not w20514;
w20517 <= not w20515 and w20516;
w20518 <= pi0608 and not w20338;
w20519 <= not w20517 and w20518;
w20520 <= not w20513 and not w20519;
w20521 <= pi0778 and not w20520;
w20522 <= not pi0778 and w20507;
w20523 <= not w20521 and not w20522;
w20524 <= not pi0609 and not w20523;
w20525 <= not pi1155 and not w20470;
w20526 <= not w20524 and w20525;
w20527 <= not pi0660 and not w20401;
w20528 <= not w20526 and w20527;
w20529 <= not pi0609 and w20341;
w20530 <= pi0609 and not w20523;
w20531 <= pi1155 and not w20529;
w20532 <= not w20530 and w20531;
w20533 <= pi0660 and not w20405;
w20534 <= not w20532 and w20533;
w20535 <= not w20528 and not w20534;
w20536 <= pi0785 and not w20535;
w20537 <= not pi0785 and not w20523;
w20538 <= not w20536 and not w20537;
w20539 <= not pi0618 and not w20538;
w20540 <= pi0618 and w20344;
w20541 <= not pi1154 and not w20540;
w20542 <= not w20539 and w20541;
w20543 <= not pi0627 and not w20413;
w20544 <= not w20542 and w20543;
w20545 <= not pi0618 and w20344;
w20546 <= pi0618 and not w20538;
w20547 <= pi1154 and not w20545;
w20548 <= not w20546 and w20547;
w20549 <= pi0627 and not w20417;
w20550 <= not w20548 and w20549;
w20551 <= not w20544 and not w20550;
w20552 <= pi0781 and not w20551;
w20553 <= not pi0781 and not w20538;
w20554 <= not w20552 and not w20553;
w20555 <= not pi0789 and w20554;
w20556 <= pi0619 and not w20347;
w20557 <= not pi0619 and not w20554;
w20558 <= not pi1159 and not w20556;
w20559 <= not w20557 and w20558;
w20560 <= not pi0648 and not w20425;
w20561 <= not w20559 and w20560;
w20562 <= pi0619 and not w20554;
w20563 <= not pi0619 and not w20347;
w20564 <= pi1159 and not w20563;
w20565 <= not w20562 and w20564;
w20566 <= pi0648 and not w20429;
w20567 <= not w20565 and w20566;
w20568 <= pi0789 and not w20561;
w20569 <= not w20567 and w20568;
w20570 <= w15533 and not w20555;
w20571 <= not w20569 and w20570;
w20572 <= w15434 and w20349;
w20573 <= not w14193 and w20442;
w20574 <= not w20572 and not w20573;
w20575 <= pi0788 and not w20574;
w20576 <= not w17927 and not w20575;
w20577 <= not w20571 and w20576;
w20578 <= not w20469 and not w20577;
w20579 <= not w17769 and not w20578;
w20580 <= not w20463 and not w20579;
w20581 <= not pi0644 and w20580;
w20582 <= not pi0715 and not w20457;
w20583 <= not w20581 and w20582;
w20584 <= pi0644 and w20316;
w20585 <= not pi0644 and not w20450;
w20586 <= pi0715 and not w20584;
w20587 <= not w20585 and w20586;
w20588 <= not pi1160 and not w20587;
w20589 <= not w20583 and w20588;
w20590 <= not w20456 and not w20589;
w20591 <= pi0790 and not w20590;
w20592 <= pi0644 and w20455;
w20593 <= pi0790 and not w20592;
w20594 <= w20580 and not w20593;
w20595 <= not w20591 and not w20594;
w20596 <= w4989 and not w20595;
w20597 <= not pi0832 and not w20315;
w20598 <= not w20596 and w20597;
w20599 <= not pi0173 and not w489;
w20600 <= not pi0723 and w14208;
w20601 <= not w20599 and not w20600;
w20602 <= not pi0778 and not w20601;
w20603 <= not pi0625 and w20600;
w20604 <= not w20601 and not w20603;
w20605 <= pi1153 and not w20604;
w20606 <= not pi1153 and not w20599;
w20607 <= not w20603 and w20606;
w20608 <= pi0778 and not w20607;
w20609 <= not w20605 and w20608;
w20610 <= not w20602 and not w20609;
w20611 <= not w15408 and not w20610;
w20612 <= not w15410 and w20611;
w20613 <= not w15412 and w20612;
w20614 <= not w15414 and w20613;
w20615 <= not w15420 and w20614;
w20616 <= not pi0647 and w20615;
w20617 <= pi0647 and w20599;
w20618 <= not pi1157 and not w20617;
w20619 <= not w20616 and w20618;
w20620 <= pi0630 and w20619;
w20621 <= not w20496 and not w20599;
w20622 <= not w15437 and not w20621;
w20623 <= not pi0785 and not w20622;
w20624 <= w14859 and w20496;
w20625 <= w20622 and not w20624;
w20626 <= pi1155 and not w20625;
w20627 <= not pi1155 and not w20599;
w20628 <= not w20624 and w20627;
w20629 <= not w20626 and not w20628;
w20630 <= pi0785 and not w20629;
w20631 <= not w20623 and not w20630;
w20632 <= not pi0781 and not w20631;
w20633 <= not w15452 and w20631;
w20634 <= pi1154 and not w20633;
w20635 <= not w15455 and w20631;
w20636 <= not pi1154 and not w20635;
w20637 <= not w20634 and not w20636;
w20638 <= pi0781 and not w20637;
w20639 <= not w20632 and not w20638;
w20640 <= not pi0789 and not w20639;
w20641 <= not pi0619 and w489;
w20642 <= w20639 and not w20641;
w20643 <= pi1159 and not w20642;
w20644 <= pi0619 and w489;
w20645 <= w20639 and not w20644;
w20646 <= not pi1159 and not w20645;
w20647 <= not w20643 and not w20646;
w20648 <= pi0789 and not w20647;
w20649 <= not w20640 and not w20648;
w20650 <= not pi0788 and not w20649;
w20651 <= not pi0626 and w20599;
w20652 <= pi0626 and w20649;
w20653 <= pi1158 and not w20651;
w20654 <= not w20652 and w20653;
w20655 <= not pi0626 and w20649;
w20656 <= pi0626 and w20599;
w20657 <= not pi1158 and not w20656;
w20658 <= not w20655 and w20657;
w20659 <= not w20654 and not w20658;
w20660 <= pi0788 and not w20659;
w20661 <= not w20650 and not w20660;
w20662 <= not w15342 and w20661;
w20663 <= w15342 and w20599;
w20664 <= not w20662 and not w20663;
w20665 <= not w18122 and w20664;
w20666 <= pi0647 and not w20615;
w20667 <= not pi0647 and not w20599;
w20668 <= not w20666 and not w20667;
w20669 <= w15364 and not w20668;
w20670 <= not w20620 and not w20669;
w20671 <= not w20665 and w20670;
w20672 <= pi0787 and not w20671;
w20673 <= w15434 and w20613;
w20674 <= not w14193 and w20659;
w20675 <= not w20673 and not w20674;
w20676 <= pi0788 and not w20675;
w20677 <= pi0618 and w20611;
w20678 <= not w14731 and not w20601;
w20679 <= pi0625 and w20678;
w20680 <= w20621 and not w20678;
w20681 <= not w20679 and not w20680;
w20682 <= w20606 and not w20681;
w20683 <= not pi0608 and not w20605;
w20684 <= not w20682 and w20683;
w20685 <= pi1153 and w20621;
w20686 <= not w20679 and w20685;
w20687 <= pi0608 and not w20607;
w20688 <= not w20686 and w20687;
w20689 <= not w20684 and not w20688;
w20690 <= pi0778 and not w20689;
w20691 <= not pi0778 and not w20680;
w20692 <= not w20690 and not w20691;
w20693 <= not pi0609 and not w20692;
w20694 <= pi0609 and not w20610;
w20695 <= not pi1155 and not w20694;
w20696 <= not w20693 and w20695;
w20697 <= not pi0660 and not w20626;
w20698 <= not w20696 and w20697;
w20699 <= pi0609 and not w20692;
w20700 <= not pi0609 and not w20610;
w20701 <= pi1155 and not w20700;
w20702 <= not w20699 and w20701;
w20703 <= pi0660 and not w20628;
w20704 <= not w20702 and w20703;
w20705 <= not w20698 and not w20704;
w20706 <= pi0785 and not w20705;
w20707 <= not pi0785 and not w20692;
w20708 <= not w20706 and not w20707;
w20709 <= not pi0618 and not w20708;
w20710 <= not pi1154 and not w20677;
w20711 <= not w20709 and w20710;
w20712 <= not pi0627 and not w20634;
w20713 <= not w20711 and w20712;
w20714 <= not pi0618 and w20611;
w20715 <= pi0618 and not w20708;
w20716 <= pi1154 and not w20714;
w20717 <= not w20715 and w20716;
w20718 <= pi0627 and not w20636;
w20719 <= not w20717 and w20718;
w20720 <= not w20713 and not w20719;
w20721 <= pi0781 and not w20720;
w20722 <= not pi0781 and not w20708;
w20723 <= not w20721 and not w20722;
w20724 <= not pi0789 and w20723;
w20725 <= not pi0619 and not w20723;
w20726 <= pi0619 and w20612;
w20727 <= not pi1159 and not w20726;
w20728 <= not w20725 and w20727;
w20729 <= not pi0648 and not w20643;
w20730 <= not w20728 and w20729;
w20731 <= not pi0619 and w20612;
w20732 <= pi0619 and not w20723;
w20733 <= pi1159 and not w20731;
w20734 <= not w20732 and w20733;
w20735 <= pi0648 and not w20646;
w20736 <= not w20734 and w20735;
w20737 <= pi0789 and not w20730;
w20738 <= not w20736 and w20737;
w20739 <= w15533 and not w20724;
w20740 <= not w20738 and w20739;
w20741 <= not w20676 and not w20740;
w20742 <= not w17927 and not w20741;
w20743 <= w15417 and w20661;
w20744 <= w18414 and w20614;
w20745 <= not w20743 and not w20744;
w20746 <= not pi0629 and not w20745;
w20747 <= w18418 and w20614;
w20748 <= w15416 and w20661;
w20749 <= not w20747 and not w20748;
w20750 <= pi0629 and not w20749;
w20751 <= not w20746 and not w20750;
w20752 <= pi0792 and not w20751;
w20753 <= not w17769 and not w20752;
w20754 <= not w20742 and w20753;
w20755 <= not w20672 and not w20754;
w20756 <= not pi0790 and w20755;
w20757 <= not pi0787 and not w20615;
w20758 <= pi1157 and not w20668;
w20759 <= not w20619 and not w20758;
w20760 <= pi0787 and not w20759;
w20761 <= not w20757 and not w20760;
w20762 <= not pi0644 and w20761;
w20763 <= pi0644 and w20755;
w20764 <= pi0715 and not w20762;
w20765 <= not w20763 and w20764;
w20766 <= not w15367 and not w20664;
w20767 <= w15367 and w20599;
w20768 <= not w20766 and not w20767;
w20769 <= pi0644 and not w20768;
w20770 <= not pi0644 and w20599;
w20771 <= not pi0715 and not w20770;
w20772 <= not w20769 and w20771;
w20773 <= pi1160 and not w20772;
w20774 <= not w20765 and w20773;
w20775 <= not pi0644 and not w20768;
w20776 <= pi0644 and w20599;
w20777 <= pi0715 and not w20776;
w20778 <= not w20775 and w20777;
w20779 <= pi0644 and w20761;
w20780 <= not pi0644 and w20755;
w20781 <= not pi0715 and not w20779;
w20782 <= not w20780 and w20781;
w20783 <= not pi1160 and not w20778;
w20784 <= not w20782 and w20783;
w20785 <= not w20774 and not w20784;
w20786 <= pi0790 and not w20785;
w20787 <= pi0832 and not w20756;
w20788 <= not w20786 and w20787;
w20789 <= not w20598 and not w20788;
w20790 <= pi0174 and not w14622;
w20791 <= w14198 and not w20790;
w20792 <= w14638 and not w20790;
w20793 <= pi0696 and w134;
w20794 <= not w20790 and not w20793;
w20795 <= not pi0174 and not w14204;
w20796 <= w17462 and not w20795;
w20797 <= not pi0174 and w15639;
w20798 <= pi0174 and not w15635;
w20799 <= not pi0038 and not w20797;
w20800 <= not w20798 and w20799;
w20801 <= w20793 and not w20796;
w20802 <= not w20800 and w20801;
w20803 <= not w20794 and not w20802;
w20804 <= not pi0778 and w20803;
w20805 <= not pi0625 and not w20790;
w20806 <= pi0625 and not w20803;
w20807 <= pi1153 and not w20805;
w20808 <= not w20806 and w20807;
w20809 <= not pi0625 and not w20803;
w20810 <= pi0625 and not w20790;
w20811 <= not pi1153 and not w20810;
w20812 <= not w20809 and w20811;
w20813 <= not w20808 and not w20812;
w20814 <= pi0778 and not w20813;
w20815 <= not w20804 and not w20814;
w20816 <= not w14638 and w20815;
w20817 <= not w20792 and not w20816;
w20818 <= not w14202 and w20817;
w20819 <= w14202 and w20790;
w20820 <= not w20818 and not w20819;
w20821 <= not w14198 and w20820;
w20822 <= not w20791 and not w20821;
w20823 <= not w14194 and w20822;
w20824 <= w14194 and w20790;
w20825 <= not w20823 and not w20824;
w20826 <= not pi0792 and not w20825;
w20827 <= not pi0628 and not w20790;
w20828 <= pi0628 and w20825;
w20829 <= pi1156 and not w20827;
w20830 <= not w20828 and w20829;
w20831 <= pi0628 and not w20790;
w20832 <= not pi0628 and w20825;
w20833 <= not pi1156 and not w20831;
w20834 <= not w20832 and w20833;
w20835 <= not w20830 and not w20834;
w20836 <= pi0792 and not w20835;
w20837 <= not w20826 and not w20836;
w20838 <= not pi0787 and not w20837;
w20839 <= not pi0647 and not w20790;
w20840 <= pi0647 and w20837;
w20841 <= pi1157 and not w20839;
w20842 <= not w20840 and w20841;
w20843 <= pi0647 and not w20790;
w20844 <= not pi0647 and w20837;
w20845 <= not pi1157 and not w20843;
w20846 <= not w20844 and w20845;
w20847 <= not w20842 and not w20846;
w20848 <= pi0787 and not w20847;
w20849 <= not w20838 and not w20848;
w20850 <= not pi0644 and w20849;
w20851 <= not pi0619 and not w20790;
w20852 <= w14680 and not w20790;
w20853 <= pi0174 and not w134;
w20854 <= pi0759 and w14782;
w20855 <= not w19033 and not w20854;
w20856 <= pi0039 and not w20855;
w20857 <= not pi0759 and w14521;
w20858 <= pi0759 and w14702;
w20859 <= not pi0039 and not w20857;
w20860 <= not w20858 and w20859;
w20861 <= not w20856 and not w20860;
w20862 <= pi0174 and not w20861;
w20863 <= not pi0174 and pi0759;
w20864 <= w14838 and w20863;
w20865 <= not w20862 and not w20864;
w20866 <= not pi0038 and not w20865;
w20867 <= pi0759 and w14731;
w20868 <= w14204 and not w20867;
w20869 <= pi0038 and not w20795;
w20870 <= not w20868 and w20869;
w20871 <= not w20866 and not w20870;
w20872 <= w134 and not w20871;
w20873 <= not w20853 and not w20872;
w20874 <= not w14680 and w20873;
w20875 <= not w20852 and not w20874;
w20876 <= not pi0785 and w20875;
w20877 <= not pi0609 and not w20790;
w20878 <= pi0609 and not w20875;
w20879 <= pi1155 and not w20877;
w20880 <= not w20878 and w20879;
w20881 <= not pi0609 and not w20875;
w20882 <= pi0609 and not w20790;
w20883 <= not pi1155 and not w20882;
w20884 <= not w20881 and w20883;
w20885 <= not w20880 and not w20884;
w20886 <= pi0785 and not w20885;
w20887 <= not w20876 and not w20886;
w20888 <= not pi0781 and not w20887;
w20889 <= not pi0618 and not w20790;
w20890 <= pi0618 and w20887;
w20891 <= pi1154 and not w20889;
w20892 <= not w20890 and w20891;
w20893 <= pi0618 and not w20790;
w20894 <= not pi0618 and w20887;
w20895 <= not pi1154 and not w20893;
w20896 <= not w20894 and w20895;
w20897 <= not w20892 and not w20896;
w20898 <= pi0781 and not w20897;
w20899 <= not w20888 and not w20898;
w20900 <= pi0619 and w20899;
w20901 <= pi1159 and not w20851;
w20902 <= not w20900 and w20901;
w20903 <= not pi0696 and w20871;
w20904 <= not pi0174 and not w15168;
w20905 <= pi0174 and w15109;
w20906 <= pi0759 and not w20905;
w20907 <= not w20904 and w20906;
w20908 <= pi0174 and not w14967;
w20909 <= not pi0174 and not w15048;
w20910 <= not pi0759 and not w20909;
w20911 <= not w20908 and w20910;
w20912 <= pi0039 and not w20907;
w20913 <= not w20911 and w20912;
w20914 <= not pi0174 and w15194;
w20915 <= pi0174 and w15192;
w20916 <= pi0759 and not w20914;
w20917 <= not w20915 and w20916;
w20918 <= not pi0174 and not w15188;
w20919 <= pi0174 and not w15175;
w20920 <= not pi0759 and not w20918;
w20921 <= not w20919 and w20920;
w20922 <= not pi0039 and not w20917;
w20923 <= not w20921 and w20922;
w20924 <= not pi0038 and not w20923;
w20925 <= not w20913 and w20924;
w20926 <= pi0696 and not w17033;
w20927 <= not w20870 and w20926;
w20928 <= not w20925 and w20927;
w20929 <= w134 and not w20928;
w20930 <= not w20903 and w20929;
w20931 <= not w20853 and not w20930;
w20932 <= not pi0625 and w20931;
w20933 <= pi0625 and w20873;
w20934 <= not pi1153 and not w20933;
w20935 <= not w20932 and w20934;
w20936 <= not pi0608 and not w20808;
w20937 <= not w20935 and w20936;
w20938 <= not pi0625 and w20873;
w20939 <= pi0625 and w20931;
w20940 <= pi1153 and not w20938;
w20941 <= not w20939 and w20940;
w20942 <= pi0608 and not w20812;
w20943 <= not w20941 and w20942;
w20944 <= not w20937 and not w20943;
w20945 <= pi0778 and not w20944;
w20946 <= not pi0778 and w20931;
w20947 <= not w20945 and not w20946;
w20948 <= not pi0609 and not w20947;
w20949 <= pi0609 and w20815;
w20950 <= not pi1155 and not w20949;
w20951 <= not w20948 and w20950;
w20952 <= not pi0660 and not w20880;
w20953 <= not w20951 and w20952;
w20954 <= not pi0609 and w20815;
w20955 <= pi0609 and not w20947;
w20956 <= pi1155 and not w20954;
w20957 <= not w20955 and w20956;
w20958 <= pi0660 and not w20884;
w20959 <= not w20957 and w20958;
w20960 <= not w20953 and not w20959;
w20961 <= pi0785 and not w20960;
w20962 <= not pi0785 and not w20947;
w20963 <= not w20961 and not w20962;
w20964 <= not pi0618 and not w20963;
w20965 <= pi0618 and not w20817;
w20966 <= not pi1154 and not w20965;
w20967 <= not w20964 and w20966;
w20968 <= not pi0627 and not w20892;
w20969 <= not w20967 and w20968;
w20970 <= pi0618 and not w20963;
w20971 <= not pi0618 and not w20817;
w20972 <= pi1154 and not w20971;
w20973 <= not w20970 and w20972;
w20974 <= pi0627 and not w20896;
w20975 <= not w20973 and w20974;
w20976 <= not w20969 and not w20975;
w20977 <= pi0781 and not w20976;
w20978 <= not pi0781 and not w20963;
w20979 <= not w20977 and not w20978;
w20980 <= not pi0619 and not w20979;
w20981 <= pi0619 and w20820;
w20982 <= not pi1159 and not w20981;
w20983 <= not w20980 and w20982;
w20984 <= not pi0648 and not w20902;
w20985 <= not w20983 and w20984;
w20986 <= pi0619 and not w20790;
w20987 <= not pi0619 and w20899;
w20988 <= not pi1159 and not w20986;
w20989 <= not w20987 and w20988;
w20990 <= not pi0619 and w20820;
w20991 <= pi0619 and not w20979;
w20992 <= pi1159 and not w20990;
w20993 <= not w20991 and w20992;
w20994 <= pi0648 and not w20989;
w20995 <= not w20993 and w20994;
w20996 <= not w20985 and not w20995;
w20997 <= pi0789 and not w20996;
w20998 <= not pi0789 and not w20979;
w20999 <= not w20997 and not w20998;
w21000 <= not pi0788 and w20999;
w21001 <= not pi0626 and w20999;
w21002 <= pi0626 and w20822;
w21003 <= not pi0641 and not w21002;
w21004 <= not w21001 and w21003;
w21005 <= not pi0789 and not w20899;
w21006 <= not w20902 and not w20989;
w21007 <= pi0789 and not w21006;
w21008 <= not w21005 and not w21007;
w21009 <= not pi0626 and not w21008;
w21010 <= pi0626 and w20790;
w21011 <= pi0641 and not w21010;
w21012 <= not w21009 and w21011;
w21013 <= not pi1158 and not w21012;
w21014 <= not w21004 and w21013;
w21015 <= pi0626 and w20999;
w21016 <= not pi0626 and w20822;
w21017 <= pi0641 and not w21016;
w21018 <= not w21015 and w21017;
w21019 <= pi0626 and not w21008;
w21020 <= not pi0626 and w20790;
w21021 <= not pi0641 and not w21020;
w21022 <= not w21019 and w21021;
w21023 <= pi1158 and not w21022;
w21024 <= not w21018 and w21023;
w21025 <= not w21014 and not w21024;
w21026 <= pi0788 and not w21025;
w21027 <= not w21000 and not w21026;
w21028 <= not pi0628 and w21027;
w21029 <= not w15532 and not w21008;
w21030 <= w15532 and w20790;
w21031 <= not w21029 and not w21030;
w21032 <= pi0628 and w21031;
w21033 <= not pi1156 and not w21032;
w21034 <= not w21028 and w21033;
w21035 <= not pi0629 and not w20830;
w21036 <= not w21034 and w21035;
w21037 <= pi0628 and w21027;
w21038 <= not pi0628 and w21031;
w21039 <= pi1156 and not w21038;
w21040 <= not w21037 and w21039;
w21041 <= pi0629 and not w20834;
w21042 <= not w21040 and w21041;
w21043 <= not w21036 and not w21042;
w21044 <= pi0792 and not w21043;
w21045 <= not pi0792 and w21027;
w21046 <= not w21044 and not w21045;
w21047 <= not pi0647 and not w21046;
w21048 <= not w15342 and not w21031;
w21049 <= w15342 and w20790;
w21050 <= not w21048 and not w21049;
w21051 <= pi0647 and w21050;
w21052 <= not pi1157 and not w21051;
w21053 <= not w21047 and w21052;
w21054 <= not pi0630 and not w20842;
w21055 <= not w21053 and w21054;
w21056 <= pi0647 and not w21046;
w21057 <= not pi0647 and w21050;
w21058 <= pi1157 and not w21057;
w21059 <= not w21056 and w21058;
w21060 <= pi0630 and not w20846;
w21061 <= not w21059 and w21060;
w21062 <= not w21055 and not w21061;
w21063 <= pi0787 and not w21062;
w21064 <= not pi0787 and not w21046;
w21065 <= not w21063 and not w21064;
w21066 <= pi0644 and not w21065;
w21067 <= pi0715 and not w20850;
w21068 <= not w21066 and w21067;
w21069 <= w15367 and not w20790;
w21070 <= not w15367 and w21050;
w21071 <= not w21069 and not w21070;
w21072 <= pi0644 and not w21071;
w21073 <= not pi0644 and not w20790;
w21074 <= not pi0715 and not w21073;
w21075 <= not w21072 and w21074;
w21076 <= pi1160 and not w21075;
w21077 <= not w21068 and w21076;
w21078 <= not pi0644 and not w21065;
w21079 <= pi0644 and w20849;
w21080 <= not pi0715 and not w21079;
w21081 <= not w21078 and w21080;
w21082 <= not pi0644 and not w21071;
w21083 <= pi0644 and not w20790;
w21084 <= pi0715 and not w21083;
w21085 <= not w21082 and w21084;
w21086 <= not pi1160 and not w21085;
w21087 <= not w21081 and w21086;
w21088 <= pi0790 and not w21077;
w21089 <= not w21087 and w21088;
w21090 <= not pi0790 and w21065;
w21091 <= w3868 and not w21090;
w21092 <= not w21089 and w21091;
w21093 <= not pi0174 and not w3868;
w21094 <= not pi0057 and not w21093;
w21095 <= not w21092 and w21094;
w21096 <= pi0057 and pi0174;
w21097 <= not pi0832 and not w21096;
w21098 <= not w21095 and w21097;
w21099 <= pi0174 and not w489;
w21100 <= pi0759 and w14807;
w21101 <= w14854 and w21100;
w21102 <= pi1155 and not w21099;
w21103 <= not w21101 and w21102;
w21104 <= pi0696 and w14208;
w21105 <= not w21099 and not w21104;
w21106 <= not pi0778 and w21105;
w21107 <= pi0625 and w21104;
w21108 <= not w21105 and not w21107;
w21109 <= not pi1153 and not w21108;
w21110 <= pi1153 and not w21099;
w21111 <= not w21107 and w21110;
w21112 <= not w21109 and not w21111;
w21113 <= pi0778 and not w21112;
w21114 <= not w21106 and not w21113;
w21115 <= pi0609 and w21114;
w21116 <= not w21099 and not w21100;
w21117 <= pi0696 and w15032;
w21118 <= w21116 and not w21117;
w21119 <= pi0625 and w21117;
w21120 <= not w21118 and not w21119;
w21121 <= not pi1153 and not w21120;
w21122 <= not pi0608 and not w21111;
w21123 <= not w21121 and w21122;
w21124 <= pi1153 and w21116;
w21125 <= not w21119 and w21124;
w21126 <= pi0608 and not w21109;
w21127 <= not w21125 and w21126;
w21128 <= not w21123 and not w21127;
w21129 <= pi0778 and not w21128;
w21130 <= not pi0778 and not w21118;
w21131 <= not w21129 and not w21130;
w21132 <= not pi0609 and not w21131;
w21133 <= not pi1155 and not w21115;
w21134 <= not w21132 and w21133;
w21135 <= not pi0660 and not w21103;
w21136 <= not w21134 and w21135;
w21137 <= w14859 and w21100;
w21138 <= not pi1155 and not w21099;
w21139 <= not w21137 and w21138;
w21140 <= not pi0609 and w21114;
w21141 <= pi0609 and not w21131;
w21142 <= pi1155 and not w21140;
w21143 <= not w21141 and w21142;
w21144 <= pi0660 and not w21139;
w21145 <= not w21143 and w21144;
w21146 <= not w21136 and not w21145;
w21147 <= pi0785 and not w21146;
w21148 <= not pi0785 and not w21131;
w21149 <= not w21147 and not w21148;
w21150 <= not pi0781 and not w21149;
w21151 <= not w17788 and w21100;
w21152 <= w17833 and w21151;
w21153 <= pi1154 and not w21099;
w21154 <= not w21152 and w21153;
w21155 <= not w14638 and w21114;
w21156 <= not w21099 and not w21155;
w21157 <= pi0618 and not w21156;
w21158 <= not pi0618 and not w21149;
w21159 <= not pi1154 and not w21157;
w21160 <= not w21158 and w21159;
w21161 <= not pi0627 and not w21154;
w21162 <= not w21160 and w21161;
w21163 <= w17882 and w21151;
w21164 <= not pi1154 and not w21099;
w21165 <= not w21163 and w21164;
w21166 <= not pi0618 and not w21156;
w21167 <= pi0618 and not w21149;
w21168 <= pi1154 and not w21166;
w21169 <= not w21167 and w21168;
w21170 <= pi0627 and not w21165;
w21171 <= not w21169 and w21170;
w21172 <= not w21162 and not w21171;
w21173 <= pi0781 and not w21172;
w21174 <= pi0648 and w17791;
w21175 <= not pi0648 and w17792;
w21176 <= not w21174 and not w21175;
w21177 <= w14197 and w21176;
w21178 <= pi0789 and not w21177;
w21179 <= not w21150 and not w21178;
w21180 <= not w21173 and w21179;
w21181 <= not w17798 and w21151;
w21182 <= w17908 and w21181;
w21183 <= w14196 and not w21182;
w21184 <= w16713 and w21114;
w21185 <= not w21176 and not w21184;
w21186 <= w17898 and w21181;
w21187 <= w14195 and not w21186;
w21188 <= not w21183 and not w21187;
w21189 <= not w21185 and w21188;
w21190 <= pi0789 and not w21099;
w21191 <= not w21189 and w21190;
w21192 <= w15533 and not w21191;
w21193 <= not w21180 and w21192;
w21194 <= w17800 and w21151;
w21195 <= not pi0626 and w21194;
w21196 <= not w21099 and not w21195;
w21197 <= not pi1158 and not w21196;
w21198 <= not w14198 and w21184;
w21199 <= not w21099 and not w21198;
w21200 <= w15428 and not w21199;
w21201 <= pi0641 and not w21197;
w21202 <= not w21200 and w21201;
w21203 <= w15429 and not w21199;
w21204 <= pi0626 and w21194;
w21205 <= not w21099 and not w21204;
w21206 <= pi1158 and not w21205;
w21207 <= not pi0641 and not w21206;
w21208 <= not w21203 and w21207;
w21209 <= pi0788 and not w21202;
w21210 <= not w21208 and w21209;
w21211 <= not w17927 and not w21210;
w21212 <= not w21193 and w21211;
w21213 <= not w15532 and w21194;
w21214 <= not pi0629 and w21213;
w21215 <= pi0628 and not w21214;
w21216 <= w16714 and w21114;
w21217 <= pi0629 and not w21216;
w21218 <= not w21215 and not w21217;
w21219 <= not pi1156 and not w21218;
w21220 <= not pi0628 and not w21213;
w21221 <= pi0629 and not w21220;
w21222 <= pi0628 and w21216;
w21223 <= pi1156 and not w21221;
w21224 <= not w21222 and w21223;
w21225 <= not w21219 and not w21224;
w21226 <= pi0792 and not w21099;
w21227 <= not w21225 and w21226;
w21228 <= not w21212 and not w21227;
w21229 <= not w17769 and not w21228;
w21230 <= not w15342 and w21213;
w21231 <= not pi0630 and w21230;
w21232 <= pi0647 and not w21231;
w21233 <= not w16705 and w21216;
w21234 <= pi0630 and not w21233;
w21235 <= not w21232 and not w21234;
w21236 <= not pi1157 and not w21235;
w21237 <= pi0630 and w21230;
w21238 <= not pi0630 and not w21233;
w21239 <= pi0647 and not w21238;
w21240 <= pi1157 and not w21237;
w21241 <= not w21239 and w21240;
w21242 <= not w21236 and not w21241;
w21243 <= pi0787 and not w21099;
w21244 <= not w21242 and w21243;
w21245 <= not w21229 and not w21244;
w21246 <= not pi0790 and w21245;
w21247 <= not w15342 and not w15367;
w21248 <= w21213 and w21247;
w21249 <= pi0644 and w21248;
w21250 <= not pi0715 and not w21099;
w21251 <= not w21249 and w21250;
w21252 <= not w16905 and w21233;
w21253 <= not w21099 and not w21252;
w21254 <= not pi0644 and not w21253;
w21255 <= pi0644 and w21245;
w21256 <= pi0715 and not w21254;
w21257 <= not w21255 and w21256;
w21258 <= pi1160 and not w21251;
w21259 <= not w21257 and w21258;
w21260 <= not pi0644 and w21248;
w21261 <= pi0715 and not w21099;
w21262 <= not w21260 and w21261;
w21263 <= not pi0644 and w21245;
w21264 <= pi0644 and not w21253;
w21265 <= not pi0715 and not w21264;
w21266 <= not w21263 and w21265;
w21267 <= not pi1160 and not w21262;
w21268 <= not w21266 and w21267;
w21269 <= not w21259 and not w21268;
w21270 <= pi0790 and not w21269;
w21271 <= pi0832 and not w21246;
w21272 <= not w21270 and w21271;
w21273 <= not w21098 and not w21272;
w21274 <= not pi0175 and not w489;
w21275 <= pi0700 and w14208;
w21276 <= not w21274 and not w21275;
w21277 <= not pi0778 and not w21276;
w21278 <= not pi0625 and w21275;
w21279 <= not w21276 and not w21278;
w21280 <= pi1153 and not w21279;
w21281 <= not pi1153 and not w21274;
w21282 <= not w21278 and w21281;
w21283 <= pi0778 and not w21282;
w21284 <= not w21280 and w21283;
w21285 <= not w21277 and not w21284;
w21286 <= not w15408 and not w21285;
w21287 <= not w15410 and w21286;
w21288 <= not w15412 and w21287;
w21289 <= not w15414 and w21288;
w21290 <= not w15420 and w21289;
w21291 <= not pi0647 and w21290;
w21292 <= pi0647 and w21274;
w21293 <= not pi1157 and not w21292;
w21294 <= not w21291 and w21293;
w21295 <= pi0630 and w21294;
w21296 <= pi0766 and w14807;
w21297 <= not w21274 and not w21296;
w21298 <= not w15437 and not w21297;
w21299 <= not pi0785 and not w21298;
w21300 <= w14859 and w21296;
w21301 <= w21298 and not w21300;
w21302 <= pi1155 and not w21301;
w21303 <= not pi1155 and not w21274;
w21304 <= not w21300 and w21303;
w21305 <= not w21302 and not w21304;
w21306 <= pi0785 and not w21305;
w21307 <= not w21299 and not w21306;
w21308 <= not pi0781 and not w21307;
w21309 <= not w15452 and w21307;
w21310 <= pi1154 and not w21309;
w21311 <= not w15455 and w21307;
w21312 <= not pi1154 and not w21311;
w21313 <= not w21310 and not w21312;
w21314 <= pi0781 and not w21313;
w21315 <= not w21308 and not w21314;
w21316 <= not pi0789 and not w21315;
w21317 <= not w20641 and w21315;
w21318 <= pi1159 and not w21317;
w21319 <= not w20644 and w21315;
w21320 <= not pi1159 and not w21319;
w21321 <= not w21318 and not w21320;
w21322 <= pi0789 and not w21321;
w21323 <= not w21316 and not w21322;
w21324 <= not w15532 and w21323;
w21325 <= w15532 and w21274;
w21326 <= not w21324 and not w21325;
w21327 <= not w15342 and not w21326;
w21328 <= w15342 and w21274;
w21329 <= not w21327 and not w21328;
w21330 <= not w18122 and w21329;
w21331 <= pi0647 and not w21290;
w21332 <= not pi0647 and not w21274;
w21333 <= not w21331 and not w21332;
w21334 <= w15364 and not w21333;
w21335 <= not w21295 and not w21334;
w21336 <= not w21330 and w21335;
w21337 <= pi0787 and not w21336;
w21338 <= w15434 and w21288;
w21339 <= not pi0626 and not w21323;
w21340 <= pi0626 and not w21274;
w21341 <= w14192 and not w21340;
w21342 <= not w21339 and w21341;
w21343 <= pi0626 and not w21323;
w21344 <= not pi0626 and not w21274;
w21345 <= w14191 and not w21344;
w21346 <= not w21343 and w21345;
w21347 <= not w21338 and not w21342;
w21348 <= not w21346 and w21347;
w21349 <= pi0788 and not w21348;
w21350 <= pi0618 and w21286;
w21351 <= not w14731 and not w21276;
w21352 <= pi0625 and w21351;
w21353 <= w21297 and not w21351;
w21354 <= not w21352 and not w21353;
w21355 <= w21281 and not w21354;
w21356 <= not pi0608 and not w21280;
w21357 <= not w21355 and w21356;
w21358 <= pi1153 and w21297;
w21359 <= not w21352 and w21358;
w21360 <= pi0608 and not w21282;
w21361 <= not w21359 and w21360;
w21362 <= not w21357 and not w21361;
w21363 <= pi0778 and not w21362;
w21364 <= not pi0778 and not w21353;
w21365 <= not w21363 and not w21364;
w21366 <= not pi0609 and not w21365;
w21367 <= pi0609 and not w21285;
w21368 <= not pi1155 and not w21367;
w21369 <= not w21366 and w21368;
w21370 <= not pi0660 and not w21302;
w21371 <= not w21369 and w21370;
w21372 <= pi0609 and not w21365;
w21373 <= not pi0609 and not w21285;
w21374 <= pi1155 and not w21373;
w21375 <= not w21372 and w21374;
w21376 <= pi0660 and not w21304;
w21377 <= not w21375 and w21376;
w21378 <= not w21371 and not w21377;
w21379 <= pi0785 and not w21378;
w21380 <= not pi0785 and not w21365;
w21381 <= not w21379 and not w21380;
w21382 <= not pi0618 and not w21381;
w21383 <= not pi1154 and not w21350;
w21384 <= not w21382 and w21383;
w21385 <= not pi0627 and not w21310;
w21386 <= not w21384 and w21385;
w21387 <= not pi0618 and w21286;
w21388 <= pi0618 and not w21381;
w21389 <= pi1154 and not w21387;
w21390 <= not w21388 and w21389;
w21391 <= pi0627 and not w21312;
w21392 <= not w21390 and w21391;
w21393 <= not w21386 and not w21392;
w21394 <= pi0781 and not w21393;
w21395 <= not pi0781 and not w21381;
w21396 <= not w21394 and not w21395;
w21397 <= not pi0789 and w21396;
w21398 <= not pi0619 and not w21396;
w21399 <= pi0619 and w21287;
w21400 <= not pi1159 and not w21399;
w21401 <= not w21398 and w21400;
w21402 <= not pi0648 and not w21318;
w21403 <= not w21401 and w21402;
w21404 <= pi0619 and not w21396;
w21405 <= not pi0619 and w21287;
w21406 <= pi1159 and not w21405;
w21407 <= not w21404 and w21406;
w21408 <= pi0648 and not w21320;
w21409 <= not w21407 and w21408;
w21410 <= pi0789 and not w21403;
w21411 <= not w21409 and w21410;
w21412 <= w15533 and not w21397;
w21413 <= not w21411 and w21412;
w21414 <= not w21349 and not w21413;
w21415 <= not w17927 and not w21414;
w21416 <= w15417 and not w21326;
w21417 <= w18414 and w21289;
w21418 <= not w21416 and not w21417;
w21419 <= not pi0629 and not w21418;
w21420 <= w18418 and w21289;
w21421 <= w15416 and not w21326;
w21422 <= not w21420 and not w21421;
w21423 <= pi0629 and not w21422;
w21424 <= not w21419 and not w21423;
w21425 <= pi0792 and not w21424;
w21426 <= not w17769 and not w21425;
w21427 <= not w21415 and w21426;
w21428 <= not w21337 and not w21427;
w21429 <= not pi0790 and w21428;
w21430 <= not pi0787 and not w21290;
w21431 <= pi1157 and not w21333;
w21432 <= not w21294 and not w21431;
w21433 <= pi0787 and not w21432;
w21434 <= not w21430 and not w21433;
w21435 <= not pi0644 and w21434;
w21436 <= pi0644 and w21428;
w21437 <= pi0715 and not w21435;
w21438 <= not w21436 and w21437;
w21439 <= not w15367 and not w21329;
w21440 <= w15367 and w21274;
w21441 <= not w21439 and not w21440;
w21442 <= pi0644 and not w21441;
w21443 <= not pi0644 and w21274;
w21444 <= not pi0715 and not w21443;
w21445 <= not w21442 and w21444;
w21446 <= pi1160 and not w21445;
w21447 <= not w21438 and w21446;
w21448 <= not pi0644 and not w21441;
w21449 <= pi0644 and w21274;
w21450 <= pi0715 and not w21449;
w21451 <= not w21448 and w21450;
w21452 <= pi0644 and w21434;
w21453 <= not pi0644 and w21428;
w21454 <= not pi0715 and not w21452;
w21455 <= not w21453 and w21454;
w21456 <= not pi1160 and not w21451;
w21457 <= not w21455 and w21456;
w21458 <= not w21447 and not w21457;
w21459 <= pi0790 and not w21458;
w21460 <= pi0832 and not w21429;
w21461 <= not w21459 and w21460;
w21462 <= not pi0175 and not w4989;
w21463 <= not pi0175 and not w14622;
w21464 <= w14198 and not w21463;
w21465 <= pi0175 and not w134;
w21466 <= not pi0175 and not w14204;
w21467 <= w14210 and not w21466;
w21468 <= not pi0175 and w15635;
w21469 <= pi0175 and not w15639;
w21470 <= not pi0038 and not w21469;
w21471 <= not w21468 and w21470;
w21472 <= pi0700 and not w21467;
w21473 <= not w21471 and w21472;
w21474 <= not pi0175 and not pi0700;
w21475 <= not w14615 and w21474;
w21476 <= w134 and not w21475;
w21477 <= not w21473 and w21476;
w21478 <= not w21465 and not w21477;
w21479 <= not pi0778 and not w21478;
w21480 <= not pi0625 and w21463;
w21481 <= pi0625 and w21478;
w21482 <= pi1153 and not w21480;
w21483 <= not w21481 and w21482;
w21484 <= not pi0625 and w21478;
w21485 <= pi0625 and w21463;
w21486 <= not pi1153 and not w21485;
w21487 <= not w21484 and w21486;
w21488 <= not w21483 and not w21487;
w21489 <= pi0778 and not w21488;
w21490 <= not w21479 and not w21489;
w21491 <= not w14638 and not w21490;
w21492 <= w14638 and not w21463;
w21493 <= not w21491 and not w21492;
w21494 <= not w14202 and w21493;
w21495 <= w14202 and w21463;
w21496 <= not w21494 and not w21495;
w21497 <= not w14198 and w21496;
w21498 <= not w21464 and not w21497;
w21499 <= not w14194 and w21498;
w21500 <= w14194 and w21463;
w21501 <= not w21499 and not w21500;
w21502 <= not pi0628 and not w21501;
w21503 <= pi0628 and w21463;
w21504 <= not w21502 and not w21503;
w21505 <= not pi1156 and not w21504;
w21506 <= pi0628 and not w21501;
w21507 <= not pi0628 and w21463;
w21508 <= not w21506 and not w21507;
w21509 <= pi1156 and not w21508;
w21510 <= not w21505 and not w21509;
w21511 <= pi0792 and not w21510;
w21512 <= not pi0792 and not w21501;
w21513 <= not w21511 and not w21512;
w21514 <= not pi0647 and not w21513;
w21515 <= pi0647 and w21463;
w21516 <= not w21514 and not w21515;
w21517 <= not pi1157 and not w21516;
w21518 <= pi0647 and not w21513;
w21519 <= not pi0647 and w21463;
w21520 <= not w21518 and not w21519;
w21521 <= pi1157 and not w21520;
w21522 <= not w21517 and not w21521;
w21523 <= pi0787 and not w21522;
w21524 <= not pi0787 and not w21513;
w21525 <= not w21523 and not w21524;
w21526 <= not pi0644 and not w21525;
w21527 <= pi0715 and not w21526;
w21528 <= not pi0766 and w14609;
w21529 <= pi0175 and w14836;
w21530 <= not w21528 and not w21529;
w21531 <= pi0039 and not w21530;
w21532 <= pi0766 and not w14797;
w21533 <= pi0175 and not w21532;
w21534 <= not pi0175 and pi0766;
w21535 <= w14784 and w21534;
w21536 <= not w19062 and not w21533;
w21537 <= not w21535 and w21536;
w21538 <= not w21531 and w21537;
w21539 <= not pi0038 and not w21538;
w21540 <= pi0766 and w14843;
w21541 <= pi0038 and not w21466;
w21542 <= not w21540 and w21541;
w21543 <= not w21539 and not w21542;
w21544 <= w134 and not w21543;
w21545 <= not w21465 and not w21544;
w21546 <= not w14680 and not w21545;
w21547 <= w14680 and not w21463;
w21548 <= not w21546 and not w21547;
w21549 <= not pi0785 and not w21548;
w21550 <= not w14854 and not w21463;
w21551 <= pi0609 and w21546;
w21552 <= not w21550 and not w21551;
w21553 <= pi1155 and not w21552;
w21554 <= not w14859 and not w21463;
w21555 <= not pi0609 and w21546;
w21556 <= not w21554 and not w21555;
w21557 <= not pi1155 and not w21556;
w21558 <= not w21553 and not w21557;
w21559 <= pi0785 and not w21558;
w21560 <= not w21549 and not w21559;
w21561 <= not pi0781 and not w21560;
w21562 <= not pi0618 and w21463;
w21563 <= pi0618 and w21560;
w21564 <= pi1154 and not w21562;
w21565 <= not w21563 and w21564;
w21566 <= not pi0618 and w21560;
w21567 <= pi0618 and w21463;
w21568 <= not pi1154 and not w21567;
w21569 <= not w21566 and w21568;
w21570 <= not w21565 and not w21569;
w21571 <= pi0781 and not w21570;
w21572 <= not w21561 and not w21571;
w21573 <= not pi0789 and not w21572;
w21574 <= not pi0619 and w21463;
w21575 <= pi0619 and w21572;
w21576 <= pi1159 and not w21574;
w21577 <= not w21575 and w21576;
w21578 <= not pi0619 and w21572;
w21579 <= pi0619 and w21463;
w21580 <= not pi1159 and not w21579;
w21581 <= not w21578 and w21580;
w21582 <= not w21577 and not w21581;
w21583 <= pi0789 and not w21582;
w21584 <= not w21573 and not w21583;
w21585 <= not w15532 and w21584;
w21586 <= w15532 and w21463;
w21587 <= not w21585 and not w21586;
w21588 <= not w15342 and not w21587;
w21589 <= w15342 and w21463;
w21590 <= not w21588 and not w21589;
w21591 <= not w15367 and not w21590;
w21592 <= w15367 and w21463;
w21593 <= not w21591 and not w21592;
w21594 <= pi0644 and not w21593;
w21595 <= not pi0644 and w21463;
w21596 <= not pi0715 and not w21595;
w21597 <= not w21594 and w21596;
w21598 <= pi1160 and not w21597;
w21599 <= not w21527 and w21598;
w21600 <= pi0644 and not w21525;
w21601 <= not pi0715 and not w21600;
w21602 <= not pi0644 and not w21593;
w21603 <= pi0644 and w21463;
w21604 <= pi0715 and not w21603;
w21605 <= not w21602 and w21604;
w21606 <= not pi1160 and not w21605;
w21607 <= not w21601 and w21606;
w21608 <= not w21599 and not w21607;
w21609 <= pi0790 and not w21608;
w21610 <= w15340 and w21504;
w21611 <= not w18133 and w21587;
w21612 <= w15339 and w21508;
w21613 <= not w21610 and not w21612;
w21614 <= not w21611 and w21613;
w21615 <= pi0792 and not w21614;
w21616 <= pi0609 and w21490;
w21617 <= not pi0700 and w21543;
w21618 <= w14230 and not w14899;
w21619 <= not pi0766 and w21618;
w21620 <= not w15053 and not w21619;
w21621 <= not pi0039 and not w21620;
w21622 <= not pi0175 and not w21621;
w21623 <= not w15032 and not w21296;
w21624 <= pi0175 and not w21623;
w21625 <= w3847 and w21624;
w21626 <= pi0038 and not w21625;
w21627 <= not w21622 and w21626;
w21628 <= not pi0175 and not w15192;
w21629 <= pi0175 and not w15194;
w21630 <= pi0766 and not w21629;
w21631 <= not w21628 and w21630;
w21632 <= not pi0175 and w15175;
w21633 <= pi0175 and w15188;
w21634 <= not pi0766 and not w21632;
w21635 <= not w21633 and w21634;
w21636 <= not pi0039 and not w21631;
w21637 <= not w21635 and w21636;
w21638 <= pi0175 and w15168;
w21639 <= not pi0175 and not w15109;
w21640 <= pi0766 and not w21639;
w21641 <= not w21638 and w21640;
w21642 <= not pi0175 and w14967;
w21643 <= pi0175 and w15048;
w21644 <= not pi0766 and not w21643;
w21645 <= not w21642 and w21644;
w21646 <= pi0039 and not w21641;
w21647 <= not w21645 and w21646;
w21648 <= not pi0038 and not w21637;
w21649 <= not w21647 and w21648;
w21650 <= pi0700 and not w21627;
w21651 <= not w21649 and w21650;
w21652 <= w134 and not w21651;
w21653 <= not w21617 and w21652;
w21654 <= not w21465 and not w21653;
w21655 <= not pi0625 and w21654;
w21656 <= pi0625 and w21545;
w21657 <= not pi1153 and not w21656;
w21658 <= not w21655 and w21657;
w21659 <= not pi0608 and not w21483;
w21660 <= not w21658 and w21659;
w21661 <= not pi0625 and w21545;
w21662 <= pi0625 and w21654;
w21663 <= pi1153 and not w21661;
w21664 <= not w21662 and w21663;
w21665 <= pi0608 and not w21487;
w21666 <= not w21664 and w21665;
w21667 <= not w21660 and not w21666;
w21668 <= pi0778 and not w21667;
w21669 <= not pi0778 and w21654;
w21670 <= not w21668 and not w21669;
w21671 <= not pi0609 and not w21670;
w21672 <= not pi1155 and not w21616;
w21673 <= not w21671 and w21672;
w21674 <= not pi0660 and not w21553;
w21675 <= not w21673 and w21674;
w21676 <= not pi0609 and w21490;
w21677 <= pi0609 and not w21670;
w21678 <= pi1155 and not w21676;
w21679 <= not w21677 and w21678;
w21680 <= pi0660 and not w21557;
w21681 <= not w21679 and w21680;
w21682 <= not w21675 and not w21681;
w21683 <= pi0785 and not w21682;
w21684 <= not pi0785 and not w21670;
w21685 <= not w21683 and not w21684;
w21686 <= not pi0618 and not w21685;
w21687 <= pi0618 and w21493;
w21688 <= not pi1154 and not w21687;
w21689 <= not w21686 and w21688;
w21690 <= not pi0627 and not w21565;
w21691 <= not w21689 and w21690;
w21692 <= not pi0618 and w21493;
w21693 <= pi0618 and not w21685;
w21694 <= pi1154 and not w21692;
w21695 <= not w21693 and w21694;
w21696 <= pi0627 and not w21569;
w21697 <= not w21695 and w21696;
w21698 <= not w21691 and not w21697;
w21699 <= pi0781 and not w21698;
w21700 <= not pi0781 and not w21685;
w21701 <= not w21699 and not w21700;
w21702 <= not pi0789 and w21701;
w21703 <= pi0619 and not w21496;
w21704 <= not pi0619 and not w21701;
w21705 <= not pi1159 and not w21703;
w21706 <= not w21704 and w21705;
w21707 <= not pi0648 and not w21577;
w21708 <= not w21706 and w21707;
w21709 <= not pi0619 and not w21496;
w21710 <= pi0619 and not w21701;
w21711 <= pi1159 and not w21709;
w21712 <= not w21710 and w21711;
w21713 <= pi0648 and not w21581;
w21714 <= not w21712 and w21713;
w21715 <= pi0789 and not w21708;
w21716 <= not w21714 and w21715;
w21717 <= w15533 and not w21702;
w21718 <= not w21716 and w21717;
w21719 <= w15434 and w21498;
w21720 <= not pi0626 and not w21584;
w21721 <= pi0626 and not w21463;
w21722 <= w14192 and not w21721;
w21723 <= not w21720 and w21722;
w21724 <= pi0626 and not w21584;
w21725 <= not pi0626 and not w21463;
w21726 <= w14191 and not w21725;
w21727 <= not w21724 and w21726;
w21728 <= not w21719 and not w21723;
w21729 <= not w21727 and w21728;
w21730 <= pi0788 and not w21729;
w21731 <= not w17927 and not w21730;
w21732 <= not w21718 and w21731;
w21733 <= not w21615 and not w21732;
w21734 <= not w17769 and not w21733;
w21735 <= w15365 and w21516;
w21736 <= not w18122 and w21590;
w21737 <= w15364 and w21520;
w21738 <= not w21735 and not w21736;
w21739 <= not w21737 and w21738;
w21740 <= pi0787 and not w21739;
w21741 <= not pi0644 and w21606;
w21742 <= pi0644 and w21598;
w21743 <= pi0790 and not w21741;
w21744 <= not w21742 and w21743;
w21745 <= not w21734 and not w21740;
w21746 <= not w21744 and w21745;
w21747 <= not w21609 and not w21746;
w21748 <= w4989 and not w21747;
w21749 <= not pi0832 and not w21462;
w21750 <= not w21748 and w21749;
w21751 <= not w21461 and not w21750;
w21752 <= not pi0176 and not w489;
w21753 <= not pi0704 and w14208;
w21754 <= not w21752 and not w21753;
w21755 <= not pi0778 and w21754;
w21756 <= not pi0625 and w21753;
w21757 <= not w21754 and not w21756;
w21758 <= pi1153 and not w21757;
w21759 <= not pi1153 and not w21752;
w21760 <= not w21756 and w21759;
w21761 <= not w21758 and not w21760;
w21762 <= pi0778 and not w21761;
w21763 <= not w21755 and not w21762;
w21764 <= not w15408 and w21763;
w21765 <= not w15410 and w21764;
w21766 <= not w15412 and w21765;
w21767 <= not w15414 and w21766;
w21768 <= not w15420 and w21767;
w21769 <= not pi0647 and w21768;
w21770 <= pi0647 and w21752;
w21771 <= not pi1157 and not w21770;
w21772 <= not w21769 and w21771;
w21773 <= pi0630 and w21772;
w21774 <= not pi0742 and w14807;
w21775 <= not w21752 and not w21774;
w21776 <= not w15437 and not w21775;
w21777 <= not pi0785 and not w21776;
w21778 <= not w15442 and not w21775;
w21779 <= pi1155 and not w21778;
w21780 <= not w15445 and w21776;
w21781 <= not pi1155 and not w21780;
w21782 <= not w21779 and not w21781;
w21783 <= pi0785 and not w21782;
w21784 <= not w21777 and not w21783;
w21785 <= not pi0781 and not w21784;
w21786 <= not w15452 and w21784;
w21787 <= pi1154 and not w21786;
w21788 <= not w15455 and w21784;
w21789 <= not pi1154 and not w21788;
w21790 <= not w21787 and not w21789;
w21791 <= pi0781 and not w21790;
w21792 <= not w21785 and not w21791;
w21793 <= not pi0789 and not w21792;
w21794 <= not pi0619 and w21752;
w21795 <= pi0619 and w21792;
w21796 <= pi1159 and not w21794;
w21797 <= not w21795 and w21796;
w21798 <= not pi0619 and w21792;
w21799 <= pi0619 and w21752;
w21800 <= not pi1159 and not w21799;
w21801 <= not w21798 and w21800;
w21802 <= not w21797 and not w21801;
w21803 <= pi0789 and not w21802;
w21804 <= not w21793 and not w21803;
w21805 <= not w15532 and w21804;
w21806 <= w15532 and w21752;
w21807 <= not w21805 and not w21806;
w21808 <= not w15342 and not w21807;
w21809 <= w15342 and w21752;
w21810 <= not w21808 and not w21809;
w21811 <= not w18122 and w21810;
w21812 <= pi0647 and not w21768;
w21813 <= not pi0647 and not w21752;
w21814 <= not w21812 and not w21813;
w21815 <= w15364 and not w21814;
w21816 <= not w21773 and not w21815;
w21817 <= not w21811 and w21816;
w21818 <= pi0787 and not w21817;
w21819 <= w15434 and w21766;
w21820 <= not pi0626 and not w21804;
w21821 <= pi0626 and not w21752;
w21822 <= w14192 and not w21821;
w21823 <= not w21820 and w21822;
w21824 <= pi0626 and not w21804;
w21825 <= not pi0626 and not w21752;
w21826 <= w14191 and not w21825;
w21827 <= not w21824 and w21826;
w21828 <= not w21819 and not w21823;
w21829 <= not w21827 and w21828;
w21830 <= pi0788 and not w21829;
w21831 <= pi0618 and w21764;
w21832 <= pi0609 and w21763;
w21833 <= not w14731 and not w21754;
w21834 <= pi0625 and w21833;
w21835 <= w21775 and not w21833;
w21836 <= not w21834 and not w21835;
w21837 <= w21759 and not w21836;
w21838 <= not pi0608 and not w21758;
w21839 <= not w21837 and w21838;
w21840 <= pi1153 and w21775;
w21841 <= not w21834 and w21840;
w21842 <= pi0608 and not w21760;
w21843 <= not w21841 and w21842;
w21844 <= not w21839 and not w21843;
w21845 <= pi0778 and not w21844;
w21846 <= not pi0778 and not w21835;
w21847 <= not w21845 and not w21846;
w21848 <= not pi0609 and not w21847;
w21849 <= not pi1155 and not w21832;
w21850 <= not w21848 and w21849;
w21851 <= not pi0660 and not w21779;
w21852 <= not w21850 and w21851;
w21853 <= not pi0609 and w21763;
w21854 <= pi0609 and not w21847;
w21855 <= pi1155 and not w21853;
w21856 <= not w21854 and w21855;
w21857 <= pi0660 and not w21781;
w21858 <= not w21856 and w21857;
w21859 <= not w21852 and not w21858;
w21860 <= pi0785 and not w21859;
w21861 <= not pi0785 and not w21847;
w21862 <= not w21860 and not w21861;
w21863 <= not pi0618 and not w21862;
w21864 <= not pi1154 and not w21831;
w21865 <= not w21863 and w21864;
w21866 <= not pi0627 and not w21787;
w21867 <= not w21865 and w21866;
w21868 <= not pi0618 and w21764;
w21869 <= pi0618 and not w21862;
w21870 <= pi1154 and not w21868;
w21871 <= not w21869 and w21870;
w21872 <= pi0627 and not w21789;
w21873 <= not w21871 and w21872;
w21874 <= not w21867 and not w21873;
w21875 <= pi0781 and not w21874;
w21876 <= not pi0781 and not w21862;
w21877 <= not w21875 and not w21876;
w21878 <= not pi0789 and w21877;
w21879 <= not pi0619 and not w21877;
w21880 <= pi0619 and w21765;
w21881 <= not pi1159 and not w21880;
w21882 <= not w21879 and w21881;
w21883 <= not pi0648 and not w21797;
w21884 <= not w21882 and w21883;
w21885 <= pi0619 and not w21877;
w21886 <= not pi0619 and w21765;
w21887 <= pi1159 and not w21886;
w21888 <= not w21885 and w21887;
w21889 <= pi0648 and not w21801;
w21890 <= not w21888 and w21889;
w21891 <= pi0789 and not w21884;
w21892 <= not w21890 and w21891;
w21893 <= w15533 and not w21878;
w21894 <= not w21892 and w21893;
w21895 <= not w21830 and not w21894;
w21896 <= not w17927 and not w21895;
w21897 <= w15417 and not w21807;
w21898 <= w18414 and w21767;
w21899 <= not w21897 and not w21898;
w21900 <= not pi0629 and not w21899;
w21901 <= w18418 and w21767;
w21902 <= w15416 and not w21807;
w21903 <= not w21901 and not w21902;
w21904 <= pi0629 and not w21903;
w21905 <= not w21900 and not w21904;
w21906 <= pi0792 and not w21905;
w21907 <= not w17769 and not w21906;
w21908 <= not w21896 and w21907;
w21909 <= not w21818 and not w21908;
w21910 <= not pi0790 and w21909;
w21911 <= not pi0787 and not w21768;
w21912 <= pi1157 and not w21814;
w21913 <= not w21772 and not w21912;
w21914 <= pi0787 and not w21913;
w21915 <= not w21911 and not w21914;
w21916 <= not pi0644 and w21915;
w21917 <= pi0644 and w21909;
w21918 <= pi0715 and not w21916;
w21919 <= not w21917 and w21918;
w21920 <= not w15367 and not w21810;
w21921 <= w15367 and w21752;
w21922 <= not w21920 and not w21921;
w21923 <= pi0644 and not w21922;
w21924 <= not pi0644 and w21752;
w21925 <= not pi0715 and not w21924;
w21926 <= not w21923 and w21925;
w21927 <= pi1160 and not w21926;
w21928 <= not w21919 and w21927;
w21929 <= not pi0644 and not w21922;
w21930 <= pi0644 and w21752;
w21931 <= pi0715 and not w21930;
w21932 <= not w21929 and w21931;
w21933 <= pi0644 and w21915;
w21934 <= not pi0644 and w21909;
w21935 <= not pi0715 and not w21933;
w21936 <= not w21934 and w21935;
w21937 <= not pi1160 and not w21932;
w21938 <= not w21936 and w21937;
w21939 <= not w21928 and not w21938;
w21940 <= pi0790 and not w21939;
w21941 <= pi0832 and not w21910;
w21942 <= not w21940 and w21941;
w21943 <= not pi0176 and not w4989;
w21944 <= not pi0176 and not w14622;
w21945 <= w14198 and not w21944;
w21946 <= not pi0038 and w15639;
w21947 <= w134 and not w14210;
w21948 <= not w21946 and w21947;
w21949 <= pi0176 and not w21948;
w21950 <= not pi0038 and w15635;
w21951 <= not w17462 and not w21950;
w21952 <= not pi0176 and w21951;
w21953 <= not pi0704 and not w21952;
w21954 <= not pi0176 and not w14615;
w21955 <= pi0704 and w21954;
w21956 <= w134 and not w21955;
w21957 <= not w21953 and w21956;
w21958 <= not w21949 and not w21957;
w21959 <= not pi0778 and not w21958;
w21960 <= not pi0625 and w21944;
w21961 <= pi0625 and w21958;
w21962 <= pi1153 and not w21960;
w21963 <= not w21961 and w21962;
w21964 <= not pi0625 and w21958;
w21965 <= pi0625 and w21944;
w21966 <= not pi1153 and not w21965;
w21967 <= not w21964 and w21966;
w21968 <= not w21963 and not w21967;
w21969 <= pi0778 and not w21968;
w21970 <= not w21959 and not w21969;
w21971 <= not w14638 and not w21970;
w21972 <= w14638 and not w21944;
w21973 <= not w21971 and not w21972;
w21974 <= not w14202 and w21973;
w21975 <= w14202 and w21944;
w21976 <= not w21974 and not w21975;
w21977 <= not w14198 and w21976;
w21978 <= not w21945 and not w21977;
w21979 <= not w14194 and w21978;
w21980 <= w14194 and w21944;
w21981 <= not w21979 and not w21980;
w21982 <= not pi0628 and not w21981;
w21983 <= pi0628 and w21944;
w21984 <= not w21982 and not w21983;
w21985 <= not pi1156 and not w21984;
w21986 <= pi0628 and not w21981;
w21987 <= not pi0628 and w21944;
w21988 <= not w21986 and not w21987;
w21989 <= pi1156 and not w21988;
w21990 <= not w21985 and not w21989;
w21991 <= pi0792 and not w21990;
w21992 <= not pi0792 and not w21981;
w21993 <= not w21991 and not w21992;
w21994 <= not pi0647 and not w21993;
w21995 <= pi0647 and w21944;
w21996 <= not w21994 and not w21995;
w21997 <= not pi1157 and not w21996;
w21998 <= pi0647 and not w21993;
w21999 <= not pi0647 and w21944;
w22000 <= not w21998 and not w21999;
w22001 <= pi1157 and not w22000;
w22002 <= not w21997 and not w22001;
w22003 <= pi0787 and not w22002;
w22004 <= not pi0787 and not w21993;
w22005 <= not w22003 and not w22004;
w22006 <= not pi0644 and not w22005;
w22007 <= pi0715 and not w22006;
w22008 <= pi0176 and not w134;
w22009 <= not pi0176 and w17002;
w22010 <= not w16996 and not w16997;
w22011 <= pi0176 and w22010;
w22012 <= not w22009 and not w22011;
w22013 <= not pi0742 and not w22012;
w22014 <= pi0742 and not w21954;
w22015 <= not w22013 and not w22014;
w22016 <= w134 and not w22015;
w22017 <= not w22008 and not w22016;
w22018 <= not w14680 and not w22017;
w22019 <= w14680 and not w21944;
w22020 <= not w22018 and not w22019;
w22021 <= not pi0785 and not w22020;
w22022 <= not w14854 and not w21944;
w22023 <= pi0609 and w22018;
w22024 <= not w22022 and not w22023;
w22025 <= pi1155 and not w22024;
w22026 <= not w14859 and not w21944;
w22027 <= not pi0609 and w22018;
w22028 <= not w22026 and not w22027;
w22029 <= not pi1155 and not w22028;
w22030 <= not w22025 and not w22029;
w22031 <= pi0785 and not w22030;
w22032 <= not w22021 and not w22031;
w22033 <= not pi0781 and not w22032;
w22034 <= not pi0618 and w21944;
w22035 <= pi0618 and w22032;
w22036 <= pi1154 and not w22034;
w22037 <= not w22035 and w22036;
w22038 <= not pi0618 and w22032;
w22039 <= pi0618 and w21944;
w22040 <= not pi1154 and not w22039;
w22041 <= not w22038 and w22040;
w22042 <= not w22037 and not w22041;
w22043 <= pi0781 and not w22042;
w22044 <= not w22033 and not w22043;
w22045 <= not pi0789 and not w22044;
w22046 <= not pi0619 and w21944;
w22047 <= pi0619 and w22044;
w22048 <= pi1159 and not w22046;
w22049 <= not w22047 and w22048;
w22050 <= not pi0619 and w22044;
w22051 <= pi0619 and w21944;
w22052 <= not pi1159 and not w22051;
w22053 <= not w22050 and w22052;
w22054 <= not w22049 and not w22053;
w22055 <= pi0789 and not w22054;
w22056 <= not w22045 and not w22055;
w22057 <= not w15532 and w22056;
w22058 <= w15532 and w21944;
w22059 <= not w22057 and not w22058;
w22060 <= not w15342 and not w22059;
w22061 <= w15342 and w21944;
w22062 <= not w22060 and not w22061;
w22063 <= not w15367 and not w22062;
w22064 <= w15367 and w21944;
w22065 <= not w22063 and not w22064;
w22066 <= pi0644 and not w22065;
w22067 <= not pi0644 and w21944;
w22068 <= not pi0715 and not w22067;
w22069 <= not w22066 and w22068;
w22070 <= pi1160 and not w22069;
w22071 <= not w22007 and w22070;
w22072 <= pi0644 and not w22005;
w22073 <= not pi0715 and not w22072;
w22074 <= not pi0644 and not w22065;
w22075 <= pi0644 and w21944;
w22076 <= pi0715 and not w22075;
w22077 <= not w22074 and w22076;
w22078 <= not pi1160 and not w22077;
w22079 <= not w22073 and w22078;
w22080 <= not w22071 and not w22079;
w22081 <= pi0790 and not w22080;
w22082 <= w15365 and w21996;
w22083 <= not w18122 and w22062;
w22084 <= w15364 and w22000;
w22085 <= not w22082 and not w22083;
w22086 <= not w22084 and w22085;
w22087 <= pi0787 and not w22086;
w22088 <= w15340 and w21984;
w22089 <= not w18133 and w22059;
w22090 <= w15339 and w21988;
w22091 <= not w22088 and not w22090;
w22092 <= not w22089 and w22091;
w22093 <= pi0792 and not w22092;
w22094 <= w15434 and w21978;
w22095 <= not pi0626 and not w22056;
w22096 <= pi0626 and not w21944;
w22097 <= w14192 and not w22096;
w22098 <= not w22095 and w22097;
w22099 <= pi0626 and not w22056;
w22100 <= not pi0626 and not w21944;
w22101 <= w14191 and not w22100;
w22102 <= not w22099 and w22101;
w22103 <= not w22094 and not w22098;
w22104 <= not w22102 and w22103;
w22105 <= pi0788 and not w22104;
w22106 <= pi0609 and w21970;
w22107 <= not pi0176 and not w17051;
w22108 <= pi0176 and w17059;
w22109 <= not pi0742 and not w22107;
w22110 <= not w22108 and w22109;
w22111 <= not pi0176 and w17040;
w22112 <= not w17031 and not w17033;
w22113 <= pi0176 and not w22112;
w22114 <= pi0742 and not w22113;
w22115 <= not w22111 and w22114;
w22116 <= not pi0704 and not w22110;
w22117 <= not w22115 and w22116;
w22118 <= pi0704 and w22015;
w22119 <= w134 and not w22117;
w22120 <= not w22118 and w22119;
w22121 <= not w22008 and not w22120;
w22122 <= not pi0625 and w22121;
w22123 <= pi0625 and w22017;
w22124 <= not pi1153 and not w22123;
w22125 <= not w22122 and w22124;
w22126 <= not pi0608 and not w21963;
w22127 <= not w22125 and w22126;
w22128 <= not pi0625 and w22017;
w22129 <= pi0625 and w22121;
w22130 <= pi1153 and not w22128;
w22131 <= not w22129 and w22130;
w22132 <= pi0608 and not w21967;
w22133 <= not w22131 and w22132;
w22134 <= not w22127 and not w22133;
w22135 <= pi0778 and not w22134;
w22136 <= not pi0778 and w22121;
w22137 <= not w22135 and not w22136;
w22138 <= not pi0609 and not w22137;
w22139 <= not pi1155 and not w22106;
w22140 <= not w22138 and w22139;
w22141 <= not pi0660 and not w22025;
w22142 <= not w22140 and w22141;
w22143 <= not pi0609 and w21970;
w22144 <= pi0609 and not w22137;
w22145 <= pi1155 and not w22143;
w22146 <= not w22144 and w22145;
w22147 <= pi0660 and not w22029;
w22148 <= not w22146 and w22147;
w22149 <= not w22142 and not w22148;
w22150 <= pi0785 and not w22149;
w22151 <= not pi0785 and not w22137;
w22152 <= not w22150 and not w22151;
w22153 <= not pi0618 and not w22152;
w22154 <= pi0618 and w21973;
w22155 <= not pi1154 and not w22154;
w22156 <= not w22153 and w22155;
w22157 <= not pi0627 and not w22037;
w22158 <= not w22156 and w22157;
w22159 <= not pi0618 and w21973;
w22160 <= pi0618 and not w22152;
w22161 <= pi1154 and not w22159;
w22162 <= not w22160 and w22161;
w22163 <= pi0627 and not w22041;
w22164 <= not w22162 and w22163;
w22165 <= not w22158 and not w22164;
w22166 <= pi0781 and not w22165;
w22167 <= not pi0781 and not w22152;
w22168 <= not w22166 and not w22167;
w22169 <= not pi0789 and w22168;
w22170 <= pi0619 and not w21976;
w22171 <= not pi0619 and not w22168;
w22172 <= not pi1159 and not w22170;
w22173 <= not w22171 and w22172;
w22174 <= not pi0648 and not w22049;
w22175 <= not w22173 and w22174;
w22176 <= pi0619 and not w22168;
w22177 <= not pi0619 and not w21976;
w22178 <= pi1159 and not w22177;
w22179 <= not w22176 and w22178;
w22180 <= pi0648 and not w22053;
w22181 <= not w22179 and w22180;
w22182 <= pi0789 and not w22175;
w22183 <= not w22181 and w22182;
w22184 <= w15533 and not w22169;
w22185 <= not w22183 and w22184;
w22186 <= not w22105 and not w22185;
w22187 <= not w22093 and not w22186;
w22188 <= w17927 and w22092;
w22189 <= not w17769 and not w22188;
w22190 <= not w22187 and w22189;
w22191 <= not pi0644 and w22078;
w22192 <= pi0644 and w22070;
w22193 <= pi0790 and not w22191;
w22194 <= not w22192 and w22193;
w22195 <= not w22087 and not w22190;
w22196 <= not w22194 and w22195;
w22197 <= not w22081 and not w22196;
w22198 <= w4989 and not w22197;
w22199 <= not pi0832 and not w21943;
w22200 <= not w22198 and w22199;
w22201 <= not w21942 and not w22200;
w22202 <= not pi0177 and not w14622;
w22203 <= w14198 and not w22202;
w22204 <= pi0177 and not w134;
w22205 <= not pi0177 and w15635;
w22206 <= pi0177 and not w15639;
w22207 <= not pi0038 and not w22206;
w22208 <= not w22205 and w22207;
w22209 <= not pi0177 and not w14204;
w22210 <= w14210 and not w22209;
w22211 <= not pi0686 and not w22210;
w22212 <= not w22208 and w22211;
w22213 <= not pi0177 and pi0686;
w22214 <= not w14615 and w22213;
w22215 <= w134 and not w22214;
w22216 <= not w22212 and w22215;
w22217 <= not w22204 and not w22216;
w22218 <= not pi0778 and not w22217;
w22219 <= not pi0625 and w22202;
w22220 <= pi0625 and w22217;
w22221 <= pi1153 and not w22219;
w22222 <= not w22220 and w22221;
w22223 <= not pi0625 and w22217;
w22224 <= pi0625 and w22202;
w22225 <= not pi1153 and not w22224;
w22226 <= not w22223 and w22225;
w22227 <= not w22222 and not w22226;
w22228 <= pi0778 and not w22227;
w22229 <= not w22218 and not w22228;
w22230 <= not w14638 and not w22229;
w22231 <= w14638 and not w22202;
w22232 <= not w22230 and not w22231;
w22233 <= not w14202 and w22232;
w22234 <= w14202 and w22202;
w22235 <= not w22233 and not w22234;
w22236 <= not w14198 and w22235;
w22237 <= not w22203 and not w22236;
w22238 <= not w14194 and w22237;
w22239 <= w14194 and w22202;
w22240 <= not w22238 and not w22239;
w22241 <= not pi0792 and w22240;
w22242 <= not pi0628 and w22202;
w22243 <= pi0628 and not w22240;
w22244 <= pi1156 and not w22242;
w22245 <= not w22243 and w22244;
w22246 <= pi0628 and w22202;
w22247 <= not pi0628 and not w22240;
w22248 <= not pi1156 and not w22246;
w22249 <= not w22247 and w22248;
w22250 <= not w22245 and not w22249;
w22251 <= pi0792 and not w22250;
w22252 <= not w22241 and not w22251;
w22253 <= not pi0787 and not w22252;
w22254 <= not pi0647 and w22202;
w22255 <= pi0647 and w22252;
w22256 <= pi1157 and not w22254;
w22257 <= not w22255 and w22256;
w22258 <= not pi0647 and w22252;
w22259 <= pi0647 and w22202;
w22260 <= not pi1157 and not w22259;
w22261 <= not w22258 and w22260;
w22262 <= not w22257 and not w22261;
w22263 <= pi0787 and not w22262;
w22264 <= not w22253 and not w22263;
w22265 <= not pi0644 and w22264;
w22266 <= not pi0619 and w22202;
w22267 <= not pi0757 and not w17002;
w22268 <= not w19209 and not w22267;
w22269 <= not pi0177 and not w22268;
w22270 <= not pi0177 and not w16996;
w22271 <= not pi0757 and not w22270;
w22272 <= not w22010 and w22271;
w22273 <= not w22269 and not w22272;
w22274 <= w134 and w22273;
w22275 <= not w22204 and not w22274;
w22276 <= not w14680 and not w22275;
w22277 <= w14680 and not w22202;
w22278 <= not w22276 and not w22277;
w22279 <= not pi0785 and not w22278;
w22280 <= not w14854 and not w22202;
w22281 <= pi0609 and w22276;
w22282 <= not w22280 and not w22281;
w22283 <= pi1155 and not w22282;
w22284 <= not w14859 and not w22202;
w22285 <= not pi0609 and w22276;
w22286 <= not w22284 and not w22285;
w22287 <= not pi1155 and not w22286;
w22288 <= not w22283 and not w22287;
w22289 <= pi0785 and not w22288;
w22290 <= not w22279 and not w22289;
w22291 <= not pi0781 and not w22290;
w22292 <= not pi0618 and w22202;
w22293 <= pi0618 and w22290;
w22294 <= pi1154 and not w22292;
w22295 <= not w22293 and w22294;
w22296 <= not pi0618 and w22290;
w22297 <= pi0618 and w22202;
w22298 <= not pi1154 and not w22297;
w22299 <= not w22296 and w22298;
w22300 <= not w22295 and not w22299;
w22301 <= pi0781 and not w22300;
w22302 <= not w22291 and not w22301;
w22303 <= pi0619 and w22302;
w22304 <= pi1159 and not w22266;
w22305 <= not w22303 and w22304;
w22306 <= w15739 and not w22209;
w22307 <= not pi0177 and w17038;
w22308 <= pi0177 and w17030;
w22309 <= not pi0038 and not w22308;
w22310 <= not w22307 and w22309;
w22311 <= pi0757 and not w22306;
w22312 <= not w22310 and w22311;
w22313 <= not pi0177 and not w17048;
w22314 <= pi0177 and w17053;
w22315 <= pi0038 and not w22314;
w22316 <= not w22313 and w22315;
w22317 <= not w17045 and not w17047;
w22318 <= not pi0177 and not w22317;
w22319 <= pi0177 and w17057;
w22320 <= not pi0038 and not w22318;
w22321 <= not w22319 and w22320;
w22322 <= not pi0757 and not w22316;
w22323 <= not w22321 and w22322;
w22324 <= not w22312 and not w22323;
w22325 <= not pi0686 and not w22324;
w22326 <= pi0686 and not w22273;
w22327 <= w134 and not w22325;
w22328 <= not w22326 and w22327;
w22329 <= not w22204 and not w22328;
w22330 <= not pi0625 and w22329;
w22331 <= pi0625 and w22275;
w22332 <= not pi1153 and not w22331;
w22333 <= not w22330 and w22332;
w22334 <= not pi0608 and not w22222;
w22335 <= not w22333 and w22334;
w22336 <= not pi0625 and w22275;
w22337 <= pi0625 and w22329;
w22338 <= pi1153 and not w22336;
w22339 <= not w22337 and w22338;
w22340 <= pi0608 and not w22226;
w22341 <= not w22339 and w22340;
w22342 <= not w22335 and not w22341;
w22343 <= pi0778 and not w22342;
w22344 <= not pi0778 and w22329;
w22345 <= not w22343 and not w22344;
w22346 <= not pi0609 and not w22345;
w22347 <= pi0609 and w22229;
w22348 <= not pi1155 and not w22347;
w22349 <= not w22346 and w22348;
w22350 <= not pi0660 and not w22283;
w22351 <= not w22349 and w22350;
w22352 <= not pi0609 and w22229;
w22353 <= pi0609 and not w22345;
w22354 <= pi1155 and not w22352;
w22355 <= not w22353 and w22354;
w22356 <= pi0660 and not w22287;
w22357 <= not w22355 and w22356;
w22358 <= not w22351 and not w22357;
w22359 <= pi0785 and not w22358;
w22360 <= not pi0785 and not w22345;
w22361 <= not w22359 and not w22360;
w22362 <= not pi0618 and not w22361;
w22363 <= pi0618 and w22232;
w22364 <= not pi1154 and not w22363;
w22365 <= not w22362 and w22364;
w22366 <= not pi0627 and not w22295;
w22367 <= not w22365 and w22366;
w22368 <= not pi0618 and w22232;
w22369 <= pi0618 and not w22361;
w22370 <= pi1154 and not w22368;
w22371 <= not w22369 and w22370;
w22372 <= pi0627 and not w22299;
w22373 <= not w22371 and w22372;
w22374 <= not w22367 and not w22373;
w22375 <= pi0781 and not w22374;
w22376 <= not pi0781 and not w22361;
w22377 <= not w22375 and not w22376;
w22378 <= not pi0619 and not w22377;
w22379 <= pi0619 and not w22235;
w22380 <= not pi1159 and not w22379;
w22381 <= not w22378 and w22380;
w22382 <= not pi0648 and not w22305;
w22383 <= not w22381 and w22382;
w22384 <= not pi0619 and w22302;
w22385 <= pi0619 and w22202;
w22386 <= not pi1159 and not w22385;
w22387 <= not w22384 and w22386;
w22388 <= pi0619 and not w22377;
w22389 <= not pi0619 and not w22235;
w22390 <= pi1159 and not w22389;
w22391 <= not w22388 and w22390;
w22392 <= pi0648 and not w22387;
w22393 <= not w22391 and w22392;
w22394 <= not w22383 and not w22393;
w22395 <= pi0789 and not w22394;
w22396 <= not pi0789 and not w22377;
w22397 <= not w22395 and not w22396;
w22398 <= not pi0788 and w22397;
w22399 <= not pi0626 and w22397;
w22400 <= pi0626 and not w22237;
w22401 <= not pi0641 and not w22400;
w22402 <= not w22399 and w22401;
w22403 <= not pi0789 and not w22302;
w22404 <= not w22305 and not w22387;
w22405 <= pi0789 and not w22404;
w22406 <= not w22403 and not w22405;
w22407 <= not pi0626 and not w22406;
w22408 <= pi0626 and not w22202;
w22409 <= pi0641 and not w22408;
w22410 <= not w22407 and w22409;
w22411 <= not pi1158 and not w22410;
w22412 <= not w22402 and w22411;
w22413 <= pi0626 and w22397;
w22414 <= not pi0626 and not w22237;
w22415 <= pi0641 and not w22414;
w22416 <= not w22413 and w22415;
w22417 <= pi0626 and not w22406;
w22418 <= not pi0626 and not w22202;
w22419 <= not pi0641 and not w22418;
w22420 <= not w22417 and w22419;
w22421 <= pi1158 and not w22420;
w22422 <= not w22416 and w22421;
w22423 <= not w22412 and not w22422;
w22424 <= pi0788 and not w22423;
w22425 <= not w22398 and not w22424;
w22426 <= not pi0628 and w22425;
w22427 <= not w15532 and w22406;
w22428 <= w15532 and w22202;
w22429 <= not w22427 and not w22428;
w22430 <= pi0628 and not w22429;
w22431 <= not pi1156 and not w22430;
w22432 <= not w22426 and w22431;
w22433 <= not pi0629 and not w22245;
w22434 <= not w22432 and w22433;
w22435 <= pi0628 and w22425;
w22436 <= not pi0628 and not w22429;
w22437 <= pi1156 and not w22436;
w22438 <= not w22435 and w22437;
w22439 <= pi0629 and not w22249;
w22440 <= not w22438 and w22439;
w22441 <= not w22434 and not w22440;
w22442 <= pi0792 and not w22441;
w22443 <= not pi0792 and w22425;
w22444 <= not w22442 and not w22443;
w22445 <= not pi0647 and not w22444;
w22446 <= not w15342 and not w22429;
w22447 <= w15342 and w22202;
w22448 <= not w22446 and not w22447;
w22449 <= pi0647 and not w22448;
w22450 <= not pi1157 and not w22449;
w22451 <= not w22445 and w22450;
w22452 <= not pi0630 and not w22257;
w22453 <= not w22451 and w22452;
w22454 <= pi0647 and not w22444;
w22455 <= not pi0647 and not w22448;
w22456 <= pi1157 and not w22455;
w22457 <= not w22454 and w22456;
w22458 <= pi0630 and not w22261;
w22459 <= not w22457 and w22458;
w22460 <= not w22453 and not w22459;
w22461 <= pi0787 and not w22460;
w22462 <= not pi0787 and not w22444;
w22463 <= not w22461 and not w22462;
w22464 <= pi0644 and not w22463;
w22465 <= pi0715 and not w22265;
w22466 <= not w22464 and w22465;
w22467 <= w15367 and not w22202;
w22468 <= not w15367 and w22448;
w22469 <= not w22467 and not w22468;
w22470 <= pi0644 and w22469;
w22471 <= not pi0644 and w22202;
w22472 <= not pi0715 and not w22471;
w22473 <= not w22470 and w22472;
w22474 <= pi1160 and not w22473;
w22475 <= not w22466 and w22474;
w22476 <= not pi0644 and not w22463;
w22477 <= pi0644 and w22264;
w22478 <= not pi0715 and not w22477;
w22479 <= not w22476 and w22478;
w22480 <= not pi0644 and w22469;
w22481 <= pi0644 and w22202;
w22482 <= pi0715 and not w22481;
w22483 <= not w22480 and w22482;
w22484 <= not pi1160 and not w22483;
w22485 <= not w22479 and w22484;
w22486 <= pi0790 and not w22475;
w22487 <= not w22485 and w22486;
w22488 <= not pi0790 and w22463;
w22489 <= w4989 and not w22488;
w22490 <= not w22487 and w22489;
w22491 <= not pi0177 and not w4989;
w22492 <= not pi0832 and not w22491;
w22493 <= not w22490 and w22492;
w22494 <= not pi0177 and not w489;
w22495 <= not pi0686 and w14208;
w22496 <= not w22494 and not w22495;
w22497 <= not pi0778 and w22496;
w22498 <= not pi0625 and w22495;
w22499 <= not w22496 and not w22498;
w22500 <= pi1153 and not w22499;
w22501 <= not pi1153 and not w22494;
w22502 <= not w22498 and w22501;
w22503 <= not w22500 and not w22502;
w22504 <= pi0778 and not w22503;
w22505 <= not w22497 and not w22504;
w22506 <= not w15408 and w22505;
w22507 <= not w15410 and w22506;
w22508 <= not w15412 and w22507;
w22509 <= not w15414 and w22508;
w22510 <= not w15420 and w22509;
w22511 <= not pi0647 and w22510;
w22512 <= pi0647 and w22494;
w22513 <= not pi1157 and not w22512;
w22514 <= not w22511 and w22513;
w22515 <= pi0630 and w22514;
w22516 <= not pi0757 and w14807;
w22517 <= not w22494 and not w22516;
w22518 <= not w15437 and not w22517;
w22519 <= not pi0785 and not w22518;
w22520 <= not w15442 and not w22517;
w22521 <= pi1155 and not w22520;
w22522 <= not w15445 and w22518;
w22523 <= not pi1155 and not w22522;
w22524 <= not w22521 and not w22523;
w22525 <= pi0785 and not w22524;
w22526 <= not w22519 and not w22525;
w22527 <= not pi0781 and not w22526;
w22528 <= not w15452 and w22526;
w22529 <= pi1154 and not w22528;
w22530 <= not w15455 and w22526;
w22531 <= not pi1154 and not w22530;
w22532 <= not w22529 and not w22531;
w22533 <= pi0781 and not w22532;
w22534 <= not w22527 and not w22533;
w22535 <= not pi0789 and not w22534;
w22536 <= not pi0619 and w22494;
w22537 <= pi0619 and w22534;
w22538 <= pi1159 and not w22536;
w22539 <= not w22537 and w22538;
w22540 <= not pi0619 and w22534;
w22541 <= pi0619 and w22494;
w22542 <= not pi1159 and not w22541;
w22543 <= not w22540 and w22542;
w22544 <= not w22539 and not w22543;
w22545 <= pi0789 and not w22544;
w22546 <= not w22535 and not w22545;
w22547 <= not w15532 and w22546;
w22548 <= w15532 and w22494;
w22549 <= not w22547 and not w22548;
w22550 <= not w15342 and not w22549;
w22551 <= w15342 and w22494;
w22552 <= not w22550 and not w22551;
w22553 <= not w18122 and w22552;
w22554 <= pi0647 and not w22510;
w22555 <= not pi0647 and not w22494;
w22556 <= not w22554 and not w22555;
w22557 <= w15364 and not w22556;
w22558 <= not w22515 and not w22557;
w22559 <= not w22553 and w22558;
w22560 <= pi0787 and not w22559;
w22561 <= w15434 and w22508;
w22562 <= not pi0626 and not w22546;
w22563 <= pi0626 and not w22494;
w22564 <= w14192 and not w22563;
w22565 <= not w22562 and w22564;
w22566 <= pi0626 and not w22546;
w22567 <= not pi0626 and not w22494;
w22568 <= w14191 and not w22567;
w22569 <= not w22566 and w22568;
w22570 <= not w22561 and not w22565;
w22571 <= not w22569 and w22570;
w22572 <= pi0788 and not w22571;
w22573 <= pi0618 and w22506;
w22574 <= pi0609 and w22505;
w22575 <= not w14731 and not w22496;
w22576 <= pi0625 and w22575;
w22577 <= w22517 and not w22575;
w22578 <= not w22576 and not w22577;
w22579 <= w22501 and not w22578;
w22580 <= not pi0608 and not w22500;
w22581 <= not w22579 and w22580;
w22582 <= pi1153 and w22517;
w22583 <= not w22576 and w22582;
w22584 <= pi0608 and not w22502;
w22585 <= not w22583 and w22584;
w22586 <= not w22581 and not w22585;
w22587 <= pi0778 and not w22586;
w22588 <= not pi0778 and not w22577;
w22589 <= not w22587 and not w22588;
w22590 <= not pi0609 and not w22589;
w22591 <= not pi1155 and not w22574;
w22592 <= not w22590 and w22591;
w22593 <= not pi0660 and not w22521;
w22594 <= not w22592 and w22593;
w22595 <= not pi0609 and w22505;
w22596 <= pi0609 and not w22589;
w22597 <= pi1155 and not w22595;
w22598 <= not w22596 and w22597;
w22599 <= pi0660 and not w22523;
w22600 <= not w22598 and w22599;
w22601 <= not w22594 and not w22600;
w22602 <= pi0785 and not w22601;
w22603 <= not pi0785 and not w22589;
w22604 <= not w22602 and not w22603;
w22605 <= not pi0618 and not w22604;
w22606 <= not pi1154 and not w22573;
w22607 <= not w22605 and w22606;
w22608 <= not pi0627 and not w22529;
w22609 <= not w22607 and w22608;
w22610 <= not pi0618 and w22506;
w22611 <= pi0618 and not w22604;
w22612 <= pi1154 and not w22610;
w22613 <= not w22611 and w22612;
w22614 <= pi0627 and not w22531;
w22615 <= not w22613 and w22614;
w22616 <= not w22609 and not w22615;
w22617 <= pi0781 and not w22616;
w22618 <= not pi0781 and not w22604;
w22619 <= not w22617 and not w22618;
w22620 <= not pi0789 and w22619;
w22621 <= not pi0619 and not w22619;
w22622 <= pi0619 and w22507;
w22623 <= not pi1159 and not w22622;
w22624 <= not w22621 and w22623;
w22625 <= not pi0648 and not w22539;
w22626 <= not w22624 and w22625;
w22627 <= pi0619 and not w22619;
w22628 <= not pi0619 and w22507;
w22629 <= pi1159 and not w22628;
w22630 <= not w22627 and w22629;
w22631 <= pi0648 and not w22543;
w22632 <= not w22630 and w22631;
w22633 <= pi0789 and not w22626;
w22634 <= not w22632 and w22633;
w22635 <= w15533 and not w22620;
w22636 <= not w22634 and w22635;
w22637 <= not w22572 and not w22636;
w22638 <= not w17927 and not w22637;
w22639 <= w15417 and not w22549;
w22640 <= w18414 and w22509;
w22641 <= not w22639 and not w22640;
w22642 <= not pi0629 and not w22641;
w22643 <= w18418 and w22509;
w22644 <= w15416 and not w22549;
w22645 <= not w22643 and not w22644;
w22646 <= pi0629 and not w22645;
w22647 <= not w22642 and not w22646;
w22648 <= pi0792 and not w22647;
w22649 <= not w17769 and not w22648;
w22650 <= not w22638 and w22649;
w22651 <= not w22560 and not w22650;
w22652 <= not pi0790 and w22651;
w22653 <= not pi0787 and not w22510;
w22654 <= pi1157 and not w22556;
w22655 <= not w22514 and not w22654;
w22656 <= pi0787 and not w22655;
w22657 <= not w22653 and not w22656;
w22658 <= not pi0644 and w22657;
w22659 <= pi0644 and w22651;
w22660 <= pi0715 and not w22658;
w22661 <= not w22659 and w22660;
w22662 <= not w15367 and not w22552;
w22663 <= w15367 and w22494;
w22664 <= not w22662 and not w22663;
w22665 <= pi0644 and not w22664;
w22666 <= not pi0644 and w22494;
w22667 <= not pi0715 and not w22666;
w22668 <= not w22665 and w22667;
w22669 <= pi1160 and not w22668;
w22670 <= not w22661 and w22669;
w22671 <= not pi0644 and not w22664;
w22672 <= pi0644 and w22494;
w22673 <= pi0715 and not w22672;
w22674 <= not w22671 and w22673;
w22675 <= pi0644 and w22657;
w22676 <= not pi0644 and w22651;
w22677 <= not pi0715 and not w22675;
w22678 <= not w22676 and w22677;
w22679 <= not pi1160 and not w22674;
w22680 <= not w22678 and w22679;
w22681 <= not w22670 and not w22680;
w22682 <= pi0790 and not w22681;
w22683 <= pi0832 and not w22652;
w22684 <= not w22682 and w22683;
w22685 <= not w22493 and not w22684;
w22686 <= not pi0178 and not w489;
w22687 <= not pi0688 and w14208;
w22688 <= not w22686 and not w22687;
w22689 <= not pi0778 and not w22688;
w22690 <= not pi0625 and w22687;
w22691 <= not w22688 and not w22690;
w22692 <= pi1153 and not w22691;
w22693 <= not pi1153 and not w22686;
w22694 <= not w22690 and w22693;
w22695 <= pi0778 and not w22694;
w22696 <= not w22692 and w22695;
w22697 <= not w22689 and not w22696;
w22698 <= not w15408 and not w22697;
w22699 <= not w15410 and w22698;
w22700 <= not w15412 and w22699;
w22701 <= not w15414 and w22700;
w22702 <= not w15420 and w22701;
w22703 <= not pi0647 and w22702;
w22704 <= pi0647 and w22686;
w22705 <= not pi1157 and not w22704;
w22706 <= not w22703 and w22705;
w22707 <= pi0630 and w22706;
w22708 <= not pi0760 and w14807;
w22709 <= not w22686 and not w22708;
w22710 <= not w15437 and not w22709;
w22711 <= not pi0785 and not w22710;
w22712 <= w14859 and w22708;
w22713 <= w22710 and not w22712;
w22714 <= pi1155 and not w22713;
w22715 <= not pi1155 and not w22686;
w22716 <= not w22712 and w22715;
w22717 <= not w22714 and not w22716;
w22718 <= pi0785 and not w22717;
w22719 <= not w22711 and not w22718;
w22720 <= not pi0781 and not w22719;
w22721 <= not w15452 and w22719;
w22722 <= pi1154 and not w22721;
w22723 <= not w15455 and w22719;
w22724 <= not pi1154 and not w22723;
w22725 <= not w22722 and not w22724;
w22726 <= pi0781 and not w22725;
w22727 <= not w22720 and not w22726;
w22728 <= not pi0789 and not w22727;
w22729 <= not w20641 and w22727;
w22730 <= pi1159 and not w22729;
w22731 <= not w20644 and w22727;
w22732 <= not pi1159 and not w22731;
w22733 <= not w22730 and not w22732;
w22734 <= pi0789 and not w22733;
w22735 <= not w22728 and not w22734;
w22736 <= not w15532 and w22735;
w22737 <= w15532 and w22686;
w22738 <= not w22736 and not w22737;
w22739 <= not w15342 and not w22738;
w22740 <= w15342 and w22686;
w22741 <= not w22739 and not w22740;
w22742 <= not w18122 and w22741;
w22743 <= pi0647 and not w22702;
w22744 <= not pi0647 and not w22686;
w22745 <= not w22743 and not w22744;
w22746 <= w15364 and not w22745;
w22747 <= not w22707 and not w22746;
w22748 <= not w22742 and w22747;
w22749 <= pi0787 and not w22748;
w22750 <= w15434 and w22700;
w22751 <= not pi0626 and not w22735;
w22752 <= pi0626 and not w22686;
w22753 <= w14192 and not w22752;
w22754 <= not w22751 and w22753;
w22755 <= pi0626 and not w22735;
w22756 <= not pi0626 and not w22686;
w22757 <= w14191 and not w22756;
w22758 <= not w22755 and w22757;
w22759 <= not w22750 and not w22754;
w22760 <= not w22758 and w22759;
w22761 <= pi0788 and not w22760;
w22762 <= pi0618 and w22698;
w22763 <= not w14731 and not w22688;
w22764 <= pi0625 and w22763;
w22765 <= w22709 and not w22763;
w22766 <= not w22764 and not w22765;
w22767 <= w22693 and not w22766;
w22768 <= not pi0608 and not w22692;
w22769 <= not w22767 and w22768;
w22770 <= pi1153 and w22709;
w22771 <= not w22764 and w22770;
w22772 <= pi0608 and not w22694;
w22773 <= not w22771 and w22772;
w22774 <= not w22769 and not w22773;
w22775 <= pi0778 and not w22774;
w22776 <= not pi0778 and not w22765;
w22777 <= not w22775 and not w22776;
w22778 <= not pi0609 and not w22777;
w22779 <= pi0609 and not w22697;
w22780 <= not pi1155 and not w22779;
w22781 <= not w22778 and w22780;
w22782 <= not pi0660 and not w22714;
w22783 <= not w22781 and w22782;
w22784 <= pi0609 and not w22777;
w22785 <= not pi0609 and not w22697;
w22786 <= pi1155 and not w22785;
w22787 <= not w22784 and w22786;
w22788 <= pi0660 and not w22716;
w22789 <= not w22787 and w22788;
w22790 <= not w22783 and not w22789;
w22791 <= pi0785 and not w22790;
w22792 <= not pi0785 and not w22777;
w22793 <= not w22791 and not w22792;
w22794 <= not pi0618 and not w22793;
w22795 <= not pi1154 and not w22762;
w22796 <= not w22794 and w22795;
w22797 <= not pi0627 and not w22722;
w22798 <= not w22796 and w22797;
w22799 <= not pi0618 and w22698;
w22800 <= pi0618 and not w22793;
w22801 <= pi1154 and not w22799;
w22802 <= not w22800 and w22801;
w22803 <= pi0627 and not w22724;
w22804 <= not w22802 and w22803;
w22805 <= not w22798 and not w22804;
w22806 <= pi0781 and not w22805;
w22807 <= not pi0781 and not w22793;
w22808 <= not w22806 and not w22807;
w22809 <= not pi0789 and w22808;
w22810 <= not pi0619 and not w22808;
w22811 <= pi0619 and w22699;
w22812 <= not pi1159 and not w22811;
w22813 <= not w22810 and w22812;
w22814 <= not pi0648 and not w22730;
w22815 <= not w22813 and w22814;
w22816 <= pi0619 and not w22808;
w22817 <= not pi0619 and w22699;
w22818 <= pi1159 and not w22817;
w22819 <= not w22816 and w22818;
w22820 <= pi0648 and not w22732;
w22821 <= not w22819 and w22820;
w22822 <= pi0789 and not w22815;
w22823 <= not w22821 and w22822;
w22824 <= w15533 and not w22809;
w22825 <= not w22823 and w22824;
w22826 <= not w22761 and not w22825;
w22827 <= not w17927 and not w22826;
w22828 <= w15417 and not w22738;
w22829 <= w18414 and w22701;
w22830 <= not w22828 and not w22829;
w22831 <= not pi0629 and not w22830;
w22832 <= w18418 and w22701;
w22833 <= w15416 and not w22738;
w22834 <= not w22832 and not w22833;
w22835 <= pi0629 and not w22834;
w22836 <= not w22831 and not w22835;
w22837 <= pi0792 and not w22836;
w22838 <= not w17769 and not w22837;
w22839 <= not w22827 and w22838;
w22840 <= not w22749 and not w22839;
w22841 <= not pi0790 and w22840;
w22842 <= not pi0787 and not w22702;
w22843 <= pi1157 and not w22745;
w22844 <= not w22706 and not w22843;
w22845 <= pi0787 and not w22844;
w22846 <= not w22842 and not w22845;
w22847 <= not pi0644 and w22846;
w22848 <= pi0644 and w22840;
w22849 <= pi0715 and not w22847;
w22850 <= not w22848 and w22849;
w22851 <= not w15367 and not w22741;
w22852 <= w15367 and w22686;
w22853 <= not w22851 and not w22852;
w22854 <= pi0644 and not w22853;
w22855 <= not pi0644 and w22686;
w22856 <= not pi0715 and not w22855;
w22857 <= not w22854 and w22856;
w22858 <= pi1160 and not w22857;
w22859 <= not w22850 and w22858;
w22860 <= not pi0644 and not w22853;
w22861 <= pi0644 and w22686;
w22862 <= pi0715 and not w22861;
w22863 <= not w22860 and w22862;
w22864 <= pi0644 and w22846;
w22865 <= not pi0644 and w22840;
w22866 <= not pi0715 and not w22864;
w22867 <= not w22865 and w22866;
w22868 <= not pi1160 and not w22863;
w22869 <= not w22867 and w22868;
w22870 <= not w22859 and not w22869;
w22871 <= pi0790 and not w22870;
w22872 <= pi0832 and not w22841;
w22873 <= not w22871 and w22872;
w22874 <= not pi0178 and not w4989;
w22875 <= not pi0178 and not w14622;
w22876 <= w14198 and not w22875;
w22877 <= not pi0688 and w134;
w22878 <= w22875 and not w22877;
w22879 <= not pi0178 and not w14204;
w22880 <= w14210 and not w22879;
w22881 <= pi0178 and not w15639;
w22882 <= not pi0038 and not w22881;
w22883 <= w134 and not w22882;
w22884 <= not pi0178 and w15635;
w22885 <= not w22883 and not w22884;
w22886 <= not pi0688 and not w22880;
w22887 <= not w22885 and w22886;
w22888 <= not w22878 and not w22887;
w22889 <= not pi0778 and w22888;
w22890 <= not pi0625 and w22875;
w22891 <= pi0625 and not w22888;
w22892 <= pi1153 and not w22890;
w22893 <= not w22891 and w22892;
w22894 <= pi0625 and w22875;
w22895 <= not pi0625 and not w22888;
w22896 <= not pi1153 and not w22894;
w22897 <= not w22895 and w22896;
w22898 <= not w22893 and not w22897;
w22899 <= pi0778 and not w22898;
w22900 <= not w22889 and not w22899;
w22901 <= not w14638 and not w22900;
w22902 <= w14638 and not w22875;
w22903 <= not w22901 and not w22902;
w22904 <= not w14202 and w22903;
w22905 <= w14202 and w22875;
w22906 <= not w22904 and not w22905;
w22907 <= not w14198 and w22906;
w22908 <= not w22876 and not w22907;
w22909 <= not w14194 and w22908;
w22910 <= w14194 and w22875;
w22911 <= not w22909 and not w22910;
w22912 <= not pi0792 and w22911;
w22913 <= pi0628 and not w22911;
w22914 <= not pi0628 and w22875;
w22915 <= pi1156 and not w22914;
w22916 <= not w22913 and w22915;
w22917 <= pi0628 and w22875;
w22918 <= not pi0628 and not w22911;
w22919 <= not pi1156 and not w22917;
w22920 <= not w22918 and w22919;
w22921 <= not w22916 and not w22920;
w22922 <= pi0792 and not w22921;
w22923 <= not w22912 and not w22922;
w22924 <= not pi0647 and not w22923;
w22925 <= pi0647 and not w22875;
w22926 <= not w22924 and not w22925;
w22927 <= not pi1157 and w22926;
w22928 <= pi0647 and not w22923;
w22929 <= not pi0647 and not w22875;
w22930 <= not w22928 and not w22929;
w22931 <= pi1157 and w22930;
w22932 <= not w22927 and not w22931;
w22933 <= pi0787 and not w22932;
w22934 <= not pi0787 and w22923;
w22935 <= not w22933 and not w22934;
w22936 <= not pi0644 and not w22935;
w22937 <= pi0715 and not w22936;
w22938 <= pi0178 and not w134;
w22939 <= not pi0760 and w14843;
w22940 <= not w22879 and not w22939;
w22941 <= pi0038 and not w22940;
w22942 <= not pi0178 and w14784;
w22943 <= pi0178 and not w14838;
w22944 <= not pi0760 and not w22943;
w22945 <= not w22942 and w22944;
w22946 <= not pi0178 and pi0760;
w22947 <= not w14611 and w22946;
w22948 <= not w22945 and not w22947;
w22949 <= not pi0038 and not w22948;
w22950 <= not w22941 and not w22949;
w22951 <= w134 and w22950;
w22952 <= not w22938 and not w22951;
w22953 <= not w14680 and not w22952;
w22954 <= w14680 and not w22875;
w22955 <= not w22953 and not w22954;
w22956 <= not pi0785 and not w22955;
w22957 <= not w14854 and not w22875;
w22958 <= pi0609 and w22953;
w22959 <= not w22957 and not w22958;
w22960 <= pi1155 and not w22959;
w22961 <= not w14859 and not w22875;
w22962 <= not pi0609 and w22953;
w22963 <= not w22961 and not w22962;
w22964 <= not pi1155 and not w22963;
w22965 <= not w22960 and not w22964;
w22966 <= pi0785 and not w22965;
w22967 <= not w22956 and not w22966;
w22968 <= not pi0781 and not w22967;
w22969 <= not pi0618 and w22875;
w22970 <= pi0618 and w22967;
w22971 <= pi1154 and not w22969;
w22972 <= not w22970 and w22971;
w22973 <= not pi0618 and w22967;
w22974 <= pi0618 and w22875;
w22975 <= not pi1154 and not w22974;
w22976 <= not w22973 and w22975;
w22977 <= not w22972 and not w22976;
w22978 <= pi0781 and not w22977;
w22979 <= not w22968 and not w22978;
w22980 <= not pi0789 and not w22979;
w22981 <= not pi0619 and w22875;
w22982 <= pi0619 and w22979;
w22983 <= pi1159 and not w22981;
w22984 <= not w22982 and w22983;
w22985 <= not pi0619 and w22979;
w22986 <= pi0619 and w22875;
w22987 <= not pi1159 and not w22986;
w22988 <= not w22985 and w22987;
w22989 <= not w22984 and not w22988;
w22990 <= pi0789 and not w22989;
w22991 <= not w22980 and not w22990;
w22992 <= not w15532 and w22991;
w22993 <= w15532 and w22875;
w22994 <= not w22992 and not w22993;
w22995 <= not w15342 and not w22994;
w22996 <= w15342 and w22875;
w22997 <= not w22995 and not w22996;
w22998 <= not w15367 and not w22997;
w22999 <= w15367 and w22875;
w23000 <= not w22998 and not w22999;
w23001 <= pi0644 and not w23000;
w23002 <= not pi0644 and w22875;
w23003 <= not pi0715 and not w23002;
w23004 <= not w23001 and w23003;
w23005 <= pi1160 and not w23004;
w23006 <= not w22937 and w23005;
w23007 <= pi0644 and not w22935;
w23008 <= not pi0715 and not w23007;
w23009 <= not pi0644 and not w23000;
w23010 <= pi0644 and w22875;
w23011 <= pi0715 and not w23010;
w23012 <= not w23009 and w23011;
w23013 <= not pi1160 and not w23012;
w23014 <= not w23008 and w23013;
w23015 <= not w23006 and not w23014;
w23016 <= pi0790 and not w23015;
w23017 <= not pi0629 and w22916;
w23018 <= not w18133 and w22994;
w23019 <= pi0629 and w22920;
w23020 <= not w23017 and not w23019;
w23021 <= not w23018 and w23020;
w23022 <= pi0792 and not w23021;
w23023 <= pi0609 and w22900;
w23024 <= pi0178 and not w15188;
w23025 <= not pi0178 and not w15175;
w23026 <= pi0760 and not w23024;
w23027 <= not w23025 and w23026;
w23028 <= not pi0178 and w15192;
w23029 <= pi0178 and w15194;
w23030 <= not pi0760 and not w23029;
w23031 <= not w23028 and w23030;
w23032 <= not w23027 and not w23031;
w23033 <= not pi0039 and not w23032;
w23034 <= pi0178 and w15168;
w23035 <= not pi0178 and not w15109;
w23036 <= not pi0760 and not w23035;
w23037 <= not w23034 and w23036;
w23038 <= not pi0178 and w14967;
w23039 <= pi0178 and w15048;
w23040 <= pi0760 and not w23039;
w23041 <= not w23038 and w23040;
w23042 <= pi0039 and not w23037;
w23043 <= not w23041 and w23042;
w23044 <= not pi0038 and not w23033;
w23045 <= not w23043 and w23044;
w23046 <= not pi0760 and not w15053;
w23047 <= w17034 and not w23046;
w23048 <= not pi0178 and not w23047;
w23049 <= not w15032 and not w22708;
w23050 <= pi0178 and not w23049;
w23051 <= w3847 and w23050;
w23052 <= pi0038 and not w23051;
w23053 <= not w23048 and w23052;
w23054 <= not pi0688 and not w23053;
w23055 <= not w23045 and w23054;
w23056 <= pi0688 and not w22950;
w23057 <= w134 and not w23055;
w23058 <= not w23056 and w23057;
w23059 <= not w22938 and not w23058;
w23060 <= not pi0625 and w23059;
w23061 <= pi0625 and w22952;
w23062 <= not pi1153 and not w23061;
w23063 <= not w23060 and w23062;
w23064 <= not pi0608 and not w22893;
w23065 <= not w23063 and w23064;
w23066 <= not pi0625 and w22952;
w23067 <= pi0625 and w23059;
w23068 <= pi1153 and not w23066;
w23069 <= not w23067 and w23068;
w23070 <= pi0608 and not w22897;
w23071 <= not w23069 and w23070;
w23072 <= not w23065 and not w23071;
w23073 <= pi0778 and not w23072;
w23074 <= not pi0778 and w23059;
w23075 <= not w23073 and not w23074;
w23076 <= not pi0609 and not w23075;
w23077 <= not pi1155 and not w23023;
w23078 <= not w23076 and w23077;
w23079 <= not pi0660 and not w22960;
w23080 <= not w23078 and w23079;
w23081 <= not pi0609 and w22900;
w23082 <= pi0609 and not w23075;
w23083 <= pi1155 and not w23081;
w23084 <= not w23082 and w23083;
w23085 <= pi0660 and not w22964;
w23086 <= not w23084 and w23085;
w23087 <= not w23080 and not w23086;
w23088 <= pi0785 and not w23087;
w23089 <= not pi0785 and not w23075;
w23090 <= not w23088 and not w23089;
w23091 <= not pi0618 and not w23090;
w23092 <= pi0618 and w22903;
w23093 <= not pi1154 and not w23092;
w23094 <= not w23091 and w23093;
w23095 <= not pi0627 and not w22972;
w23096 <= not w23094 and w23095;
w23097 <= not pi0618 and w22903;
w23098 <= pi0618 and not w23090;
w23099 <= pi1154 and not w23097;
w23100 <= not w23098 and w23099;
w23101 <= pi0627 and not w22976;
w23102 <= not w23100 and w23101;
w23103 <= not w23096 and not w23102;
w23104 <= pi0781 and not w23103;
w23105 <= not pi0781 and not w23090;
w23106 <= not w23104 and not w23105;
w23107 <= not pi0789 and w23106;
w23108 <= pi0619 and not w22906;
w23109 <= not pi0619 and not w23106;
w23110 <= not pi1159 and not w23108;
w23111 <= not w23109 and w23110;
w23112 <= not pi0648 and not w22984;
w23113 <= not w23111 and w23112;
w23114 <= not pi0619 and not w22906;
w23115 <= pi0619 and not w23106;
w23116 <= pi1159 and not w23114;
w23117 <= not w23115 and w23116;
w23118 <= pi0648 and not w22988;
w23119 <= not w23117 and w23118;
w23120 <= pi0789 and not w23113;
w23121 <= not w23119 and w23120;
w23122 <= w15533 and not w23107;
w23123 <= not w23121 and w23122;
w23124 <= w15434 and w22908;
w23125 <= not pi0626 and not w22991;
w23126 <= pi0626 and not w22875;
w23127 <= w14192 and not w23126;
w23128 <= not w23125 and w23127;
w23129 <= pi0626 and not w22991;
w23130 <= not pi0626 and not w22875;
w23131 <= w14191 and not w23130;
w23132 <= not w23129 and w23131;
w23133 <= not w23124 and not w23128;
w23134 <= not w23132 and w23133;
w23135 <= pi0788 and not w23134;
w23136 <= not w17927 and not w23135;
w23137 <= not w23123 and w23136;
w23138 <= not w23022 and not w23137;
w23139 <= not w17769 and not w23138;
w23140 <= w15365 and not w22926;
w23141 <= not w18122 and w22997;
w23142 <= w15364 and not w22930;
w23143 <= not w23140 and not w23142;
w23144 <= not w23141 and w23143;
w23145 <= pi0787 and not w23144;
w23146 <= not pi0644 and w23013;
w23147 <= pi0644 and w23005;
w23148 <= pi0790 and not w23146;
w23149 <= not w23147 and w23148;
w23150 <= not w23139 and not w23145;
w23151 <= not w23149 and w23150;
w23152 <= not w23016 and not w23151;
w23153 <= w4989 and not w23152;
w23154 <= not pi0832 and not w22874;
w23155 <= not w23153 and w23154;
w23156 <= not w22873 and not w23155;
w23157 <= not pi0179 and not w14622;
w23158 <= w14198 and not w23157;
w23159 <= not pi0724 and w134;
w23160 <= w23157 and not w23159;
w23161 <= not pi0179 and not w14204;
w23162 <= w14210 and not w23161;
w23163 <= not pi0179 and w15635;
w23164 <= pi0179 and not w15639;
w23165 <= not pi0038 and not w23164;
w23166 <= w134 and not w23165;
w23167 <= not w23163 and not w23166;
w23168 <= not pi0724 and not w23162;
w23169 <= not w23167 and w23168;
w23170 <= not w23160 and not w23169;
w23171 <= not pi0778 and w23170;
w23172 <= not pi0625 and w23157;
w23173 <= pi0625 and not w23170;
w23174 <= pi1153 and not w23172;
w23175 <= not w23173 and w23174;
w23176 <= pi0625 and w23157;
w23177 <= not pi0625 and not w23170;
w23178 <= not pi1153 and not w23176;
w23179 <= not w23177 and w23178;
w23180 <= not w23175 and not w23179;
w23181 <= pi0778 and not w23180;
w23182 <= not w23171 and not w23181;
w23183 <= not w14638 and not w23182;
w23184 <= w14638 and not w23157;
w23185 <= not w23183 and not w23184;
w23186 <= not w14202 and w23185;
w23187 <= w14202 and w23157;
w23188 <= not w23186 and not w23187;
w23189 <= not w14198 and w23188;
w23190 <= not w23158 and not w23189;
w23191 <= not w14194 and w23190;
w23192 <= w14194 and w23157;
w23193 <= not w23191 and not w23192;
w23194 <= not pi0792 and w23193;
w23195 <= not pi0628 and w23157;
w23196 <= pi0628 and not w23193;
w23197 <= pi1156 and not w23195;
w23198 <= not w23196 and w23197;
w23199 <= pi0628 and w23157;
w23200 <= not pi0628 and not w23193;
w23201 <= not pi1156 and not w23199;
w23202 <= not w23200 and w23201;
w23203 <= not w23198 and not w23202;
w23204 <= pi0792 and not w23203;
w23205 <= not w23194 and not w23204;
w23206 <= not pi0787 and not w23205;
w23207 <= not pi0647 and w23157;
w23208 <= pi0647 and w23205;
w23209 <= pi1157 and not w23207;
w23210 <= not w23208 and w23209;
w23211 <= not pi0647 and w23205;
w23212 <= pi0647 and w23157;
w23213 <= not pi1157 and not w23212;
w23214 <= not w23211 and w23213;
w23215 <= not w23210 and not w23214;
w23216 <= pi0787 and not w23215;
w23217 <= not w23206 and not w23216;
w23218 <= not pi0644 and w23217;
w23219 <= not pi0618 and w23157;
w23220 <= pi0179 and not w134;
w23221 <= not pi0741 and not w22010;
w23222 <= pi0179 and not w23221;
w23223 <= not pi0179 and not pi0741;
w23224 <= not w16996 and w23223;
w23225 <= w17002 and w23224;
w23226 <= not w23222 and not w23225;
w23227 <= not w19237 and w23226;
w23228 <= w134 and not w23227;
w23229 <= not w23220 and not w23228;
w23230 <= not w14680 and not w23229;
w23231 <= w14680 and not w23157;
w23232 <= not w23230 and not w23231;
w23233 <= not pi0785 and not w23232;
w23234 <= not w14854 and not w23157;
w23235 <= pi0609 and w23230;
w23236 <= not w23234 and not w23235;
w23237 <= pi1155 and not w23236;
w23238 <= not w14859 and not w23157;
w23239 <= not pi0609 and w23230;
w23240 <= not w23238 and not w23239;
w23241 <= not pi1155 and not w23240;
w23242 <= not w23237 and not w23241;
w23243 <= pi0785 and not w23242;
w23244 <= not w23233 and not w23243;
w23245 <= pi0618 and w23244;
w23246 <= pi1154 and not w23219;
w23247 <= not w23245 and w23246;
w23248 <= w15739 and not w23161;
w23249 <= not pi0179 and w14967;
w23250 <= pi0179 and w15048;
w23251 <= pi0039 and not w23250;
w23252 <= not w23249 and w23251;
w23253 <= not pi0179 and w15175;
w23254 <= pi0179 and w15188;
w23255 <= not pi0039 and not w23253;
w23256 <= not w23254 and w23255;
w23257 <= not w23252 and not w23256;
w23258 <= not pi0038 and not w23257;
w23259 <= not w23248 and not w23258;
w23260 <= pi0741 and not w23259;
w23261 <= not pi0179 and not w17051;
w23262 <= pi0179 and w17059;
w23263 <= not pi0741 and not w23261;
w23264 <= not w23262 and w23263;
w23265 <= not pi0724 and not w23264;
w23266 <= not w23260 and w23265;
w23267 <= pi0724 and w23227;
w23268 <= w134 and not w23267;
w23269 <= not w23266 and w23268;
w23270 <= not w23220 and not w23269;
w23271 <= not pi0625 and w23270;
w23272 <= pi0625 and w23229;
w23273 <= not pi1153 and not w23272;
w23274 <= not w23271 and w23273;
w23275 <= not pi0608 and not w23175;
w23276 <= not w23274 and w23275;
w23277 <= not pi0625 and w23229;
w23278 <= pi0625 and w23270;
w23279 <= pi1153 and not w23277;
w23280 <= not w23278 and w23279;
w23281 <= pi0608 and not w23179;
w23282 <= not w23280 and w23281;
w23283 <= not w23276 and not w23282;
w23284 <= pi0778 and not w23283;
w23285 <= not pi0778 and w23270;
w23286 <= not w23284 and not w23285;
w23287 <= not pi0609 and not w23286;
w23288 <= pi0609 and w23182;
w23289 <= not pi1155 and not w23288;
w23290 <= not w23287 and w23289;
w23291 <= not pi0660 and not w23237;
w23292 <= not w23290 and w23291;
w23293 <= not pi0609 and w23182;
w23294 <= pi0609 and not w23286;
w23295 <= pi1155 and not w23293;
w23296 <= not w23294 and w23295;
w23297 <= pi0660 and not w23241;
w23298 <= not w23296 and w23297;
w23299 <= not w23292 and not w23298;
w23300 <= pi0785 and not w23299;
w23301 <= not pi0785 and not w23286;
w23302 <= not w23300 and not w23301;
w23303 <= not pi0618 and not w23302;
w23304 <= pi0618 and w23185;
w23305 <= not pi1154 and not w23304;
w23306 <= not w23303 and w23305;
w23307 <= not pi0627 and not w23247;
w23308 <= not w23306 and w23307;
w23309 <= not pi0618 and w23244;
w23310 <= pi0618 and w23157;
w23311 <= not pi1154 and not w23310;
w23312 <= not w23309 and w23311;
w23313 <= not pi0618 and w23185;
w23314 <= pi0618 and not w23302;
w23315 <= pi1154 and not w23313;
w23316 <= not w23314 and w23315;
w23317 <= pi0627 and not w23312;
w23318 <= not w23316 and w23317;
w23319 <= not w23308 and not w23318;
w23320 <= pi0781 and not w23319;
w23321 <= not pi0781 and not w23302;
w23322 <= not w23320 and not w23321;
w23323 <= not pi0619 and not w23322;
w23324 <= pi0619 and not w23188;
w23325 <= not pi1159 and not w23324;
w23326 <= not w23323 and w23325;
w23327 <= not pi0619 and w23157;
w23328 <= not pi0781 and not w23244;
w23329 <= not w23247 and not w23312;
w23330 <= pi0781 and not w23329;
w23331 <= not w23328 and not w23330;
w23332 <= pi0619 and w23331;
w23333 <= pi1159 and not w23327;
w23334 <= not w23332 and w23333;
w23335 <= not pi0648 and not w23334;
w23336 <= not w23326 and w23335;
w23337 <= pi0619 and not w23322;
w23338 <= not pi0619 and not w23188;
w23339 <= pi1159 and not w23338;
w23340 <= not w23337 and w23339;
w23341 <= not pi0619 and w23331;
w23342 <= pi0619 and w23157;
w23343 <= not pi1159 and not w23342;
w23344 <= not w23341 and w23343;
w23345 <= pi0648 and not w23344;
w23346 <= not w23340 and w23345;
w23347 <= not w23336 and not w23346;
w23348 <= pi0789 and not w23347;
w23349 <= not pi0789 and not w23322;
w23350 <= not w23348 and not w23349;
w23351 <= not pi0788 and w23350;
w23352 <= not pi0626 and w23350;
w23353 <= pi0626 and not w23190;
w23354 <= not pi0641 and not w23353;
w23355 <= not w23352 and w23354;
w23356 <= not pi0789 and not w23331;
w23357 <= not w23334 and not w23344;
w23358 <= pi0789 and not w23357;
w23359 <= not w23356 and not w23358;
w23360 <= not pi0626 and not w23359;
w23361 <= pi0626 and not w23157;
w23362 <= pi0641 and not w23361;
w23363 <= not w23360 and w23362;
w23364 <= not pi1158 and not w23363;
w23365 <= not w23355 and w23364;
w23366 <= pi0626 and w23350;
w23367 <= not pi0626 and not w23190;
w23368 <= pi0641 and not w23367;
w23369 <= not w23366 and w23368;
w23370 <= pi0626 and not w23359;
w23371 <= not pi0626 and not w23157;
w23372 <= not pi0641 and not w23371;
w23373 <= not w23370 and w23372;
w23374 <= pi1158 and not w23373;
w23375 <= not w23369 and w23374;
w23376 <= not w23365 and not w23375;
w23377 <= pi0788 and not w23376;
w23378 <= not w23351 and not w23377;
w23379 <= not pi0628 and w23378;
w23380 <= not w15532 and w23359;
w23381 <= w15532 and w23157;
w23382 <= not w23380 and not w23381;
w23383 <= pi0628 and not w23382;
w23384 <= not pi1156 and not w23383;
w23385 <= not w23379 and w23384;
w23386 <= not pi0629 and not w23198;
w23387 <= not w23385 and w23386;
w23388 <= pi0628 and w23378;
w23389 <= not pi0628 and not w23382;
w23390 <= pi1156 and not w23389;
w23391 <= not w23388 and w23390;
w23392 <= pi0629 and not w23202;
w23393 <= not w23391 and w23392;
w23394 <= not w23387 and not w23393;
w23395 <= pi0792 and not w23394;
w23396 <= not pi0792 and w23378;
w23397 <= not w23395 and not w23396;
w23398 <= not pi0647 and not w23397;
w23399 <= not w15342 and not w23382;
w23400 <= w15342 and w23157;
w23401 <= not w23399 and not w23400;
w23402 <= pi0647 and not w23401;
w23403 <= not pi1157 and not w23402;
w23404 <= not w23398 and w23403;
w23405 <= not pi0630 and not w23210;
w23406 <= not w23404 and w23405;
w23407 <= pi0647 and not w23397;
w23408 <= not pi0647 and not w23401;
w23409 <= pi1157 and not w23408;
w23410 <= not w23407 and w23409;
w23411 <= pi0630 and not w23214;
w23412 <= not w23410 and w23411;
w23413 <= not w23406 and not w23412;
w23414 <= pi0787 and not w23413;
w23415 <= not pi0787 and not w23397;
w23416 <= not w23414 and not w23415;
w23417 <= pi0644 and not w23416;
w23418 <= pi0715 and not w23218;
w23419 <= not w23417 and w23418;
w23420 <= w15367 and not w23157;
w23421 <= not w15367 and w23401;
w23422 <= not w23420 and not w23421;
w23423 <= pi0644 and w23422;
w23424 <= not pi0644 and w23157;
w23425 <= not pi0715 and not w23424;
w23426 <= not w23423 and w23425;
w23427 <= pi1160 and not w23426;
w23428 <= not w23419 and w23427;
w23429 <= not pi0644 and not w23416;
w23430 <= pi0644 and w23217;
w23431 <= not pi0715 and not w23430;
w23432 <= not w23429 and w23431;
w23433 <= not pi0644 and w23422;
w23434 <= pi0644 and w23157;
w23435 <= pi0715 and not w23434;
w23436 <= not w23433 and w23435;
w23437 <= not pi1160 and not w23436;
w23438 <= not w23432 and w23437;
w23439 <= pi0790 and not w23428;
w23440 <= not w23438 and w23439;
w23441 <= not pi0790 and w23416;
w23442 <= w4989 and not w23441;
w23443 <= not w23440 and w23442;
w23444 <= not pi0179 and not w4989;
w23445 <= not pi0832 and not w23444;
w23446 <= not w23443 and w23445;
w23447 <= not pi0179 and not w489;
w23448 <= not pi0724 and w14208;
w23449 <= not w23447 and not w23448;
w23450 <= not pi0778 and w23449;
w23451 <= not pi0625 and w23448;
w23452 <= not w23449 and not w23451;
w23453 <= pi1153 and not w23452;
w23454 <= not pi1153 and not w23447;
w23455 <= not w23451 and w23454;
w23456 <= not w23453 and not w23455;
w23457 <= pi0778 and not w23456;
w23458 <= not w23450 and not w23457;
w23459 <= not w15408 and w23458;
w23460 <= not w15410 and w23459;
w23461 <= not w15412 and w23460;
w23462 <= not w15414 and w23461;
w23463 <= not w15420 and w23462;
w23464 <= not pi0647 and w23463;
w23465 <= pi0647 and w23447;
w23466 <= not pi1157 and not w23465;
w23467 <= not w23464 and w23466;
w23468 <= pi0630 and w23467;
w23469 <= not pi0741 and w14807;
w23470 <= not w23447 and not w23469;
w23471 <= not w15437 and not w23470;
w23472 <= not pi0785 and not w23471;
w23473 <= not w15442 and not w23470;
w23474 <= pi1155 and not w23473;
w23475 <= not w15445 and w23471;
w23476 <= not pi1155 and not w23475;
w23477 <= not w23474 and not w23476;
w23478 <= pi0785 and not w23477;
w23479 <= not w23472 and not w23478;
w23480 <= not pi0781 and not w23479;
w23481 <= not w15452 and w23479;
w23482 <= pi1154 and not w23481;
w23483 <= not w15455 and w23479;
w23484 <= not pi1154 and not w23483;
w23485 <= not w23482 and not w23484;
w23486 <= pi0781 and not w23485;
w23487 <= not w23480 and not w23486;
w23488 <= not pi0789 and not w23487;
w23489 <= not pi0619 and w23447;
w23490 <= pi0619 and w23487;
w23491 <= pi1159 and not w23489;
w23492 <= not w23490 and w23491;
w23493 <= not pi0619 and w23487;
w23494 <= pi0619 and w23447;
w23495 <= not pi1159 and not w23494;
w23496 <= not w23493 and w23495;
w23497 <= not w23492 and not w23496;
w23498 <= pi0789 and not w23497;
w23499 <= not w23488 and not w23498;
w23500 <= not w15532 and w23499;
w23501 <= w15532 and w23447;
w23502 <= not w23500 and not w23501;
w23503 <= not w15342 and not w23502;
w23504 <= w15342 and w23447;
w23505 <= not w23503 and not w23504;
w23506 <= not w18122 and w23505;
w23507 <= pi0647 and not w23463;
w23508 <= not pi0647 and not w23447;
w23509 <= not w23507 and not w23508;
w23510 <= w15364 and not w23509;
w23511 <= not w23468 and not w23510;
w23512 <= not w23506 and w23511;
w23513 <= pi0787 and not w23512;
w23514 <= w15434 and w23461;
w23515 <= not pi0626 and not w23499;
w23516 <= pi0626 and not w23447;
w23517 <= w14192 and not w23516;
w23518 <= not w23515 and w23517;
w23519 <= pi0626 and not w23499;
w23520 <= not pi0626 and not w23447;
w23521 <= w14191 and not w23520;
w23522 <= not w23519 and w23521;
w23523 <= not w23514 and not w23518;
w23524 <= not w23522 and w23523;
w23525 <= pi0788 and not w23524;
w23526 <= pi0618 and w23459;
w23527 <= pi0609 and w23458;
w23528 <= not w14731 and not w23449;
w23529 <= pi0625 and w23528;
w23530 <= w23470 and not w23528;
w23531 <= not w23529 and not w23530;
w23532 <= w23454 and not w23531;
w23533 <= not pi0608 and not w23453;
w23534 <= not w23532 and w23533;
w23535 <= pi1153 and w23470;
w23536 <= not w23529 and w23535;
w23537 <= pi0608 and not w23455;
w23538 <= not w23536 and w23537;
w23539 <= not w23534 and not w23538;
w23540 <= pi0778 and not w23539;
w23541 <= not pi0778 and not w23530;
w23542 <= not w23540 and not w23541;
w23543 <= not pi0609 and not w23542;
w23544 <= not pi1155 and not w23527;
w23545 <= not w23543 and w23544;
w23546 <= not pi0660 and not w23474;
w23547 <= not w23545 and w23546;
w23548 <= not pi0609 and w23458;
w23549 <= pi0609 and not w23542;
w23550 <= pi1155 and not w23548;
w23551 <= not w23549 and w23550;
w23552 <= pi0660 and not w23476;
w23553 <= not w23551 and w23552;
w23554 <= not w23547 and not w23553;
w23555 <= pi0785 and not w23554;
w23556 <= not pi0785 and not w23542;
w23557 <= not w23555 and not w23556;
w23558 <= not pi0618 and not w23557;
w23559 <= not pi1154 and not w23526;
w23560 <= not w23558 and w23559;
w23561 <= not pi0627 and not w23482;
w23562 <= not w23560 and w23561;
w23563 <= not pi0618 and w23459;
w23564 <= pi0618 and not w23557;
w23565 <= pi1154 and not w23563;
w23566 <= not w23564 and w23565;
w23567 <= pi0627 and not w23484;
w23568 <= not w23566 and w23567;
w23569 <= not w23562 and not w23568;
w23570 <= pi0781 and not w23569;
w23571 <= not pi0781 and not w23557;
w23572 <= not w23570 and not w23571;
w23573 <= not pi0789 and w23572;
w23574 <= not pi0619 and not w23572;
w23575 <= pi0619 and w23460;
w23576 <= not pi1159 and not w23575;
w23577 <= not w23574 and w23576;
w23578 <= not pi0648 and not w23492;
w23579 <= not w23577 and w23578;
w23580 <= pi0619 and not w23572;
w23581 <= not pi0619 and w23460;
w23582 <= pi1159 and not w23581;
w23583 <= not w23580 and w23582;
w23584 <= pi0648 and not w23496;
w23585 <= not w23583 and w23584;
w23586 <= pi0789 and not w23579;
w23587 <= not w23585 and w23586;
w23588 <= w15533 and not w23573;
w23589 <= not w23587 and w23588;
w23590 <= not w23525 and not w23589;
w23591 <= not w17927 and not w23590;
w23592 <= w15417 and not w23502;
w23593 <= w18414 and w23462;
w23594 <= not w23592 and not w23593;
w23595 <= not pi0629 and not w23594;
w23596 <= w18418 and w23462;
w23597 <= w15416 and not w23502;
w23598 <= not w23596 and not w23597;
w23599 <= pi0629 and not w23598;
w23600 <= not w23595 and not w23599;
w23601 <= pi0792 and not w23600;
w23602 <= not w17769 and not w23601;
w23603 <= not w23591 and w23602;
w23604 <= not w23513 and not w23603;
w23605 <= not pi0790 and w23604;
w23606 <= not pi0787 and not w23463;
w23607 <= pi1157 and not w23509;
w23608 <= not w23467 and not w23607;
w23609 <= pi0787 and not w23608;
w23610 <= not w23606 and not w23609;
w23611 <= not pi0644 and w23610;
w23612 <= pi0644 and w23604;
w23613 <= pi0715 and not w23611;
w23614 <= not w23612 and w23613;
w23615 <= not w15367 and not w23505;
w23616 <= w15367 and w23447;
w23617 <= not w23615 and not w23616;
w23618 <= pi0644 and not w23617;
w23619 <= not pi0644 and w23447;
w23620 <= not pi0715 and not w23619;
w23621 <= not w23618 and w23620;
w23622 <= pi1160 and not w23621;
w23623 <= not w23614 and w23622;
w23624 <= not pi0644 and not w23617;
w23625 <= pi0644 and w23447;
w23626 <= pi0715 and not w23625;
w23627 <= not w23624 and w23626;
w23628 <= pi0644 and w23610;
w23629 <= not pi0644 and w23604;
w23630 <= not pi0715 and not w23628;
w23631 <= not w23629 and w23630;
w23632 <= not pi1160 and not w23627;
w23633 <= not w23631 and w23632;
w23634 <= not w23623 and not w23633;
w23635 <= pi0790 and not w23634;
w23636 <= pi0832 and not w23605;
w23637 <= not w23635 and w23636;
w23638 <= not w23446 and not w23637;
w23639 <= not pi0180 and not w489;
w23640 <= not pi0702 and w14208;
w23641 <= not w23639 and not w23640;
w23642 <= not pi0778 and not w23641;
w23643 <= not pi0625 and w23640;
w23644 <= not w23641 and not w23643;
w23645 <= pi1153 and not w23644;
w23646 <= not pi1153 and not w23639;
w23647 <= not w23643 and w23646;
w23648 <= pi0778 and not w23647;
w23649 <= not w23645 and w23648;
w23650 <= not w23642 and not w23649;
w23651 <= not w15408 and not w23650;
w23652 <= not w15410 and w23651;
w23653 <= not w15412 and w23652;
w23654 <= not w15414 and w23653;
w23655 <= not w15420 and w23654;
w23656 <= not pi0647 and w23655;
w23657 <= pi0647 and w23639;
w23658 <= not pi1157 and not w23657;
w23659 <= not w23656 and w23658;
w23660 <= pi0630 and w23659;
w23661 <= not pi0753 and w14807;
w23662 <= not w23639 and not w23661;
w23663 <= not w15437 and not w23662;
w23664 <= not pi0785 and not w23663;
w23665 <= w14859 and w23661;
w23666 <= w23663 and not w23665;
w23667 <= pi1155 and not w23666;
w23668 <= not pi1155 and not w23639;
w23669 <= not w23665 and w23668;
w23670 <= not w23667 and not w23669;
w23671 <= pi0785 and not w23670;
w23672 <= not w23664 and not w23671;
w23673 <= not pi0781 and not w23672;
w23674 <= not w15452 and w23672;
w23675 <= pi1154 and not w23674;
w23676 <= not w15455 and w23672;
w23677 <= not pi1154 and not w23676;
w23678 <= not w23675 and not w23677;
w23679 <= pi0781 and not w23678;
w23680 <= not w23673 and not w23679;
w23681 <= not pi0789 and not w23680;
w23682 <= not w20641 and w23680;
w23683 <= pi1159 and not w23682;
w23684 <= not w20644 and w23680;
w23685 <= not pi1159 and not w23684;
w23686 <= not w23683 and not w23685;
w23687 <= pi0789 and not w23686;
w23688 <= not w23681 and not w23687;
w23689 <= not w15532 and w23688;
w23690 <= w15532 and w23639;
w23691 <= not w23689 and not w23690;
w23692 <= not w15342 and not w23691;
w23693 <= w15342 and w23639;
w23694 <= not w23692 and not w23693;
w23695 <= not w18122 and w23694;
w23696 <= pi0647 and not w23655;
w23697 <= not pi0647 and not w23639;
w23698 <= not w23696 and not w23697;
w23699 <= w15364 and not w23698;
w23700 <= not w23660 and not w23699;
w23701 <= not w23695 and w23700;
w23702 <= pi0787 and not w23701;
w23703 <= w15434 and w23653;
w23704 <= not pi0626 and not w23688;
w23705 <= pi0626 and not w23639;
w23706 <= w14192 and not w23705;
w23707 <= not w23704 and w23706;
w23708 <= pi0626 and not w23688;
w23709 <= not pi0626 and not w23639;
w23710 <= w14191 and not w23709;
w23711 <= not w23708 and w23710;
w23712 <= not w23703 and not w23707;
w23713 <= not w23711 and w23712;
w23714 <= pi0788 and not w23713;
w23715 <= pi0618 and w23651;
w23716 <= not w14731 and not w23641;
w23717 <= pi0625 and w23716;
w23718 <= w23662 and not w23716;
w23719 <= not w23717 and not w23718;
w23720 <= w23646 and not w23719;
w23721 <= not pi0608 and not w23645;
w23722 <= not w23720 and w23721;
w23723 <= pi1153 and w23662;
w23724 <= not w23717 and w23723;
w23725 <= pi0608 and not w23647;
w23726 <= not w23724 and w23725;
w23727 <= not w23722 and not w23726;
w23728 <= pi0778 and not w23727;
w23729 <= not pi0778 and not w23718;
w23730 <= not w23728 and not w23729;
w23731 <= not pi0609 and not w23730;
w23732 <= pi0609 and not w23650;
w23733 <= not pi1155 and not w23732;
w23734 <= not w23731 and w23733;
w23735 <= not pi0660 and not w23667;
w23736 <= not w23734 and w23735;
w23737 <= pi0609 and not w23730;
w23738 <= not pi0609 and not w23650;
w23739 <= pi1155 and not w23738;
w23740 <= not w23737 and w23739;
w23741 <= pi0660 and not w23669;
w23742 <= not w23740 and w23741;
w23743 <= not w23736 and not w23742;
w23744 <= pi0785 and not w23743;
w23745 <= not pi0785 and not w23730;
w23746 <= not w23744 and not w23745;
w23747 <= not pi0618 and not w23746;
w23748 <= not pi1154 and not w23715;
w23749 <= not w23747 and w23748;
w23750 <= not pi0627 and not w23675;
w23751 <= not w23749 and w23750;
w23752 <= not pi0618 and w23651;
w23753 <= pi0618 and not w23746;
w23754 <= pi1154 and not w23752;
w23755 <= not w23753 and w23754;
w23756 <= pi0627 and not w23677;
w23757 <= not w23755 and w23756;
w23758 <= not w23751 and not w23757;
w23759 <= pi0781 and not w23758;
w23760 <= not pi0781 and not w23746;
w23761 <= not w23759 and not w23760;
w23762 <= not pi0789 and w23761;
w23763 <= not pi0619 and not w23761;
w23764 <= pi0619 and w23652;
w23765 <= not pi1159 and not w23764;
w23766 <= not w23763 and w23765;
w23767 <= not pi0648 and not w23683;
w23768 <= not w23766 and w23767;
w23769 <= pi0619 and not w23761;
w23770 <= not pi0619 and w23652;
w23771 <= pi1159 and not w23770;
w23772 <= not w23769 and w23771;
w23773 <= pi0648 and not w23685;
w23774 <= not w23772 and w23773;
w23775 <= pi0789 and not w23768;
w23776 <= not w23774 and w23775;
w23777 <= w15533 and not w23762;
w23778 <= not w23776 and w23777;
w23779 <= not w23714 and not w23778;
w23780 <= not w17927 and not w23779;
w23781 <= w15417 and not w23691;
w23782 <= w18414 and w23654;
w23783 <= not w23781 and not w23782;
w23784 <= not pi0629 and not w23783;
w23785 <= w18418 and w23654;
w23786 <= w15416 and not w23691;
w23787 <= not w23785 and not w23786;
w23788 <= pi0629 and not w23787;
w23789 <= not w23784 and not w23788;
w23790 <= pi0792 and not w23789;
w23791 <= not w17769 and not w23790;
w23792 <= not w23780 and w23791;
w23793 <= not w23702 and not w23792;
w23794 <= not pi0790 and w23793;
w23795 <= not pi0787 and not w23655;
w23796 <= pi1157 and not w23698;
w23797 <= not w23659 and not w23796;
w23798 <= pi0787 and not w23797;
w23799 <= not w23795 and not w23798;
w23800 <= not pi0644 and w23799;
w23801 <= pi0644 and w23793;
w23802 <= pi0715 and not w23800;
w23803 <= not w23801 and w23802;
w23804 <= not w15367 and not w23694;
w23805 <= w15367 and w23639;
w23806 <= not w23804 and not w23805;
w23807 <= pi0644 and not w23806;
w23808 <= not pi0644 and w23639;
w23809 <= not pi0715 and not w23808;
w23810 <= not w23807 and w23809;
w23811 <= pi1160 and not w23810;
w23812 <= not w23803 and w23811;
w23813 <= not pi0644 and not w23806;
w23814 <= pi0644 and w23639;
w23815 <= pi0715 and not w23814;
w23816 <= not w23813 and w23815;
w23817 <= pi0644 and w23799;
w23818 <= not pi0644 and w23793;
w23819 <= not pi0715 and not w23817;
w23820 <= not w23818 and w23819;
w23821 <= not pi1160 and not w23816;
w23822 <= not w23820 and w23821;
w23823 <= not w23812 and not w23822;
w23824 <= pi0790 and not w23823;
w23825 <= pi0832 and not w23794;
w23826 <= not w23824 and w23825;
w23827 <= not pi0180 and not w4989;
w23828 <= not pi0180 and not w14622;
w23829 <= w14198 and not w23828;
w23830 <= not pi0702 and w134;
w23831 <= w23828 and not w23830;
w23832 <= not pi0180 and not w14204;
w23833 <= w14210 and not w23832;
w23834 <= pi0180 and not w15639;
w23835 <= not pi0038 and not w23834;
w23836 <= w134 and not w23835;
w23837 <= not pi0180 and w15635;
w23838 <= not w23836 and not w23837;
w23839 <= not pi0702 and not w23833;
w23840 <= not w23838 and w23839;
w23841 <= not w23831 and not w23840;
w23842 <= not pi0778 and w23841;
w23843 <= not pi0625 and w23828;
w23844 <= pi0625 and not w23841;
w23845 <= pi1153 and not w23843;
w23846 <= not w23844 and w23845;
w23847 <= pi0625 and w23828;
w23848 <= not pi0625 and not w23841;
w23849 <= not pi1153 and not w23847;
w23850 <= not w23848 and w23849;
w23851 <= not w23846 and not w23850;
w23852 <= pi0778 and not w23851;
w23853 <= not w23842 and not w23852;
w23854 <= not w14638 and not w23853;
w23855 <= w14638 and not w23828;
w23856 <= not w23854 and not w23855;
w23857 <= not w14202 and w23856;
w23858 <= w14202 and w23828;
w23859 <= not w23857 and not w23858;
w23860 <= not w14198 and w23859;
w23861 <= not w23829 and not w23860;
w23862 <= not w14194 and w23861;
w23863 <= w14194 and w23828;
w23864 <= not w23862 and not w23863;
w23865 <= not pi0792 and w23864;
w23866 <= pi0628 and not w23864;
w23867 <= not pi0628 and w23828;
w23868 <= pi1156 and not w23867;
w23869 <= not w23866 and w23868;
w23870 <= pi0628 and w23828;
w23871 <= not pi0628 and not w23864;
w23872 <= not pi1156 and not w23870;
w23873 <= not w23871 and w23872;
w23874 <= not w23869 and not w23873;
w23875 <= pi0792 and not w23874;
w23876 <= not w23865 and not w23875;
w23877 <= not pi0647 and not w23876;
w23878 <= pi0647 and not w23828;
w23879 <= not w23877 and not w23878;
w23880 <= not pi1157 and w23879;
w23881 <= pi0647 and not w23876;
w23882 <= not pi0647 and not w23828;
w23883 <= not w23881 and not w23882;
w23884 <= pi1157 and w23883;
w23885 <= not w23880 and not w23884;
w23886 <= pi0787 and not w23885;
w23887 <= not pi0787 and w23876;
w23888 <= not w23886 and not w23887;
w23889 <= not pi0644 and not w23888;
w23890 <= pi0715 and not w23889;
w23891 <= pi0180 and not w134;
w23892 <= pi0180 and pi0753;
w23893 <= pi0753 and w14609;
w23894 <= pi0180 and w14836;
w23895 <= not w23893 and not w23894;
w23896 <= pi0039 and not w23895;
w23897 <= pi0180 and not w14796;
w23898 <= not w19319 and not w23897;
w23899 <= not pi0039 and not w23898;
w23900 <= not pi0180 and not pi0753;
w23901 <= w14784 and w23900;
w23902 <= not w23892 and not w23899;
w23903 <= not w23901 and w23902;
w23904 <= not w23896 and w23903;
w23905 <= not pi0038 and not w23904;
w23906 <= not pi0753 and w14843;
w23907 <= pi0038 and not w23832;
w23908 <= not w23906 and w23907;
w23909 <= not w23905 and not w23908;
w23910 <= w134 and not w23909;
w23911 <= not w23891 and not w23910;
w23912 <= not w14680 and not w23911;
w23913 <= w14680 and not w23828;
w23914 <= not w23912 and not w23913;
w23915 <= not pi0785 and not w23914;
w23916 <= not w14854 and not w23828;
w23917 <= pi0609 and w23912;
w23918 <= not w23916 and not w23917;
w23919 <= pi1155 and not w23918;
w23920 <= not w14859 and not w23828;
w23921 <= not pi0609 and w23912;
w23922 <= not w23920 and not w23921;
w23923 <= not pi1155 and not w23922;
w23924 <= not w23919 and not w23923;
w23925 <= pi0785 and not w23924;
w23926 <= not w23915 and not w23925;
w23927 <= not pi0781 and not w23926;
w23928 <= not pi0618 and w23828;
w23929 <= pi0618 and w23926;
w23930 <= pi1154 and not w23928;
w23931 <= not w23929 and w23930;
w23932 <= not pi0618 and w23926;
w23933 <= pi0618 and w23828;
w23934 <= not pi1154 and not w23933;
w23935 <= not w23932 and w23934;
w23936 <= not w23931 and not w23935;
w23937 <= pi0781 and not w23936;
w23938 <= not w23927 and not w23937;
w23939 <= not pi0789 and not w23938;
w23940 <= not pi0619 and w23828;
w23941 <= pi0619 and w23938;
w23942 <= pi1159 and not w23940;
w23943 <= not w23941 and w23942;
w23944 <= not pi0619 and w23938;
w23945 <= pi0619 and w23828;
w23946 <= not pi1159 and not w23945;
w23947 <= not w23944 and w23946;
w23948 <= not w23943 and not w23947;
w23949 <= pi0789 and not w23948;
w23950 <= not w23939 and not w23949;
w23951 <= not w15532 and w23950;
w23952 <= w15532 and w23828;
w23953 <= not w23951 and not w23952;
w23954 <= not w15342 and not w23953;
w23955 <= w15342 and w23828;
w23956 <= not w23954 and not w23955;
w23957 <= not w15367 and not w23956;
w23958 <= w15367 and w23828;
w23959 <= not w23957 and not w23958;
w23960 <= pi0644 and not w23959;
w23961 <= not pi0644 and w23828;
w23962 <= not pi0715 and not w23961;
w23963 <= not w23960 and w23962;
w23964 <= pi1160 and not w23963;
w23965 <= not w23890 and w23964;
w23966 <= pi0644 and not w23888;
w23967 <= not pi0715 and not w23966;
w23968 <= not pi0644 and not w23959;
w23969 <= pi0644 and w23828;
w23970 <= pi0715 and not w23969;
w23971 <= not w23968 and w23970;
w23972 <= not pi1160 and not w23971;
w23973 <= not w23967 and w23972;
w23974 <= not w23965 and not w23973;
w23975 <= pi0790 and not w23974;
w23976 <= not pi0629 and w23869;
w23977 <= not w18133 and w23953;
w23978 <= pi0629 and w23873;
w23979 <= not w23976 and not w23978;
w23980 <= not w23977 and w23979;
w23981 <= pi0792 and not w23980;
w23982 <= pi0609 and w23853;
w23983 <= pi0180 and not w15188;
w23984 <= not pi0180 and not w15175;
w23985 <= pi0753 and not w23983;
w23986 <= not w23984 and w23985;
w23987 <= not pi0180 and w15192;
w23988 <= pi0180 and w15194;
w23989 <= not pi0753 and not w23988;
w23990 <= not w23987 and w23989;
w23991 <= not w23986 and not w23990;
w23992 <= not pi0039 and not w23991;
w23993 <= pi0180 and w15168;
w23994 <= not pi0180 and not w15109;
w23995 <= not pi0753 and not w23994;
w23996 <= not w23993 and w23995;
w23997 <= not pi0180 and w14967;
w23998 <= pi0180 and w15048;
w23999 <= pi0753 and not w23998;
w24000 <= not w23997 and w23999;
w24001 <= pi0039 and not w23996;
w24002 <= not w24000 and w24001;
w24003 <= not pi0038 and not w23992;
w24004 <= not w24002 and w24003;
w24005 <= not w15032 and not w23661;
w24006 <= pi0180 and not w24005;
w24007 <= w3847 and w24006;
w24008 <= not pi0753 and not w15053;
w24009 <= w17034 and not w24008;
w24010 <= not pi0180 and not w24009;
w24011 <= pi0038 and not w24007;
w24012 <= not w24010 and w24011;
w24013 <= not pi0702 and not w24012;
w24014 <= not w24004 and w24013;
w24015 <= pi0702 and w23909;
w24016 <= w134 and not w24014;
w24017 <= not w24015 and w24016;
w24018 <= not w23891 and not w24017;
w24019 <= not pi0625 and w24018;
w24020 <= pi0625 and w23911;
w24021 <= not pi1153 and not w24020;
w24022 <= not w24019 and w24021;
w24023 <= not pi0608 and not w23846;
w24024 <= not w24022 and w24023;
w24025 <= not pi0625 and w23911;
w24026 <= pi0625 and w24018;
w24027 <= pi1153 and not w24025;
w24028 <= not w24026 and w24027;
w24029 <= pi0608 and not w23850;
w24030 <= not w24028 and w24029;
w24031 <= not w24024 and not w24030;
w24032 <= pi0778 and not w24031;
w24033 <= not pi0778 and w24018;
w24034 <= not w24032 and not w24033;
w24035 <= not pi0609 and not w24034;
w24036 <= not pi1155 and not w23982;
w24037 <= not w24035 and w24036;
w24038 <= not pi0660 and not w23919;
w24039 <= not w24037 and w24038;
w24040 <= not pi0609 and w23853;
w24041 <= pi0609 and not w24034;
w24042 <= pi1155 and not w24040;
w24043 <= not w24041 and w24042;
w24044 <= pi0660 and not w23923;
w24045 <= not w24043 and w24044;
w24046 <= not w24039 and not w24045;
w24047 <= pi0785 and not w24046;
w24048 <= not pi0785 and not w24034;
w24049 <= not w24047 and not w24048;
w24050 <= not pi0618 and not w24049;
w24051 <= pi0618 and w23856;
w24052 <= not pi1154 and not w24051;
w24053 <= not w24050 and w24052;
w24054 <= not pi0627 and not w23931;
w24055 <= not w24053 and w24054;
w24056 <= not pi0618 and w23856;
w24057 <= pi0618 and not w24049;
w24058 <= pi1154 and not w24056;
w24059 <= not w24057 and w24058;
w24060 <= pi0627 and not w23935;
w24061 <= not w24059 and w24060;
w24062 <= not w24055 and not w24061;
w24063 <= pi0781 and not w24062;
w24064 <= not pi0781 and not w24049;
w24065 <= not w24063 and not w24064;
w24066 <= not pi0789 and w24065;
w24067 <= pi0619 and not w23859;
w24068 <= not pi0619 and not w24065;
w24069 <= not pi1159 and not w24067;
w24070 <= not w24068 and w24069;
w24071 <= not pi0648 and not w23943;
w24072 <= not w24070 and w24071;
w24073 <= not pi0619 and not w23859;
w24074 <= pi0619 and not w24065;
w24075 <= pi1159 and not w24073;
w24076 <= not w24074 and w24075;
w24077 <= pi0648 and not w23947;
w24078 <= not w24076 and w24077;
w24079 <= pi0789 and not w24072;
w24080 <= not w24078 and w24079;
w24081 <= w15533 and not w24066;
w24082 <= not w24080 and w24081;
w24083 <= w15434 and w23861;
w24084 <= not pi0626 and not w23950;
w24085 <= pi0626 and not w23828;
w24086 <= w14192 and not w24085;
w24087 <= not w24084 and w24086;
w24088 <= pi0626 and not w23950;
w24089 <= not pi0626 and not w23828;
w24090 <= w14191 and not w24089;
w24091 <= not w24088 and w24090;
w24092 <= not w24083 and not w24087;
w24093 <= not w24091 and w24092;
w24094 <= pi0788 and not w24093;
w24095 <= not w17927 and not w24094;
w24096 <= not w24082 and w24095;
w24097 <= not w23981 and not w24096;
w24098 <= not w17769 and not w24097;
w24099 <= w15365 and not w23879;
w24100 <= not w18122 and w23956;
w24101 <= w15364 and not w23883;
w24102 <= not w24099 and not w24101;
w24103 <= not w24100 and w24102;
w24104 <= pi0787 and not w24103;
w24105 <= not pi0644 and w23972;
w24106 <= pi0644 and w23964;
w24107 <= pi0790 and not w24105;
w24108 <= not w24106 and w24107;
w24109 <= not w24098 and not w24104;
w24110 <= not w24108 and w24109;
w24111 <= not w23975 and not w24110;
w24112 <= w4989 and not w24111;
w24113 <= not pi0832 and not w23827;
w24114 <= not w24112 and w24113;
w24115 <= not w23826 and not w24114;
w24116 <= not pi0181 and not w489;
w24117 <= not pi0709 and w14208;
w24118 <= not w24116 and not w24117;
w24119 <= not pi0778 and not w24118;
w24120 <= not pi0625 and w24117;
w24121 <= not w24118 and not w24120;
w24122 <= pi1153 and not w24121;
w24123 <= not pi1153 and not w24116;
w24124 <= not w24120 and w24123;
w24125 <= pi0778 and not w24124;
w24126 <= not w24122 and w24125;
w24127 <= not w24119 and not w24126;
w24128 <= not w15408 and not w24127;
w24129 <= not w15410 and w24128;
w24130 <= not w15412 and w24129;
w24131 <= not w15414 and w24130;
w24132 <= not w15420 and w24131;
w24133 <= not pi0647 and w24132;
w24134 <= pi0647 and w24116;
w24135 <= not pi1157 and not w24134;
w24136 <= not w24133 and w24135;
w24137 <= pi0630 and w24136;
w24138 <= not pi0754 and w14807;
w24139 <= not w24116 and not w24138;
w24140 <= not w15437 and not w24139;
w24141 <= not pi0785 and not w24140;
w24142 <= w14859 and w24138;
w24143 <= w24140 and not w24142;
w24144 <= pi1155 and not w24143;
w24145 <= not pi1155 and not w24116;
w24146 <= not w24142 and w24145;
w24147 <= not w24144 and not w24146;
w24148 <= pi0785 and not w24147;
w24149 <= not w24141 and not w24148;
w24150 <= not pi0781 and not w24149;
w24151 <= not w15452 and w24149;
w24152 <= pi1154 and not w24151;
w24153 <= not w15455 and w24149;
w24154 <= not pi1154 and not w24153;
w24155 <= not w24152 and not w24154;
w24156 <= pi0781 and not w24155;
w24157 <= not w24150 and not w24156;
w24158 <= not pi0789 and not w24157;
w24159 <= not w20641 and w24157;
w24160 <= pi1159 and not w24159;
w24161 <= not w20644 and w24157;
w24162 <= not pi1159 and not w24161;
w24163 <= not w24160 and not w24162;
w24164 <= pi0789 and not w24163;
w24165 <= not w24158 and not w24164;
w24166 <= not w15532 and w24165;
w24167 <= w15532 and w24116;
w24168 <= not w24166 and not w24167;
w24169 <= not w15342 and not w24168;
w24170 <= w15342 and w24116;
w24171 <= not w24169 and not w24170;
w24172 <= not w18122 and w24171;
w24173 <= pi0647 and not w24132;
w24174 <= not pi0647 and not w24116;
w24175 <= not w24173 and not w24174;
w24176 <= w15364 and not w24175;
w24177 <= not w24137 and not w24176;
w24178 <= not w24172 and w24177;
w24179 <= pi0787 and not w24178;
w24180 <= w15434 and w24130;
w24181 <= not pi0626 and not w24165;
w24182 <= pi0626 and not w24116;
w24183 <= w14192 and not w24182;
w24184 <= not w24181 and w24183;
w24185 <= pi0626 and not w24165;
w24186 <= not pi0626 and not w24116;
w24187 <= w14191 and not w24186;
w24188 <= not w24185 and w24187;
w24189 <= not w24180 and not w24184;
w24190 <= not w24188 and w24189;
w24191 <= pi0788 and not w24190;
w24192 <= pi0618 and w24128;
w24193 <= not w14731 and not w24118;
w24194 <= pi0625 and w24193;
w24195 <= w24139 and not w24193;
w24196 <= not w24194 and not w24195;
w24197 <= w24123 and not w24196;
w24198 <= not pi0608 and not w24122;
w24199 <= not w24197 and w24198;
w24200 <= pi1153 and w24139;
w24201 <= not w24194 and w24200;
w24202 <= pi0608 and not w24124;
w24203 <= not w24201 and w24202;
w24204 <= not w24199 and not w24203;
w24205 <= pi0778 and not w24204;
w24206 <= not pi0778 and not w24195;
w24207 <= not w24205 and not w24206;
w24208 <= not pi0609 and not w24207;
w24209 <= pi0609 and not w24127;
w24210 <= not pi1155 and not w24209;
w24211 <= not w24208 and w24210;
w24212 <= not pi0660 and not w24144;
w24213 <= not w24211 and w24212;
w24214 <= pi0609 and not w24207;
w24215 <= not pi0609 and not w24127;
w24216 <= pi1155 and not w24215;
w24217 <= not w24214 and w24216;
w24218 <= pi0660 and not w24146;
w24219 <= not w24217 and w24218;
w24220 <= not w24213 and not w24219;
w24221 <= pi0785 and not w24220;
w24222 <= not pi0785 and not w24207;
w24223 <= not w24221 and not w24222;
w24224 <= not pi0618 and not w24223;
w24225 <= not pi1154 and not w24192;
w24226 <= not w24224 and w24225;
w24227 <= not pi0627 and not w24152;
w24228 <= not w24226 and w24227;
w24229 <= not pi0618 and w24128;
w24230 <= pi0618 and not w24223;
w24231 <= pi1154 and not w24229;
w24232 <= not w24230 and w24231;
w24233 <= pi0627 and not w24154;
w24234 <= not w24232 and w24233;
w24235 <= not w24228 and not w24234;
w24236 <= pi0781 and not w24235;
w24237 <= not pi0781 and not w24223;
w24238 <= not w24236 and not w24237;
w24239 <= not pi0789 and w24238;
w24240 <= not pi0619 and not w24238;
w24241 <= pi0619 and w24129;
w24242 <= not pi1159 and not w24241;
w24243 <= not w24240 and w24242;
w24244 <= not pi0648 and not w24160;
w24245 <= not w24243 and w24244;
w24246 <= pi0619 and not w24238;
w24247 <= not pi0619 and w24129;
w24248 <= pi1159 and not w24247;
w24249 <= not w24246 and w24248;
w24250 <= pi0648 and not w24162;
w24251 <= not w24249 and w24250;
w24252 <= pi0789 and not w24245;
w24253 <= not w24251 and w24252;
w24254 <= w15533 and not w24239;
w24255 <= not w24253 and w24254;
w24256 <= not w24191 and not w24255;
w24257 <= not w17927 and not w24256;
w24258 <= w15417 and not w24168;
w24259 <= w18414 and w24131;
w24260 <= not w24258 and not w24259;
w24261 <= not pi0629 and not w24260;
w24262 <= w18418 and w24131;
w24263 <= w15416 and not w24168;
w24264 <= not w24262 and not w24263;
w24265 <= pi0629 and not w24264;
w24266 <= not w24261 and not w24265;
w24267 <= pi0792 and not w24266;
w24268 <= not w17769 and not w24267;
w24269 <= not w24257 and w24268;
w24270 <= not w24179 and not w24269;
w24271 <= not pi0790 and w24270;
w24272 <= not pi0787 and not w24132;
w24273 <= pi1157 and not w24175;
w24274 <= not w24136 and not w24273;
w24275 <= pi0787 and not w24274;
w24276 <= not w24272 and not w24275;
w24277 <= not pi0644 and w24276;
w24278 <= pi0644 and w24270;
w24279 <= pi0715 and not w24277;
w24280 <= not w24278 and w24279;
w24281 <= not w15367 and not w24171;
w24282 <= w15367 and w24116;
w24283 <= not w24281 and not w24282;
w24284 <= pi0644 and not w24283;
w24285 <= not pi0644 and w24116;
w24286 <= not pi0715 and not w24285;
w24287 <= not w24284 and w24286;
w24288 <= pi1160 and not w24287;
w24289 <= not w24280 and w24288;
w24290 <= not pi0644 and not w24283;
w24291 <= pi0644 and w24116;
w24292 <= pi0715 and not w24291;
w24293 <= not w24290 and w24292;
w24294 <= pi0644 and w24276;
w24295 <= not pi0644 and w24270;
w24296 <= not pi0715 and not w24294;
w24297 <= not w24295 and w24296;
w24298 <= not pi1160 and not w24293;
w24299 <= not w24297 and w24298;
w24300 <= not w24289 and not w24299;
w24301 <= pi0790 and not w24300;
w24302 <= pi0832 and not w24271;
w24303 <= not w24301 and w24302;
w24304 <= not pi0181 and not w4989;
w24305 <= not pi0181 and not w14622;
w24306 <= w14198 and not w24305;
w24307 <= not pi0709 and w134;
w24308 <= w24305 and not w24307;
w24309 <= not pi0181 and not w14204;
w24310 <= w14210 and not w24309;
w24311 <= pi0181 and not w15639;
w24312 <= not pi0038 and not w24311;
w24313 <= w134 and not w24312;
w24314 <= not pi0181 and w15635;
w24315 <= not w24313 and not w24314;
w24316 <= not pi0709 and not w24310;
w24317 <= not w24315 and w24316;
w24318 <= not w24308 and not w24317;
w24319 <= not pi0778 and w24318;
w24320 <= not pi0625 and w24305;
w24321 <= pi0625 and not w24318;
w24322 <= pi1153 and not w24320;
w24323 <= not w24321 and w24322;
w24324 <= pi0625 and w24305;
w24325 <= not pi0625 and not w24318;
w24326 <= not pi1153 and not w24324;
w24327 <= not w24325 and w24326;
w24328 <= not w24323 and not w24327;
w24329 <= pi0778 and not w24328;
w24330 <= not w24319 and not w24329;
w24331 <= not w14638 and not w24330;
w24332 <= w14638 and not w24305;
w24333 <= not w24331 and not w24332;
w24334 <= not w14202 and w24333;
w24335 <= w14202 and w24305;
w24336 <= not w24334 and not w24335;
w24337 <= not w14198 and w24336;
w24338 <= not w24306 and not w24337;
w24339 <= not w14194 and w24338;
w24340 <= w14194 and w24305;
w24341 <= not w24339 and not w24340;
w24342 <= not pi0792 and w24341;
w24343 <= pi0628 and not w24341;
w24344 <= not pi0628 and w24305;
w24345 <= pi1156 and not w24344;
w24346 <= not w24343 and w24345;
w24347 <= pi0628 and w24305;
w24348 <= not pi0628 and not w24341;
w24349 <= not pi1156 and not w24347;
w24350 <= not w24348 and w24349;
w24351 <= not w24346 and not w24350;
w24352 <= pi0792 and not w24351;
w24353 <= not w24342 and not w24352;
w24354 <= not pi0647 and not w24353;
w24355 <= pi0647 and not w24305;
w24356 <= not w24354 and not w24355;
w24357 <= not pi1157 and w24356;
w24358 <= pi0647 and not w24353;
w24359 <= not pi0647 and not w24305;
w24360 <= not w24358 and not w24359;
w24361 <= pi1157 and w24360;
w24362 <= not w24357 and not w24361;
w24363 <= pi0787 and not w24362;
w24364 <= not pi0787 and w24353;
w24365 <= not w24363 and not w24364;
w24366 <= not pi0644 and not w24365;
w24367 <= pi0715 and not w24366;
w24368 <= pi0181 and not w134;
w24369 <= pi0181 and pi0754;
w24370 <= pi0754 and w14609;
w24371 <= pi0181 and w14836;
w24372 <= not w24370 and not w24371;
w24373 <= pi0039 and not w24372;
w24374 <= pi0181 and not w14796;
w24375 <= not w19375 and not w24374;
w24376 <= not pi0039 and not w24375;
w24377 <= not pi0181 and not pi0754;
w24378 <= w14784 and w24377;
w24379 <= not w24369 and not w24376;
w24380 <= not w24378 and w24379;
w24381 <= not w24373 and w24380;
w24382 <= not pi0038 and not w24381;
w24383 <= not pi0754 and w14843;
w24384 <= pi0038 and not w24309;
w24385 <= not w24383 and w24384;
w24386 <= not w24382 and not w24385;
w24387 <= w134 and not w24386;
w24388 <= not w24368 and not w24387;
w24389 <= not w14680 and not w24388;
w24390 <= w14680 and not w24305;
w24391 <= not w24389 and not w24390;
w24392 <= not pi0785 and not w24391;
w24393 <= not w14854 and not w24305;
w24394 <= pi0609 and w24389;
w24395 <= not w24393 and not w24394;
w24396 <= pi1155 and not w24395;
w24397 <= not w14859 and not w24305;
w24398 <= not pi0609 and w24389;
w24399 <= not w24397 and not w24398;
w24400 <= not pi1155 and not w24399;
w24401 <= not w24396 and not w24400;
w24402 <= pi0785 and not w24401;
w24403 <= not w24392 and not w24402;
w24404 <= not pi0781 and not w24403;
w24405 <= not pi0618 and w24305;
w24406 <= pi0618 and w24403;
w24407 <= pi1154 and not w24405;
w24408 <= not w24406 and w24407;
w24409 <= not pi0618 and w24403;
w24410 <= pi0618 and w24305;
w24411 <= not pi1154 and not w24410;
w24412 <= not w24409 and w24411;
w24413 <= not w24408 and not w24412;
w24414 <= pi0781 and not w24413;
w24415 <= not w24404 and not w24414;
w24416 <= not pi0789 and not w24415;
w24417 <= not pi0619 and w24305;
w24418 <= pi0619 and w24415;
w24419 <= pi1159 and not w24417;
w24420 <= not w24418 and w24419;
w24421 <= not pi0619 and w24415;
w24422 <= pi0619 and w24305;
w24423 <= not pi1159 and not w24422;
w24424 <= not w24421 and w24423;
w24425 <= not w24420 and not w24424;
w24426 <= pi0789 and not w24425;
w24427 <= not w24416 and not w24426;
w24428 <= not w15532 and w24427;
w24429 <= w15532 and w24305;
w24430 <= not w24428 and not w24429;
w24431 <= not w15342 and not w24430;
w24432 <= w15342 and w24305;
w24433 <= not w24431 and not w24432;
w24434 <= not w15367 and not w24433;
w24435 <= w15367 and w24305;
w24436 <= not w24434 and not w24435;
w24437 <= pi0644 and not w24436;
w24438 <= not pi0644 and w24305;
w24439 <= not pi0715 and not w24438;
w24440 <= not w24437 and w24439;
w24441 <= pi1160 and not w24440;
w24442 <= not w24367 and w24441;
w24443 <= pi0644 and not w24365;
w24444 <= not pi0715 and not w24443;
w24445 <= not pi0644 and not w24436;
w24446 <= pi0644 and w24305;
w24447 <= pi0715 and not w24446;
w24448 <= not w24445 and w24447;
w24449 <= not pi1160 and not w24448;
w24450 <= not w24444 and w24449;
w24451 <= not w24442 and not w24450;
w24452 <= pi0790 and not w24451;
w24453 <= not pi0629 and w24346;
w24454 <= not w18133 and w24430;
w24455 <= pi0629 and w24350;
w24456 <= not w24453 and not w24455;
w24457 <= not w24454 and w24456;
w24458 <= pi0792 and not w24457;
w24459 <= pi0609 and w24330;
w24460 <= pi0181 and not w15188;
w24461 <= not pi0181 and not w15175;
w24462 <= pi0754 and not w24460;
w24463 <= not w24461 and w24462;
w24464 <= not pi0181 and w15192;
w24465 <= pi0181 and w15194;
w24466 <= not pi0754 and not w24465;
w24467 <= not w24464 and w24466;
w24468 <= not w24463 and not w24467;
w24469 <= not pi0039 and not w24468;
w24470 <= pi0181 and w15168;
w24471 <= not pi0181 and not w15109;
w24472 <= not pi0754 and not w24471;
w24473 <= not w24470 and w24472;
w24474 <= not pi0181 and w14967;
w24475 <= pi0181 and w15048;
w24476 <= pi0754 and not w24475;
w24477 <= not w24474 and w24476;
w24478 <= pi0039 and not w24473;
w24479 <= not w24477 and w24478;
w24480 <= not pi0038 and not w24469;
w24481 <= not w24479 and w24480;
w24482 <= not w15032 and not w24138;
w24483 <= pi0181 and not w24482;
w24484 <= w3847 and w24483;
w24485 <= not pi0754 and not w15053;
w24486 <= w17034 and not w24485;
w24487 <= not pi0181 and not w24486;
w24488 <= pi0038 and not w24484;
w24489 <= not w24487 and w24488;
w24490 <= not pi0709 and not w24489;
w24491 <= not w24481 and w24490;
w24492 <= pi0709 and w24386;
w24493 <= w134 and not w24491;
w24494 <= not w24492 and w24493;
w24495 <= not w24368 and not w24494;
w24496 <= not pi0625 and w24495;
w24497 <= pi0625 and w24388;
w24498 <= not pi1153 and not w24497;
w24499 <= not w24496 and w24498;
w24500 <= not pi0608 and not w24323;
w24501 <= not w24499 and w24500;
w24502 <= not pi0625 and w24388;
w24503 <= pi0625 and w24495;
w24504 <= pi1153 and not w24502;
w24505 <= not w24503 and w24504;
w24506 <= pi0608 and not w24327;
w24507 <= not w24505 and w24506;
w24508 <= not w24501 and not w24507;
w24509 <= pi0778 and not w24508;
w24510 <= not pi0778 and w24495;
w24511 <= not w24509 and not w24510;
w24512 <= not pi0609 and not w24511;
w24513 <= not pi1155 and not w24459;
w24514 <= not w24512 and w24513;
w24515 <= not pi0660 and not w24396;
w24516 <= not w24514 and w24515;
w24517 <= not pi0609 and w24330;
w24518 <= pi0609 and not w24511;
w24519 <= pi1155 and not w24517;
w24520 <= not w24518 and w24519;
w24521 <= pi0660 and not w24400;
w24522 <= not w24520 and w24521;
w24523 <= not w24516 and not w24522;
w24524 <= pi0785 and not w24523;
w24525 <= not pi0785 and not w24511;
w24526 <= not w24524 and not w24525;
w24527 <= not pi0618 and not w24526;
w24528 <= pi0618 and w24333;
w24529 <= not pi1154 and not w24528;
w24530 <= not w24527 and w24529;
w24531 <= not pi0627 and not w24408;
w24532 <= not w24530 and w24531;
w24533 <= not pi0618 and w24333;
w24534 <= pi0618 and not w24526;
w24535 <= pi1154 and not w24533;
w24536 <= not w24534 and w24535;
w24537 <= pi0627 and not w24412;
w24538 <= not w24536 and w24537;
w24539 <= not w24532 and not w24538;
w24540 <= pi0781 and not w24539;
w24541 <= not pi0781 and not w24526;
w24542 <= not w24540 and not w24541;
w24543 <= not pi0789 and w24542;
w24544 <= pi0619 and not w24336;
w24545 <= not pi0619 and not w24542;
w24546 <= not pi1159 and not w24544;
w24547 <= not w24545 and w24546;
w24548 <= not pi0648 and not w24420;
w24549 <= not w24547 and w24548;
w24550 <= not pi0619 and not w24336;
w24551 <= pi0619 and not w24542;
w24552 <= pi1159 and not w24550;
w24553 <= not w24551 and w24552;
w24554 <= pi0648 and not w24424;
w24555 <= not w24553 and w24554;
w24556 <= pi0789 and not w24549;
w24557 <= not w24555 and w24556;
w24558 <= w15533 and not w24543;
w24559 <= not w24557 and w24558;
w24560 <= w15434 and w24338;
w24561 <= not pi0626 and not w24427;
w24562 <= pi0626 and not w24305;
w24563 <= w14192 and not w24562;
w24564 <= not w24561 and w24563;
w24565 <= pi0626 and not w24427;
w24566 <= not pi0626 and not w24305;
w24567 <= w14191 and not w24566;
w24568 <= not w24565 and w24567;
w24569 <= not w24560 and not w24564;
w24570 <= not w24568 and w24569;
w24571 <= pi0788 and not w24570;
w24572 <= not w17927 and not w24571;
w24573 <= not w24559 and w24572;
w24574 <= not w24458 and not w24573;
w24575 <= not w17769 and not w24574;
w24576 <= w15365 and not w24356;
w24577 <= not w18122 and w24433;
w24578 <= w15364 and not w24360;
w24579 <= not w24576 and not w24578;
w24580 <= not w24577 and w24579;
w24581 <= pi0787 and not w24580;
w24582 <= not pi0644 and w24449;
w24583 <= pi0644 and w24441;
w24584 <= pi0790 and not w24582;
w24585 <= not w24583 and w24584;
w24586 <= not w24575 and not w24581;
w24587 <= not w24585 and w24586;
w24588 <= not w24452 and not w24587;
w24589 <= w4989 and not w24588;
w24590 <= not pi0832 and not w24304;
w24591 <= not w24589 and w24590;
w24592 <= not w24303 and not w24591;
w24593 <= not pi0182 and not w489;
w24594 <= not pi0734 and w14208;
w24595 <= not w24593 and not w24594;
w24596 <= not pi0778 and not w24595;
w24597 <= not pi0625 and w24594;
w24598 <= not w24595 and not w24597;
w24599 <= pi1153 and not w24598;
w24600 <= not pi1153 and not w24593;
w24601 <= not w24597 and w24600;
w24602 <= pi0778 and not w24601;
w24603 <= not w24599 and w24602;
w24604 <= not w24596 and not w24603;
w24605 <= not w15408 and not w24604;
w24606 <= not w15410 and w24605;
w24607 <= not w15412 and w24606;
w24608 <= not w15414 and w24607;
w24609 <= not w15420 and w24608;
w24610 <= not pi0647 and w24609;
w24611 <= pi0647 and w24593;
w24612 <= not pi1157 and not w24611;
w24613 <= not w24610 and w24612;
w24614 <= pi0630 and w24613;
w24615 <= not pi0756 and w14807;
w24616 <= not w24593 and not w24615;
w24617 <= not w15437 and not w24616;
w24618 <= not pi0785 and not w24617;
w24619 <= w14859 and w24615;
w24620 <= w24617 and not w24619;
w24621 <= pi1155 and not w24620;
w24622 <= not pi1155 and not w24593;
w24623 <= not w24619 and w24622;
w24624 <= not w24621 and not w24623;
w24625 <= pi0785 and not w24624;
w24626 <= not w24618 and not w24625;
w24627 <= not pi0781 and not w24626;
w24628 <= not w15452 and w24626;
w24629 <= pi1154 and not w24628;
w24630 <= not w15455 and w24626;
w24631 <= not pi1154 and not w24630;
w24632 <= not w24629 and not w24631;
w24633 <= pi0781 and not w24632;
w24634 <= not w24627 and not w24633;
w24635 <= not pi0789 and not w24634;
w24636 <= not w20641 and w24634;
w24637 <= pi1159 and not w24636;
w24638 <= not w20644 and w24634;
w24639 <= not pi1159 and not w24638;
w24640 <= not w24637 and not w24639;
w24641 <= pi0789 and not w24640;
w24642 <= not w24635 and not w24641;
w24643 <= not w15532 and w24642;
w24644 <= w15532 and w24593;
w24645 <= not w24643 and not w24644;
w24646 <= not w15342 and not w24645;
w24647 <= w15342 and w24593;
w24648 <= not w24646 and not w24647;
w24649 <= not w18122 and w24648;
w24650 <= pi0647 and not w24609;
w24651 <= not pi0647 and not w24593;
w24652 <= not w24650 and not w24651;
w24653 <= w15364 and not w24652;
w24654 <= not w24614 and not w24653;
w24655 <= not w24649 and w24654;
w24656 <= pi0787 and not w24655;
w24657 <= w15434 and w24607;
w24658 <= not pi0626 and not w24642;
w24659 <= pi0626 and not w24593;
w24660 <= w14192 and not w24659;
w24661 <= not w24658 and w24660;
w24662 <= pi0626 and not w24642;
w24663 <= not pi0626 and not w24593;
w24664 <= w14191 and not w24663;
w24665 <= not w24662 and w24664;
w24666 <= not w24657 and not w24661;
w24667 <= not w24665 and w24666;
w24668 <= pi0788 and not w24667;
w24669 <= pi0618 and w24605;
w24670 <= not w14731 and not w24595;
w24671 <= pi0625 and w24670;
w24672 <= w24616 and not w24670;
w24673 <= not w24671 and not w24672;
w24674 <= w24600 and not w24673;
w24675 <= not pi0608 and not w24599;
w24676 <= not w24674 and w24675;
w24677 <= pi1153 and w24616;
w24678 <= not w24671 and w24677;
w24679 <= pi0608 and not w24601;
w24680 <= not w24678 and w24679;
w24681 <= not w24676 and not w24680;
w24682 <= pi0778 and not w24681;
w24683 <= not pi0778 and not w24672;
w24684 <= not w24682 and not w24683;
w24685 <= not pi0609 and not w24684;
w24686 <= pi0609 and not w24604;
w24687 <= not pi1155 and not w24686;
w24688 <= not w24685 and w24687;
w24689 <= not pi0660 and not w24621;
w24690 <= not w24688 and w24689;
w24691 <= pi0609 and not w24684;
w24692 <= not pi0609 and not w24604;
w24693 <= pi1155 and not w24692;
w24694 <= not w24691 and w24693;
w24695 <= pi0660 and not w24623;
w24696 <= not w24694 and w24695;
w24697 <= not w24690 and not w24696;
w24698 <= pi0785 and not w24697;
w24699 <= not pi0785 and not w24684;
w24700 <= not w24698 and not w24699;
w24701 <= not pi0618 and not w24700;
w24702 <= not pi1154 and not w24669;
w24703 <= not w24701 and w24702;
w24704 <= not pi0627 and not w24629;
w24705 <= not w24703 and w24704;
w24706 <= not pi0618 and w24605;
w24707 <= pi0618 and not w24700;
w24708 <= pi1154 and not w24706;
w24709 <= not w24707 and w24708;
w24710 <= pi0627 and not w24631;
w24711 <= not w24709 and w24710;
w24712 <= not w24705 and not w24711;
w24713 <= pi0781 and not w24712;
w24714 <= not pi0781 and not w24700;
w24715 <= not w24713 and not w24714;
w24716 <= not pi0789 and w24715;
w24717 <= not pi0619 and not w24715;
w24718 <= pi0619 and w24606;
w24719 <= not pi1159 and not w24718;
w24720 <= not w24717 and w24719;
w24721 <= not pi0648 and not w24637;
w24722 <= not w24720 and w24721;
w24723 <= pi0619 and not w24715;
w24724 <= not pi0619 and w24606;
w24725 <= pi1159 and not w24724;
w24726 <= not w24723 and w24725;
w24727 <= pi0648 and not w24639;
w24728 <= not w24726 and w24727;
w24729 <= pi0789 and not w24722;
w24730 <= not w24728 and w24729;
w24731 <= w15533 and not w24716;
w24732 <= not w24730 and w24731;
w24733 <= not w24668 and not w24732;
w24734 <= not w17927 and not w24733;
w24735 <= w15417 and not w24645;
w24736 <= w18414 and w24608;
w24737 <= not w24735 and not w24736;
w24738 <= not pi0629 and not w24737;
w24739 <= w18418 and w24608;
w24740 <= w15416 and not w24645;
w24741 <= not w24739 and not w24740;
w24742 <= pi0629 and not w24741;
w24743 <= not w24738 and not w24742;
w24744 <= pi0792 and not w24743;
w24745 <= not w17769 and not w24744;
w24746 <= not w24734 and w24745;
w24747 <= not w24656 and not w24746;
w24748 <= not pi0790 and w24747;
w24749 <= not pi0787 and not w24609;
w24750 <= pi1157 and not w24652;
w24751 <= not w24613 and not w24750;
w24752 <= pi0787 and not w24751;
w24753 <= not w24749 and not w24752;
w24754 <= not pi0644 and w24753;
w24755 <= pi0644 and w24747;
w24756 <= pi0715 and not w24754;
w24757 <= not w24755 and w24756;
w24758 <= not w15367 and not w24648;
w24759 <= w15367 and w24593;
w24760 <= not w24758 and not w24759;
w24761 <= pi0644 and not w24760;
w24762 <= not pi0644 and w24593;
w24763 <= not pi0715 and not w24762;
w24764 <= not w24761 and w24763;
w24765 <= pi1160 and not w24764;
w24766 <= not w24757 and w24765;
w24767 <= not pi0644 and not w24760;
w24768 <= pi0644 and w24593;
w24769 <= pi0715 and not w24768;
w24770 <= not w24767 and w24769;
w24771 <= pi0644 and w24753;
w24772 <= not pi0644 and w24747;
w24773 <= not pi0715 and not w24771;
w24774 <= not w24772 and w24773;
w24775 <= not pi1160 and not w24770;
w24776 <= not w24774 and w24775;
w24777 <= not w24766 and not w24776;
w24778 <= pi0790 and not w24777;
w24779 <= pi0832 and not w24748;
w24780 <= not w24778 and w24779;
w24781 <= not pi0182 and not w4989;
w24782 <= not pi0182 and not w14622;
w24783 <= w14198 and not w24782;
w24784 <= not pi0734 and w134;
w24785 <= w24782 and not w24784;
w24786 <= not pi0182 and not w14204;
w24787 <= w14210 and not w24786;
w24788 <= pi0182 and not w15639;
w24789 <= not pi0038 and not w24788;
w24790 <= w134 and not w24789;
w24791 <= not pi0182 and w15635;
w24792 <= not w24790 and not w24791;
w24793 <= not pi0734 and not w24787;
w24794 <= not w24792 and w24793;
w24795 <= not w24785 and not w24794;
w24796 <= not pi0778 and w24795;
w24797 <= not pi0625 and w24782;
w24798 <= pi0625 and not w24795;
w24799 <= pi1153 and not w24797;
w24800 <= not w24798 and w24799;
w24801 <= pi0625 and w24782;
w24802 <= not pi0625 and not w24795;
w24803 <= not pi1153 and not w24801;
w24804 <= not w24802 and w24803;
w24805 <= not w24800 and not w24804;
w24806 <= pi0778 and not w24805;
w24807 <= not w24796 and not w24806;
w24808 <= not w14638 and not w24807;
w24809 <= w14638 and not w24782;
w24810 <= not w24808 and not w24809;
w24811 <= not w14202 and w24810;
w24812 <= w14202 and w24782;
w24813 <= not w24811 and not w24812;
w24814 <= not w14198 and w24813;
w24815 <= not w24783 and not w24814;
w24816 <= not w14194 and w24815;
w24817 <= w14194 and w24782;
w24818 <= not w24816 and not w24817;
w24819 <= not pi0792 and w24818;
w24820 <= pi0628 and not w24818;
w24821 <= not pi0628 and w24782;
w24822 <= pi1156 and not w24821;
w24823 <= not w24820 and w24822;
w24824 <= pi0628 and w24782;
w24825 <= not pi0628 and not w24818;
w24826 <= not pi1156 and not w24824;
w24827 <= not w24825 and w24826;
w24828 <= not w24823 and not w24827;
w24829 <= pi0792 and not w24828;
w24830 <= not w24819 and not w24829;
w24831 <= not pi0647 and not w24830;
w24832 <= pi0647 and not w24782;
w24833 <= not w24831 and not w24832;
w24834 <= not pi1157 and w24833;
w24835 <= pi0647 and not w24830;
w24836 <= not pi0647 and not w24782;
w24837 <= not w24835 and not w24836;
w24838 <= pi1157 and w24837;
w24839 <= not w24834 and not w24838;
w24840 <= pi0787 and not w24839;
w24841 <= not pi0787 and w24830;
w24842 <= not w24840 and not w24841;
w24843 <= not pi0644 and not w24842;
w24844 <= pi0715 and not w24843;
w24845 <= pi0182 and not w134;
w24846 <= not pi0756 and w14843;
w24847 <= not w24786 and not w24846;
w24848 <= pi0038 and not w24847;
w24849 <= not pi0182 and w14784;
w24850 <= pi0182 and not w14838;
w24851 <= not pi0756 and not w24850;
w24852 <= not w24849 and w24851;
w24853 <= not pi0182 and pi0756;
w24854 <= not w14611 and w24853;
w24855 <= not w24852 and not w24854;
w24856 <= not pi0038 and not w24855;
w24857 <= not w24848 and not w24856;
w24858 <= w134 and w24857;
w24859 <= not w24845 and not w24858;
w24860 <= not w14680 and not w24859;
w24861 <= w14680 and not w24782;
w24862 <= not w24860 and not w24861;
w24863 <= not pi0785 and not w24862;
w24864 <= not w14854 and not w24782;
w24865 <= pi0609 and w24860;
w24866 <= not w24864 and not w24865;
w24867 <= pi1155 and not w24866;
w24868 <= not w14859 and not w24782;
w24869 <= not pi0609 and w24860;
w24870 <= not w24868 and not w24869;
w24871 <= not pi1155 and not w24870;
w24872 <= not w24867 and not w24871;
w24873 <= pi0785 and not w24872;
w24874 <= not w24863 and not w24873;
w24875 <= not pi0781 and not w24874;
w24876 <= not pi0618 and w24782;
w24877 <= pi0618 and w24874;
w24878 <= pi1154 and not w24876;
w24879 <= not w24877 and w24878;
w24880 <= not pi0618 and w24874;
w24881 <= pi0618 and w24782;
w24882 <= not pi1154 and not w24881;
w24883 <= not w24880 and w24882;
w24884 <= not w24879 and not w24883;
w24885 <= pi0781 and not w24884;
w24886 <= not w24875 and not w24885;
w24887 <= not pi0789 and not w24886;
w24888 <= not pi0619 and w24782;
w24889 <= pi0619 and w24886;
w24890 <= pi1159 and not w24888;
w24891 <= not w24889 and w24890;
w24892 <= not pi0619 and w24886;
w24893 <= pi0619 and w24782;
w24894 <= not pi1159 and not w24893;
w24895 <= not w24892 and w24894;
w24896 <= not w24891 and not w24895;
w24897 <= pi0789 and not w24896;
w24898 <= not w24887 and not w24897;
w24899 <= not w15532 and w24898;
w24900 <= w15532 and w24782;
w24901 <= not w24899 and not w24900;
w24902 <= not w15342 and not w24901;
w24903 <= w15342 and w24782;
w24904 <= not w24902 and not w24903;
w24905 <= not w15367 and not w24904;
w24906 <= w15367 and w24782;
w24907 <= not w24905 and not w24906;
w24908 <= pi0644 and not w24907;
w24909 <= not pi0644 and w24782;
w24910 <= not pi0715 and not w24909;
w24911 <= not w24908 and w24910;
w24912 <= pi1160 and not w24911;
w24913 <= not w24844 and w24912;
w24914 <= pi0644 and not w24842;
w24915 <= not pi0715 and not w24914;
w24916 <= not pi0644 and not w24907;
w24917 <= pi0644 and w24782;
w24918 <= pi0715 and not w24917;
w24919 <= not w24916 and w24918;
w24920 <= not pi1160 and not w24919;
w24921 <= not w24915 and w24920;
w24922 <= not w24913 and not w24921;
w24923 <= pi0790 and not w24922;
w24924 <= not pi0629 and w24823;
w24925 <= not w18133 and w24901;
w24926 <= pi0629 and w24827;
w24927 <= not w24924 and not w24926;
w24928 <= not w24925 and w24927;
w24929 <= pi0792 and not w24928;
w24930 <= pi0609 and w24807;
w24931 <= pi0182 and not w15188;
w24932 <= not pi0182 and not w15175;
w24933 <= pi0756 and not w24931;
w24934 <= not w24932 and w24933;
w24935 <= not pi0182 and w15192;
w24936 <= pi0182 and w15194;
w24937 <= not pi0756 and not w24936;
w24938 <= not w24935 and w24937;
w24939 <= not w24934 and not w24938;
w24940 <= not pi0039 and not w24939;
w24941 <= pi0182 and w15168;
w24942 <= not pi0182 and not w15109;
w24943 <= not pi0756 and not w24942;
w24944 <= not w24941 and w24943;
w24945 <= not pi0182 and w14967;
w24946 <= pi0182 and w15048;
w24947 <= pi0756 and not w24946;
w24948 <= not w24945 and w24947;
w24949 <= pi0039 and not w24944;
w24950 <= not w24948 and w24949;
w24951 <= not pi0038 and not w24940;
w24952 <= not w24950 and w24951;
w24953 <= not pi0756 and not w15053;
w24954 <= w17034 and not w24953;
w24955 <= not pi0182 and not w24954;
w24956 <= not w15032 and not w24615;
w24957 <= pi0182 and not w24956;
w24958 <= w3847 and w24957;
w24959 <= pi0038 and not w24958;
w24960 <= not w24955 and w24959;
w24961 <= not pi0734 and not w24960;
w24962 <= not w24952 and w24961;
w24963 <= pi0734 and not w24857;
w24964 <= w134 and not w24962;
w24965 <= not w24963 and w24964;
w24966 <= not w24845 and not w24965;
w24967 <= not pi0625 and w24966;
w24968 <= pi0625 and w24859;
w24969 <= not pi1153 and not w24968;
w24970 <= not w24967 and w24969;
w24971 <= not pi0608 and not w24800;
w24972 <= not w24970 and w24971;
w24973 <= not pi0625 and w24859;
w24974 <= pi0625 and w24966;
w24975 <= pi1153 and not w24973;
w24976 <= not w24974 and w24975;
w24977 <= pi0608 and not w24804;
w24978 <= not w24976 and w24977;
w24979 <= not w24972 and not w24978;
w24980 <= pi0778 and not w24979;
w24981 <= not pi0778 and w24966;
w24982 <= not w24980 and not w24981;
w24983 <= not pi0609 and not w24982;
w24984 <= not pi1155 and not w24930;
w24985 <= not w24983 and w24984;
w24986 <= not pi0660 and not w24867;
w24987 <= not w24985 and w24986;
w24988 <= not pi0609 and w24807;
w24989 <= pi0609 and not w24982;
w24990 <= pi1155 and not w24988;
w24991 <= not w24989 and w24990;
w24992 <= pi0660 and not w24871;
w24993 <= not w24991 and w24992;
w24994 <= not w24987 and not w24993;
w24995 <= pi0785 and not w24994;
w24996 <= not pi0785 and not w24982;
w24997 <= not w24995 and not w24996;
w24998 <= not pi0618 and not w24997;
w24999 <= pi0618 and w24810;
w25000 <= not pi1154 and not w24999;
w25001 <= not w24998 and w25000;
w25002 <= not pi0627 and not w24879;
w25003 <= not w25001 and w25002;
w25004 <= not pi0618 and w24810;
w25005 <= pi0618 and not w24997;
w25006 <= pi1154 and not w25004;
w25007 <= not w25005 and w25006;
w25008 <= pi0627 and not w24883;
w25009 <= not w25007 and w25008;
w25010 <= not w25003 and not w25009;
w25011 <= pi0781 and not w25010;
w25012 <= not pi0781 and not w24997;
w25013 <= not w25011 and not w25012;
w25014 <= not pi0789 and w25013;
w25015 <= pi0619 and not w24813;
w25016 <= not pi0619 and not w25013;
w25017 <= not pi1159 and not w25015;
w25018 <= not w25016 and w25017;
w25019 <= not pi0648 and not w24891;
w25020 <= not w25018 and w25019;
w25021 <= not pi0619 and not w24813;
w25022 <= pi0619 and not w25013;
w25023 <= pi1159 and not w25021;
w25024 <= not w25022 and w25023;
w25025 <= pi0648 and not w24895;
w25026 <= not w25024 and w25025;
w25027 <= pi0789 and not w25020;
w25028 <= not w25026 and w25027;
w25029 <= w15533 and not w25014;
w25030 <= not w25028 and w25029;
w25031 <= w15434 and w24815;
w25032 <= not pi0626 and not w24898;
w25033 <= pi0626 and not w24782;
w25034 <= w14192 and not w25033;
w25035 <= not w25032 and w25034;
w25036 <= pi0626 and not w24898;
w25037 <= not pi0626 and not w24782;
w25038 <= w14191 and not w25037;
w25039 <= not w25036 and w25038;
w25040 <= not w25031 and not w25035;
w25041 <= not w25039 and w25040;
w25042 <= pi0788 and not w25041;
w25043 <= not w17927 and not w25042;
w25044 <= not w25030 and w25043;
w25045 <= not w24929 and not w25044;
w25046 <= not w17769 and not w25045;
w25047 <= w15365 and not w24833;
w25048 <= not w18122 and w24904;
w25049 <= w15364 and not w24837;
w25050 <= not w25047 and not w25049;
w25051 <= not w25048 and w25050;
w25052 <= pi0787 and not w25051;
w25053 <= not pi0644 and w24920;
w25054 <= pi0644 and w24912;
w25055 <= pi0790 and not w25053;
w25056 <= not w25054 and w25055;
w25057 <= not w25046 and not w25052;
w25058 <= not w25056 and w25057;
w25059 <= not w24923 and not w25058;
w25060 <= w4989 and not w25059;
w25061 <= not pi0832 and not w24781;
w25062 <= not w25060 and w25061;
w25063 <= not w24780 and not w25062;
w25064 <= not pi0183 and not w489;
w25065 <= not pi0725 and w14208;
w25066 <= not w25064 and not w25065;
w25067 <= not pi0778 and not w25066;
w25068 <= not pi0625 and w25065;
w25069 <= not w25066 and not w25068;
w25070 <= pi1153 and not w25069;
w25071 <= not pi1153 and not w25064;
w25072 <= not w25068 and w25071;
w25073 <= pi0778 and not w25072;
w25074 <= not w25070 and w25073;
w25075 <= not w25067 and not w25074;
w25076 <= not w15408 and not w25075;
w25077 <= not w15410 and w25076;
w25078 <= not w15412 and w25077;
w25079 <= not w15414 and w25078;
w25080 <= not w15420 and w25079;
w25081 <= not pi0647 and w25080;
w25082 <= pi0647 and w25064;
w25083 <= not pi1157 and not w25082;
w25084 <= not w25081 and w25083;
w25085 <= pi0630 and w25084;
w25086 <= not pi0755 and w14807;
w25087 <= not w25064 and not w25086;
w25088 <= not w15437 and not w25087;
w25089 <= not pi0785 and not w25088;
w25090 <= w14859 and w25086;
w25091 <= w25088 and not w25090;
w25092 <= pi1155 and not w25091;
w25093 <= not pi1155 and not w25064;
w25094 <= not w25090 and w25093;
w25095 <= not w25092 and not w25094;
w25096 <= pi0785 and not w25095;
w25097 <= not w25089 and not w25096;
w25098 <= not pi0781 and not w25097;
w25099 <= not w15452 and w25097;
w25100 <= pi1154 and not w25099;
w25101 <= not w15455 and w25097;
w25102 <= not pi1154 and not w25101;
w25103 <= not w25100 and not w25102;
w25104 <= pi0781 and not w25103;
w25105 <= not w25098 and not w25104;
w25106 <= not pi0789 and not w25105;
w25107 <= not w20641 and w25105;
w25108 <= pi1159 and not w25107;
w25109 <= not w20644 and w25105;
w25110 <= not pi1159 and not w25109;
w25111 <= not w25108 and not w25110;
w25112 <= pi0789 and not w25111;
w25113 <= not w25106 and not w25112;
w25114 <= not w15532 and w25113;
w25115 <= w15532 and w25064;
w25116 <= not w25114 and not w25115;
w25117 <= not w15342 and not w25116;
w25118 <= w15342 and w25064;
w25119 <= not w25117 and not w25118;
w25120 <= not w18122 and w25119;
w25121 <= pi0647 and not w25080;
w25122 <= not pi0647 and not w25064;
w25123 <= not w25121 and not w25122;
w25124 <= w15364 and not w25123;
w25125 <= not w25085 and not w25124;
w25126 <= not w25120 and w25125;
w25127 <= pi0787 and not w25126;
w25128 <= w15434 and w25078;
w25129 <= not pi0626 and not w25113;
w25130 <= pi0626 and not w25064;
w25131 <= w14192 and not w25130;
w25132 <= not w25129 and w25131;
w25133 <= pi0626 and not w25113;
w25134 <= not pi0626 and not w25064;
w25135 <= w14191 and not w25134;
w25136 <= not w25133 and w25135;
w25137 <= not w25128 and not w25132;
w25138 <= not w25136 and w25137;
w25139 <= pi0788 and not w25138;
w25140 <= pi0618 and w25076;
w25141 <= not w14731 and not w25066;
w25142 <= pi0625 and w25141;
w25143 <= w25087 and not w25141;
w25144 <= not w25142 and not w25143;
w25145 <= w25071 and not w25144;
w25146 <= not pi0608 and not w25070;
w25147 <= not w25145 and w25146;
w25148 <= pi1153 and w25087;
w25149 <= not w25142 and w25148;
w25150 <= pi0608 and not w25072;
w25151 <= not w25149 and w25150;
w25152 <= not w25147 and not w25151;
w25153 <= pi0778 and not w25152;
w25154 <= not pi0778 and not w25143;
w25155 <= not w25153 and not w25154;
w25156 <= not pi0609 and not w25155;
w25157 <= pi0609 and not w25075;
w25158 <= not pi1155 and not w25157;
w25159 <= not w25156 and w25158;
w25160 <= not pi0660 and not w25092;
w25161 <= not w25159 and w25160;
w25162 <= pi0609 and not w25155;
w25163 <= not pi0609 and not w25075;
w25164 <= pi1155 and not w25163;
w25165 <= not w25162 and w25164;
w25166 <= pi0660 and not w25094;
w25167 <= not w25165 and w25166;
w25168 <= not w25161 and not w25167;
w25169 <= pi0785 and not w25168;
w25170 <= not pi0785 and not w25155;
w25171 <= not w25169 and not w25170;
w25172 <= not pi0618 and not w25171;
w25173 <= not pi1154 and not w25140;
w25174 <= not w25172 and w25173;
w25175 <= not pi0627 and not w25100;
w25176 <= not w25174 and w25175;
w25177 <= not pi0618 and w25076;
w25178 <= pi0618 and not w25171;
w25179 <= pi1154 and not w25177;
w25180 <= not w25178 and w25179;
w25181 <= pi0627 and not w25102;
w25182 <= not w25180 and w25181;
w25183 <= not w25176 and not w25182;
w25184 <= pi0781 and not w25183;
w25185 <= not pi0781 and not w25171;
w25186 <= not w25184 and not w25185;
w25187 <= not pi0789 and w25186;
w25188 <= not pi0619 and not w25186;
w25189 <= pi0619 and w25077;
w25190 <= not pi1159 and not w25189;
w25191 <= not w25188 and w25190;
w25192 <= not pi0648 and not w25108;
w25193 <= not w25191 and w25192;
w25194 <= pi0619 and not w25186;
w25195 <= not pi0619 and w25077;
w25196 <= pi1159 and not w25195;
w25197 <= not w25194 and w25196;
w25198 <= pi0648 and not w25110;
w25199 <= not w25197 and w25198;
w25200 <= pi0789 and not w25193;
w25201 <= not w25199 and w25200;
w25202 <= w15533 and not w25187;
w25203 <= not w25201 and w25202;
w25204 <= not w25139 and not w25203;
w25205 <= not w17927 and not w25204;
w25206 <= w15417 and not w25116;
w25207 <= w18414 and w25079;
w25208 <= not w25206 and not w25207;
w25209 <= not pi0629 and not w25208;
w25210 <= w18418 and w25079;
w25211 <= w15416 and not w25116;
w25212 <= not w25210 and not w25211;
w25213 <= pi0629 and not w25212;
w25214 <= not w25209 and not w25213;
w25215 <= pi0792 and not w25214;
w25216 <= not w17769 and not w25215;
w25217 <= not w25205 and w25216;
w25218 <= not w25127 and not w25217;
w25219 <= not pi0790 and w25218;
w25220 <= not pi0787 and not w25080;
w25221 <= pi1157 and not w25123;
w25222 <= not w25084 and not w25221;
w25223 <= pi0787 and not w25222;
w25224 <= not w25220 and not w25223;
w25225 <= not pi0644 and w25224;
w25226 <= pi0644 and w25218;
w25227 <= pi0715 and not w25225;
w25228 <= not w25226 and w25227;
w25229 <= not w15367 and not w25119;
w25230 <= w15367 and w25064;
w25231 <= not w25229 and not w25230;
w25232 <= pi0644 and not w25231;
w25233 <= not pi0644 and w25064;
w25234 <= not pi0715 and not w25233;
w25235 <= not w25232 and w25234;
w25236 <= pi1160 and not w25235;
w25237 <= not w25228 and w25236;
w25238 <= not pi0644 and not w25231;
w25239 <= pi0644 and w25064;
w25240 <= pi0715 and not w25239;
w25241 <= not w25238 and w25240;
w25242 <= pi0644 and w25224;
w25243 <= not pi0644 and w25218;
w25244 <= not pi0715 and not w25242;
w25245 <= not w25243 and w25244;
w25246 <= not pi1160 and not w25241;
w25247 <= not w25245 and w25246;
w25248 <= not w25237 and not w25247;
w25249 <= pi0790 and not w25248;
w25250 <= pi0832 and not w25219;
w25251 <= not w25249 and w25250;
w25252 <= not pi0183 and not w4989;
w25253 <= not pi0183 and not w14622;
w25254 <= w14198 and not w25253;
w25255 <= not pi0725 and w134;
w25256 <= w25253 and not w25255;
w25257 <= not pi0183 and not w14204;
w25258 <= w14210 and not w25257;
w25259 <= pi0183 and not w15639;
w25260 <= not pi0038 and not w25259;
w25261 <= w134 and not w25260;
w25262 <= not pi0183 and w15635;
w25263 <= not w25261 and not w25262;
w25264 <= not pi0725 and not w25258;
w25265 <= not w25263 and w25264;
w25266 <= not w25256 and not w25265;
w25267 <= not pi0778 and w25266;
w25268 <= not pi0625 and w25253;
w25269 <= pi0625 and not w25266;
w25270 <= pi1153 and not w25268;
w25271 <= not w25269 and w25270;
w25272 <= pi0625 and w25253;
w25273 <= not pi0625 and not w25266;
w25274 <= not pi1153 and not w25272;
w25275 <= not w25273 and w25274;
w25276 <= not w25271 and not w25275;
w25277 <= pi0778 and not w25276;
w25278 <= not w25267 and not w25277;
w25279 <= not w14638 and not w25278;
w25280 <= w14638 and not w25253;
w25281 <= not w25279 and not w25280;
w25282 <= not w14202 and w25281;
w25283 <= w14202 and w25253;
w25284 <= not w25282 and not w25283;
w25285 <= not w14198 and w25284;
w25286 <= not w25254 and not w25285;
w25287 <= not w14194 and w25286;
w25288 <= w14194 and w25253;
w25289 <= not w25287 and not w25288;
w25290 <= not pi0792 and w25289;
w25291 <= pi0628 and not w25289;
w25292 <= not pi0628 and w25253;
w25293 <= pi1156 and not w25292;
w25294 <= not w25291 and w25293;
w25295 <= pi0628 and w25253;
w25296 <= not pi0628 and not w25289;
w25297 <= not pi1156 and not w25295;
w25298 <= not w25296 and w25297;
w25299 <= not w25294 and not w25298;
w25300 <= pi0792 and not w25299;
w25301 <= not w25290 and not w25300;
w25302 <= not pi0647 and not w25301;
w25303 <= pi0647 and not w25253;
w25304 <= not w25302 and not w25303;
w25305 <= not pi1157 and w25304;
w25306 <= pi0647 and not w25301;
w25307 <= not pi0647 and not w25253;
w25308 <= not w25306 and not w25307;
w25309 <= pi1157 and w25308;
w25310 <= not w25305 and not w25309;
w25311 <= pi0787 and not w25310;
w25312 <= not pi0787 and w25301;
w25313 <= not w25311 and not w25312;
w25314 <= not pi0644 and not w25313;
w25315 <= pi0715 and not w25314;
w25316 <= pi0183 and not w134;
w25317 <= not pi0755 and w14843;
w25318 <= not w25257 and not w25317;
w25319 <= pi0038 and not w25318;
w25320 <= not pi0183 and w14784;
w25321 <= pi0183 and not w14838;
w25322 <= not pi0755 and not w25321;
w25323 <= not w25320 and w25322;
w25324 <= not pi0183 and pi0755;
w25325 <= not w14611 and w25324;
w25326 <= not w25323 and not w25325;
w25327 <= not pi0038 and not w25326;
w25328 <= not w25319 and not w25327;
w25329 <= w134 and w25328;
w25330 <= not w25316 and not w25329;
w25331 <= not w14680 and not w25330;
w25332 <= w14680 and not w25253;
w25333 <= not w25331 and not w25332;
w25334 <= not pi0785 and not w25333;
w25335 <= not w14854 and not w25253;
w25336 <= pi0609 and w25331;
w25337 <= not w25335 and not w25336;
w25338 <= pi1155 and not w25337;
w25339 <= not w14859 and not w25253;
w25340 <= not pi0609 and w25331;
w25341 <= not w25339 and not w25340;
w25342 <= not pi1155 and not w25341;
w25343 <= not w25338 and not w25342;
w25344 <= pi0785 and not w25343;
w25345 <= not w25334 and not w25344;
w25346 <= not pi0781 and not w25345;
w25347 <= not pi0618 and w25253;
w25348 <= pi0618 and w25345;
w25349 <= pi1154 and not w25347;
w25350 <= not w25348 and w25349;
w25351 <= not pi0618 and w25345;
w25352 <= pi0618 and w25253;
w25353 <= not pi1154 and not w25352;
w25354 <= not w25351 and w25353;
w25355 <= not w25350 and not w25354;
w25356 <= pi0781 and not w25355;
w25357 <= not w25346 and not w25356;
w25358 <= not pi0789 and not w25357;
w25359 <= not pi0619 and w25253;
w25360 <= pi0619 and w25357;
w25361 <= pi1159 and not w25359;
w25362 <= not w25360 and w25361;
w25363 <= not pi0619 and w25357;
w25364 <= pi0619 and w25253;
w25365 <= not pi1159 and not w25364;
w25366 <= not w25363 and w25365;
w25367 <= not w25362 and not w25366;
w25368 <= pi0789 and not w25367;
w25369 <= not w25358 and not w25368;
w25370 <= not w15532 and w25369;
w25371 <= w15532 and w25253;
w25372 <= not w25370 and not w25371;
w25373 <= not w15342 and not w25372;
w25374 <= w15342 and w25253;
w25375 <= not w25373 and not w25374;
w25376 <= not w15367 and not w25375;
w25377 <= w15367 and w25253;
w25378 <= not w25376 and not w25377;
w25379 <= pi0644 and not w25378;
w25380 <= not pi0644 and w25253;
w25381 <= not pi0715 and not w25380;
w25382 <= not w25379 and w25381;
w25383 <= pi1160 and not w25382;
w25384 <= not w25315 and w25383;
w25385 <= pi0644 and not w25313;
w25386 <= not pi0715 and not w25385;
w25387 <= not pi0644 and not w25378;
w25388 <= pi0644 and w25253;
w25389 <= pi0715 and not w25388;
w25390 <= not w25387 and w25389;
w25391 <= not pi1160 and not w25390;
w25392 <= not w25386 and w25391;
w25393 <= not w25384 and not w25392;
w25394 <= pi0790 and not w25393;
w25395 <= not pi0629 and w25294;
w25396 <= not w18133 and w25372;
w25397 <= pi0629 and w25298;
w25398 <= not w25395 and not w25397;
w25399 <= not w25396 and w25398;
w25400 <= pi0792 and not w25399;
w25401 <= pi0609 and w25278;
w25402 <= pi0183 and not w15188;
w25403 <= not pi0183 and not w15175;
w25404 <= pi0755 and not w25402;
w25405 <= not w25403 and w25404;
w25406 <= not pi0183 and w15192;
w25407 <= pi0183 and w15194;
w25408 <= not pi0755 and not w25407;
w25409 <= not w25406 and w25408;
w25410 <= not w25405 and not w25409;
w25411 <= not pi0039 and not w25410;
w25412 <= pi0183 and w15168;
w25413 <= not pi0183 and not w15109;
w25414 <= not pi0755 and not w25413;
w25415 <= not w25412 and w25414;
w25416 <= not pi0183 and w14967;
w25417 <= pi0183 and w15048;
w25418 <= pi0755 and not w25417;
w25419 <= not w25416 and w25418;
w25420 <= pi0039 and not w25415;
w25421 <= not w25419 and w25420;
w25422 <= not pi0038 and not w25411;
w25423 <= not w25421 and w25422;
w25424 <= not pi0755 and not w15053;
w25425 <= w17034 and not w25424;
w25426 <= not pi0183 and not w25425;
w25427 <= not w15032 and not w25086;
w25428 <= pi0183 and not w25427;
w25429 <= w3847 and w25428;
w25430 <= pi0038 and not w25429;
w25431 <= not w25426 and w25430;
w25432 <= not pi0725 and not w25431;
w25433 <= not w25423 and w25432;
w25434 <= pi0725 and not w25328;
w25435 <= w134 and not w25433;
w25436 <= not w25434 and w25435;
w25437 <= not w25316 and not w25436;
w25438 <= not pi0625 and w25437;
w25439 <= pi0625 and w25330;
w25440 <= not pi1153 and not w25439;
w25441 <= not w25438 and w25440;
w25442 <= not pi0608 and not w25271;
w25443 <= not w25441 and w25442;
w25444 <= not pi0625 and w25330;
w25445 <= pi0625 and w25437;
w25446 <= pi1153 and not w25444;
w25447 <= not w25445 and w25446;
w25448 <= pi0608 and not w25275;
w25449 <= not w25447 and w25448;
w25450 <= not w25443 and not w25449;
w25451 <= pi0778 and not w25450;
w25452 <= not pi0778 and w25437;
w25453 <= not w25451 and not w25452;
w25454 <= not pi0609 and not w25453;
w25455 <= not pi1155 and not w25401;
w25456 <= not w25454 and w25455;
w25457 <= not pi0660 and not w25338;
w25458 <= not w25456 and w25457;
w25459 <= not pi0609 and w25278;
w25460 <= pi0609 and not w25453;
w25461 <= pi1155 and not w25459;
w25462 <= not w25460 and w25461;
w25463 <= pi0660 and not w25342;
w25464 <= not w25462 and w25463;
w25465 <= not w25458 and not w25464;
w25466 <= pi0785 and not w25465;
w25467 <= not pi0785 and not w25453;
w25468 <= not w25466 and not w25467;
w25469 <= not pi0618 and not w25468;
w25470 <= pi0618 and w25281;
w25471 <= not pi1154 and not w25470;
w25472 <= not w25469 and w25471;
w25473 <= not pi0627 and not w25350;
w25474 <= not w25472 and w25473;
w25475 <= not pi0618 and w25281;
w25476 <= pi0618 and not w25468;
w25477 <= pi1154 and not w25475;
w25478 <= not w25476 and w25477;
w25479 <= pi0627 and not w25354;
w25480 <= not w25478 and w25479;
w25481 <= not w25474 and not w25480;
w25482 <= pi0781 and not w25481;
w25483 <= not pi0781 and not w25468;
w25484 <= not w25482 and not w25483;
w25485 <= not pi0789 and w25484;
w25486 <= pi0619 and not w25284;
w25487 <= not pi0619 and not w25484;
w25488 <= not pi1159 and not w25486;
w25489 <= not w25487 and w25488;
w25490 <= not pi0648 and not w25362;
w25491 <= not w25489 and w25490;
w25492 <= not pi0619 and not w25284;
w25493 <= pi0619 and not w25484;
w25494 <= pi1159 and not w25492;
w25495 <= not w25493 and w25494;
w25496 <= pi0648 and not w25366;
w25497 <= not w25495 and w25496;
w25498 <= pi0789 and not w25491;
w25499 <= not w25497 and w25498;
w25500 <= w15533 and not w25485;
w25501 <= not w25499 and w25500;
w25502 <= w15434 and w25286;
w25503 <= not pi0626 and not w25369;
w25504 <= pi0626 and not w25253;
w25505 <= w14192 and not w25504;
w25506 <= not w25503 and w25505;
w25507 <= pi0626 and not w25369;
w25508 <= not pi0626 and not w25253;
w25509 <= w14191 and not w25508;
w25510 <= not w25507 and w25509;
w25511 <= not w25502 and not w25506;
w25512 <= not w25510 and w25511;
w25513 <= pi0788 and not w25512;
w25514 <= not w17927 and not w25513;
w25515 <= not w25501 and w25514;
w25516 <= not w25400 and not w25515;
w25517 <= not w17769 and not w25516;
w25518 <= w15365 and not w25304;
w25519 <= not w18122 and w25375;
w25520 <= w15364 and not w25308;
w25521 <= not w25518 and not w25520;
w25522 <= not w25519 and w25521;
w25523 <= pi0787 and not w25522;
w25524 <= not pi0644 and w25391;
w25525 <= pi0644 and w25383;
w25526 <= pi0790 and not w25524;
w25527 <= not w25525 and w25526;
w25528 <= not w25517 and not w25523;
w25529 <= not w25527 and w25528;
w25530 <= not w25394 and not w25529;
w25531 <= w4989 and not w25530;
w25532 <= not pi0832 and not w25252;
w25533 <= not w25531 and w25532;
w25534 <= not w25251 and not w25533;
w25535 <= not pi0184 and not w489;
w25536 <= not pi0737 and w14208;
w25537 <= not w25535 and not w25536;
w25538 <= not pi0778 and not w25537;
w25539 <= not pi0625 and w25536;
w25540 <= not w25537 and not w25539;
w25541 <= pi1153 and not w25540;
w25542 <= not pi1153 and not w25535;
w25543 <= not w25539 and w25542;
w25544 <= pi0778 and not w25543;
w25545 <= not w25541 and w25544;
w25546 <= not w25538 and not w25545;
w25547 <= not w15408 and not w25546;
w25548 <= not w15410 and w25547;
w25549 <= not w15412 and w25548;
w25550 <= not w15414 and w25549;
w25551 <= not w15420 and w25550;
w25552 <= not pi0647 and w25551;
w25553 <= pi0647 and w25535;
w25554 <= not pi1157 and not w25553;
w25555 <= not w25552 and w25554;
w25556 <= pi0630 and w25555;
w25557 <= not pi0777 and w14807;
w25558 <= not w25535 and not w25557;
w25559 <= not w15437 and not w25558;
w25560 <= not pi0785 and not w25559;
w25561 <= w14859 and w25557;
w25562 <= w25559 and not w25561;
w25563 <= pi1155 and not w25562;
w25564 <= not pi1155 and not w25535;
w25565 <= not w25561 and w25564;
w25566 <= not w25563 and not w25565;
w25567 <= pi0785 and not w25566;
w25568 <= not w25560 and not w25567;
w25569 <= not pi0781 and not w25568;
w25570 <= not w15452 and w25568;
w25571 <= pi1154 and not w25570;
w25572 <= not w15455 and w25568;
w25573 <= not pi1154 and not w25572;
w25574 <= not w25571 and not w25573;
w25575 <= pi0781 and not w25574;
w25576 <= not w25569 and not w25575;
w25577 <= not pi0789 and not w25576;
w25578 <= not w20641 and w25576;
w25579 <= pi1159 and not w25578;
w25580 <= not w20644 and w25576;
w25581 <= not pi1159 and not w25580;
w25582 <= not w25579 and not w25581;
w25583 <= pi0789 and not w25582;
w25584 <= not w25577 and not w25583;
w25585 <= not w15532 and w25584;
w25586 <= w15532 and w25535;
w25587 <= not w25585 and not w25586;
w25588 <= not w15342 and not w25587;
w25589 <= w15342 and w25535;
w25590 <= not w25588 and not w25589;
w25591 <= not w18122 and w25590;
w25592 <= pi0647 and not w25551;
w25593 <= not pi0647 and not w25535;
w25594 <= not w25592 and not w25593;
w25595 <= w15364 and not w25594;
w25596 <= not w25556 and not w25595;
w25597 <= not w25591 and w25596;
w25598 <= pi0787 and not w25597;
w25599 <= w15434 and w25549;
w25600 <= not pi0626 and not w25584;
w25601 <= pi0626 and not w25535;
w25602 <= w14192 and not w25601;
w25603 <= not w25600 and w25602;
w25604 <= pi0626 and not w25584;
w25605 <= not pi0626 and not w25535;
w25606 <= w14191 and not w25605;
w25607 <= not w25604 and w25606;
w25608 <= not w25599 and not w25603;
w25609 <= not w25607 and w25608;
w25610 <= pi0788 and not w25609;
w25611 <= pi0618 and w25547;
w25612 <= not w14731 and not w25537;
w25613 <= pi0625 and w25612;
w25614 <= w25558 and not w25612;
w25615 <= not w25613 and not w25614;
w25616 <= w25542 and not w25615;
w25617 <= not pi0608 and not w25541;
w25618 <= not w25616 and w25617;
w25619 <= pi1153 and w25558;
w25620 <= not w25613 and w25619;
w25621 <= pi0608 and not w25543;
w25622 <= not w25620 and w25621;
w25623 <= not w25618 and not w25622;
w25624 <= pi0778 and not w25623;
w25625 <= not pi0778 and not w25614;
w25626 <= not w25624 and not w25625;
w25627 <= not pi0609 and not w25626;
w25628 <= pi0609 and not w25546;
w25629 <= not pi1155 and not w25628;
w25630 <= not w25627 and w25629;
w25631 <= not pi0660 and not w25563;
w25632 <= not w25630 and w25631;
w25633 <= pi0609 and not w25626;
w25634 <= not pi0609 and not w25546;
w25635 <= pi1155 and not w25634;
w25636 <= not w25633 and w25635;
w25637 <= pi0660 and not w25565;
w25638 <= not w25636 and w25637;
w25639 <= not w25632 and not w25638;
w25640 <= pi0785 and not w25639;
w25641 <= not pi0785 and not w25626;
w25642 <= not w25640 and not w25641;
w25643 <= not pi0618 and not w25642;
w25644 <= not pi1154 and not w25611;
w25645 <= not w25643 and w25644;
w25646 <= not pi0627 and not w25571;
w25647 <= not w25645 and w25646;
w25648 <= not pi0618 and w25547;
w25649 <= pi0618 and not w25642;
w25650 <= pi1154 and not w25648;
w25651 <= not w25649 and w25650;
w25652 <= pi0627 and not w25573;
w25653 <= not w25651 and w25652;
w25654 <= not w25647 and not w25653;
w25655 <= pi0781 and not w25654;
w25656 <= not pi0781 and not w25642;
w25657 <= not w25655 and not w25656;
w25658 <= not pi0789 and w25657;
w25659 <= not pi0619 and not w25657;
w25660 <= pi0619 and w25548;
w25661 <= not pi1159 and not w25660;
w25662 <= not w25659 and w25661;
w25663 <= not pi0648 and not w25579;
w25664 <= not w25662 and w25663;
w25665 <= pi0619 and not w25657;
w25666 <= not pi0619 and w25548;
w25667 <= pi1159 and not w25666;
w25668 <= not w25665 and w25667;
w25669 <= pi0648 and not w25581;
w25670 <= not w25668 and w25669;
w25671 <= pi0789 and not w25664;
w25672 <= not w25670 and w25671;
w25673 <= w15533 and not w25658;
w25674 <= not w25672 and w25673;
w25675 <= not w25610 and not w25674;
w25676 <= not w17927 and not w25675;
w25677 <= w15417 and not w25587;
w25678 <= w18414 and w25550;
w25679 <= not w25677 and not w25678;
w25680 <= not pi0629 and not w25679;
w25681 <= w18418 and w25550;
w25682 <= w15416 and not w25587;
w25683 <= not w25681 and not w25682;
w25684 <= pi0629 and not w25683;
w25685 <= not w25680 and not w25684;
w25686 <= pi0792 and not w25685;
w25687 <= not w17769 and not w25686;
w25688 <= not w25676 and w25687;
w25689 <= not w25598 and not w25688;
w25690 <= not pi0790 and w25689;
w25691 <= not pi0787 and not w25551;
w25692 <= pi1157 and not w25594;
w25693 <= not w25555 and not w25692;
w25694 <= pi0787 and not w25693;
w25695 <= not w25691 and not w25694;
w25696 <= not pi0644 and w25695;
w25697 <= pi0644 and w25689;
w25698 <= pi0715 and not w25696;
w25699 <= not w25697 and w25698;
w25700 <= not w15367 and not w25590;
w25701 <= w15367 and w25535;
w25702 <= not w25700 and not w25701;
w25703 <= pi0644 and not w25702;
w25704 <= not pi0644 and w25535;
w25705 <= not pi0715 and not w25704;
w25706 <= not w25703 and w25705;
w25707 <= pi1160 and not w25706;
w25708 <= not w25699 and w25707;
w25709 <= not pi0644 and not w25702;
w25710 <= pi0644 and w25535;
w25711 <= pi0715 and not w25710;
w25712 <= not w25709 and w25711;
w25713 <= pi0644 and w25695;
w25714 <= not pi0644 and w25689;
w25715 <= not pi0715 and not w25713;
w25716 <= not w25714 and w25715;
w25717 <= not pi1160 and not w25712;
w25718 <= not w25716 and w25717;
w25719 <= not w25708 and not w25718;
w25720 <= pi0790 and not w25719;
w25721 <= pi0832 and not w25690;
w25722 <= not w25720 and w25721;
w25723 <= not pi0184 and not w4989;
w25724 <= not pi0184 and not w14622;
w25725 <= w14198 and not w25724;
w25726 <= not pi0737 and w134;
w25727 <= w25724 and not w25726;
w25728 <= not pi0184 and not w14204;
w25729 <= w14210 and not w25728;
w25730 <= pi0184 and not w15639;
w25731 <= not pi0038 and not w25730;
w25732 <= w134 and not w25731;
w25733 <= not pi0184 and w15635;
w25734 <= not w25732 and not w25733;
w25735 <= not pi0737 and not w25729;
w25736 <= not w25734 and w25735;
w25737 <= not w25727 and not w25736;
w25738 <= not pi0778 and w25737;
w25739 <= not pi0625 and w25724;
w25740 <= pi0625 and not w25737;
w25741 <= pi1153 and not w25739;
w25742 <= not w25740 and w25741;
w25743 <= pi0625 and w25724;
w25744 <= not pi0625 and not w25737;
w25745 <= not pi1153 and not w25743;
w25746 <= not w25744 and w25745;
w25747 <= not w25742 and not w25746;
w25748 <= pi0778 and not w25747;
w25749 <= not w25738 and not w25748;
w25750 <= not w14638 and not w25749;
w25751 <= w14638 and not w25724;
w25752 <= not w25750 and not w25751;
w25753 <= not w14202 and w25752;
w25754 <= w14202 and w25724;
w25755 <= not w25753 and not w25754;
w25756 <= not w14198 and w25755;
w25757 <= not w25725 and not w25756;
w25758 <= not w14194 and w25757;
w25759 <= w14194 and w25724;
w25760 <= not w25758 and not w25759;
w25761 <= not pi0792 and w25760;
w25762 <= pi0628 and not w25760;
w25763 <= not pi0628 and w25724;
w25764 <= pi1156 and not w25763;
w25765 <= not w25762 and w25764;
w25766 <= pi0628 and w25724;
w25767 <= not pi0628 and not w25760;
w25768 <= not pi1156 and not w25766;
w25769 <= not w25767 and w25768;
w25770 <= not w25765 and not w25769;
w25771 <= pi0792 and not w25770;
w25772 <= not w25761 and not w25771;
w25773 <= not pi0647 and not w25772;
w25774 <= pi0647 and not w25724;
w25775 <= not w25773 and not w25774;
w25776 <= not pi1157 and w25775;
w25777 <= pi0647 and not w25772;
w25778 <= not pi0647 and not w25724;
w25779 <= not w25777 and not w25778;
w25780 <= pi1157 and w25779;
w25781 <= not w25776 and not w25780;
w25782 <= pi0787 and not w25781;
w25783 <= not pi0787 and w25772;
w25784 <= not w25782 and not w25783;
w25785 <= not pi0644 and not w25784;
w25786 <= pi0715 and not w25785;
w25787 <= pi0184 and not w134;
w25788 <= not pi0777 and w14843;
w25789 <= not w25728 and not w25788;
w25790 <= pi0038 and not w25789;
w25791 <= not pi0184 and w14784;
w25792 <= pi0184 and not w14838;
w25793 <= not pi0777 and not w25792;
w25794 <= not w25791 and w25793;
w25795 <= not pi0184 and pi0777;
w25796 <= not w14611 and w25795;
w25797 <= not w25794 and not w25796;
w25798 <= not pi0038 and not w25797;
w25799 <= not w25790 and not w25798;
w25800 <= w134 and w25799;
w25801 <= not w25787 and not w25800;
w25802 <= not w14680 and not w25801;
w25803 <= w14680 and not w25724;
w25804 <= not w25802 and not w25803;
w25805 <= not pi0785 and not w25804;
w25806 <= not w14854 and not w25724;
w25807 <= pi0609 and w25802;
w25808 <= not w25806 and not w25807;
w25809 <= pi1155 and not w25808;
w25810 <= not w14859 and not w25724;
w25811 <= not pi0609 and w25802;
w25812 <= not w25810 and not w25811;
w25813 <= not pi1155 and not w25812;
w25814 <= not w25809 and not w25813;
w25815 <= pi0785 and not w25814;
w25816 <= not w25805 and not w25815;
w25817 <= not pi0781 and not w25816;
w25818 <= not pi0618 and w25724;
w25819 <= pi0618 and w25816;
w25820 <= pi1154 and not w25818;
w25821 <= not w25819 and w25820;
w25822 <= not pi0618 and w25816;
w25823 <= pi0618 and w25724;
w25824 <= not pi1154 and not w25823;
w25825 <= not w25822 and w25824;
w25826 <= not w25821 and not w25825;
w25827 <= pi0781 and not w25826;
w25828 <= not w25817 and not w25827;
w25829 <= not pi0789 and not w25828;
w25830 <= not pi0619 and w25724;
w25831 <= pi0619 and w25828;
w25832 <= pi1159 and not w25830;
w25833 <= not w25831 and w25832;
w25834 <= not pi0619 and w25828;
w25835 <= pi0619 and w25724;
w25836 <= not pi1159 and not w25835;
w25837 <= not w25834 and w25836;
w25838 <= not w25833 and not w25837;
w25839 <= pi0789 and not w25838;
w25840 <= not w25829 and not w25839;
w25841 <= not w15532 and w25840;
w25842 <= w15532 and w25724;
w25843 <= not w25841 and not w25842;
w25844 <= not w15342 and not w25843;
w25845 <= w15342 and w25724;
w25846 <= not w25844 and not w25845;
w25847 <= not w15367 and not w25846;
w25848 <= w15367 and w25724;
w25849 <= not w25847 and not w25848;
w25850 <= pi0644 and not w25849;
w25851 <= not pi0644 and w25724;
w25852 <= not pi0715 and not w25851;
w25853 <= not w25850 and w25852;
w25854 <= pi1160 and not w25853;
w25855 <= not w25786 and w25854;
w25856 <= pi0644 and not w25784;
w25857 <= not pi0715 and not w25856;
w25858 <= not pi0644 and not w25849;
w25859 <= pi0644 and w25724;
w25860 <= pi0715 and not w25859;
w25861 <= not w25858 and w25860;
w25862 <= not pi1160 and not w25861;
w25863 <= not w25857 and w25862;
w25864 <= not w25855 and not w25863;
w25865 <= pi0790 and not w25864;
w25866 <= not pi0629 and w25765;
w25867 <= not w18133 and w25843;
w25868 <= pi0629 and w25769;
w25869 <= not w25866 and not w25868;
w25870 <= not w25867 and w25869;
w25871 <= pi0792 and not w25870;
w25872 <= pi0609 and w25749;
w25873 <= pi0184 and not w15188;
w25874 <= not pi0184 and not w15175;
w25875 <= pi0777 and not w25873;
w25876 <= not w25874 and w25875;
w25877 <= not pi0184 and w15192;
w25878 <= pi0184 and w15194;
w25879 <= not pi0777 and not w25878;
w25880 <= not w25877 and w25879;
w25881 <= not w25876 and not w25880;
w25882 <= not pi0039 and not w25881;
w25883 <= pi0184 and w15168;
w25884 <= not pi0184 and not w15109;
w25885 <= not pi0777 and not w25884;
w25886 <= not w25883 and w25885;
w25887 <= not pi0184 and w14967;
w25888 <= pi0184 and w15048;
w25889 <= pi0777 and not w25888;
w25890 <= not w25887 and w25889;
w25891 <= pi0039 and not w25886;
w25892 <= not w25890 and w25891;
w25893 <= not pi0038 and not w25882;
w25894 <= not w25892 and w25893;
w25895 <= not pi0777 and not w15053;
w25896 <= w17034 and not w25895;
w25897 <= not pi0184 and not w25896;
w25898 <= not w15032 and not w25557;
w25899 <= pi0184 and not w25898;
w25900 <= w3847 and w25899;
w25901 <= pi0038 and not w25900;
w25902 <= not w25897 and w25901;
w25903 <= not pi0737 and not w25902;
w25904 <= not w25894 and w25903;
w25905 <= pi0737 and not w25799;
w25906 <= w134 and not w25904;
w25907 <= not w25905 and w25906;
w25908 <= not w25787 and not w25907;
w25909 <= not pi0625 and w25908;
w25910 <= pi0625 and w25801;
w25911 <= not pi1153 and not w25910;
w25912 <= not w25909 and w25911;
w25913 <= not pi0608 and not w25742;
w25914 <= not w25912 and w25913;
w25915 <= not pi0625 and w25801;
w25916 <= pi0625 and w25908;
w25917 <= pi1153 and not w25915;
w25918 <= not w25916 and w25917;
w25919 <= pi0608 and not w25746;
w25920 <= not w25918 and w25919;
w25921 <= not w25914 and not w25920;
w25922 <= pi0778 and not w25921;
w25923 <= not pi0778 and w25908;
w25924 <= not w25922 and not w25923;
w25925 <= not pi0609 and not w25924;
w25926 <= not pi1155 and not w25872;
w25927 <= not w25925 and w25926;
w25928 <= not pi0660 and not w25809;
w25929 <= not w25927 and w25928;
w25930 <= not pi0609 and w25749;
w25931 <= pi0609 and not w25924;
w25932 <= pi1155 and not w25930;
w25933 <= not w25931 and w25932;
w25934 <= pi0660 and not w25813;
w25935 <= not w25933 and w25934;
w25936 <= not w25929 and not w25935;
w25937 <= pi0785 and not w25936;
w25938 <= not pi0785 and not w25924;
w25939 <= not w25937 and not w25938;
w25940 <= not pi0618 and not w25939;
w25941 <= pi0618 and w25752;
w25942 <= not pi1154 and not w25941;
w25943 <= not w25940 and w25942;
w25944 <= not pi0627 and not w25821;
w25945 <= not w25943 and w25944;
w25946 <= not pi0618 and w25752;
w25947 <= pi0618 and not w25939;
w25948 <= pi1154 and not w25946;
w25949 <= not w25947 and w25948;
w25950 <= pi0627 and not w25825;
w25951 <= not w25949 and w25950;
w25952 <= not w25945 and not w25951;
w25953 <= pi0781 and not w25952;
w25954 <= not pi0781 and not w25939;
w25955 <= not w25953 and not w25954;
w25956 <= not pi0789 and w25955;
w25957 <= pi0619 and not w25755;
w25958 <= not pi0619 and not w25955;
w25959 <= not pi1159 and not w25957;
w25960 <= not w25958 and w25959;
w25961 <= not pi0648 and not w25833;
w25962 <= not w25960 and w25961;
w25963 <= not pi0619 and not w25755;
w25964 <= pi0619 and not w25955;
w25965 <= pi1159 and not w25963;
w25966 <= not w25964 and w25965;
w25967 <= pi0648 and not w25837;
w25968 <= not w25966 and w25967;
w25969 <= pi0789 and not w25962;
w25970 <= not w25968 and w25969;
w25971 <= w15533 and not w25956;
w25972 <= not w25970 and w25971;
w25973 <= w15434 and w25757;
w25974 <= not pi0626 and not w25840;
w25975 <= pi0626 and not w25724;
w25976 <= w14192 and not w25975;
w25977 <= not w25974 and w25976;
w25978 <= pi0626 and not w25840;
w25979 <= not pi0626 and not w25724;
w25980 <= w14191 and not w25979;
w25981 <= not w25978 and w25980;
w25982 <= not w25973 and not w25977;
w25983 <= not w25981 and w25982;
w25984 <= pi0788 and not w25983;
w25985 <= not w17927 and not w25984;
w25986 <= not w25972 and w25985;
w25987 <= not w25871 and not w25986;
w25988 <= not w17769 and not w25987;
w25989 <= w15365 and not w25775;
w25990 <= not w18122 and w25846;
w25991 <= w15364 and not w25779;
w25992 <= not w25989 and not w25991;
w25993 <= not w25990 and w25992;
w25994 <= pi0787 and not w25993;
w25995 <= not pi0644 and w25862;
w25996 <= pi0644 and w25854;
w25997 <= pi0790 and not w25995;
w25998 <= not w25996 and w25997;
w25999 <= not w25988 and not w25994;
w26000 <= not w25998 and w25999;
w26001 <= not w25865 and not w26000;
w26002 <= w4989 and not w26001;
w26003 <= not pi0832 and not w25723;
w26004 <= not w26002 and w26003;
w26005 <= not w25722 and not w26004;
w26006 <= not pi0185 and not w489;
w26007 <= not pi0701 and w14208;
w26008 <= not w26006 and not w26007;
w26009 <= not pi0778 and not w26008;
w26010 <= not pi0625 and w26007;
w26011 <= not w26008 and not w26010;
w26012 <= pi1153 and not w26011;
w26013 <= not pi1153 and not w26006;
w26014 <= not w26010 and w26013;
w26015 <= pi0778 and not w26014;
w26016 <= not w26012 and w26015;
w26017 <= not w26009 and not w26016;
w26018 <= not w15408 and not w26017;
w26019 <= not w15410 and w26018;
w26020 <= not w15412 and w26019;
w26021 <= not w15414 and w26020;
w26022 <= not w15420 and w26021;
w26023 <= not pi0647 and w26022;
w26024 <= pi0647 and w26006;
w26025 <= not pi1157 and not w26024;
w26026 <= not w26023 and w26025;
w26027 <= pi0630 and w26026;
w26028 <= not pi0751 and w14807;
w26029 <= not w26006 and not w26028;
w26030 <= not w15437 and not w26029;
w26031 <= not pi0785 and not w26030;
w26032 <= w14859 and w26028;
w26033 <= w26030 and not w26032;
w26034 <= pi1155 and not w26033;
w26035 <= not pi1155 and not w26006;
w26036 <= not w26032 and w26035;
w26037 <= not w26034 and not w26036;
w26038 <= pi0785 and not w26037;
w26039 <= not w26031 and not w26038;
w26040 <= not pi0781 and not w26039;
w26041 <= not w15452 and w26039;
w26042 <= pi1154 and not w26041;
w26043 <= not w15455 and w26039;
w26044 <= not pi1154 and not w26043;
w26045 <= not w26042 and not w26044;
w26046 <= pi0781 and not w26045;
w26047 <= not w26040 and not w26046;
w26048 <= not pi0789 and not w26047;
w26049 <= not w20641 and w26047;
w26050 <= pi1159 and not w26049;
w26051 <= not w20644 and w26047;
w26052 <= not pi1159 and not w26051;
w26053 <= not w26050 and not w26052;
w26054 <= pi0789 and not w26053;
w26055 <= not w26048 and not w26054;
w26056 <= not w15532 and w26055;
w26057 <= w15532 and w26006;
w26058 <= not w26056 and not w26057;
w26059 <= not w15342 and not w26058;
w26060 <= w15342 and w26006;
w26061 <= not w26059 and not w26060;
w26062 <= not w18122 and w26061;
w26063 <= pi0647 and not w26022;
w26064 <= not pi0647 and not w26006;
w26065 <= not w26063 and not w26064;
w26066 <= w15364 and not w26065;
w26067 <= not w26027 and not w26066;
w26068 <= not w26062 and w26067;
w26069 <= pi0787 and not w26068;
w26070 <= w15434 and w26020;
w26071 <= not pi0626 and not w26055;
w26072 <= pi0626 and not w26006;
w26073 <= w14192 and not w26072;
w26074 <= not w26071 and w26073;
w26075 <= pi0626 and not w26055;
w26076 <= not pi0626 and not w26006;
w26077 <= w14191 and not w26076;
w26078 <= not w26075 and w26077;
w26079 <= not w26070 and not w26074;
w26080 <= not w26078 and w26079;
w26081 <= pi0788 and not w26080;
w26082 <= pi0618 and w26018;
w26083 <= not w14731 and not w26008;
w26084 <= pi0625 and w26083;
w26085 <= w26029 and not w26083;
w26086 <= not w26084 and not w26085;
w26087 <= w26013 and not w26086;
w26088 <= not pi0608 and not w26012;
w26089 <= not w26087 and w26088;
w26090 <= pi1153 and w26029;
w26091 <= not w26084 and w26090;
w26092 <= pi0608 and not w26014;
w26093 <= not w26091 and w26092;
w26094 <= not w26089 and not w26093;
w26095 <= pi0778 and not w26094;
w26096 <= not pi0778 and not w26085;
w26097 <= not w26095 and not w26096;
w26098 <= not pi0609 and not w26097;
w26099 <= pi0609 and not w26017;
w26100 <= not pi1155 and not w26099;
w26101 <= not w26098 and w26100;
w26102 <= not pi0660 and not w26034;
w26103 <= not w26101 and w26102;
w26104 <= pi0609 and not w26097;
w26105 <= not pi0609 and not w26017;
w26106 <= pi1155 and not w26105;
w26107 <= not w26104 and w26106;
w26108 <= pi0660 and not w26036;
w26109 <= not w26107 and w26108;
w26110 <= not w26103 and not w26109;
w26111 <= pi0785 and not w26110;
w26112 <= not pi0785 and not w26097;
w26113 <= not w26111 and not w26112;
w26114 <= not pi0618 and not w26113;
w26115 <= not pi1154 and not w26082;
w26116 <= not w26114 and w26115;
w26117 <= not pi0627 and not w26042;
w26118 <= not w26116 and w26117;
w26119 <= not pi0618 and w26018;
w26120 <= pi0618 and not w26113;
w26121 <= pi1154 and not w26119;
w26122 <= not w26120 and w26121;
w26123 <= pi0627 and not w26044;
w26124 <= not w26122 and w26123;
w26125 <= not w26118 and not w26124;
w26126 <= pi0781 and not w26125;
w26127 <= not pi0781 and not w26113;
w26128 <= not w26126 and not w26127;
w26129 <= not pi0789 and w26128;
w26130 <= not pi0619 and not w26128;
w26131 <= pi0619 and w26019;
w26132 <= not pi1159 and not w26131;
w26133 <= not w26130 and w26132;
w26134 <= not pi0648 and not w26050;
w26135 <= not w26133 and w26134;
w26136 <= pi0619 and not w26128;
w26137 <= not pi0619 and w26019;
w26138 <= pi1159 and not w26137;
w26139 <= not w26136 and w26138;
w26140 <= pi0648 and not w26052;
w26141 <= not w26139 and w26140;
w26142 <= pi0789 and not w26135;
w26143 <= not w26141 and w26142;
w26144 <= w15533 and not w26129;
w26145 <= not w26143 and w26144;
w26146 <= not w26081 and not w26145;
w26147 <= not w17927 and not w26146;
w26148 <= w15417 and not w26058;
w26149 <= w18414 and w26021;
w26150 <= not w26148 and not w26149;
w26151 <= not pi0629 and not w26150;
w26152 <= w18418 and w26021;
w26153 <= w15416 and not w26058;
w26154 <= not w26152 and not w26153;
w26155 <= pi0629 and not w26154;
w26156 <= not w26151 and not w26155;
w26157 <= pi0792 and not w26156;
w26158 <= not w17769 and not w26157;
w26159 <= not w26147 and w26158;
w26160 <= not w26069 and not w26159;
w26161 <= not pi0790 and w26160;
w26162 <= not pi0787 and not w26022;
w26163 <= pi1157 and not w26065;
w26164 <= not w26026 and not w26163;
w26165 <= pi0787 and not w26164;
w26166 <= not w26162 and not w26165;
w26167 <= not pi0644 and w26166;
w26168 <= pi0644 and w26160;
w26169 <= pi0715 and not w26167;
w26170 <= not w26168 and w26169;
w26171 <= not w15367 and not w26061;
w26172 <= w15367 and w26006;
w26173 <= not w26171 and not w26172;
w26174 <= pi0644 and not w26173;
w26175 <= not pi0644 and w26006;
w26176 <= not pi0715 and not w26175;
w26177 <= not w26174 and w26176;
w26178 <= pi1160 and not w26177;
w26179 <= not w26170 and w26178;
w26180 <= not pi0644 and not w26173;
w26181 <= pi0644 and w26006;
w26182 <= pi0715 and not w26181;
w26183 <= not w26180 and w26182;
w26184 <= pi0644 and w26166;
w26185 <= not pi0644 and w26160;
w26186 <= not pi0715 and not w26184;
w26187 <= not w26185 and w26186;
w26188 <= not pi1160 and not w26183;
w26189 <= not w26187 and w26188;
w26190 <= not w26179 and not w26189;
w26191 <= pi0790 and not w26190;
w26192 <= pi0832 and not w26161;
w26193 <= not w26191 and w26192;
w26194 <= not pi0185 and not w4989;
w26195 <= not pi0185 and not w14622;
w26196 <= w14198 and not w26195;
w26197 <= not pi0701 and w134;
w26198 <= w26195 and not w26197;
w26199 <= not pi0185 and not w14204;
w26200 <= w14210 and not w26199;
w26201 <= pi0185 and not w15639;
w26202 <= not pi0038 and not w26201;
w26203 <= w134 and not w26202;
w26204 <= not pi0185 and w15635;
w26205 <= not w26203 and not w26204;
w26206 <= not pi0701 and not w26200;
w26207 <= not w26205 and w26206;
w26208 <= not w26198 and not w26207;
w26209 <= not pi0778 and w26208;
w26210 <= not pi0625 and w26195;
w26211 <= pi0625 and not w26208;
w26212 <= pi1153 and not w26210;
w26213 <= not w26211 and w26212;
w26214 <= pi0625 and w26195;
w26215 <= not pi0625 and not w26208;
w26216 <= not pi1153 and not w26214;
w26217 <= not w26215 and w26216;
w26218 <= not w26213 and not w26217;
w26219 <= pi0778 and not w26218;
w26220 <= not w26209 and not w26219;
w26221 <= not w14638 and not w26220;
w26222 <= w14638 and not w26195;
w26223 <= not w26221 and not w26222;
w26224 <= not w14202 and w26223;
w26225 <= w14202 and w26195;
w26226 <= not w26224 and not w26225;
w26227 <= not w14198 and w26226;
w26228 <= not w26196 and not w26227;
w26229 <= not w14194 and w26228;
w26230 <= w14194 and w26195;
w26231 <= not w26229 and not w26230;
w26232 <= not pi0792 and w26231;
w26233 <= pi0628 and not w26231;
w26234 <= not pi0628 and w26195;
w26235 <= pi1156 and not w26234;
w26236 <= not w26233 and w26235;
w26237 <= pi0628 and w26195;
w26238 <= not pi0628 and not w26231;
w26239 <= not pi1156 and not w26237;
w26240 <= not w26238 and w26239;
w26241 <= not w26236 and not w26240;
w26242 <= pi0792 and not w26241;
w26243 <= not w26232 and not w26242;
w26244 <= not pi0647 and not w26243;
w26245 <= pi0647 and not w26195;
w26246 <= not w26244 and not w26245;
w26247 <= not pi1157 and w26246;
w26248 <= pi0647 and not w26243;
w26249 <= not pi0647 and not w26195;
w26250 <= not w26248 and not w26249;
w26251 <= pi1157 and w26250;
w26252 <= not w26247 and not w26251;
w26253 <= pi0787 and not w26252;
w26254 <= not pi0787 and w26243;
w26255 <= not w26253 and not w26254;
w26256 <= not pi0644 and not w26255;
w26257 <= pi0715 and not w26256;
w26258 <= pi0185 and not w134;
w26259 <= pi0185 and pi0751;
w26260 <= pi0751 and w14609;
w26261 <= pi0185 and w14836;
w26262 <= not w26260 and not w26261;
w26263 <= pi0039 and not w26262;
w26264 <= pi0185 and not w14796;
w26265 <= not w18822 and not w26264;
w26266 <= not pi0039 and not w26265;
w26267 <= not pi0185 and not pi0751;
w26268 <= w14784 and w26267;
w26269 <= not w26259 and not w26266;
w26270 <= not w26268 and w26269;
w26271 <= not w26263 and w26270;
w26272 <= not pi0038 and not w26271;
w26273 <= not pi0751 and w14843;
w26274 <= pi0038 and not w26199;
w26275 <= not w26273 and w26274;
w26276 <= not w26272 and not w26275;
w26277 <= w134 and not w26276;
w26278 <= not w26258 and not w26277;
w26279 <= not w14680 and not w26278;
w26280 <= w14680 and not w26195;
w26281 <= not w26279 and not w26280;
w26282 <= not pi0785 and not w26281;
w26283 <= not w14854 and not w26195;
w26284 <= pi0609 and w26279;
w26285 <= not w26283 and not w26284;
w26286 <= pi1155 and not w26285;
w26287 <= not w14859 and not w26195;
w26288 <= not pi0609 and w26279;
w26289 <= not w26287 and not w26288;
w26290 <= not pi1155 and not w26289;
w26291 <= not w26286 and not w26290;
w26292 <= pi0785 and not w26291;
w26293 <= not w26282 and not w26292;
w26294 <= not pi0781 and not w26293;
w26295 <= not pi0618 and w26195;
w26296 <= pi0618 and w26293;
w26297 <= pi1154 and not w26295;
w26298 <= not w26296 and w26297;
w26299 <= not pi0618 and w26293;
w26300 <= pi0618 and w26195;
w26301 <= not pi1154 and not w26300;
w26302 <= not w26299 and w26301;
w26303 <= not w26298 and not w26302;
w26304 <= pi0781 and not w26303;
w26305 <= not w26294 and not w26304;
w26306 <= not pi0789 and not w26305;
w26307 <= not pi0619 and w26195;
w26308 <= pi0619 and w26305;
w26309 <= pi1159 and not w26307;
w26310 <= not w26308 and w26309;
w26311 <= not pi0619 and w26305;
w26312 <= pi0619 and w26195;
w26313 <= not pi1159 and not w26312;
w26314 <= not w26311 and w26313;
w26315 <= not w26310 and not w26314;
w26316 <= pi0789 and not w26315;
w26317 <= not w26306 and not w26316;
w26318 <= not w15532 and w26317;
w26319 <= w15532 and w26195;
w26320 <= not w26318 and not w26319;
w26321 <= not w15342 and not w26320;
w26322 <= w15342 and w26195;
w26323 <= not w26321 and not w26322;
w26324 <= not w15367 and not w26323;
w26325 <= w15367 and w26195;
w26326 <= not w26324 and not w26325;
w26327 <= pi0644 and not w26326;
w26328 <= not pi0644 and w26195;
w26329 <= not pi0715 and not w26328;
w26330 <= not w26327 and w26329;
w26331 <= pi1160 and not w26330;
w26332 <= not w26257 and w26331;
w26333 <= pi0644 and not w26255;
w26334 <= not pi0715 and not w26333;
w26335 <= not pi0644 and not w26326;
w26336 <= pi0644 and w26195;
w26337 <= pi0715 and not w26336;
w26338 <= not w26335 and w26337;
w26339 <= not pi1160 and not w26338;
w26340 <= not w26334 and w26339;
w26341 <= not w26332 and not w26340;
w26342 <= pi0790 and not w26341;
w26343 <= not pi0629 and w26236;
w26344 <= not w18133 and w26320;
w26345 <= pi0629 and w26240;
w26346 <= not w26343 and not w26345;
w26347 <= not w26344 and w26346;
w26348 <= pi0792 and not w26347;
w26349 <= pi0609 and w26220;
w26350 <= pi0185 and not w15188;
w26351 <= not pi0185 and not w15175;
w26352 <= pi0751 and not w26350;
w26353 <= not w26351 and w26352;
w26354 <= not pi0185 and w15192;
w26355 <= pi0185 and w15194;
w26356 <= not pi0751 and not w26355;
w26357 <= not w26354 and w26356;
w26358 <= not w26353 and not w26357;
w26359 <= not pi0039 and not w26358;
w26360 <= pi0185 and w15168;
w26361 <= not pi0185 and not w15109;
w26362 <= not pi0751 and not w26361;
w26363 <= not w26360 and w26362;
w26364 <= not pi0185 and w14967;
w26365 <= pi0185 and w15048;
w26366 <= pi0751 and not w26365;
w26367 <= not w26364 and w26366;
w26368 <= pi0039 and not w26363;
w26369 <= not w26367 and w26368;
w26370 <= not pi0038 and not w26359;
w26371 <= not w26369 and w26370;
w26372 <= not w15032 and not w26028;
w26373 <= pi0185 and not w26372;
w26374 <= w3847 and w26373;
w26375 <= not pi0751 and not w15053;
w26376 <= w17034 and not w26375;
w26377 <= not pi0185 and not w26376;
w26378 <= pi0038 and not w26374;
w26379 <= not w26377 and w26378;
w26380 <= not pi0701 and not w26379;
w26381 <= not w26371 and w26380;
w26382 <= pi0701 and w26276;
w26383 <= w134 and not w26381;
w26384 <= not w26382 and w26383;
w26385 <= not w26258 and not w26384;
w26386 <= not pi0625 and w26385;
w26387 <= pi0625 and w26278;
w26388 <= not pi1153 and not w26387;
w26389 <= not w26386 and w26388;
w26390 <= not pi0608 and not w26213;
w26391 <= not w26389 and w26390;
w26392 <= not pi0625 and w26278;
w26393 <= pi0625 and w26385;
w26394 <= pi1153 and not w26392;
w26395 <= not w26393 and w26394;
w26396 <= pi0608 and not w26217;
w26397 <= not w26395 and w26396;
w26398 <= not w26391 and not w26397;
w26399 <= pi0778 and not w26398;
w26400 <= not pi0778 and w26385;
w26401 <= not w26399 and not w26400;
w26402 <= not pi0609 and not w26401;
w26403 <= not pi1155 and not w26349;
w26404 <= not w26402 and w26403;
w26405 <= not pi0660 and not w26286;
w26406 <= not w26404 and w26405;
w26407 <= not pi0609 and w26220;
w26408 <= pi0609 and not w26401;
w26409 <= pi1155 and not w26407;
w26410 <= not w26408 and w26409;
w26411 <= pi0660 and not w26290;
w26412 <= not w26410 and w26411;
w26413 <= not w26406 and not w26412;
w26414 <= pi0785 and not w26413;
w26415 <= not pi0785 and not w26401;
w26416 <= not w26414 and not w26415;
w26417 <= not pi0618 and not w26416;
w26418 <= pi0618 and w26223;
w26419 <= not pi1154 and not w26418;
w26420 <= not w26417 and w26419;
w26421 <= not pi0627 and not w26298;
w26422 <= not w26420 and w26421;
w26423 <= not pi0618 and w26223;
w26424 <= pi0618 and not w26416;
w26425 <= pi1154 and not w26423;
w26426 <= not w26424 and w26425;
w26427 <= pi0627 and not w26302;
w26428 <= not w26426 and w26427;
w26429 <= not w26422 and not w26428;
w26430 <= pi0781 and not w26429;
w26431 <= not pi0781 and not w26416;
w26432 <= not w26430 and not w26431;
w26433 <= not pi0789 and w26432;
w26434 <= pi0619 and not w26226;
w26435 <= not pi0619 and not w26432;
w26436 <= not pi1159 and not w26434;
w26437 <= not w26435 and w26436;
w26438 <= not pi0648 and not w26310;
w26439 <= not w26437 and w26438;
w26440 <= not pi0619 and not w26226;
w26441 <= pi0619 and not w26432;
w26442 <= pi1159 and not w26440;
w26443 <= not w26441 and w26442;
w26444 <= pi0648 and not w26314;
w26445 <= not w26443 and w26444;
w26446 <= pi0789 and not w26439;
w26447 <= not w26445 and w26446;
w26448 <= w15533 and not w26433;
w26449 <= not w26447 and w26448;
w26450 <= w15434 and w26228;
w26451 <= not pi0626 and not w26317;
w26452 <= pi0626 and not w26195;
w26453 <= w14192 and not w26452;
w26454 <= not w26451 and w26453;
w26455 <= pi0626 and not w26317;
w26456 <= not pi0626 and not w26195;
w26457 <= w14191 and not w26456;
w26458 <= not w26455 and w26457;
w26459 <= not w26450 and not w26454;
w26460 <= not w26458 and w26459;
w26461 <= pi0788 and not w26460;
w26462 <= not w17927 and not w26461;
w26463 <= not w26449 and w26462;
w26464 <= not w26348 and not w26463;
w26465 <= not w17769 and not w26464;
w26466 <= w15365 and not w26246;
w26467 <= not w18122 and w26323;
w26468 <= w15364 and not w26250;
w26469 <= not w26466 and not w26468;
w26470 <= not w26467 and w26469;
w26471 <= pi0787 and not w26470;
w26472 <= not pi0644 and w26339;
w26473 <= pi0644 and w26331;
w26474 <= pi0790 and not w26472;
w26475 <= not w26473 and w26474;
w26476 <= not w26465 and not w26471;
w26477 <= not w26475 and w26476;
w26478 <= not w26342 and not w26477;
w26479 <= w4989 and not w26478;
w26480 <= not pi0832 and not w26194;
w26481 <= not w26479 and w26480;
w26482 <= not w26193 and not w26481;
w26483 <= not pi0186 and not w14622;
w26484 <= w14198 and not w26483;
w26485 <= pi0186 and not w134;
w26486 <= not pi0186 and not w14615;
w26487 <= not pi0703 and w26486;
w26488 <= not pi0186 and not w14204;
w26489 <= w14210 and not w26488;
w26490 <= not pi0186 and w15635;
w26491 <= pi0186 and not w15639;
w26492 <= not pi0038 and not w26491;
w26493 <= not w26490 and w26492;
w26494 <= pi0703 and not w26489;
w26495 <= not w26493 and w26494;
w26496 <= w134 and not w26487;
w26497 <= not w26495 and w26496;
w26498 <= not w26485 and not w26497;
w26499 <= not pi0778 and not w26498;
w26500 <= not pi0625 and w26483;
w26501 <= pi0625 and w26498;
w26502 <= pi1153 and not w26500;
w26503 <= not w26501 and w26502;
w26504 <= not pi0625 and w26498;
w26505 <= pi0625 and w26483;
w26506 <= not pi1153 and not w26505;
w26507 <= not w26504 and w26506;
w26508 <= not w26503 and not w26507;
w26509 <= pi0778 and not w26508;
w26510 <= not w26499 and not w26509;
w26511 <= not w14638 and not w26510;
w26512 <= w14638 and not w26483;
w26513 <= not w26511 and not w26512;
w26514 <= not w14202 and w26513;
w26515 <= w14202 and w26483;
w26516 <= not w26514 and not w26515;
w26517 <= not w14198 and w26516;
w26518 <= not w26484 and not w26517;
w26519 <= not w14194 and w26518;
w26520 <= w14194 and w26483;
w26521 <= not w26519 and not w26520;
w26522 <= not pi0792 and w26521;
w26523 <= not pi0628 and w26483;
w26524 <= pi0628 and not w26521;
w26525 <= pi1156 and not w26523;
w26526 <= not w26524 and w26525;
w26527 <= pi0628 and w26483;
w26528 <= not pi0628 and not w26521;
w26529 <= not pi1156 and not w26527;
w26530 <= not w26528 and w26529;
w26531 <= not w26526 and not w26530;
w26532 <= pi0792 and not w26531;
w26533 <= not w26522 and not w26532;
w26534 <= not pi0787 and not w26533;
w26535 <= not pi0647 and w26483;
w26536 <= pi0647 and w26533;
w26537 <= pi1157 and not w26535;
w26538 <= not w26536 and w26537;
w26539 <= not pi0647 and w26533;
w26540 <= pi0647 and w26483;
w26541 <= not pi1157 and not w26540;
w26542 <= not w26539 and w26541;
w26543 <= not w26538 and not w26542;
w26544 <= pi0787 and not w26543;
w26545 <= not w26534 and not w26544;
w26546 <= not pi0644 and w26545;
w26547 <= not pi0618 and w26483;
w26548 <= pi0752 and not w26486;
w26549 <= pi0186 and not w16997;
w26550 <= not pi0186 and not pi0752;
w26551 <= w17002 and w26550;
w26552 <= not w26549 and not w26551;
w26553 <= not w16996 and not w26552;
w26554 <= not w26548 and not w26553;
w26555 <= w134 and not w26554;
w26556 <= not w26485 and not w26555;
w26557 <= not w14680 and not w26556;
w26558 <= w14680 and not w26483;
w26559 <= not w26557 and not w26558;
w26560 <= not pi0785 and not w26559;
w26561 <= not w14854 and not w26483;
w26562 <= pi0609 and w26557;
w26563 <= not w26561 and not w26562;
w26564 <= pi1155 and not w26563;
w26565 <= not w14859 and not w26483;
w26566 <= not pi0609 and w26557;
w26567 <= not w26565 and not w26566;
w26568 <= not pi1155 and not w26567;
w26569 <= not w26564 and not w26568;
w26570 <= pi0785 and not w26569;
w26571 <= not w26560 and not w26570;
w26572 <= pi0618 and w26571;
w26573 <= pi1154 and not w26547;
w26574 <= not w26572 and w26573;
w26575 <= pi0186 and w17031;
w26576 <= not pi0186 and w17040;
w26577 <= pi0752 and not w17033;
w26578 <= not w26575 and w26577;
w26579 <= not w26576 and w26578;
w26580 <= not pi0186 and not w17051;
w26581 <= pi0186 and w17059;
w26582 <= not pi0752 and not w26580;
w26583 <= not w26581 and w26582;
w26584 <= pi0703 and not w26583;
w26585 <= not w26579 and w26584;
w26586 <= not pi0703 and w26554;
w26587 <= w134 and not w26585;
w26588 <= not w26586 and w26587;
w26589 <= not w26485 and not w26588;
w26590 <= not pi0625 and w26589;
w26591 <= pi0625 and w26556;
w26592 <= not pi1153 and not w26591;
w26593 <= not w26590 and w26592;
w26594 <= not pi0608 and not w26503;
w26595 <= not w26593 and w26594;
w26596 <= not pi0625 and w26556;
w26597 <= pi0625 and w26589;
w26598 <= pi1153 and not w26596;
w26599 <= not w26597 and w26598;
w26600 <= pi0608 and not w26507;
w26601 <= not w26599 and w26600;
w26602 <= not w26595 and not w26601;
w26603 <= pi0778 and not w26602;
w26604 <= not pi0778 and w26589;
w26605 <= not w26603 and not w26604;
w26606 <= not pi0609 and not w26605;
w26607 <= pi0609 and w26510;
w26608 <= not pi1155 and not w26607;
w26609 <= not w26606 and w26608;
w26610 <= not pi0660 and not w26564;
w26611 <= not w26609 and w26610;
w26612 <= not pi0609 and w26510;
w26613 <= pi0609 and not w26605;
w26614 <= pi1155 and not w26612;
w26615 <= not w26613 and w26614;
w26616 <= pi0660 and not w26568;
w26617 <= not w26615 and w26616;
w26618 <= not w26611 and not w26617;
w26619 <= pi0785 and not w26618;
w26620 <= not pi0785 and not w26605;
w26621 <= not w26619 and not w26620;
w26622 <= not pi0618 and not w26621;
w26623 <= pi0618 and w26513;
w26624 <= not pi1154 and not w26623;
w26625 <= not w26622 and w26624;
w26626 <= not pi0627 and not w26574;
w26627 <= not w26625 and w26626;
w26628 <= not pi0618 and w26571;
w26629 <= pi0618 and w26483;
w26630 <= not pi1154 and not w26629;
w26631 <= not w26628 and w26630;
w26632 <= not pi0618 and w26513;
w26633 <= pi0618 and not w26621;
w26634 <= pi1154 and not w26632;
w26635 <= not w26633 and w26634;
w26636 <= pi0627 and not w26631;
w26637 <= not w26635 and w26636;
w26638 <= not w26627 and not w26637;
w26639 <= pi0781 and not w26638;
w26640 <= not pi0781 and not w26621;
w26641 <= not w26639 and not w26640;
w26642 <= not pi0619 and not w26641;
w26643 <= pi0619 and not w26516;
w26644 <= not pi1159 and not w26643;
w26645 <= not w26642 and w26644;
w26646 <= not pi0619 and w26483;
w26647 <= not pi0781 and not w26571;
w26648 <= not w26574 and not w26631;
w26649 <= pi0781 and not w26648;
w26650 <= not w26647 and not w26649;
w26651 <= pi0619 and w26650;
w26652 <= pi1159 and not w26646;
w26653 <= not w26651 and w26652;
w26654 <= not pi0648 and not w26653;
w26655 <= not w26645 and w26654;
w26656 <= pi0619 and not w26641;
w26657 <= not pi0619 and not w26516;
w26658 <= pi1159 and not w26657;
w26659 <= not w26656 and w26658;
w26660 <= not pi0619 and w26650;
w26661 <= pi0619 and w26483;
w26662 <= not pi1159 and not w26661;
w26663 <= not w26660 and w26662;
w26664 <= pi0648 and not w26663;
w26665 <= not w26659 and w26664;
w26666 <= not w26655 and not w26665;
w26667 <= pi0789 and not w26666;
w26668 <= not pi0789 and not w26641;
w26669 <= not w26667 and not w26668;
w26670 <= not pi0788 and w26669;
w26671 <= not pi0626 and w26669;
w26672 <= pi0626 and not w26518;
w26673 <= not pi0641 and not w26672;
w26674 <= not w26671 and w26673;
w26675 <= not pi0789 and not w26650;
w26676 <= not w26653 and not w26663;
w26677 <= pi0789 and not w26676;
w26678 <= not w26675 and not w26677;
w26679 <= not pi0626 and not w26678;
w26680 <= pi0626 and not w26483;
w26681 <= pi0641 and not w26680;
w26682 <= not w26679 and w26681;
w26683 <= not pi1158 and not w26682;
w26684 <= not w26674 and w26683;
w26685 <= pi0626 and w26669;
w26686 <= not pi0626 and not w26518;
w26687 <= pi0641 and not w26686;
w26688 <= not w26685 and w26687;
w26689 <= pi0626 and not w26678;
w26690 <= not pi0626 and not w26483;
w26691 <= not pi0641 and not w26690;
w26692 <= not w26689 and w26691;
w26693 <= pi1158 and not w26692;
w26694 <= not w26688 and w26693;
w26695 <= not w26684 and not w26694;
w26696 <= pi0788 and not w26695;
w26697 <= not w26670 and not w26696;
w26698 <= not pi0628 and w26697;
w26699 <= not w15532 and w26678;
w26700 <= w15532 and w26483;
w26701 <= not w26699 and not w26700;
w26702 <= pi0628 and not w26701;
w26703 <= not pi1156 and not w26702;
w26704 <= not w26698 and w26703;
w26705 <= not pi0629 and not w26526;
w26706 <= not w26704 and w26705;
w26707 <= pi0628 and w26697;
w26708 <= not pi0628 and not w26701;
w26709 <= pi1156 and not w26708;
w26710 <= not w26707 and w26709;
w26711 <= pi0629 and not w26530;
w26712 <= not w26710 and w26711;
w26713 <= not w26706 and not w26712;
w26714 <= pi0792 and not w26713;
w26715 <= not pi0792 and w26697;
w26716 <= not w26714 and not w26715;
w26717 <= not pi0647 and not w26716;
w26718 <= not w15342 and not w26701;
w26719 <= w15342 and w26483;
w26720 <= not w26718 and not w26719;
w26721 <= pi0647 and not w26720;
w26722 <= not pi1157 and not w26721;
w26723 <= not w26717 and w26722;
w26724 <= not pi0630 and not w26538;
w26725 <= not w26723 and w26724;
w26726 <= pi0647 and not w26716;
w26727 <= not pi0647 and not w26720;
w26728 <= pi1157 and not w26727;
w26729 <= not w26726 and w26728;
w26730 <= pi0630 and not w26542;
w26731 <= not w26729 and w26730;
w26732 <= not w26725 and not w26731;
w26733 <= pi0787 and not w26732;
w26734 <= not pi0787 and not w26716;
w26735 <= not w26733 and not w26734;
w26736 <= pi0644 and not w26735;
w26737 <= pi0715 and not w26546;
w26738 <= not w26736 and w26737;
w26739 <= w15367 and not w26483;
w26740 <= not w15367 and w26720;
w26741 <= not w26739 and not w26740;
w26742 <= pi0644 and w26741;
w26743 <= not pi0644 and w26483;
w26744 <= not pi0715 and not w26743;
w26745 <= not w26742 and w26744;
w26746 <= pi1160 and not w26745;
w26747 <= not w26738 and w26746;
w26748 <= not pi0644 and not w26735;
w26749 <= pi0644 and w26545;
w26750 <= not pi0715 and not w26749;
w26751 <= not w26748 and w26750;
w26752 <= not pi0644 and w26741;
w26753 <= pi0644 and w26483;
w26754 <= pi0715 and not w26753;
w26755 <= not w26752 and w26754;
w26756 <= not pi1160 and not w26755;
w26757 <= not w26751 and w26756;
w26758 <= pi0790 and not w26747;
w26759 <= not w26757 and w26758;
w26760 <= not pi0790 and w26735;
w26761 <= w4989 and not w26760;
w26762 <= not w26759 and w26761;
w26763 <= not pi0186 and not w4989;
w26764 <= not pi0832 and not w26763;
w26765 <= not w26762 and w26764;
w26766 <= not pi0186 and not w489;
w26767 <= pi0703 and w14208;
w26768 <= not w26766 and not w26767;
w26769 <= not pi0778 and w26768;
w26770 <= not pi0625 and w26767;
w26771 <= not w26768 and not w26770;
w26772 <= pi1153 and not w26771;
w26773 <= not pi1153 and not w26766;
w26774 <= not w26770 and w26773;
w26775 <= not w26772 and not w26774;
w26776 <= pi0778 and not w26775;
w26777 <= not w26769 and not w26776;
w26778 <= not w15408 and w26777;
w26779 <= not w15410 and w26778;
w26780 <= not w15412 and w26779;
w26781 <= not w15414 and w26780;
w26782 <= not w15420 and w26781;
w26783 <= not pi0647 and w26782;
w26784 <= pi0647 and w26766;
w26785 <= not pi1157 and not w26784;
w26786 <= not w26783 and w26785;
w26787 <= pi0630 and w26786;
w26788 <= not pi0752 and w14807;
w26789 <= not w26766 and not w26788;
w26790 <= not w15437 and not w26789;
w26791 <= not pi0785 and not w26790;
w26792 <= not w15442 and not w26789;
w26793 <= pi1155 and not w26792;
w26794 <= not w15445 and w26790;
w26795 <= not pi1155 and not w26794;
w26796 <= not w26793 and not w26795;
w26797 <= pi0785 and not w26796;
w26798 <= not w26791 and not w26797;
w26799 <= not pi0781 and not w26798;
w26800 <= not w15452 and w26798;
w26801 <= pi1154 and not w26800;
w26802 <= not w15455 and w26798;
w26803 <= not pi1154 and not w26802;
w26804 <= not w26801 and not w26803;
w26805 <= pi0781 and not w26804;
w26806 <= not w26799 and not w26805;
w26807 <= not pi0789 and not w26806;
w26808 <= not pi0619 and w26766;
w26809 <= pi0619 and w26806;
w26810 <= pi1159 and not w26808;
w26811 <= not w26809 and w26810;
w26812 <= not pi0619 and w26806;
w26813 <= pi0619 and w26766;
w26814 <= not pi1159 and not w26813;
w26815 <= not w26812 and w26814;
w26816 <= not w26811 and not w26815;
w26817 <= pi0789 and not w26816;
w26818 <= not w26807 and not w26817;
w26819 <= not w15532 and w26818;
w26820 <= w15532 and w26766;
w26821 <= not w26819 and not w26820;
w26822 <= not w15342 and not w26821;
w26823 <= w15342 and w26766;
w26824 <= not w26822 and not w26823;
w26825 <= not w18122 and w26824;
w26826 <= pi0647 and not w26782;
w26827 <= not pi0647 and not w26766;
w26828 <= not w26826 and not w26827;
w26829 <= w15364 and not w26828;
w26830 <= not w26787 and not w26829;
w26831 <= not w26825 and w26830;
w26832 <= pi0787 and not w26831;
w26833 <= w15434 and w26780;
w26834 <= not pi0626 and not w26818;
w26835 <= pi0626 and not w26766;
w26836 <= w14192 and not w26835;
w26837 <= not w26834 and w26836;
w26838 <= pi0626 and not w26818;
w26839 <= not pi0626 and not w26766;
w26840 <= w14191 and not w26839;
w26841 <= not w26838 and w26840;
w26842 <= not w26833 and not w26837;
w26843 <= not w26841 and w26842;
w26844 <= pi0788 and not w26843;
w26845 <= pi0618 and w26778;
w26846 <= pi0609 and w26777;
w26847 <= not w14731 and not w26768;
w26848 <= pi0625 and w26847;
w26849 <= w26789 and not w26847;
w26850 <= not w26848 and not w26849;
w26851 <= w26773 and not w26850;
w26852 <= not pi0608 and not w26772;
w26853 <= not w26851 and w26852;
w26854 <= pi1153 and w26789;
w26855 <= not w26848 and w26854;
w26856 <= pi0608 and not w26774;
w26857 <= not w26855 and w26856;
w26858 <= not w26853 and not w26857;
w26859 <= pi0778 and not w26858;
w26860 <= not pi0778 and not w26849;
w26861 <= not w26859 and not w26860;
w26862 <= not pi0609 and not w26861;
w26863 <= not pi1155 and not w26846;
w26864 <= not w26862 and w26863;
w26865 <= not pi0660 and not w26793;
w26866 <= not w26864 and w26865;
w26867 <= not pi0609 and w26777;
w26868 <= pi0609 and not w26861;
w26869 <= pi1155 and not w26867;
w26870 <= not w26868 and w26869;
w26871 <= pi0660 and not w26795;
w26872 <= not w26870 and w26871;
w26873 <= not w26866 and not w26872;
w26874 <= pi0785 and not w26873;
w26875 <= not pi0785 and not w26861;
w26876 <= not w26874 and not w26875;
w26877 <= not pi0618 and not w26876;
w26878 <= not pi1154 and not w26845;
w26879 <= not w26877 and w26878;
w26880 <= not pi0627 and not w26801;
w26881 <= not w26879 and w26880;
w26882 <= not pi0618 and w26778;
w26883 <= pi0618 and not w26876;
w26884 <= pi1154 and not w26882;
w26885 <= not w26883 and w26884;
w26886 <= pi0627 and not w26803;
w26887 <= not w26885 and w26886;
w26888 <= not w26881 and not w26887;
w26889 <= pi0781 and not w26888;
w26890 <= not pi0781 and not w26876;
w26891 <= not w26889 and not w26890;
w26892 <= not pi0789 and w26891;
w26893 <= not pi0619 and not w26891;
w26894 <= pi0619 and w26779;
w26895 <= not pi1159 and not w26894;
w26896 <= not w26893 and w26895;
w26897 <= not pi0648 and not w26811;
w26898 <= not w26896 and w26897;
w26899 <= pi0619 and not w26891;
w26900 <= not pi0619 and w26779;
w26901 <= pi1159 and not w26900;
w26902 <= not w26899 and w26901;
w26903 <= pi0648 and not w26815;
w26904 <= not w26902 and w26903;
w26905 <= pi0789 and not w26898;
w26906 <= not w26904 and w26905;
w26907 <= w15533 and not w26892;
w26908 <= not w26906 and w26907;
w26909 <= not w26844 and not w26908;
w26910 <= not w17927 and not w26909;
w26911 <= w15417 and not w26821;
w26912 <= w18414 and w26781;
w26913 <= not w26911 and not w26912;
w26914 <= not pi0629 and not w26913;
w26915 <= w18418 and w26781;
w26916 <= w15416 and not w26821;
w26917 <= not w26915 and not w26916;
w26918 <= pi0629 and not w26917;
w26919 <= not w26914 and not w26918;
w26920 <= pi0792 and not w26919;
w26921 <= not w17769 and not w26920;
w26922 <= not w26910 and w26921;
w26923 <= not w26832 and not w26922;
w26924 <= not pi0790 and w26923;
w26925 <= not pi0787 and not w26782;
w26926 <= pi1157 and not w26828;
w26927 <= not w26786 and not w26926;
w26928 <= pi0787 and not w26927;
w26929 <= not w26925 and not w26928;
w26930 <= not pi0644 and w26929;
w26931 <= pi0644 and w26923;
w26932 <= pi0715 and not w26930;
w26933 <= not w26931 and w26932;
w26934 <= not w15367 and not w26824;
w26935 <= w15367 and w26766;
w26936 <= not w26934 and not w26935;
w26937 <= pi0644 and not w26936;
w26938 <= not pi0644 and w26766;
w26939 <= not pi0715 and not w26938;
w26940 <= not w26937 and w26939;
w26941 <= pi1160 and not w26940;
w26942 <= not w26933 and w26941;
w26943 <= not pi0644 and not w26936;
w26944 <= pi0644 and w26766;
w26945 <= pi0715 and not w26944;
w26946 <= not w26943 and w26945;
w26947 <= pi0644 and w26929;
w26948 <= not pi0644 and w26923;
w26949 <= not pi0715 and not w26947;
w26950 <= not w26948 and w26949;
w26951 <= not pi1160 and not w26946;
w26952 <= not w26950 and w26951;
w26953 <= not w26942 and not w26952;
w26954 <= pi0790 and not w26953;
w26955 <= pi0832 and not w26924;
w26956 <= not w26954 and w26955;
w26957 <= not w26765 and not w26956;
w26958 <= not pi0187 and not w14622;
w26959 <= w14198 and not w26958;
w26960 <= pi0187 and not w134;
w26961 <= not pi0187 and not pi0726;
w26962 <= not w14615 and w26961;
w26963 <= not pi0187 and not w14204;
w26964 <= w14210 and not w26963;
w26965 <= not pi0187 and w15635;
w26966 <= pi0187 and not w15639;
w26967 <= not pi0038 and not w26966;
w26968 <= not w26965 and w26967;
w26969 <= pi0726 and not w26964;
w26970 <= not w26968 and w26969;
w26971 <= w134 and not w26962;
w26972 <= not w26970 and w26971;
w26973 <= not w26960 and not w26972;
w26974 <= not pi0778 and not w26973;
w26975 <= not pi0625 and w26958;
w26976 <= pi0625 and w26973;
w26977 <= pi1153 and not w26975;
w26978 <= not w26976 and w26977;
w26979 <= not pi0625 and w26973;
w26980 <= pi0625 and w26958;
w26981 <= not pi1153 and not w26980;
w26982 <= not w26979 and w26981;
w26983 <= not w26978 and not w26982;
w26984 <= pi0778 and not w26983;
w26985 <= not w26974 and not w26984;
w26986 <= not w14638 and not w26985;
w26987 <= w14638 and not w26958;
w26988 <= not w26986 and not w26987;
w26989 <= not w14202 and w26988;
w26990 <= w14202 and w26958;
w26991 <= not w26989 and not w26990;
w26992 <= not w14198 and w26991;
w26993 <= not w26959 and not w26992;
w26994 <= not w14194 and w26993;
w26995 <= w14194 and w26958;
w26996 <= not w26994 and not w26995;
w26997 <= not pi0792 and w26996;
w26998 <= not pi0628 and w26958;
w26999 <= pi0628 and not w26996;
w27000 <= pi1156 and not w26998;
w27001 <= not w26999 and w27000;
w27002 <= pi0628 and w26958;
w27003 <= not pi0628 and not w26996;
w27004 <= not pi1156 and not w27002;
w27005 <= not w27003 and w27004;
w27006 <= not w27001 and not w27005;
w27007 <= pi0792 and not w27006;
w27008 <= not w26997 and not w27007;
w27009 <= not pi0787 and not w27008;
w27010 <= not pi0647 and w26958;
w27011 <= pi0647 and w27008;
w27012 <= pi1157 and not w27010;
w27013 <= not w27011 and w27012;
w27014 <= not pi0647 and w27008;
w27015 <= pi0647 and w26958;
w27016 <= not pi1157 and not w27015;
w27017 <= not w27014 and w27016;
w27018 <= not w27013 and not w27017;
w27019 <= pi0787 and not w27018;
w27020 <= not w27009 and not w27019;
w27021 <= not pi0644 and w27020;
w27022 <= not pi0618 and w26958;
w27023 <= not pi0770 and not w17002;
w27024 <= not w18575 and not w27023;
w27025 <= not pi0187 and not w27024;
w27026 <= not pi0187 and not w16996;
w27027 <= not pi0770 and not w27026;
w27028 <= not w22010 and w27027;
w27029 <= not w27025 and not w27028;
w27030 <= w134 and w27029;
w27031 <= not w26960 and not w27030;
w27032 <= not w14680 and not w27031;
w27033 <= w14680 and not w26958;
w27034 <= not w27032 and not w27033;
w27035 <= not pi0785 and not w27034;
w27036 <= not w14854 and not w26958;
w27037 <= pi0609 and w27032;
w27038 <= not w27036 and not w27037;
w27039 <= pi1155 and not w27038;
w27040 <= not w14859 and not w26958;
w27041 <= not pi0609 and w27032;
w27042 <= not w27040 and not w27041;
w27043 <= not pi1155 and not w27042;
w27044 <= not w27039 and not w27043;
w27045 <= pi0785 and not w27044;
w27046 <= not w27035 and not w27045;
w27047 <= pi0618 and w27046;
w27048 <= pi1154 and not w27022;
w27049 <= not w27047 and w27048;
w27050 <= pi0187 and w17031;
w27051 <= not pi0187 and w17040;
w27052 <= pi0770 and not w17033;
w27053 <= not w27050 and w27052;
w27054 <= not w27051 and w27053;
w27055 <= not pi0187 and not w17051;
w27056 <= pi0187 and w17059;
w27057 <= not pi0770 and not w27055;
w27058 <= not w27056 and w27057;
w27059 <= pi0726 and not w27058;
w27060 <= not w27054 and w27059;
w27061 <= not pi0726 and not w27029;
w27062 <= w134 and not w27060;
w27063 <= not w27061 and w27062;
w27064 <= not w26960 and not w27063;
w27065 <= not pi0625 and w27064;
w27066 <= pi0625 and w27031;
w27067 <= not pi1153 and not w27066;
w27068 <= not w27065 and w27067;
w27069 <= not pi0608 and not w26978;
w27070 <= not w27068 and w27069;
w27071 <= not pi0625 and w27031;
w27072 <= pi0625 and w27064;
w27073 <= pi1153 and not w27071;
w27074 <= not w27072 and w27073;
w27075 <= pi0608 and not w26982;
w27076 <= not w27074 and w27075;
w27077 <= not w27070 and not w27076;
w27078 <= pi0778 and not w27077;
w27079 <= not pi0778 and w27064;
w27080 <= not w27078 and not w27079;
w27081 <= not pi0609 and not w27080;
w27082 <= pi0609 and w26985;
w27083 <= not pi1155 and not w27082;
w27084 <= not w27081 and w27083;
w27085 <= not pi0660 and not w27039;
w27086 <= not w27084 and w27085;
w27087 <= not pi0609 and w26985;
w27088 <= pi0609 and not w27080;
w27089 <= pi1155 and not w27087;
w27090 <= not w27088 and w27089;
w27091 <= pi0660 and not w27043;
w27092 <= not w27090 and w27091;
w27093 <= not w27086 and not w27092;
w27094 <= pi0785 and not w27093;
w27095 <= not pi0785 and not w27080;
w27096 <= not w27094 and not w27095;
w27097 <= not pi0618 and not w27096;
w27098 <= pi0618 and w26988;
w27099 <= not pi1154 and not w27098;
w27100 <= not w27097 and w27099;
w27101 <= not pi0627 and not w27049;
w27102 <= not w27100 and w27101;
w27103 <= not pi0618 and w27046;
w27104 <= pi0618 and w26958;
w27105 <= not pi1154 and not w27104;
w27106 <= not w27103 and w27105;
w27107 <= not pi0618 and w26988;
w27108 <= pi0618 and not w27096;
w27109 <= pi1154 and not w27107;
w27110 <= not w27108 and w27109;
w27111 <= pi0627 and not w27106;
w27112 <= not w27110 and w27111;
w27113 <= not w27102 and not w27112;
w27114 <= pi0781 and not w27113;
w27115 <= not pi0781 and not w27096;
w27116 <= not w27114 and not w27115;
w27117 <= not pi0619 and not w27116;
w27118 <= pi0619 and not w26991;
w27119 <= not pi1159 and not w27118;
w27120 <= not w27117 and w27119;
w27121 <= not pi0619 and w26958;
w27122 <= not pi0781 and not w27046;
w27123 <= not w27049 and not w27106;
w27124 <= pi0781 and not w27123;
w27125 <= not w27122 and not w27124;
w27126 <= pi0619 and w27125;
w27127 <= pi1159 and not w27121;
w27128 <= not w27126 and w27127;
w27129 <= not pi0648 and not w27128;
w27130 <= not w27120 and w27129;
w27131 <= pi0619 and not w27116;
w27132 <= not pi0619 and not w26991;
w27133 <= pi1159 and not w27132;
w27134 <= not w27131 and w27133;
w27135 <= not pi0619 and w27125;
w27136 <= pi0619 and w26958;
w27137 <= not pi1159 and not w27136;
w27138 <= not w27135 and w27137;
w27139 <= pi0648 and not w27138;
w27140 <= not w27134 and w27139;
w27141 <= not w27130 and not w27140;
w27142 <= pi0789 and not w27141;
w27143 <= not pi0789 and not w27116;
w27144 <= not w27142 and not w27143;
w27145 <= not pi0788 and w27144;
w27146 <= not pi0626 and w27144;
w27147 <= pi0626 and not w26993;
w27148 <= not pi0641 and not w27147;
w27149 <= not w27146 and w27148;
w27150 <= not pi0789 and not w27125;
w27151 <= not w27128 and not w27138;
w27152 <= pi0789 and not w27151;
w27153 <= not w27150 and not w27152;
w27154 <= not pi0626 and not w27153;
w27155 <= pi0626 and not w26958;
w27156 <= pi0641 and not w27155;
w27157 <= not w27154 and w27156;
w27158 <= not pi1158 and not w27157;
w27159 <= not w27149 and w27158;
w27160 <= pi0626 and w27144;
w27161 <= not pi0626 and not w26993;
w27162 <= pi0641 and not w27161;
w27163 <= not w27160 and w27162;
w27164 <= pi0626 and not w27153;
w27165 <= not pi0626 and not w26958;
w27166 <= not pi0641 and not w27165;
w27167 <= not w27164 and w27166;
w27168 <= pi1158 and not w27167;
w27169 <= not w27163 and w27168;
w27170 <= not w27159 and not w27169;
w27171 <= pi0788 and not w27170;
w27172 <= not w27145 and not w27171;
w27173 <= not pi0628 and w27172;
w27174 <= not w15532 and w27153;
w27175 <= w15532 and w26958;
w27176 <= not w27174 and not w27175;
w27177 <= pi0628 and not w27176;
w27178 <= not pi1156 and not w27177;
w27179 <= not w27173 and w27178;
w27180 <= not pi0629 and not w27001;
w27181 <= not w27179 and w27180;
w27182 <= pi0628 and w27172;
w27183 <= not pi0628 and not w27176;
w27184 <= pi1156 and not w27183;
w27185 <= not w27182 and w27184;
w27186 <= pi0629 and not w27005;
w27187 <= not w27185 and w27186;
w27188 <= not w27181 and not w27187;
w27189 <= pi0792 and not w27188;
w27190 <= not pi0792 and w27172;
w27191 <= not w27189 and not w27190;
w27192 <= not pi0647 and not w27191;
w27193 <= not w15342 and not w27176;
w27194 <= w15342 and w26958;
w27195 <= not w27193 and not w27194;
w27196 <= pi0647 and not w27195;
w27197 <= not pi1157 and not w27196;
w27198 <= not w27192 and w27197;
w27199 <= not pi0630 and not w27013;
w27200 <= not w27198 and w27199;
w27201 <= pi0647 and not w27191;
w27202 <= not pi0647 and not w27195;
w27203 <= pi1157 and not w27202;
w27204 <= not w27201 and w27203;
w27205 <= pi0630 and not w27017;
w27206 <= not w27204 and w27205;
w27207 <= not w27200 and not w27206;
w27208 <= pi0787 and not w27207;
w27209 <= not pi0787 and not w27191;
w27210 <= not w27208 and not w27209;
w27211 <= pi0644 and not w27210;
w27212 <= pi0715 and not w27021;
w27213 <= not w27211 and w27212;
w27214 <= w15367 and not w26958;
w27215 <= not w15367 and w27195;
w27216 <= not w27214 and not w27215;
w27217 <= pi0644 and w27216;
w27218 <= not pi0644 and w26958;
w27219 <= not pi0715 and not w27218;
w27220 <= not w27217 and w27219;
w27221 <= pi1160 and not w27220;
w27222 <= not w27213 and w27221;
w27223 <= not pi0644 and not w27210;
w27224 <= pi0644 and w27020;
w27225 <= not pi0715 and not w27224;
w27226 <= not w27223 and w27225;
w27227 <= not pi0644 and w27216;
w27228 <= pi0644 and w26958;
w27229 <= pi0715 and not w27228;
w27230 <= not w27227 and w27229;
w27231 <= not pi1160 and not w27230;
w27232 <= not w27226 and w27231;
w27233 <= pi0790 and not w27222;
w27234 <= not w27232 and w27233;
w27235 <= not pi0790 and w27210;
w27236 <= w4989 and not w27235;
w27237 <= not w27234 and w27236;
w27238 <= not pi0187 and not w4989;
w27239 <= not pi0832 and not w27238;
w27240 <= not w27237 and w27239;
w27241 <= not pi0187 and not w489;
w27242 <= pi0726 and w14208;
w27243 <= not w27241 and not w27242;
w27244 <= not pi0778 and w27243;
w27245 <= not pi0625 and w27242;
w27246 <= not w27243 and not w27245;
w27247 <= pi1153 and not w27246;
w27248 <= not pi1153 and not w27241;
w27249 <= not w27245 and w27248;
w27250 <= not w27247 and not w27249;
w27251 <= pi0778 and not w27250;
w27252 <= not w27244 and not w27251;
w27253 <= not w15408 and w27252;
w27254 <= not w15410 and w27253;
w27255 <= not w15412 and w27254;
w27256 <= not w15414 and w27255;
w27257 <= not w15420 and w27256;
w27258 <= not pi0647 and w27257;
w27259 <= pi0647 and w27241;
w27260 <= not pi1157 and not w27259;
w27261 <= not w27258 and w27260;
w27262 <= pi0630 and w27261;
w27263 <= not pi0770 and w14807;
w27264 <= not w27241 and not w27263;
w27265 <= not w15437 and not w27264;
w27266 <= not pi0785 and not w27265;
w27267 <= not w15442 and not w27264;
w27268 <= pi1155 and not w27267;
w27269 <= not w15445 and w27265;
w27270 <= not pi1155 and not w27269;
w27271 <= not w27268 and not w27270;
w27272 <= pi0785 and not w27271;
w27273 <= not w27266 and not w27272;
w27274 <= not pi0781 and not w27273;
w27275 <= not w15452 and w27273;
w27276 <= pi1154 and not w27275;
w27277 <= not w15455 and w27273;
w27278 <= not pi1154 and not w27277;
w27279 <= not w27276 and not w27278;
w27280 <= pi0781 and not w27279;
w27281 <= not w27274 and not w27280;
w27282 <= not pi0789 and not w27281;
w27283 <= not pi0619 and w27241;
w27284 <= pi0619 and w27281;
w27285 <= pi1159 and not w27283;
w27286 <= not w27284 and w27285;
w27287 <= not pi0619 and w27281;
w27288 <= pi0619 and w27241;
w27289 <= not pi1159 and not w27288;
w27290 <= not w27287 and w27289;
w27291 <= not w27286 and not w27290;
w27292 <= pi0789 and not w27291;
w27293 <= not w27282 and not w27292;
w27294 <= not w15532 and w27293;
w27295 <= w15532 and w27241;
w27296 <= not w27294 and not w27295;
w27297 <= not w15342 and not w27296;
w27298 <= w15342 and w27241;
w27299 <= not w27297 and not w27298;
w27300 <= not w18122 and w27299;
w27301 <= pi0647 and not w27257;
w27302 <= not pi0647 and not w27241;
w27303 <= not w27301 and not w27302;
w27304 <= w15364 and not w27303;
w27305 <= not w27262 and not w27304;
w27306 <= not w27300 and w27305;
w27307 <= pi0787 and not w27306;
w27308 <= w15434 and w27255;
w27309 <= not pi0626 and not w27293;
w27310 <= pi0626 and not w27241;
w27311 <= w14192 and not w27310;
w27312 <= not w27309 and w27311;
w27313 <= pi0626 and not w27293;
w27314 <= not pi0626 and not w27241;
w27315 <= w14191 and not w27314;
w27316 <= not w27313 and w27315;
w27317 <= not w27308 and not w27312;
w27318 <= not w27316 and w27317;
w27319 <= pi0788 and not w27318;
w27320 <= pi0618 and w27253;
w27321 <= pi0609 and w27252;
w27322 <= not w14731 and not w27243;
w27323 <= pi0625 and w27322;
w27324 <= w27264 and not w27322;
w27325 <= not w27323 and not w27324;
w27326 <= w27248 and not w27325;
w27327 <= not pi0608 and not w27247;
w27328 <= not w27326 and w27327;
w27329 <= pi1153 and w27264;
w27330 <= not w27323 and w27329;
w27331 <= pi0608 and not w27249;
w27332 <= not w27330 and w27331;
w27333 <= not w27328 and not w27332;
w27334 <= pi0778 and not w27333;
w27335 <= not pi0778 and not w27324;
w27336 <= not w27334 and not w27335;
w27337 <= not pi0609 and not w27336;
w27338 <= not pi1155 and not w27321;
w27339 <= not w27337 and w27338;
w27340 <= not pi0660 and not w27268;
w27341 <= not w27339 and w27340;
w27342 <= not pi0609 and w27252;
w27343 <= pi0609 and not w27336;
w27344 <= pi1155 and not w27342;
w27345 <= not w27343 and w27344;
w27346 <= pi0660 and not w27270;
w27347 <= not w27345 and w27346;
w27348 <= not w27341 and not w27347;
w27349 <= pi0785 and not w27348;
w27350 <= not pi0785 and not w27336;
w27351 <= not w27349 and not w27350;
w27352 <= not pi0618 and not w27351;
w27353 <= not pi1154 and not w27320;
w27354 <= not w27352 and w27353;
w27355 <= not pi0627 and not w27276;
w27356 <= not w27354 and w27355;
w27357 <= not pi0618 and w27253;
w27358 <= pi0618 and not w27351;
w27359 <= pi1154 and not w27357;
w27360 <= not w27358 and w27359;
w27361 <= pi0627 and not w27278;
w27362 <= not w27360 and w27361;
w27363 <= not w27356 and not w27362;
w27364 <= pi0781 and not w27363;
w27365 <= not pi0781 and not w27351;
w27366 <= not w27364 and not w27365;
w27367 <= not pi0789 and w27366;
w27368 <= not pi0619 and not w27366;
w27369 <= pi0619 and w27254;
w27370 <= not pi1159 and not w27369;
w27371 <= not w27368 and w27370;
w27372 <= not pi0648 and not w27286;
w27373 <= not w27371 and w27372;
w27374 <= pi0619 and not w27366;
w27375 <= not pi0619 and w27254;
w27376 <= pi1159 and not w27375;
w27377 <= not w27374 and w27376;
w27378 <= pi0648 and not w27290;
w27379 <= not w27377 and w27378;
w27380 <= pi0789 and not w27373;
w27381 <= not w27379 and w27380;
w27382 <= w15533 and not w27367;
w27383 <= not w27381 and w27382;
w27384 <= not w27319 and not w27383;
w27385 <= not w17927 and not w27384;
w27386 <= w15417 and not w27296;
w27387 <= w18414 and w27256;
w27388 <= not w27386 and not w27387;
w27389 <= not pi0629 and not w27388;
w27390 <= w18418 and w27256;
w27391 <= w15416 and not w27296;
w27392 <= not w27390 and not w27391;
w27393 <= pi0629 and not w27392;
w27394 <= not w27389 and not w27393;
w27395 <= pi0792 and not w27394;
w27396 <= not w17769 and not w27395;
w27397 <= not w27385 and w27396;
w27398 <= not w27307 and not w27397;
w27399 <= not pi0790 and w27398;
w27400 <= not pi0787 and not w27257;
w27401 <= pi1157 and not w27303;
w27402 <= not w27261 and not w27401;
w27403 <= pi0787 and not w27402;
w27404 <= not w27400 and not w27403;
w27405 <= not pi0644 and w27404;
w27406 <= pi0644 and w27398;
w27407 <= pi0715 and not w27405;
w27408 <= not w27406 and w27407;
w27409 <= not w15367 and not w27299;
w27410 <= w15367 and w27241;
w27411 <= not w27409 and not w27410;
w27412 <= pi0644 and not w27411;
w27413 <= not pi0644 and w27241;
w27414 <= not pi0715 and not w27413;
w27415 <= not w27412 and w27414;
w27416 <= pi1160 and not w27415;
w27417 <= not w27408 and w27416;
w27418 <= not pi0644 and not w27411;
w27419 <= pi0644 and w27241;
w27420 <= pi0715 and not w27419;
w27421 <= not w27418 and w27420;
w27422 <= pi0644 and w27404;
w27423 <= not pi0644 and w27398;
w27424 <= not pi0715 and not w27422;
w27425 <= not w27423 and w27424;
w27426 <= not pi1160 and not w27421;
w27427 <= not w27425 and w27426;
w27428 <= not w27417 and not w27427;
w27429 <= pi0790 and not w27428;
w27430 <= pi0832 and not w27399;
w27431 <= not w27429 and w27430;
w27432 <= not w27240 and not w27431;
w27433 <= not pi0188 and not w14622;
w27434 <= w14198 and not w27433;
w27435 <= pi0188 and not w134;
w27436 <= not pi0188 and not pi0705;
w27437 <= not w14615 and w27436;
w27438 <= not pi0188 and not w14204;
w27439 <= w14210 and not w27438;
w27440 <= not pi0188 and w15635;
w27441 <= pi0188 and not w15639;
w27442 <= not pi0038 and not w27441;
w27443 <= not w27440 and w27442;
w27444 <= pi0705 and not w27439;
w27445 <= not w27443 and w27444;
w27446 <= w134 and not w27437;
w27447 <= not w27445 and w27446;
w27448 <= not w27435 and not w27447;
w27449 <= not pi0778 and not w27448;
w27450 <= not pi0625 and w27433;
w27451 <= pi0625 and w27448;
w27452 <= pi1153 and not w27450;
w27453 <= not w27451 and w27452;
w27454 <= not pi0625 and w27448;
w27455 <= pi0625 and w27433;
w27456 <= not pi1153 and not w27455;
w27457 <= not w27454 and w27456;
w27458 <= not w27453 and not w27457;
w27459 <= pi0778 and not w27458;
w27460 <= not w27449 and not w27459;
w27461 <= not w14638 and not w27460;
w27462 <= w14638 and not w27433;
w27463 <= not w27461 and not w27462;
w27464 <= not w14202 and w27463;
w27465 <= w14202 and w27433;
w27466 <= not w27464 and not w27465;
w27467 <= not w14198 and w27466;
w27468 <= not w27434 and not w27467;
w27469 <= not w14194 and w27468;
w27470 <= w14194 and w27433;
w27471 <= not w27469 and not w27470;
w27472 <= not pi0792 and w27471;
w27473 <= not pi0628 and w27433;
w27474 <= pi0628 and not w27471;
w27475 <= pi1156 and not w27473;
w27476 <= not w27474 and w27475;
w27477 <= pi0628 and w27433;
w27478 <= not pi0628 and not w27471;
w27479 <= not pi1156 and not w27477;
w27480 <= not w27478 and w27479;
w27481 <= not w27476 and not w27480;
w27482 <= pi0792 and not w27481;
w27483 <= not w27472 and not w27482;
w27484 <= not pi0787 and not w27483;
w27485 <= not pi0647 and w27433;
w27486 <= pi0647 and w27483;
w27487 <= pi1157 and not w27485;
w27488 <= not w27486 and w27487;
w27489 <= not pi0647 and w27483;
w27490 <= pi0647 and w27433;
w27491 <= not pi1157 and not w27490;
w27492 <= not w27489 and w27491;
w27493 <= not w27488 and not w27492;
w27494 <= pi0787 and not w27493;
w27495 <= not w27484 and not w27494;
w27496 <= not pi0644 and w27495;
w27497 <= not pi0618 and w27433;
w27498 <= not pi0768 and not w17002;
w27499 <= not w19876 and not w27498;
w27500 <= not pi0188 and not w27499;
w27501 <= not pi0188 and not w16996;
w27502 <= not pi0768 and not w27501;
w27503 <= not w22010 and w27502;
w27504 <= not w27500 and not w27503;
w27505 <= w134 and w27504;
w27506 <= not w27435 and not w27505;
w27507 <= not w14680 and not w27506;
w27508 <= w14680 and not w27433;
w27509 <= not w27507 and not w27508;
w27510 <= not pi0785 and not w27509;
w27511 <= not w14854 and not w27433;
w27512 <= pi0609 and w27507;
w27513 <= not w27511 and not w27512;
w27514 <= pi1155 and not w27513;
w27515 <= not w14859 and not w27433;
w27516 <= not pi0609 and w27507;
w27517 <= not w27515 and not w27516;
w27518 <= not pi1155 and not w27517;
w27519 <= not w27514 and not w27518;
w27520 <= pi0785 and not w27519;
w27521 <= not w27510 and not w27520;
w27522 <= pi0618 and w27521;
w27523 <= pi1154 and not w27497;
w27524 <= not w27522 and w27523;
w27525 <= pi0188 and w17031;
w27526 <= not pi0188 and w17040;
w27527 <= pi0768 and not w17033;
w27528 <= not w27525 and w27527;
w27529 <= not w27526 and w27528;
w27530 <= not pi0188 and not w17051;
w27531 <= pi0188 and w17059;
w27532 <= not pi0768 and not w27530;
w27533 <= not w27531 and w27532;
w27534 <= pi0705 and not w27533;
w27535 <= not w27529 and w27534;
w27536 <= not pi0705 and not w27504;
w27537 <= w134 and not w27535;
w27538 <= not w27536 and w27537;
w27539 <= not w27435 and not w27538;
w27540 <= not pi0625 and w27539;
w27541 <= pi0625 and w27506;
w27542 <= not pi1153 and not w27541;
w27543 <= not w27540 and w27542;
w27544 <= not pi0608 and not w27453;
w27545 <= not w27543 and w27544;
w27546 <= not pi0625 and w27506;
w27547 <= pi0625 and w27539;
w27548 <= pi1153 and not w27546;
w27549 <= not w27547 and w27548;
w27550 <= pi0608 and not w27457;
w27551 <= not w27549 and w27550;
w27552 <= not w27545 and not w27551;
w27553 <= pi0778 and not w27552;
w27554 <= not pi0778 and w27539;
w27555 <= not w27553 and not w27554;
w27556 <= not pi0609 and not w27555;
w27557 <= pi0609 and w27460;
w27558 <= not pi1155 and not w27557;
w27559 <= not w27556 and w27558;
w27560 <= not pi0660 and not w27514;
w27561 <= not w27559 and w27560;
w27562 <= not pi0609 and w27460;
w27563 <= pi0609 and not w27555;
w27564 <= pi1155 and not w27562;
w27565 <= not w27563 and w27564;
w27566 <= pi0660 and not w27518;
w27567 <= not w27565 and w27566;
w27568 <= not w27561 and not w27567;
w27569 <= pi0785 and not w27568;
w27570 <= not pi0785 and not w27555;
w27571 <= not w27569 and not w27570;
w27572 <= not pi0618 and not w27571;
w27573 <= pi0618 and w27463;
w27574 <= not pi1154 and not w27573;
w27575 <= not w27572 and w27574;
w27576 <= not pi0627 and not w27524;
w27577 <= not w27575 and w27576;
w27578 <= not pi0618 and w27521;
w27579 <= pi0618 and w27433;
w27580 <= not pi1154 and not w27579;
w27581 <= not w27578 and w27580;
w27582 <= not pi0618 and w27463;
w27583 <= pi0618 and not w27571;
w27584 <= pi1154 and not w27582;
w27585 <= not w27583 and w27584;
w27586 <= pi0627 and not w27581;
w27587 <= not w27585 and w27586;
w27588 <= not w27577 and not w27587;
w27589 <= pi0781 and not w27588;
w27590 <= not pi0781 and not w27571;
w27591 <= not w27589 and not w27590;
w27592 <= not pi0619 and not w27591;
w27593 <= pi0619 and not w27466;
w27594 <= not pi1159 and not w27593;
w27595 <= not w27592 and w27594;
w27596 <= not pi0619 and w27433;
w27597 <= not pi0781 and not w27521;
w27598 <= not w27524 and not w27581;
w27599 <= pi0781 and not w27598;
w27600 <= not w27597 and not w27599;
w27601 <= pi0619 and w27600;
w27602 <= pi1159 and not w27596;
w27603 <= not w27601 and w27602;
w27604 <= not pi0648 and not w27603;
w27605 <= not w27595 and w27604;
w27606 <= pi0619 and not w27591;
w27607 <= not pi0619 and not w27466;
w27608 <= pi1159 and not w27607;
w27609 <= not w27606 and w27608;
w27610 <= not pi0619 and w27600;
w27611 <= pi0619 and w27433;
w27612 <= not pi1159 and not w27611;
w27613 <= not w27610 and w27612;
w27614 <= pi0648 and not w27613;
w27615 <= not w27609 and w27614;
w27616 <= not w27605 and not w27615;
w27617 <= pi0789 and not w27616;
w27618 <= not pi0789 and not w27591;
w27619 <= not w27617 and not w27618;
w27620 <= not pi0788 and w27619;
w27621 <= not pi0626 and w27619;
w27622 <= pi0626 and not w27468;
w27623 <= not pi0641 and not w27622;
w27624 <= not w27621 and w27623;
w27625 <= not pi0789 and not w27600;
w27626 <= not w27603 and not w27613;
w27627 <= pi0789 and not w27626;
w27628 <= not w27625 and not w27627;
w27629 <= not pi0626 and not w27628;
w27630 <= pi0626 and not w27433;
w27631 <= pi0641 and not w27630;
w27632 <= not w27629 and w27631;
w27633 <= not pi1158 and not w27632;
w27634 <= not w27624 and w27633;
w27635 <= pi0626 and w27619;
w27636 <= not pi0626 and not w27468;
w27637 <= pi0641 and not w27636;
w27638 <= not w27635 and w27637;
w27639 <= pi0626 and not w27628;
w27640 <= not pi0626 and not w27433;
w27641 <= not pi0641 and not w27640;
w27642 <= not w27639 and w27641;
w27643 <= pi1158 and not w27642;
w27644 <= not w27638 and w27643;
w27645 <= not w27634 and not w27644;
w27646 <= pi0788 and not w27645;
w27647 <= not w27620 and not w27646;
w27648 <= not pi0628 and w27647;
w27649 <= not w15532 and w27628;
w27650 <= w15532 and w27433;
w27651 <= not w27649 and not w27650;
w27652 <= pi0628 and not w27651;
w27653 <= not pi1156 and not w27652;
w27654 <= not w27648 and w27653;
w27655 <= not pi0629 and not w27476;
w27656 <= not w27654 and w27655;
w27657 <= pi0628 and w27647;
w27658 <= not pi0628 and not w27651;
w27659 <= pi1156 and not w27658;
w27660 <= not w27657 and w27659;
w27661 <= pi0629 and not w27480;
w27662 <= not w27660 and w27661;
w27663 <= not w27656 and not w27662;
w27664 <= pi0792 and not w27663;
w27665 <= not pi0792 and w27647;
w27666 <= not w27664 and not w27665;
w27667 <= not pi0647 and not w27666;
w27668 <= not w15342 and not w27651;
w27669 <= w15342 and w27433;
w27670 <= not w27668 and not w27669;
w27671 <= pi0647 and not w27670;
w27672 <= not pi1157 and not w27671;
w27673 <= not w27667 and w27672;
w27674 <= not pi0630 and not w27488;
w27675 <= not w27673 and w27674;
w27676 <= pi0647 and not w27666;
w27677 <= not pi0647 and not w27670;
w27678 <= pi1157 and not w27677;
w27679 <= not w27676 and w27678;
w27680 <= pi0630 and not w27492;
w27681 <= not w27679 and w27680;
w27682 <= not w27675 and not w27681;
w27683 <= pi0787 and not w27682;
w27684 <= not pi0787 and not w27666;
w27685 <= not w27683 and not w27684;
w27686 <= pi0644 and not w27685;
w27687 <= pi0715 and not w27496;
w27688 <= not w27686 and w27687;
w27689 <= w15367 and not w27433;
w27690 <= not w15367 and w27670;
w27691 <= not w27689 and not w27690;
w27692 <= pi0644 and w27691;
w27693 <= not pi0644 and w27433;
w27694 <= not pi0715 and not w27693;
w27695 <= not w27692 and w27694;
w27696 <= pi1160 and not w27695;
w27697 <= not w27688 and w27696;
w27698 <= not pi0644 and not w27685;
w27699 <= pi0644 and w27495;
w27700 <= not pi0715 and not w27699;
w27701 <= not w27698 and w27700;
w27702 <= not pi0644 and w27691;
w27703 <= pi0644 and w27433;
w27704 <= pi0715 and not w27703;
w27705 <= not w27702 and w27704;
w27706 <= not pi1160 and not w27705;
w27707 <= not w27701 and w27706;
w27708 <= pi0790 and not w27697;
w27709 <= not w27707 and w27708;
w27710 <= not pi0790 and w27685;
w27711 <= w4989 and not w27710;
w27712 <= not w27709 and w27711;
w27713 <= not pi0188 and not w4989;
w27714 <= not pi0832 and not w27713;
w27715 <= not w27712 and w27714;
w27716 <= not pi0188 and not w489;
w27717 <= pi0705 and w14208;
w27718 <= not w27716 and not w27717;
w27719 <= not pi0778 and w27718;
w27720 <= not pi0625 and w27717;
w27721 <= not w27718 and not w27720;
w27722 <= pi1153 and not w27721;
w27723 <= not pi1153 and not w27716;
w27724 <= not w27720 and w27723;
w27725 <= not w27722 and not w27724;
w27726 <= pi0778 and not w27725;
w27727 <= not w27719 and not w27726;
w27728 <= not w15408 and w27727;
w27729 <= not w15410 and w27728;
w27730 <= not w15412 and w27729;
w27731 <= not w15414 and w27730;
w27732 <= not w15420 and w27731;
w27733 <= not pi0647 and w27732;
w27734 <= pi0647 and w27716;
w27735 <= not pi1157 and not w27734;
w27736 <= not w27733 and w27735;
w27737 <= pi0630 and w27736;
w27738 <= not pi0768 and w14807;
w27739 <= not w27716 and not w27738;
w27740 <= not w15437 and not w27739;
w27741 <= not pi0785 and not w27740;
w27742 <= not w15442 and not w27739;
w27743 <= pi1155 and not w27742;
w27744 <= not w15445 and w27740;
w27745 <= not pi1155 and not w27744;
w27746 <= not w27743 and not w27745;
w27747 <= pi0785 and not w27746;
w27748 <= not w27741 and not w27747;
w27749 <= not pi0781 and not w27748;
w27750 <= not w15452 and w27748;
w27751 <= pi1154 and not w27750;
w27752 <= not w15455 and w27748;
w27753 <= not pi1154 and not w27752;
w27754 <= not w27751 and not w27753;
w27755 <= pi0781 and not w27754;
w27756 <= not w27749 and not w27755;
w27757 <= not pi0789 and not w27756;
w27758 <= not pi0619 and w27716;
w27759 <= pi0619 and w27756;
w27760 <= pi1159 and not w27758;
w27761 <= not w27759 and w27760;
w27762 <= not pi0619 and w27756;
w27763 <= pi0619 and w27716;
w27764 <= not pi1159 and not w27763;
w27765 <= not w27762 and w27764;
w27766 <= not w27761 and not w27765;
w27767 <= pi0789 and not w27766;
w27768 <= not w27757 and not w27767;
w27769 <= not w15532 and w27768;
w27770 <= w15532 and w27716;
w27771 <= not w27769 and not w27770;
w27772 <= not w15342 and not w27771;
w27773 <= w15342 and w27716;
w27774 <= not w27772 and not w27773;
w27775 <= not w18122 and w27774;
w27776 <= pi0647 and not w27732;
w27777 <= not pi0647 and not w27716;
w27778 <= not w27776 and not w27777;
w27779 <= w15364 and not w27778;
w27780 <= not w27737 and not w27779;
w27781 <= not w27775 and w27780;
w27782 <= pi0787 and not w27781;
w27783 <= w15434 and w27730;
w27784 <= not pi0626 and not w27768;
w27785 <= pi0626 and not w27716;
w27786 <= w14192 and not w27785;
w27787 <= not w27784 and w27786;
w27788 <= pi0626 and not w27768;
w27789 <= not pi0626 and not w27716;
w27790 <= w14191 and not w27789;
w27791 <= not w27788 and w27790;
w27792 <= not w27783 and not w27787;
w27793 <= not w27791 and w27792;
w27794 <= pi0788 and not w27793;
w27795 <= pi0618 and w27728;
w27796 <= pi0609 and w27727;
w27797 <= not w14731 and not w27718;
w27798 <= pi0625 and w27797;
w27799 <= w27739 and not w27797;
w27800 <= not w27798 and not w27799;
w27801 <= w27723 and not w27800;
w27802 <= not pi0608 and not w27722;
w27803 <= not w27801 and w27802;
w27804 <= pi1153 and w27739;
w27805 <= not w27798 and w27804;
w27806 <= pi0608 and not w27724;
w27807 <= not w27805 and w27806;
w27808 <= not w27803 and not w27807;
w27809 <= pi0778 and not w27808;
w27810 <= not pi0778 and not w27799;
w27811 <= not w27809 and not w27810;
w27812 <= not pi0609 and not w27811;
w27813 <= not pi1155 and not w27796;
w27814 <= not w27812 and w27813;
w27815 <= not pi0660 and not w27743;
w27816 <= not w27814 and w27815;
w27817 <= not pi0609 and w27727;
w27818 <= pi0609 and not w27811;
w27819 <= pi1155 and not w27817;
w27820 <= not w27818 and w27819;
w27821 <= pi0660 and not w27745;
w27822 <= not w27820 and w27821;
w27823 <= not w27816 and not w27822;
w27824 <= pi0785 and not w27823;
w27825 <= not pi0785 and not w27811;
w27826 <= not w27824 and not w27825;
w27827 <= not pi0618 and not w27826;
w27828 <= not pi1154 and not w27795;
w27829 <= not w27827 and w27828;
w27830 <= not pi0627 and not w27751;
w27831 <= not w27829 and w27830;
w27832 <= not pi0618 and w27728;
w27833 <= pi0618 and not w27826;
w27834 <= pi1154 and not w27832;
w27835 <= not w27833 and w27834;
w27836 <= pi0627 and not w27753;
w27837 <= not w27835 and w27836;
w27838 <= not w27831 and not w27837;
w27839 <= pi0781 and not w27838;
w27840 <= not pi0781 and not w27826;
w27841 <= not w27839 and not w27840;
w27842 <= not pi0789 and w27841;
w27843 <= not pi0619 and not w27841;
w27844 <= pi0619 and w27729;
w27845 <= not pi1159 and not w27844;
w27846 <= not w27843 and w27845;
w27847 <= not pi0648 and not w27761;
w27848 <= not w27846 and w27847;
w27849 <= pi0619 and not w27841;
w27850 <= not pi0619 and w27729;
w27851 <= pi1159 and not w27850;
w27852 <= not w27849 and w27851;
w27853 <= pi0648 and not w27765;
w27854 <= not w27852 and w27853;
w27855 <= pi0789 and not w27848;
w27856 <= not w27854 and w27855;
w27857 <= w15533 and not w27842;
w27858 <= not w27856 and w27857;
w27859 <= not w27794 and not w27858;
w27860 <= not w17927 and not w27859;
w27861 <= w15417 and not w27771;
w27862 <= w18414 and w27731;
w27863 <= not w27861 and not w27862;
w27864 <= not pi0629 and not w27863;
w27865 <= w18418 and w27731;
w27866 <= w15416 and not w27771;
w27867 <= not w27865 and not w27866;
w27868 <= pi0629 and not w27867;
w27869 <= not w27864 and not w27868;
w27870 <= pi0792 and not w27869;
w27871 <= not w17769 and not w27870;
w27872 <= not w27860 and w27871;
w27873 <= not w27782 and not w27872;
w27874 <= not pi0790 and w27873;
w27875 <= not pi0787 and not w27732;
w27876 <= pi1157 and not w27778;
w27877 <= not w27736 and not w27876;
w27878 <= pi0787 and not w27877;
w27879 <= not w27875 and not w27878;
w27880 <= not pi0644 and w27879;
w27881 <= pi0644 and w27873;
w27882 <= pi0715 and not w27880;
w27883 <= not w27881 and w27882;
w27884 <= not w15367 and not w27774;
w27885 <= w15367 and w27716;
w27886 <= not w27884 and not w27885;
w27887 <= pi0644 and not w27886;
w27888 <= not pi0644 and w27716;
w27889 <= not pi0715 and not w27888;
w27890 <= not w27887 and w27889;
w27891 <= pi1160 and not w27890;
w27892 <= not w27883 and w27891;
w27893 <= not pi0644 and not w27886;
w27894 <= pi0644 and w27716;
w27895 <= pi0715 and not w27894;
w27896 <= not w27893 and w27895;
w27897 <= pi0644 and w27879;
w27898 <= not pi0644 and w27873;
w27899 <= not pi0715 and not w27897;
w27900 <= not w27898 and w27899;
w27901 <= not pi1160 and not w27896;
w27902 <= not w27900 and w27901;
w27903 <= not w27892 and not w27902;
w27904 <= pi0790 and not w27903;
w27905 <= pi0832 and not w27874;
w27906 <= not w27904 and w27905;
w27907 <= not w27715 and not w27906;
w27908 <= pi0189 and not w14622;
w27909 <= w14198 and not w27908;
w27910 <= w14638 and not w27908;
w27911 <= pi0727 and w134;
w27912 <= not w27908 and not w27911;
w27913 <= not pi0189 and not w14204;
w27914 <= w17462 and not w27913;
w27915 <= not pi0189 and w15639;
w27916 <= pi0189 and not w15635;
w27917 <= not pi0038 and not w27915;
w27918 <= not w27916 and w27917;
w27919 <= w27911 and not w27914;
w27920 <= not w27918 and w27919;
w27921 <= not w27912 and not w27920;
w27922 <= not pi0778 and w27921;
w27923 <= not pi0625 and not w27908;
w27924 <= pi0625 and not w27921;
w27925 <= pi1153 and not w27923;
w27926 <= not w27924 and w27925;
w27927 <= not pi0625 and not w27921;
w27928 <= pi0625 and not w27908;
w27929 <= not pi1153 and not w27928;
w27930 <= not w27927 and w27929;
w27931 <= not w27926 and not w27930;
w27932 <= pi0778 and not w27931;
w27933 <= not w27922 and not w27932;
w27934 <= not w14638 and w27933;
w27935 <= not w27910 and not w27934;
w27936 <= not w14202 and w27935;
w27937 <= w14202 and w27908;
w27938 <= not w27936 and not w27937;
w27939 <= not w14198 and w27938;
w27940 <= not w27909 and not w27939;
w27941 <= not w14194 and w27940;
w27942 <= w14194 and w27908;
w27943 <= not w27941 and not w27942;
w27944 <= not pi0792 and not w27943;
w27945 <= not pi0628 and not w27908;
w27946 <= pi0628 and w27943;
w27947 <= pi1156 and not w27945;
w27948 <= not w27946 and w27947;
w27949 <= pi0628 and not w27908;
w27950 <= not pi0628 and w27943;
w27951 <= not pi1156 and not w27949;
w27952 <= not w27950 and w27951;
w27953 <= not w27948 and not w27952;
w27954 <= pi0792 and not w27953;
w27955 <= not w27944 and not w27954;
w27956 <= not pi0787 and not w27955;
w27957 <= not pi0647 and not w27908;
w27958 <= pi0647 and w27955;
w27959 <= pi1157 and not w27957;
w27960 <= not w27958 and w27959;
w27961 <= pi0647 and not w27908;
w27962 <= not pi0647 and w27955;
w27963 <= not pi1157 and not w27961;
w27964 <= not w27962 and w27963;
w27965 <= not w27960 and not w27964;
w27966 <= pi0787 and not w27965;
w27967 <= not w27956 and not w27966;
w27968 <= not pi0644 and w27967;
w27969 <= not pi0619 and not w27908;
w27970 <= w14680 and not w27908;
w27971 <= pi0189 and not w134;
w27972 <= pi0772 and w14782;
w27973 <= not w19804 and not w27972;
w27974 <= pi0039 and not w27973;
w27975 <= not pi0772 and w14521;
w27976 <= pi0772 and w14702;
w27977 <= not pi0039 and not w27975;
w27978 <= not w27976 and w27977;
w27979 <= not w27974 and not w27978;
w27980 <= pi0189 and not w27979;
w27981 <= not pi0189 and pi0772;
w27982 <= w14838 and w27981;
w27983 <= not w27980 and not w27982;
w27984 <= not pi0038 and not w27983;
w27985 <= pi0772 and w14731;
w27986 <= w14204 and not w27985;
w27987 <= pi0038 and not w27913;
w27988 <= not w27986 and w27987;
w27989 <= not w27984 and not w27988;
w27990 <= w134 and not w27989;
w27991 <= not w27971 and not w27990;
w27992 <= not w14680 and w27991;
w27993 <= not w27970 and not w27992;
w27994 <= not pi0785 and w27993;
w27995 <= not pi0609 and not w27908;
w27996 <= pi0609 and not w27993;
w27997 <= pi1155 and not w27995;
w27998 <= not w27996 and w27997;
w27999 <= not pi0609 and not w27993;
w28000 <= pi0609 and not w27908;
w28001 <= not pi1155 and not w28000;
w28002 <= not w27999 and w28001;
w28003 <= not w27998 and not w28002;
w28004 <= pi0785 and not w28003;
w28005 <= not w27994 and not w28004;
w28006 <= not pi0781 and not w28005;
w28007 <= not pi0618 and not w27908;
w28008 <= pi0618 and w28005;
w28009 <= pi1154 and not w28007;
w28010 <= not w28008 and w28009;
w28011 <= pi0618 and not w27908;
w28012 <= not pi0618 and w28005;
w28013 <= not pi1154 and not w28011;
w28014 <= not w28012 and w28013;
w28015 <= not w28010 and not w28014;
w28016 <= pi0781 and not w28015;
w28017 <= not w28006 and not w28016;
w28018 <= pi0619 and w28017;
w28019 <= pi1159 and not w27969;
w28020 <= not w28018 and w28019;
w28021 <= not pi0727 and w27989;
w28022 <= not pi0189 and not w15168;
w28023 <= pi0189 and w15109;
w28024 <= pi0772 and not w28023;
w28025 <= not w28022 and w28024;
w28026 <= pi0189 and not w14967;
w28027 <= not pi0189 and not w15048;
w28028 <= not pi0772 and not w28027;
w28029 <= not w28026 and w28028;
w28030 <= pi0039 and not w28025;
w28031 <= not w28029 and w28030;
w28032 <= not pi0189 and w15194;
w28033 <= pi0189 and w15192;
w28034 <= pi0772 and not w28032;
w28035 <= not w28033 and w28034;
w28036 <= not pi0189 and not w15188;
w28037 <= pi0189 and not w15175;
w28038 <= not pi0772 and not w28036;
w28039 <= not w28037 and w28038;
w28040 <= not pi0039 and not w28035;
w28041 <= not w28039 and w28040;
w28042 <= not pi0038 and not w28041;
w28043 <= not w28031 and w28042;
w28044 <= pi0727 and not w17033;
w28045 <= not w27988 and w28044;
w28046 <= not w28043 and w28045;
w28047 <= w134 and not w28046;
w28048 <= not w28021 and w28047;
w28049 <= not w27971 and not w28048;
w28050 <= not pi0625 and w28049;
w28051 <= pi0625 and w27991;
w28052 <= not pi1153 and not w28051;
w28053 <= not w28050 and w28052;
w28054 <= not pi0608 and not w27926;
w28055 <= not w28053 and w28054;
w28056 <= not pi0625 and w27991;
w28057 <= pi0625 and w28049;
w28058 <= pi1153 and not w28056;
w28059 <= not w28057 and w28058;
w28060 <= pi0608 and not w27930;
w28061 <= not w28059 and w28060;
w28062 <= not w28055 and not w28061;
w28063 <= pi0778 and not w28062;
w28064 <= not pi0778 and w28049;
w28065 <= not w28063 and not w28064;
w28066 <= not pi0609 and not w28065;
w28067 <= pi0609 and w27933;
w28068 <= not pi1155 and not w28067;
w28069 <= not w28066 and w28068;
w28070 <= not pi0660 and not w27998;
w28071 <= not w28069 and w28070;
w28072 <= not pi0609 and w27933;
w28073 <= pi0609 and not w28065;
w28074 <= pi1155 and not w28072;
w28075 <= not w28073 and w28074;
w28076 <= pi0660 and not w28002;
w28077 <= not w28075 and w28076;
w28078 <= not w28071 and not w28077;
w28079 <= pi0785 and not w28078;
w28080 <= not pi0785 and not w28065;
w28081 <= not w28079 and not w28080;
w28082 <= not pi0618 and not w28081;
w28083 <= pi0618 and not w27935;
w28084 <= not pi1154 and not w28083;
w28085 <= not w28082 and w28084;
w28086 <= not pi0627 and not w28010;
w28087 <= not w28085 and w28086;
w28088 <= pi0618 and not w28081;
w28089 <= not pi0618 and not w27935;
w28090 <= pi1154 and not w28089;
w28091 <= not w28088 and w28090;
w28092 <= pi0627 and not w28014;
w28093 <= not w28091 and w28092;
w28094 <= not w28087 and not w28093;
w28095 <= pi0781 and not w28094;
w28096 <= not pi0781 and not w28081;
w28097 <= not w28095 and not w28096;
w28098 <= not pi0619 and not w28097;
w28099 <= pi0619 and w27938;
w28100 <= not pi1159 and not w28099;
w28101 <= not w28098 and w28100;
w28102 <= not pi0648 and not w28020;
w28103 <= not w28101 and w28102;
w28104 <= pi0619 and not w27908;
w28105 <= not pi0619 and w28017;
w28106 <= not pi1159 and not w28104;
w28107 <= not w28105 and w28106;
w28108 <= not pi0619 and w27938;
w28109 <= pi0619 and not w28097;
w28110 <= pi1159 and not w28108;
w28111 <= not w28109 and w28110;
w28112 <= pi0648 and not w28107;
w28113 <= not w28111 and w28112;
w28114 <= not w28103 and not w28113;
w28115 <= pi0789 and not w28114;
w28116 <= not pi0789 and not w28097;
w28117 <= not w28115 and not w28116;
w28118 <= not pi0788 and w28117;
w28119 <= not pi0626 and w28117;
w28120 <= pi0626 and w27940;
w28121 <= not pi0641 and not w28120;
w28122 <= not w28119 and w28121;
w28123 <= not pi0789 and not w28017;
w28124 <= not w28020 and not w28107;
w28125 <= pi0789 and not w28124;
w28126 <= not w28123 and not w28125;
w28127 <= not pi0626 and not w28126;
w28128 <= pi0626 and w27908;
w28129 <= pi0641 and not w28128;
w28130 <= not w28127 and w28129;
w28131 <= not pi1158 and not w28130;
w28132 <= not w28122 and w28131;
w28133 <= pi0626 and w28117;
w28134 <= not pi0626 and w27940;
w28135 <= pi0641 and not w28134;
w28136 <= not w28133 and w28135;
w28137 <= pi0626 and not w28126;
w28138 <= not pi0626 and w27908;
w28139 <= not pi0641 and not w28138;
w28140 <= not w28137 and w28139;
w28141 <= pi1158 and not w28140;
w28142 <= not w28136 and w28141;
w28143 <= not w28132 and not w28142;
w28144 <= pi0788 and not w28143;
w28145 <= not w28118 and not w28144;
w28146 <= not pi0628 and w28145;
w28147 <= not w15532 and not w28126;
w28148 <= w15532 and w27908;
w28149 <= not w28147 and not w28148;
w28150 <= pi0628 and w28149;
w28151 <= not pi1156 and not w28150;
w28152 <= not w28146 and w28151;
w28153 <= not pi0629 and not w27948;
w28154 <= not w28152 and w28153;
w28155 <= pi0628 and w28145;
w28156 <= not pi0628 and w28149;
w28157 <= pi1156 and not w28156;
w28158 <= not w28155 and w28157;
w28159 <= pi0629 and not w27952;
w28160 <= not w28158 and w28159;
w28161 <= not w28154 and not w28160;
w28162 <= pi0792 and not w28161;
w28163 <= not pi0792 and w28145;
w28164 <= not w28162 and not w28163;
w28165 <= not pi0647 and not w28164;
w28166 <= not w15342 and not w28149;
w28167 <= w15342 and w27908;
w28168 <= not w28166 and not w28167;
w28169 <= pi0647 and w28168;
w28170 <= not pi1157 and not w28169;
w28171 <= not w28165 and w28170;
w28172 <= not pi0630 and not w27960;
w28173 <= not w28171 and w28172;
w28174 <= pi0647 and not w28164;
w28175 <= not pi0647 and w28168;
w28176 <= pi1157 and not w28175;
w28177 <= not w28174 and w28176;
w28178 <= pi0630 and not w27964;
w28179 <= not w28177 and w28178;
w28180 <= not w28173 and not w28179;
w28181 <= pi0787 and not w28180;
w28182 <= not pi0787 and not w28164;
w28183 <= not w28181 and not w28182;
w28184 <= pi0644 and not w28183;
w28185 <= pi0715 and not w27968;
w28186 <= not w28184 and w28185;
w28187 <= w15367 and not w27908;
w28188 <= not w15367 and w28168;
w28189 <= not w28187 and not w28188;
w28190 <= pi0644 and not w28189;
w28191 <= not pi0644 and not w27908;
w28192 <= not pi0715 and not w28191;
w28193 <= not w28190 and w28192;
w28194 <= pi1160 and not w28193;
w28195 <= not w28186 and w28194;
w28196 <= not pi0644 and not w28183;
w28197 <= pi0644 and w27967;
w28198 <= not pi0715 and not w28197;
w28199 <= not w28196 and w28198;
w28200 <= not pi0644 and not w28189;
w28201 <= pi0644 and not w27908;
w28202 <= pi0715 and not w28201;
w28203 <= not w28200 and w28202;
w28204 <= not pi1160 and not w28203;
w28205 <= not w28199 and w28204;
w28206 <= pi0790 and not w28195;
w28207 <= not w28205 and w28206;
w28208 <= not pi0790 and w28183;
w28209 <= w3868 and not w28208;
w28210 <= not w28207 and w28209;
w28211 <= not pi0189 and not w3868;
w28212 <= not pi0057 and not w28211;
w28213 <= not w28210 and w28212;
w28214 <= pi0057 and pi0189;
w28215 <= not pi0832 and not w28214;
w28216 <= not w28213 and w28215;
w28217 <= pi0189 and not w489;
w28218 <= pi0772 and w14807;
w28219 <= w14854 and w28218;
w28220 <= pi1155 and not w28217;
w28221 <= not w28219 and w28220;
w28222 <= pi0727 and w14208;
w28223 <= not w28217 and not w28222;
w28224 <= not pi0778 and w28223;
w28225 <= pi0625 and w28222;
w28226 <= not w28223 and not w28225;
w28227 <= not pi1153 and not w28226;
w28228 <= pi1153 and not w28217;
w28229 <= not w28225 and w28228;
w28230 <= not w28227 and not w28229;
w28231 <= pi0778 and not w28230;
w28232 <= not w28224 and not w28231;
w28233 <= pi0609 and w28232;
w28234 <= not w28217 and not w28218;
w28235 <= pi0727 and w15032;
w28236 <= w28234 and not w28235;
w28237 <= pi0625 and w28235;
w28238 <= not w28236 and not w28237;
w28239 <= not pi1153 and not w28238;
w28240 <= not pi0608 and not w28229;
w28241 <= not w28239 and w28240;
w28242 <= pi1153 and w28234;
w28243 <= not w28237 and w28242;
w28244 <= pi0608 and not w28227;
w28245 <= not w28243 and w28244;
w28246 <= not w28241 and not w28245;
w28247 <= pi0778 and not w28246;
w28248 <= not pi0778 and not w28236;
w28249 <= not w28247 and not w28248;
w28250 <= not pi0609 and not w28249;
w28251 <= not pi1155 and not w28233;
w28252 <= not w28250 and w28251;
w28253 <= not pi0660 and not w28221;
w28254 <= not w28252 and w28253;
w28255 <= w14859 and w28218;
w28256 <= not pi1155 and not w28217;
w28257 <= not w28255 and w28256;
w28258 <= not pi0609 and w28232;
w28259 <= pi0609 and not w28249;
w28260 <= pi1155 and not w28258;
w28261 <= not w28259 and w28260;
w28262 <= pi0660 and not w28257;
w28263 <= not w28261 and w28262;
w28264 <= not w28254 and not w28263;
w28265 <= pi0785 and not w28264;
w28266 <= not pi0785 and not w28249;
w28267 <= not w28265 and not w28266;
w28268 <= not pi0781 and not w28267;
w28269 <= not w17788 and w28218;
w28270 <= w17882 and w28269;
w28271 <= not pi1154 and not w28217;
w28272 <= not w28270 and w28271;
w28273 <= not w14638 and w28232;
w28274 <= not w28217 and not w28273;
w28275 <= not pi0618 and not w28274;
w28276 <= pi0618 and not w28267;
w28277 <= pi1154 and not w28275;
w28278 <= not w28276 and w28277;
w28279 <= pi0627 and not w28272;
w28280 <= not w28278 and w28279;
w28281 <= w17833 and w28269;
w28282 <= pi1154 and not w28217;
w28283 <= not w28281 and w28282;
w28284 <= pi0618 and not w28274;
w28285 <= not pi0618 and not w28267;
w28286 <= not pi1154 and not w28284;
w28287 <= not w28285 and w28286;
w28288 <= not pi0627 and not w28283;
w28289 <= not w28287 and w28288;
w28290 <= not w28280 and not w28289;
w28291 <= pi0781 and not w28290;
w28292 <= not w21178 and not w28268;
w28293 <= not w28291 and w28292;
w28294 <= not w17798 and w28269;
w28295 <= w17908 and w28294;
w28296 <= w14196 and not w28295;
w28297 <= w16713 and w28232;
w28298 <= not w21176 and not w28297;
w28299 <= w17898 and w28294;
w28300 <= w14195 and not w28299;
w28301 <= not w28296 and not w28300;
w28302 <= not w28298 and w28301;
w28303 <= pi0789 and not w28217;
w28304 <= not w28302 and w28303;
w28305 <= w15533 and not w28304;
w28306 <= not w28293 and w28305;
w28307 <= not w14198 and w28297;
w28308 <= not w28217 and not w28307;
w28309 <= w15428 and not w28308;
w28310 <= w17800 and w28269;
w28311 <= not pi0626 and w28310;
w28312 <= not w28217 and not w28311;
w28313 <= not pi1158 and not w28312;
w28314 <= pi0641 and not w28313;
w28315 <= not w28309 and w28314;
w28316 <= pi0626 and w28310;
w28317 <= not w28217 and not w28316;
w28318 <= pi1158 and not w28317;
w28319 <= w15429 and not w28308;
w28320 <= not pi0641 and not w28318;
w28321 <= not w28319 and w28320;
w28322 <= pi0788 and not w28315;
w28323 <= not w28321 and w28322;
w28324 <= not w17927 and not w28323;
w28325 <= not w28306 and w28324;
w28326 <= not w15532 and w28310;
w28327 <= not pi0629 and w28326;
w28328 <= pi0628 and not w28327;
w28329 <= w16714 and w28232;
w28330 <= pi0629 and not w28329;
w28331 <= not w28328 and not w28330;
w28332 <= not pi1156 and not w28331;
w28333 <= not pi0628 and not w28326;
w28334 <= pi0629 and not w28333;
w28335 <= pi0628 and w28329;
w28336 <= pi1156 and not w28334;
w28337 <= not w28335 and w28336;
w28338 <= not w28332 and not w28337;
w28339 <= pi0792 and not w28217;
w28340 <= not w28338 and w28339;
w28341 <= not w28325 and not w28340;
w28342 <= not w17769 and not w28341;
w28343 <= not w15342 and w28326;
w28344 <= not pi0630 and w28343;
w28345 <= pi0647 and not w28344;
w28346 <= not w16705 and w28329;
w28347 <= pi0630 and not w28346;
w28348 <= not w28345 and not w28347;
w28349 <= not pi1157 and not w28348;
w28350 <= pi0630 and w28343;
w28351 <= not pi0630 and not w28346;
w28352 <= pi0647 and not w28351;
w28353 <= pi1157 and not w28350;
w28354 <= not w28352 and w28353;
w28355 <= not w28349 and not w28354;
w28356 <= pi0787 and not w28217;
w28357 <= not w28355 and w28356;
w28358 <= not w28342 and not w28357;
w28359 <= not pi0790 and w28358;
w28360 <= not w15532 and w21247;
w28361 <= w28310 and w28360;
w28362 <= pi0644 and w28361;
w28363 <= not pi0715 and not w28217;
w28364 <= not w28362 and w28363;
w28365 <= not w16905 and w28346;
w28366 <= not w28217 and not w28365;
w28367 <= not pi0644 and not w28366;
w28368 <= pi0644 and w28358;
w28369 <= pi0715 and not w28367;
w28370 <= not w28368 and w28369;
w28371 <= pi1160 and not w28364;
w28372 <= not w28370 and w28371;
w28373 <= not pi0644 and w28361;
w28374 <= pi0715 and not w28217;
w28375 <= not w28373 and w28374;
w28376 <= not pi0644 and w28358;
w28377 <= pi0644 and not w28366;
w28378 <= not pi0715 and not w28377;
w28379 <= not w28376 and w28378;
w28380 <= not pi1160 and not w28375;
w28381 <= not w28379 and w28380;
w28382 <= not w28372 and not w28381;
w28383 <= pi0790 and not w28382;
w28384 <= pi0832 and not w28359;
w28385 <= not w28383 and w28384;
w28386 <= not w28216 and not w28385;
w28387 <= not pi0190 and not w489;
w28388 <= pi0699 and w14208;
w28389 <= not w28387 and not w28388;
w28390 <= not pi0778 and not w28389;
w28391 <= not pi0625 and w28388;
w28392 <= not w28389 and not w28391;
w28393 <= pi1153 and not w28392;
w28394 <= not pi1153 and not w28387;
w28395 <= not w28391 and w28394;
w28396 <= pi0778 and not w28395;
w28397 <= not w28393 and w28396;
w28398 <= not w28390 and not w28397;
w28399 <= not w15408 and not w28398;
w28400 <= not w15410 and w28399;
w28401 <= not w15412 and w28400;
w28402 <= not w15414 and w28401;
w28403 <= not w15420 and w28402;
w28404 <= not pi0647 and w28403;
w28405 <= pi0647 and w28387;
w28406 <= not pi1157 and not w28405;
w28407 <= not w28404 and w28406;
w28408 <= pi0630 and w28407;
w28409 <= pi0763 and w14807;
w28410 <= not w28387 and not w28409;
w28411 <= not w15437 and not w28410;
w28412 <= not pi0785 and not w28411;
w28413 <= w14859 and w28409;
w28414 <= w28411 and not w28413;
w28415 <= pi1155 and not w28414;
w28416 <= not pi1155 and not w28387;
w28417 <= not w28413 and w28416;
w28418 <= not w28415 and not w28417;
w28419 <= pi0785 and not w28418;
w28420 <= not w28412 and not w28419;
w28421 <= not pi0781 and not w28420;
w28422 <= not w15452 and w28420;
w28423 <= pi1154 and not w28422;
w28424 <= not w15455 and w28420;
w28425 <= not pi1154 and not w28424;
w28426 <= not w28423 and not w28425;
w28427 <= pi0781 and not w28426;
w28428 <= not w28421 and not w28427;
w28429 <= not pi0789 and not w28428;
w28430 <= not w20641 and w28428;
w28431 <= pi1159 and not w28430;
w28432 <= not w20644 and w28428;
w28433 <= not pi1159 and not w28432;
w28434 <= not w28431 and not w28433;
w28435 <= pi0789 and not w28434;
w28436 <= not w28429 and not w28435;
w28437 <= not w15532 and w28436;
w28438 <= w15532 and w28387;
w28439 <= not w28437 and not w28438;
w28440 <= not w15342 and not w28439;
w28441 <= w15342 and w28387;
w28442 <= not w28440 and not w28441;
w28443 <= not w18122 and w28442;
w28444 <= pi0647 and not w28403;
w28445 <= not pi0647 and not w28387;
w28446 <= not w28444 and not w28445;
w28447 <= w15364 and not w28446;
w28448 <= not w28408 and not w28447;
w28449 <= not w28443 and w28448;
w28450 <= pi0787 and not w28449;
w28451 <= w15434 and w28401;
w28452 <= not pi0626 and not w28436;
w28453 <= pi0626 and not w28387;
w28454 <= w14192 and not w28453;
w28455 <= not w28452 and w28454;
w28456 <= pi0626 and not w28436;
w28457 <= not pi0626 and not w28387;
w28458 <= w14191 and not w28457;
w28459 <= not w28456 and w28458;
w28460 <= not w28451 and not w28455;
w28461 <= not w28459 and w28460;
w28462 <= pi0788 and not w28461;
w28463 <= pi0618 and w28399;
w28464 <= not w14731 and not w28389;
w28465 <= pi0625 and w28464;
w28466 <= w28410 and not w28464;
w28467 <= not w28465 and not w28466;
w28468 <= w28394 and not w28467;
w28469 <= not pi0608 and not w28393;
w28470 <= not w28468 and w28469;
w28471 <= pi1153 and w28410;
w28472 <= not w28465 and w28471;
w28473 <= pi0608 and not w28395;
w28474 <= not w28472 and w28473;
w28475 <= not w28470 and not w28474;
w28476 <= pi0778 and not w28475;
w28477 <= not pi0778 and not w28466;
w28478 <= not w28476 and not w28477;
w28479 <= not pi0609 and not w28478;
w28480 <= pi0609 and not w28398;
w28481 <= not pi1155 and not w28480;
w28482 <= not w28479 and w28481;
w28483 <= not pi0660 and not w28415;
w28484 <= not w28482 and w28483;
w28485 <= pi0609 and not w28478;
w28486 <= not pi0609 and not w28398;
w28487 <= pi1155 and not w28486;
w28488 <= not w28485 and w28487;
w28489 <= pi0660 and not w28417;
w28490 <= not w28488 and w28489;
w28491 <= not w28484 and not w28490;
w28492 <= pi0785 and not w28491;
w28493 <= not pi0785 and not w28478;
w28494 <= not w28492 and not w28493;
w28495 <= not pi0618 and not w28494;
w28496 <= not pi1154 and not w28463;
w28497 <= not w28495 and w28496;
w28498 <= not pi0627 and not w28423;
w28499 <= not w28497 and w28498;
w28500 <= not pi0618 and w28399;
w28501 <= pi0618 and not w28494;
w28502 <= pi1154 and not w28500;
w28503 <= not w28501 and w28502;
w28504 <= pi0627 and not w28425;
w28505 <= not w28503 and w28504;
w28506 <= not w28499 and not w28505;
w28507 <= pi0781 and not w28506;
w28508 <= not pi0781 and not w28494;
w28509 <= not w28507 and not w28508;
w28510 <= not pi0789 and w28509;
w28511 <= not pi0619 and not w28509;
w28512 <= pi0619 and w28400;
w28513 <= not pi1159 and not w28512;
w28514 <= not w28511 and w28513;
w28515 <= not pi0648 and not w28431;
w28516 <= not w28514 and w28515;
w28517 <= pi0619 and not w28509;
w28518 <= not pi0619 and w28400;
w28519 <= pi1159 and not w28518;
w28520 <= not w28517 and w28519;
w28521 <= pi0648 and not w28433;
w28522 <= not w28520 and w28521;
w28523 <= pi0789 and not w28516;
w28524 <= not w28522 and w28523;
w28525 <= w15533 and not w28510;
w28526 <= not w28524 and w28525;
w28527 <= not w28462 and not w28526;
w28528 <= not w17927 and not w28527;
w28529 <= w15417 and not w28439;
w28530 <= w18414 and w28402;
w28531 <= not w28529 and not w28530;
w28532 <= not pi0629 and not w28531;
w28533 <= w18418 and w28402;
w28534 <= w15416 and not w28439;
w28535 <= not w28533 and not w28534;
w28536 <= pi0629 and not w28535;
w28537 <= not w28532 and not w28536;
w28538 <= pi0792 and not w28537;
w28539 <= not w17769 and not w28538;
w28540 <= not w28528 and w28539;
w28541 <= not w28450 and not w28540;
w28542 <= not pi0790 and w28541;
w28543 <= not pi0787 and not w28403;
w28544 <= pi1157 and not w28446;
w28545 <= not w28407 and not w28544;
w28546 <= pi0787 and not w28545;
w28547 <= not w28543 and not w28546;
w28548 <= not pi0644 and w28547;
w28549 <= pi0644 and w28541;
w28550 <= pi0715 and not w28548;
w28551 <= not w28549 and w28550;
w28552 <= not w15367 and not w28442;
w28553 <= w15367 and w28387;
w28554 <= not w28552 and not w28553;
w28555 <= pi0644 and not w28554;
w28556 <= not pi0644 and w28387;
w28557 <= not pi0715 and not w28556;
w28558 <= not w28555 and w28557;
w28559 <= pi1160 and not w28558;
w28560 <= not w28551 and w28559;
w28561 <= not pi0644 and not w28554;
w28562 <= pi0644 and w28387;
w28563 <= pi0715 and not w28562;
w28564 <= not w28561 and w28563;
w28565 <= pi0644 and w28547;
w28566 <= not pi0644 and w28541;
w28567 <= not pi0715 and not w28565;
w28568 <= not w28566 and w28567;
w28569 <= not pi1160 and not w28564;
w28570 <= not w28568 and w28569;
w28571 <= not w28560 and not w28570;
w28572 <= pi0790 and not w28571;
w28573 <= pi0832 and not w28542;
w28574 <= not w28572 and w28573;
w28575 <= not pi0190 and not w4989;
w28576 <= not pi0190 and not w14622;
w28577 <= w14198 and not w28576;
w28578 <= pi0190 and not w134;
w28579 <= not pi0190 and not w14204;
w28580 <= w14210 and not w28579;
w28581 <= not pi0190 and w15635;
w28582 <= pi0190 and not w15639;
w28583 <= not pi0038 and not w28582;
w28584 <= not w28581 and w28583;
w28585 <= pi0699 and not w28580;
w28586 <= not w28584 and w28585;
w28587 <= not pi0190 and not pi0699;
w28588 <= not w14615 and w28587;
w28589 <= w134 and not w28588;
w28590 <= not w28586 and w28589;
w28591 <= not w28578 and not w28590;
w28592 <= not pi0778 and not w28591;
w28593 <= not pi0625 and w28576;
w28594 <= pi0625 and w28591;
w28595 <= pi1153 and not w28593;
w28596 <= not w28594 and w28595;
w28597 <= not pi0625 and w28591;
w28598 <= pi0625 and w28576;
w28599 <= not pi1153 and not w28598;
w28600 <= not w28597 and w28599;
w28601 <= not w28596 and not w28600;
w28602 <= pi0778 and not w28601;
w28603 <= not w28592 and not w28602;
w28604 <= not w14638 and not w28603;
w28605 <= w14638 and not w28576;
w28606 <= not w28604 and not w28605;
w28607 <= not w14202 and w28606;
w28608 <= w14202 and w28576;
w28609 <= not w28607 and not w28608;
w28610 <= not w14198 and w28609;
w28611 <= not w28577 and not w28610;
w28612 <= not w14194 and w28611;
w28613 <= w14194 and w28576;
w28614 <= not w28612 and not w28613;
w28615 <= not pi0628 and not w28614;
w28616 <= pi0628 and w28576;
w28617 <= not w28615 and not w28616;
w28618 <= not pi1156 and not w28617;
w28619 <= pi0628 and not w28614;
w28620 <= not pi0628 and w28576;
w28621 <= not w28619 and not w28620;
w28622 <= pi1156 and not w28621;
w28623 <= not w28618 and not w28622;
w28624 <= pi0792 and not w28623;
w28625 <= not pi0792 and not w28614;
w28626 <= not w28624 and not w28625;
w28627 <= not pi0647 and not w28626;
w28628 <= pi0647 and w28576;
w28629 <= not w28627 and not w28628;
w28630 <= not pi1157 and not w28629;
w28631 <= pi0647 and not w28626;
w28632 <= not pi0647 and w28576;
w28633 <= not w28631 and not w28632;
w28634 <= pi1157 and not w28633;
w28635 <= not w28630 and not w28634;
w28636 <= pi0787 and not w28635;
w28637 <= not pi0787 and not w28626;
w28638 <= not w28636 and not w28637;
w28639 <= not pi0644 and not w28638;
w28640 <= pi0715 and not w28639;
w28641 <= not pi0763 and w14609;
w28642 <= pi0190 and w14836;
w28643 <= not w28641 and not w28642;
w28644 <= pi0039 and not w28643;
w28645 <= pi0763 and not w14797;
w28646 <= pi0190 and not w28645;
w28647 <= not pi0190 and pi0763;
w28648 <= w14784 and w28647;
w28649 <= not w19921 and not w28646;
w28650 <= not w28648 and w28649;
w28651 <= not w28644 and w28650;
w28652 <= not pi0038 and not w28651;
w28653 <= pi0763 and w14843;
w28654 <= pi0038 and not w28579;
w28655 <= not w28653 and w28654;
w28656 <= not w28652 and not w28655;
w28657 <= w134 and not w28656;
w28658 <= not w28578 and not w28657;
w28659 <= not w14680 and not w28658;
w28660 <= w14680 and not w28576;
w28661 <= not w28659 and not w28660;
w28662 <= not pi0785 and not w28661;
w28663 <= not w14854 and not w28576;
w28664 <= pi0609 and w28659;
w28665 <= not w28663 and not w28664;
w28666 <= pi1155 and not w28665;
w28667 <= not w14859 and not w28576;
w28668 <= not pi0609 and w28659;
w28669 <= not w28667 and not w28668;
w28670 <= not pi1155 and not w28669;
w28671 <= not w28666 and not w28670;
w28672 <= pi0785 and not w28671;
w28673 <= not w28662 and not w28672;
w28674 <= not pi0781 and not w28673;
w28675 <= not pi0618 and w28576;
w28676 <= pi0618 and w28673;
w28677 <= pi1154 and not w28675;
w28678 <= not w28676 and w28677;
w28679 <= not pi0618 and w28673;
w28680 <= pi0618 and w28576;
w28681 <= not pi1154 and not w28680;
w28682 <= not w28679 and w28681;
w28683 <= not w28678 and not w28682;
w28684 <= pi0781 and not w28683;
w28685 <= not w28674 and not w28684;
w28686 <= not pi0789 and not w28685;
w28687 <= not pi0619 and w28576;
w28688 <= pi0619 and w28685;
w28689 <= pi1159 and not w28687;
w28690 <= not w28688 and w28689;
w28691 <= not pi0619 and w28685;
w28692 <= pi0619 and w28576;
w28693 <= not pi1159 and not w28692;
w28694 <= not w28691 and w28693;
w28695 <= not w28690 and not w28694;
w28696 <= pi0789 and not w28695;
w28697 <= not w28686 and not w28696;
w28698 <= not w15532 and w28697;
w28699 <= w15532 and w28576;
w28700 <= not w28698 and not w28699;
w28701 <= not w15342 and not w28700;
w28702 <= w15342 and w28576;
w28703 <= not w28701 and not w28702;
w28704 <= not w15367 and not w28703;
w28705 <= w15367 and w28576;
w28706 <= not w28704 and not w28705;
w28707 <= pi0644 and not w28706;
w28708 <= not pi0644 and w28576;
w28709 <= not pi0715 and not w28708;
w28710 <= not w28707 and w28709;
w28711 <= pi1160 and not w28710;
w28712 <= not w28640 and w28711;
w28713 <= pi0644 and not w28638;
w28714 <= not pi0715 and not w28713;
w28715 <= not pi0644 and not w28706;
w28716 <= pi0644 and w28576;
w28717 <= pi0715 and not w28716;
w28718 <= not w28715 and w28717;
w28719 <= not pi1160 and not w28718;
w28720 <= not w28714 and w28719;
w28721 <= not w28712 and not w28720;
w28722 <= pi0790 and not w28721;
w28723 <= w15340 and w28617;
w28724 <= not w18133 and w28700;
w28725 <= w15339 and w28621;
w28726 <= not w28723 and not w28725;
w28727 <= not w28724 and w28726;
w28728 <= pi0792 and not w28727;
w28729 <= pi0609 and w28603;
w28730 <= not pi0699 and w28656;
w28731 <= not pi0763 and w21618;
w28732 <= not w15053 and not w28731;
w28733 <= not pi0039 and not w28732;
w28734 <= not pi0190 and not w28733;
w28735 <= not w15032 and not w28409;
w28736 <= pi0190 and not w28735;
w28737 <= w3847 and w28736;
w28738 <= pi0038 and not w28737;
w28739 <= not w28734 and w28738;
w28740 <= not pi0190 and not w15192;
w28741 <= pi0190 and not w15194;
w28742 <= pi0763 and not w28741;
w28743 <= not w28740 and w28742;
w28744 <= not pi0190 and w15175;
w28745 <= pi0190 and w15188;
w28746 <= not pi0763 and not w28744;
w28747 <= not w28745 and w28746;
w28748 <= not pi0039 and not w28743;
w28749 <= not w28747 and w28748;
w28750 <= pi0190 and w15168;
w28751 <= not pi0190 and not w15109;
w28752 <= pi0763 and not w28751;
w28753 <= not w28750 and w28752;
w28754 <= not pi0190 and w14967;
w28755 <= pi0190 and w15048;
w28756 <= not pi0763 and not w28755;
w28757 <= not w28754 and w28756;
w28758 <= pi0039 and not w28753;
w28759 <= not w28757 and w28758;
w28760 <= not pi0038 and not w28749;
w28761 <= not w28759 and w28760;
w28762 <= pi0699 and not w28739;
w28763 <= not w28761 and w28762;
w28764 <= w134 and not w28763;
w28765 <= not w28730 and w28764;
w28766 <= not w28578 and not w28765;
w28767 <= not pi0625 and w28766;
w28768 <= pi0625 and w28658;
w28769 <= not pi1153 and not w28768;
w28770 <= not w28767 and w28769;
w28771 <= not pi0608 and not w28596;
w28772 <= not w28770 and w28771;
w28773 <= not pi0625 and w28658;
w28774 <= pi0625 and w28766;
w28775 <= pi1153 and not w28773;
w28776 <= not w28774 and w28775;
w28777 <= pi0608 and not w28600;
w28778 <= not w28776 and w28777;
w28779 <= not w28772 and not w28778;
w28780 <= pi0778 and not w28779;
w28781 <= not pi0778 and w28766;
w28782 <= not w28780 and not w28781;
w28783 <= not pi0609 and not w28782;
w28784 <= not pi1155 and not w28729;
w28785 <= not w28783 and w28784;
w28786 <= not pi0660 and not w28666;
w28787 <= not w28785 and w28786;
w28788 <= not pi0609 and w28603;
w28789 <= pi0609 and not w28782;
w28790 <= pi1155 and not w28788;
w28791 <= not w28789 and w28790;
w28792 <= pi0660 and not w28670;
w28793 <= not w28791 and w28792;
w28794 <= not w28787 and not w28793;
w28795 <= pi0785 and not w28794;
w28796 <= not pi0785 and not w28782;
w28797 <= not w28795 and not w28796;
w28798 <= not pi0618 and not w28797;
w28799 <= pi0618 and w28606;
w28800 <= not pi1154 and not w28799;
w28801 <= not w28798 and w28800;
w28802 <= not pi0627 and not w28678;
w28803 <= not w28801 and w28802;
w28804 <= not pi0618 and w28606;
w28805 <= pi0618 and not w28797;
w28806 <= pi1154 and not w28804;
w28807 <= not w28805 and w28806;
w28808 <= pi0627 and not w28682;
w28809 <= not w28807 and w28808;
w28810 <= not w28803 and not w28809;
w28811 <= pi0781 and not w28810;
w28812 <= not pi0781 and not w28797;
w28813 <= not w28811 and not w28812;
w28814 <= not pi0789 and w28813;
w28815 <= pi0619 and not w28609;
w28816 <= not pi0619 and not w28813;
w28817 <= not pi1159 and not w28815;
w28818 <= not w28816 and w28817;
w28819 <= not pi0648 and not w28690;
w28820 <= not w28818 and w28819;
w28821 <= not pi0619 and not w28609;
w28822 <= pi0619 and not w28813;
w28823 <= pi1159 and not w28821;
w28824 <= not w28822 and w28823;
w28825 <= pi0648 and not w28694;
w28826 <= not w28824 and w28825;
w28827 <= pi0789 and not w28820;
w28828 <= not w28826 and w28827;
w28829 <= w15533 and not w28814;
w28830 <= not w28828 and w28829;
w28831 <= w15434 and w28611;
w28832 <= not pi0626 and not w28697;
w28833 <= pi0626 and not w28576;
w28834 <= w14192 and not w28833;
w28835 <= not w28832 and w28834;
w28836 <= pi0626 and not w28697;
w28837 <= not pi0626 and not w28576;
w28838 <= w14191 and not w28837;
w28839 <= not w28836 and w28838;
w28840 <= not w28831 and not w28835;
w28841 <= not w28839 and w28840;
w28842 <= pi0788 and not w28841;
w28843 <= not w17927 and not w28842;
w28844 <= not w28830 and w28843;
w28845 <= not w28728 and not w28844;
w28846 <= not w17769 and not w28845;
w28847 <= w15365 and w28629;
w28848 <= not w18122 and w28703;
w28849 <= w15364 and w28633;
w28850 <= not w28847 and not w28848;
w28851 <= not w28849 and w28850;
w28852 <= pi0787 and not w28851;
w28853 <= not pi0644 and w28719;
w28854 <= pi0644 and w28711;
w28855 <= pi0790 and not w28853;
w28856 <= not w28854 and w28855;
w28857 <= not w28846 and not w28852;
w28858 <= not w28856 and w28857;
w28859 <= not w28722 and not w28858;
w28860 <= w4989 and not w28859;
w28861 <= not pi0832 and not w28575;
w28862 <= not w28860 and w28861;
w28863 <= not w28574 and not w28862;
w28864 <= not pi0191 and not w489;
w28865 <= pi0729 and w14208;
w28866 <= not w28864 and not w28865;
w28867 <= not pi0778 and not w28866;
w28868 <= not pi0625 and w28865;
w28869 <= not w28866 and not w28868;
w28870 <= pi1153 and not w28869;
w28871 <= not pi1153 and not w28864;
w28872 <= not w28868 and w28871;
w28873 <= pi0778 and not w28872;
w28874 <= not w28870 and w28873;
w28875 <= not w28867 and not w28874;
w28876 <= not w15408 and not w28875;
w28877 <= not w15410 and w28876;
w28878 <= not w15412 and w28877;
w28879 <= not w15414 and w28878;
w28880 <= not w15420 and w28879;
w28881 <= not pi0647 and w28880;
w28882 <= pi0647 and w28864;
w28883 <= not pi1157 and not w28882;
w28884 <= not w28881 and w28883;
w28885 <= pi0630 and w28884;
w28886 <= pi0746 and w14807;
w28887 <= not w28864 and not w28886;
w28888 <= not w15437 and not w28887;
w28889 <= not pi0785 and not w28888;
w28890 <= w14859 and w28886;
w28891 <= w28888 and not w28890;
w28892 <= pi1155 and not w28891;
w28893 <= not pi1155 and not w28864;
w28894 <= not w28890 and w28893;
w28895 <= not w28892 and not w28894;
w28896 <= pi0785 and not w28895;
w28897 <= not w28889 and not w28896;
w28898 <= not pi0781 and not w28897;
w28899 <= not w15452 and w28897;
w28900 <= pi1154 and not w28899;
w28901 <= not w15455 and w28897;
w28902 <= not pi1154 and not w28901;
w28903 <= not w28900 and not w28902;
w28904 <= pi0781 and not w28903;
w28905 <= not w28898 and not w28904;
w28906 <= not pi0789 and not w28905;
w28907 <= not w20641 and w28905;
w28908 <= pi1159 and not w28907;
w28909 <= not w20644 and w28905;
w28910 <= not pi1159 and not w28909;
w28911 <= not w28908 and not w28910;
w28912 <= pi0789 and not w28911;
w28913 <= not w28906 and not w28912;
w28914 <= not w15532 and w28913;
w28915 <= w15532 and w28864;
w28916 <= not w28914 and not w28915;
w28917 <= not w15342 and not w28916;
w28918 <= w15342 and w28864;
w28919 <= not w28917 and not w28918;
w28920 <= not w18122 and w28919;
w28921 <= pi0647 and not w28880;
w28922 <= not pi0647 and not w28864;
w28923 <= not w28921 and not w28922;
w28924 <= w15364 and not w28923;
w28925 <= not w28885 and not w28924;
w28926 <= not w28920 and w28925;
w28927 <= pi0787 and not w28926;
w28928 <= w15434 and w28878;
w28929 <= not pi0626 and not w28913;
w28930 <= pi0626 and not w28864;
w28931 <= w14192 and not w28930;
w28932 <= not w28929 and w28931;
w28933 <= pi0626 and not w28913;
w28934 <= not pi0626 and not w28864;
w28935 <= w14191 and not w28934;
w28936 <= not w28933 and w28935;
w28937 <= not w28928 and not w28932;
w28938 <= not w28936 and w28937;
w28939 <= pi0788 and not w28938;
w28940 <= pi0618 and w28876;
w28941 <= not w14731 and not w28866;
w28942 <= pi0625 and w28941;
w28943 <= w28887 and not w28941;
w28944 <= not w28942 and not w28943;
w28945 <= w28871 and not w28944;
w28946 <= not pi0608 and not w28870;
w28947 <= not w28945 and w28946;
w28948 <= pi1153 and w28887;
w28949 <= not w28942 and w28948;
w28950 <= pi0608 and not w28872;
w28951 <= not w28949 and w28950;
w28952 <= not w28947 and not w28951;
w28953 <= pi0778 and not w28952;
w28954 <= not pi0778 and not w28943;
w28955 <= not w28953 and not w28954;
w28956 <= not pi0609 and not w28955;
w28957 <= pi0609 and not w28875;
w28958 <= not pi1155 and not w28957;
w28959 <= not w28956 and w28958;
w28960 <= not pi0660 and not w28892;
w28961 <= not w28959 and w28960;
w28962 <= pi0609 and not w28955;
w28963 <= not pi0609 and not w28875;
w28964 <= pi1155 and not w28963;
w28965 <= not w28962 and w28964;
w28966 <= pi0660 and not w28894;
w28967 <= not w28965 and w28966;
w28968 <= not w28961 and not w28967;
w28969 <= pi0785 and not w28968;
w28970 <= not pi0785 and not w28955;
w28971 <= not w28969 and not w28970;
w28972 <= not pi0618 and not w28971;
w28973 <= not pi1154 and not w28940;
w28974 <= not w28972 and w28973;
w28975 <= not pi0627 and not w28900;
w28976 <= not w28974 and w28975;
w28977 <= not pi0618 and w28876;
w28978 <= pi0618 and not w28971;
w28979 <= pi1154 and not w28977;
w28980 <= not w28978 and w28979;
w28981 <= pi0627 and not w28902;
w28982 <= not w28980 and w28981;
w28983 <= not w28976 and not w28982;
w28984 <= pi0781 and not w28983;
w28985 <= not pi0781 and not w28971;
w28986 <= not w28984 and not w28985;
w28987 <= not pi0789 and w28986;
w28988 <= not pi0619 and not w28986;
w28989 <= pi0619 and w28877;
w28990 <= not pi1159 and not w28989;
w28991 <= not w28988 and w28990;
w28992 <= not pi0648 and not w28908;
w28993 <= not w28991 and w28992;
w28994 <= pi0619 and not w28986;
w28995 <= not pi0619 and w28877;
w28996 <= pi1159 and not w28995;
w28997 <= not w28994 and w28996;
w28998 <= pi0648 and not w28910;
w28999 <= not w28997 and w28998;
w29000 <= pi0789 and not w28993;
w29001 <= not w28999 and w29000;
w29002 <= w15533 and not w28987;
w29003 <= not w29001 and w29002;
w29004 <= not w28939 and not w29003;
w29005 <= not w17927 and not w29004;
w29006 <= w15417 and not w28916;
w29007 <= w18414 and w28879;
w29008 <= not w29006 and not w29007;
w29009 <= not pi0629 and not w29008;
w29010 <= w18418 and w28879;
w29011 <= w15416 and not w28916;
w29012 <= not w29010 and not w29011;
w29013 <= pi0629 and not w29012;
w29014 <= not w29009 and not w29013;
w29015 <= pi0792 and not w29014;
w29016 <= not w17769 and not w29015;
w29017 <= not w29005 and w29016;
w29018 <= not w28927 and not w29017;
w29019 <= not pi0790 and w29018;
w29020 <= not pi0787 and not w28880;
w29021 <= pi1157 and not w28923;
w29022 <= not w28884 and not w29021;
w29023 <= pi0787 and not w29022;
w29024 <= not w29020 and not w29023;
w29025 <= not pi0644 and w29024;
w29026 <= pi0644 and w29018;
w29027 <= pi0715 and not w29025;
w29028 <= not w29026 and w29027;
w29029 <= not w15367 and not w28919;
w29030 <= w15367 and w28864;
w29031 <= not w29029 and not w29030;
w29032 <= pi0644 and not w29031;
w29033 <= not pi0644 and w28864;
w29034 <= not pi0715 and not w29033;
w29035 <= not w29032 and w29034;
w29036 <= pi1160 and not w29035;
w29037 <= not w29028 and w29036;
w29038 <= not pi0644 and not w29031;
w29039 <= pi0644 and w28864;
w29040 <= pi0715 and not w29039;
w29041 <= not w29038 and w29040;
w29042 <= pi0644 and w29024;
w29043 <= not pi0644 and w29018;
w29044 <= not pi0715 and not w29042;
w29045 <= not w29043 and w29044;
w29046 <= not pi1160 and not w29041;
w29047 <= not w29045 and w29046;
w29048 <= not w29037 and not w29047;
w29049 <= pi0790 and not w29048;
w29050 <= pi0832 and not w29019;
w29051 <= not w29049 and w29050;
w29052 <= not pi0191 and not w4989;
w29053 <= not pi0191 and not w14622;
w29054 <= w14198 and not w29053;
w29055 <= pi0191 and not w134;
w29056 <= not pi0191 and not w14204;
w29057 <= w14210 and not w29056;
w29058 <= not pi0191 and w15635;
w29059 <= pi0191 and not w15639;
w29060 <= not pi0038 and not w29059;
w29061 <= not w29058 and w29060;
w29062 <= pi0729 and not w29057;
w29063 <= not w29061 and w29062;
w29064 <= not pi0191 and not pi0729;
w29065 <= not w14615 and w29064;
w29066 <= w134 and not w29065;
w29067 <= not w29063 and w29066;
w29068 <= not w29055 and not w29067;
w29069 <= not pi0778 and not w29068;
w29070 <= not pi0625 and w29053;
w29071 <= pi0625 and w29068;
w29072 <= pi1153 and not w29070;
w29073 <= not w29071 and w29072;
w29074 <= not pi0625 and w29068;
w29075 <= pi0625 and w29053;
w29076 <= not pi1153 and not w29075;
w29077 <= not w29074 and w29076;
w29078 <= not w29073 and not w29077;
w29079 <= pi0778 and not w29078;
w29080 <= not w29069 and not w29079;
w29081 <= not w14638 and not w29080;
w29082 <= w14638 and not w29053;
w29083 <= not w29081 and not w29082;
w29084 <= not w14202 and w29083;
w29085 <= w14202 and w29053;
w29086 <= not w29084 and not w29085;
w29087 <= not w14198 and w29086;
w29088 <= not w29054 and not w29087;
w29089 <= not w14194 and w29088;
w29090 <= w14194 and w29053;
w29091 <= not w29089 and not w29090;
w29092 <= not pi0628 and not w29091;
w29093 <= pi0628 and w29053;
w29094 <= not w29092 and not w29093;
w29095 <= not pi1156 and not w29094;
w29096 <= pi0628 and not w29091;
w29097 <= not pi0628 and w29053;
w29098 <= not w29096 and not w29097;
w29099 <= pi1156 and not w29098;
w29100 <= not w29095 and not w29099;
w29101 <= pi0792 and not w29100;
w29102 <= not pi0792 and not w29091;
w29103 <= not w29101 and not w29102;
w29104 <= not pi0647 and not w29103;
w29105 <= pi0647 and w29053;
w29106 <= not w29104 and not w29105;
w29107 <= not pi1157 and not w29106;
w29108 <= pi0647 and not w29103;
w29109 <= not pi0647 and w29053;
w29110 <= not w29108 and not w29109;
w29111 <= pi1157 and not w29110;
w29112 <= not w29107 and not w29111;
w29113 <= pi0787 and not w29112;
w29114 <= not pi0787 and not w29103;
w29115 <= not w29113 and not w29114;
w29116 <= not pi0644 and not w29115;
w29117 <= pi0715 and not w29116;
w29118 <= not pi0746 and w14609;
w29119 <= pi0191 and w14836;
w29120 <= not w29118 and not w29119;
w29121 <= pi0039 and not w29120;
w29122 <= pi0746 and not w14797;
w29123 <= pi0191 and not w29122;
w29124 <= not pi0191 and pi0746;
w29125 <= w14784 and w29124;
w29126 <= not w20002 and not w29123;
w29127 <= not w29125 and w29126;
w29128 <= not w29121 and w29127;
w29129 <= not pi0038 and not w29128;
w29130 <= pi0746 and w14843;
w29131 <= pi0038 and not w29056;
w29132 <= not w29130 and w29131;
w29133 <= not w29129 and not w29132;
w29134 <= w134 and not w29133;
w29135 <= not w29055 and not w29134;
w29136 <= not w14680 and not w29135;
w29137 <= w14680 and not w29053;
w29138 <= not w29136 and not w29137;
w29139 <= not pi0785 and not w29138;
w29140 <= not w14854 and not w29053;
w29141 <= pi0609 and w29136;
w29142 <= not w29140 and not w29141;
w29143 <= pi1155 and not w29142;
w29144 <= not w14859 and not w29053;
w29145 <= not pi0609 and w29136;
w29146 <= not w29144 and not w29145;
w29147 <= not pi1155 and not w29146;
w29148 <= not w29143 and not w29147;
w29149 <= pi0785 and not w29148;
w29150 <= not w29139 and not w29149;
w29151 <= not pi0781 and not w29150;
w29152 <= not pi0618 and w29053;
w29153 <= pi0618 and w29150;
w29154 <= pi1154 and not w29152;
w29155 <= not w29153 and w29154;
w29156 <= not pi0618 and w29150;
w29157 <= pi0618 and w29053;
w29158 <= not pi1154 and not w29157;
w29159 <= not w29156 and w29158;
w29160 <= not w29155 and not w29159;
w29161 <= pi0781 and not w29160;
w29162 <= not w29151 and not w29161;
w29163 <= not pi0789 and not w29162;
w29164 <= not pi0619 and w29053;
w29165 <= pi0619 and w29162;
w29166 <= pi1159 and not w29164;
w29167 <= not w29165 and w29166;
w29168 <= not pi0619 and w29162;
w29169 <= pi0619 and w29053;
w29170 <= not pi1159 and not w29169;
w29171 <= not w29168 and w29170;
w29172 <= not w29167 and not w29171;
w29173 <= pi0789 and not w29172;
w29174 <= not w29163 and not w29173;
w29175 <= not w15532 and w29174;
w29176 <= w15532 and w29053;
w29177 <= not w29175 and not w29176;
w29178 <= not w15342 and not w29177;
w29179 <= w15342 and w29053;
w29180 <= not w29178 and not w29179;
w29181 <= not w15367 and not w29180;
w29182 <= w15367 and w29053;
w29183 <= not w29181 and not w29182;
w29184 <= pi0644 and not w29183;
w29185 <= not pi0644 and w29053;
w29186 <= not pi0715 and not w29185;
w29187 <= not w29184 and w29186;
w29188 <= pi1160 and not w29187;
w29189 <= not w29117 and w29188;
w29190 <= pi0644 and not w29115;
w29191 <= not pi0715 and not w29190;
w29192 <= not pi0644 and not w29183;
w29193 <= pi0644 and w29053;
w29194 <= pi0715 and not w29193;
w29195 <= not w29192 and w29194;
w29196 <= not pi1160 and not w29195;
w29197 <= not w29191 and w29196;
w29198 <= not w29189 and not w29197;
w29199 <= pi0790 and not w29198;
w29200 <= w15340 and w29094;
w29201 <= not w18133 and w29177;
w29202 <= w15339 and w29098;
w29203 <= not w29200 and not w29202;
w29204 <= not w29201 and w29203;
w29205 <= pi0792 and not w29204;
w29206 <= pi0609 and w29080;
w29207 <= not pi0729 and w29133;
w29208 <= not pi0746 and w21618;
w29209 <= not w15053 and not w29208;
w29210 <= not pi0039 and not w29209;
w29211 <= not pi0191 and not w29210;
w29212 <= not w15032 and not w28886;
w29213 <= pi0191 and not w29212;
w29214 <= w3847 and w29213;
w29215 <= pi0038 and not w29214;
w29216 <= not w29211 and w29215;
w29217 <= not pi0191 and not w15192;
w29218 <= pi0191 and not w15194;
w29219 <= pi0746 and not w29218;
w29220 <= not w29217 and w29219;
w29221 <= not pi0191 and w15175;
w29222 <= pi0191 and w15188;
w29223 <= not pi0746 and not w29221;
w29224 <= not w29222 and w29223;
w29225 <= not pi0039 and not w29220;
w29226 <= not w29224 and w29225;
w29227 <= pi0191 and w15168;
w29228 <= not pi0191 and not w15109;
w29229 <= pi0746 and not w29228;
w29230 <= not w29227 and w29229;
w29231 <= not pi0191 and w14967;
w29232 <= pi0191 and w15048;
w29233 <= not pi0746 and not w29232;
w29234 <= not w29231 and w29233;
w29235 <= pi0039 and not w29230;
w29236 <= not w29234 and w29235;
w29237 <= not pi0038 and not w29226;
w29238 <= not w29236 and w29237;
w29239 <= pi0729 and not w29216;
w29240 <= not w29238 and w29239;
w29241 <= w134 and not w29240;
w29242 <= not w29207 and w29241;
w29243 <= not w29055 and not w29242;
w29244 <= not pi0625 and w29243;
w29245 <= pi0625 and w29135;
w29246 <= not pi1153 and not w29245;
w29247 <= not w29244 and w29246;
w29248 <= not pi0608 and not w29073;
w29249 <= not w29247 and w29248;
w29250 <= not pi0625 and w29135;
w29251 <= pi0625 and w29243;
w29252 <= pi1153 and not w29250;
w29253 <= not w29251 and w29252;
w29254 <= pi0608 and not w29077;
w29255 <= not w29253 and w29254;
w29256 <= not w29249 and not w29255;
w29257 <= pi0778 and not w29256;
w29258 <= not pi0778 and w29243;
w29259 <= not w29257 and not w29258;
w29260 <= not pi0609 and not w29259;
w29261 <= not pi1155 and not w29206;
w29262 <= not w29260 and w29261;
w29263 <= not pi0660 and not w29143;
w29264 <= not w29262 and w29263;
w29265 <= not pi0609 and w29080;
w29266 <= pi0609 and not w29259;
w29267 <= pi1155 and not w29265;
w29268 <= not w29266 and w29267;
w29269 <= pi0660 and not w29147;
w29270 <= not w29268 and w29269;
w29271 <= not w29264 and not w29270;
w29272 <= pi0785 and not w29271;
w29273 <= not pi0785 and not w29259;
w29274 <= not w29272 and not w29273;
w29275 <= not pi0618 and not w29274;
w29276 <= pi0618 and w29083;
w29277 <= not pi1154 and not w29276;
w29278 <= not w29275 and w29277;
w29279 <= not pi0627 and not w29155;
w29280 <= not w29278 and w29279;
w29281 <= not pi0618 and w29083;
w29282 <= pi0618 and not w29274;
w29283 <= pi1154 and not w29281;
w29284 <= not w29282 and w29283;
w29285 <= pi0627 and not w29159;
w29286 <= not w29284 and w29285;
w29287 <= not w29280 and not w29286;
w29288 <= pi0781 and not w29287;
w29289 <= not pi0781 and not w29274;
w29290 <= not w29288 and not w29289;
w29291 <= not pi0789 and w29290;
w29292 <= pi0619 and not w29086;
w29293 <= not pi0619 and not w29290;
w29294 <= not pi1159 and not w29292;
w29295 <= not w29293 and w29294;
w29296 <= not pi0648 and not w29167;
w29297 <= not w29295 and w29296;
w29298 <= not pi0619 and not w29086;
w29299 <= pi0619 and not w29290;
w29300 <= pi1159 and not w29298;
w29301 <= not w29299 and w29300;
w29302 <= pi0648 and not w29171;
w29303 <= not w29301 and w29302;
w29304 <= pi0789 and not w29297;
w29305 <= not w29303 and w29304;
w29306 <= w15533 and not w29291;
w29307 <= not w29305 and w29306;
w29308 <= w15434 and w29088;
w29309 <= not pi0626 and not w29174;
w29310 <= pi0626 and not w29053;
w29311 <= w14192 and not w29310;
w29312 <= not w29309 and w29311;
w29313 <= pi0626 and not w29174;
w29314 <= not pi0626 and not w29053;
w29315 <= w14191 and not w29314;
w29316 <= not w29313 and w29315;
w29317 <= not w29308 and not w29312;
w29318 <= not w29316 and w29317;
w29319 <= pi0788 and not w29318;
w29320 <= not w17927 and not w29319;
w29321 <= not w29307 and w29320;
w29322 <= not w29205 and not w29321;
w29323 <= not w17769 and not w29322;
w29324 <= w15365 and w29106;
w29325 <= not w18122 and w29180;
w29326 <= w15364 and w29110;
w29327 <= not w29324 and not w29325;
w29328 <= not w29326 and w29327;
w29329 <= pi0787 and not w29328;
w29330 <= not pi0644 and w29196;
w29331 <= pi0644 and w29188;
w29332 <= pi0790 and not w29330;
w29333 <= not w29331 and w29332;
w29334 <= not w29323 and not w29329;
w29335 <= not w29333 and w29334;
w29336 <= not w29199 and not w29335;
w29337 <= w4989 and not w29336;
w29338 <= not pi0832 and not w29052;
w29339 <= not w29337 and w29338;
w29340 <= not w29051 and not w29339;
w29341 <= not pi0192 and not w489;
w29342 <= pi0691 and w14208;
w29343 <= not w29341 and not w29342;
w29344 <= not pi0778 and not w29343;
w29345 <= not pi0625 and w29342;
w29346 <= not w29343 and not w29345;
w29347 <= pi1153 and not w29346;
w29348 <= not pi1153 and not w29341;
w29349 <= not w29345 and w29348;
w29350 <= pi0778 and not w29349;
w29351 <= not w29347 and w29350;
w29352 <= not w29344 and not w29351;
w29353 <= not w15408 and not w29352;
w29354 <= not w15410 and w29353;
w29355 <= not w15412 and w29354;
w29356 <= not w15414 and w29355;
w29357 <= not w15420 and w29356;
w29358 <= not pi0647 and w29357;
w29359 <= pi0647 and w29341;
w29360 <= not pi1157 and not w29359;
w29361 <= not w29358 and w29360;
w29362 <= pi0630 and w29361;
w29363 <= pi0764 and w14807;
w29364 <= not w29341 and not w29363;
w29365 <= not w15437 and not w29364;
w29366 <= not pi0785 and not w29365;
w29367 <= w14859 and w29363;
w29368 <= w29365 and not w29367;
w29369 <= pi1155 and not w29368;
w29370 <= not pi1155 and not w29341;
w29371 <= not w29367 and w29370;
w29372 <= not w29369 and not w29371;
w29373 <= pi0785 and not w29372;
w29374 <= not w29366 and not w29373;
w29375 <= not pi0781 and not w29374;
w29376 <= not w15452 and w29374;
w29377 <= pi1154 and not w29376;
w29378 <= not w15455 and w29374;
w29379 <= not pi1154 and not w29378;
w29380 <= not w29377 and not w29379;
w29381 <= pi0781 and not w29380;
w29382 <= not w29375 and not w29381;
w29383 <= not pi0789 and not w29382;
w29384 <= not w20641 and w29382;
w29385 <= pi1159 and not w29384;
w29386 <= not w20644 and w29382;
w29387 <= not pi1159 and not w29386;
w29388 <= not w29385 and not w29387;
w29389 <= pi0789 and not w29388;
w29390 <= not w29383 and not w29389;
w29391 <= not w15532 and w29390;
w29392 <= w15532 and w29341;
w29393 <= not w29391 and not w29392;
w29394 <= not w15342 and not w29393;
w29395 <= w15342 and w29341;
w29396 <= not w29394 and not w29395;
w29397 <= not w18122 and w29396;
w29398 <= pi0647 and not w29357;
w29399 <= not pi0647 and not w29341;
w29400 <= not w29398 and not w29399;
w29401 <= w15364 and not w29400;
w29402 <= not w29362 and not w29401;
w29403 <= not w29397 and w29402;
w29404 <= pi0787 and not w29403;
w29405 <= w15434 and w29355;
w29406 <= not pi0626 and not w29390;
w29407 <= pi0626 and not w29341;
w29408 <= w14192 and not w29407;
w29409 <= not w29406 and w29408;
w29410 <= pi0626 and not w29390;
w29411 <= not pi0626 and not w29341;
w29412 <= w14191 and not w29411;
w29413 <= not w29410 and w29412;
w29414 <= not w29405 and not w29409;
w29415 <= not w29413 and w29414;
w29416 <= pi0788 and not w29415;
w29417 <= pi0618 and w29353;
w29418 <= not w14731 and not w29343;
w29419 <= pi0625 and w29418;
w29420 <= w29364 and not w29418;
w29421 <= not w29419 and not w29420;
w29422 <= w29348 and not w29421;
w29423 <= not pi0608 and not w29347;
w29424 <= not w29422 and w29423;
w29425 <= pi1153 and w29364;
w29426 <= not w29419 and w29425;
w29427 <= pi0608 and not w29349;
w29428 <= not w29426 and w29427;
w29429 <= not w29424 and not w29428;
w29430 <= pi0778 and not w29429;
w29431 <= not pi0778 and not w29420;
w29432 <= not w29430 and not w29431;
w29433 <= not pi0609 and not w29432;
w29434 <= pi0609 and not w29352;
w29435 <= not pi1155 and not w29434;
w29436 <= not w29433 and w29435;
w29437 <= not pi0660 and not w29369;
w29438 <= not w29436 and w29437;
w29439 <= pi0609 and not w29432;
w29440 <= not pi0609 and not w29352;
w29441 <= pi1155 and not w29440;
w29442 <= not w29439 and w29441;
w29443 <= pi0660 and not w29371;
w29444 <= not w29442 and w29443;
w29445 <= not w29438 and not w29444;
w29446 <= pi0785 and not w29445;
w29447 <= not pi0785 and not w29432;
w29448 <= not w29446 and not w29447;
w29449 <= not pi0618 and not w29448;
w29450 <= not pi1154 and not w29417;
w29451 <= not w29449 and w29450;
w29452 <= not pi0627 and not w29377;
w29453 <= not w29451 and w29452;
w29454 <= not pi0618 and w29353;
w29455 <= pi0618 and not w29448;
w29456 <= pi1154 and not w29454;
w29457 <= not w29455 and w29456;
w29458 <= pi0627 and not w29379;
w29459 <= not w29457 and w29458;
w29460 <= not w29453 and not w29459;
w29461 <= pi0781 and not w29460;
w29462 <= not pi0781 and not w29448;
w29463 <= not w29461 and not w29462;
w29464 <= not pi0789 and w29463;
w29465 <= not pi0619 and not w29463;
w29466 <= pi0619 and w29354;
w29467 <= not pi1159 and not w29466;
w29468 <= not w29465 and w29467;
w29469 <= not pi0648 and not w29385;
w29470 <= not w29468 and w29469;
w29471 <= pi0619 and not w29463;
w29472 <= not pi0619 and w29354;
w29473 <= pi1159 and not w29472;
w29474 <= not w29471 and w29473;
w29475 <= pi0648 and not w29387;
w29476 <= not w29474 and w29475;
w29477 <= pi0789 and not w29470;
w29478 <= not w29476 and w29477;
w29479 <= w15533 and not w29464;
w29480 <= not w29478 and w29479;
w29481 <= not w29416 and not w29480;
w29482 <= not w17927 and not w29481;
w29483 <= w15417 and not w29393;
w29484 <= w18414 and w29356;
w29485 <= not w29483 and not w29484;
w29486 <= not pi0629 and not w29485;
w29487 <= w18418 and w29356;
w29488 <= w15416 and not w29393;
w29489 <= not w29487 and not w29488;
w29490 <= pi0629 and not w29489;
w29491 <= not w29486 and not w29490;
w29492 <= pi0792 and not w29491;
w29493 <= not w17769 and not w29492;
w29494 <= not w29482 and w29493;
w29495 <= not w29404 and not w29494;
w29496 <= not pi0790 and w29495;
w29497 <= not pi0787 and not w29357;
w29498 <= pi1157 and not w29400;
w29499 <= not w29361 and not w29498;
w29500 <= pi0787 and not w29499;
w29501 <= not w29497 and not w29500;
w29502 <= not pi0644 and w29501;
w29503 <= pi0644 and w29495;
w29504 <= pi0715 and not w29502;
w29505 <= not w29503 and w29504;
w29506 <= not w15367 and not w29396;
w29507 <= w15367 and w29341;
w29508 <= not w29506 and not w29507;
w29509 <= pi0644 and not w29508;
w29510 <= not pi0644 and w29341;
w29511 <= not pi0715 and not w29510;
w29512 <= not w29509 and w29511;
w29513 <= pi1160 and not w29512;
w29514 <= not w29505 and w29513;
w29515 <= not pi0644 and not w29508;
w29516 <= pi0644 and w29341;
w29517 <= pi0715 and not w29516;
w29518 <= not w29515 and w29517;
w29519 <= pi0644 and w29501;
w29520 <= not pi0644 and w29495;
w29521 <= not pi0715 and not w29519;
w29522 <= not w29520 and w29521;
w29523 <= not pi1160 and not w29518;
w29524 <= not w29522 and w29523;
w29525 <= not w29514 and not w29524;
w29526 <= pi0790 and not w29525;
w29527 <= pi0832 and not w29496;
w29528 <= not w29526 and w29527;
w29529 <= not pi0192 and not w4989;
w29530 <= not pi0192 and not w14622;
w29531 <= w14198 and not w29530;
w29532 <= pi0192 and not w134;
w29533 <= not pi0192 and not w14204;
w29534 <= w14210 and not w29533;
w29535 <= not pi0192 and w15635;
w29536 <= pi0192 and not w15639;
w29537 <= not pi0038 and not w29536;
w29538 <= not w29535 and w29537;
w29539 <= pi0691 and not w29534;
w29540 <= not w29538 and w29539;
w29541 <= not pi0192 and not pi0691;
w29542 <= not w14615 and w29541;
w29543 <= w134 and not w29542;
w29544 <= not w29540 and w29543;
w29545 <= not w29532 and not w29544;
w29546 <= not pi0778 and not w29545;
w29547 <= not pi0625 and w29530;
w29548 <= pi0625 and w29545;
w29549 <= pi1153 and not w29547;
w29550 <= not w29548 and w29549;
w29551 <= not pi0625 and w29545;
w29552 <= pi0625 and w29530;
w29553 <= not pi1153 and not w29552;
w29554 <= not w29551 and w29553;
w29555 <= not w29550 and not w29554;
w29556 <= pi0778 and not w29555;
w29557 <= not w29546 and not w29556;
w29558 <= not w14638 and not w29557;
w29559 <= w14638 and not w29530;
w29560 <= not w29558 and not w29559;
w29561 <= not w14202 and w29560;
w29562 <= w14202 and w29530;
w29563 <= not w29561 and not w29562;
w29564 <= not w14198 and w29563;
w29565 <= not w29531 and not w29564;
w29566 <= not w14194 and w29565;
w29567 <= w14194 and w29530;
w29568 <= not w29566 and not w29567;
w29569 <= not pi0628 and not w29568;
w29570 <= pi0628 and w29530;
w29571 <= not w29569 and not w29570;
w29572 <= not pi1156 and not w29571;
w29573 <= pi0628 and not w29568;
w29574 <= not pi0628 and w29530;
w29575 <= not w29573 and not w29574;
w29576 <= pi1156 and not w29575;
w29577 <= not w29572 and not w29576;
w29578 <= pi0792 and not w29577;
w29579 <= not pi0792 and not w29568;
w29580 <= not w29578 and not w29579;
w29581 <= not pi0647 and not w29580;
w29582 <= pi0647 and w29530;
w29583 <= not w29581 and not w29582;
w29584 <= not pi1157 and not w29583;
w29585 <= pi0647 and not w29580;
w29586 <= not pi0647 and w29530;
w29587 <= not w29585 and not w29586;
w29588 <= pi1157 and not w29587;
w29589 <= not w29584 and not w29588;
w29590 <= pi0787 and not w29589;
w29591 <= not pi0787 and not w29580;
w29592 <= not w29590 and not w29591;
w29593 <= not pi0644 and not w29592;
w29594 <= pi0715 and not w29593;
w29595 <= not pi0764 and w14609;
w29596 <= pi0192 and w14836;
w29597 <= not w29595 and not w29596;
w29598 <= pi0039 and not w29597;
w29599 <= pi0764 and not w14797;
w29600 <= pi0192 and not w29599;
w29601 <= not pi0192 and pi0764;
w29602 <= w14784 and w29601;
w29603 <= not w20163 and not w29600;
w29604 <= not w29602 and w29603;
w29605 <= not w29598 and w29604;
w29606 <= not pi0038 and not w29605;
w29607 <= pi0764 and w14843;
w29608 <= pi0038 and not w29533;
w29609 <= not w29607 and w29608;
w29610 <= not w29606 and not w29609;
w29611 <= w134 and not w29610;
w29612 <= not w29532 and not w29611;
w29613 <= not w14680 and not w29612;
w29614 <= w14680 and not w29530;
w29615 <= not w29613 and not w29614;
w29616 <= not pi0785 and not w29615;
w29617 <= not w14854 and not w29530;
w29618 <= pi0609 and w29613;
w29619 <= not w29617 and not w29618;
w29620 <= pi1155 and not w29619;
w29621 <= not w14859 and not w29530;
w29622 <= not pi0609 and w29613;
w29623 <= not w29621 and not w29622;
w29624 <= not pi1155 and not w29623;
w29625 <= not w29620 and not w29624;
w29626 <= pi0785 and not w29625;
w29627 <= not w29616 and not w29626;
w29628 <= not pi0781 and not w29627;
w29629 <= not pi0618 and w29530;
w29630 <= pi0618 and w29627;
w29631 <= pi1154 and not w29629;
w29632 <= not w29630 and w29631;
w29633 <= not pi0618 and w29627;
w29634 <= pi0618 and w29530;
w29635 <= not pi1154 and not w29634;
w29636 <= not w29633 and w29635;
w29637 <= not w29632 and not w29636;
w29638 <= pi0781 and not w29637;
w29639 <= not w29628 and not w29638;
w29640 <= not pi0789 and not w29639;
w29641 <= not pi0619 and w29530;
w29642 <= pi0619 and w29639;
w29643 <= pi1159 and not w29641;
w29644 <= not w29642 and w29643;
w29645 <= not pi0619 and w29639;
w29646 <= pi0619 and w29530;
w29647 <= not pi1159 and not w29646;
w29648 <= not w29645 and w29647;
w29649 <= not w29644 and not w29648;
w29650 <= pi0789 and not w29649;
w29651 <= not w29640 and not w29650;
w29652 <= not w15532 and w29651;
w29653 <= w15532 and w29530;
w29654 <= not w29652 and not w29653;
w29655 <= not w15342 and not w29654;
w29656 <= w15342 and w29530;
w29657 <= not w29655 and not w29656;
w29658 <= not w15367 and not w29657;
w29659 <= w15367 and w29530;
w29660 <= not w29658 and not w29659;
w29661 <= pi0644 and not w29660;
w29662 <= not pi0644 and w29530;
w29663 <= not pi0715 and not w29662;
w29664 <= not w29661 and w29663;
w29665 <= pi1160 and not w29664;
w29666 <= not w29594 and w29665;
w29667 <= pi0644 and not w29592;
w29668 <= not pi0715 and not w29667;
w29669 <= not pi0644 and not w29660;
w29670 <= pi0644 and w29530;
w29671 <= pi0715 and not w29670;
w29672 <= not w29669 and w29671;
w29673 <= not pi1160 and not w29672;
w29674 <= not w29668 and w29673;
w29675 <= not w29666 and not w29674;
w29676 <= pi0790 and not w29675;
w29677 <= w15340 and w29571;
w29678 <= not w18133 and w29654;
w29679 <= w15339 and w29575;
w29680 <= not w29677 and not w29679;
w29681 <= not w29678 and w29680;
w29682 <= pi0792 and not w29681;
w29683 <= pi0609 and w29557;
w29684 <= not pi0691 and w29610;
w29685 <= not pi0764 and w21618;
w29686 <= not w15053 and not w29685;
w29687 <= not pi0039 and not w29686;
w29688 <= not pi0192 and not w29687;
w29689 <= not w15032 and not w29363;
w29690 <= pi0192 and not w29689;
w29691 <= w3847 and w29690;
w29692 <= pi0038 and not w29691;
w29693 <= not w29688 and w29692;
w29694 <= not pi0192 and not w15192;
w29695 <= pi0192 and not w15194;
w29696 <= pi0764 and not w29695;
w29697 <= not w29694 and w29696;
w29698 <= not pi0192 and w15175;
w29699 <= pi0192 and w15188;
w29700 <= not pi0764 and not w29698;
w29701 <= not w29699 and w29700;
w29702 <= not pi0039 and not w29697;
w29703 <= not w29701 and w29702;
w29704 <= pi0192 and w15168;
w29705 <= not pi0192 and not w15109;
w29706 <= pi0764 and not w29705;
w29707 <= not w29704 and w29706;
w29708 <= not pi0192 and w14967;
w29709 <= pi0192 and w15048;
w29710 <= not pi0764 and not w29709;
w29711 <= not w29708 and w29710;
w29712 <= pi0039 and not w29707;
w29713 <= not w29711 and w29712;
w29714 <= not pi0038 and not w29703;
w29715 <= not w29713 and w29714;
w29716 <= pi0691 and not w29693;
w29717 <= not w29715 and w29716;
w29718 <= w134 and not w29717;
w29719 <= not w29684 and w29718;
w29720 <= not w29532 and not w29719;
w29721 <= not pi0625 and w29720;
w29722 <= pi0625 and w29612;
w29723 <= not pi1153 and not w29722;
w29724 <= not w29721 and w29723;
w29725 <= not pi0608 and not w29550;
w29726 <= not w29724 and w29725;
w29727 <= not pi0625 and w29612;
w29728 <= pi0625 and w29720;
w29729 <= pi1153 and not w29727;
w29730 <= not w29728 and w29729;
w29731 <= pi0608 and not w29554;
w29732 <= not w29730 and w29731;
w29733 <= not w29726 and not w29732;
w29734 <= pi0778 and not w29733;
w29735 <= not pi0778 and w29720;
w29736 <= not w29734 and not w29735;
w29737 <= not pi0609 and not w29736;
w29738 <= not pi1155 and not w29683;
w29739 <= not w29737 and w29738;
w29740 <= not pi0660 and not w29620;
w29741 <= not w29739 and w29740;
w29742 <= not pi0609 and w29557;
w29743 <= pi0609 and not w29736;
w29744 <= pi1155 and not w29742;
w29745 <= not w29743 and w29744;
w29746 <= pi0660 and not w29624;
w29747 <= not w29745 and w29746;
w29748 <= not w29741 and not w29747;
w29749 <= pi0785 and not w29748;
w29750 <= not pi0785 and not w29736;
w29751 <= not w29749 and not w29750;
w29752 <= not pi0618 and not w29751;
w29753 <= pi0618 and w29560;
w29754 <= not pi1154 and not w29753;
w29755 <= not w29752 and w29754;
w29756 <= not pi0627 and not w29632;
w29757 <= not w29755 and w29756;
w29758 <= not pi0618 and w29560;
w29759 <= pi0618 and not w29751;
w29760 <= pi1154 and not w29758;
w29761 <= not w29759 and w29760;
w29762 <= pi0627 and not w29636;
w29763 <= not w29761 and w29762;
w29764 <= not w29757 and not w29763;
w29765 <= pi0781 and not w29764;
w29766 <= not pi0781 and not w29751;
w29767 <= not w29765 and not w29766;
w29768 <= not pi0789 and w29767;
w29769 <= pi0619 and not w29563;
w29770 <= not pi0619 and not w29767;
w29771 <= not pi1159 and not w29769;
w29772 <= not w29770 and w29771;
w29773 <= not pi0648 and not w29644;
w29774 <= not w29772 and w29773;
w29775 <= not pi0619 and not w29563;
w29776 <= pi0619 and not w29767;
w29777 <= pi1159 and not w29775;
w29778 <= not w29776 and w29777;
w29779 <= pi0648 and not w29648;
w29780 <= not w29778 and w29779;
w29781 <= pi0789 and not w29774;
w29782 <= not w29780 and w29781;
w29783 <= w15533 and not w29768;
w29784 <= not w29782 and w29783;
w29785 <= w15434 and w29565;
w29786 <= not pi0626 and not w29651;
w29787 <= pi0626 and not w29530;
w29788 <= w14192 and not w29787;
w29789 <= not w29786 and w29788;
w29790 <= pi0626 and not w29651;
w29791 <= not pi0626 and not w29530;
w29792 <= w14191 and not w29791;
w29793 <= not w29790 and w29792;
w29794 <= not w29785 and not w29789;
w29795 <= not w29793 and w29794;
w29796 <= pi0788 and not w29795;
w29797 <= not w17927 and not w29796;
w29798 <= not w29784 and w29797;
w29799 <= not w29682 and not w29798;
w29800 <= not w17769 and not w29799;
w29801 <= w15365 and w29583;
w29802 <= not w18122 and w29657;
w29803 <= w15364 and w29587;
w29804 <= not w29801 and not w29802;
w29805 <= not w29803 and w29804;
w29806 <= pi0787 and not w29805;
w29807 <= not pi0644 and w29673;
w29808 <= pi0644 and w29665;
w29809 <= pi0790 and not w29807;
w29810 <= not w29808 and w29809;
w29811 <= not w29800 and not w29806;
w29812 <= not w29810 and w29811;
w29813 <= not w29676 and not w29812;
w29814 <= w4989 and not w29813;
w29815 <= not pi0832 and not w29529;
w29816 <= not w29814 and w29815;
w29817 <= not w29528 and not w29816;
w29818 <= not pi0193 and not w489;
w29819 <= pi0690 and w14208;
w29820 <= not w29818 and not w29819;
w29821 <= not pi0778 and not w29820;
w29822 <= not pi0625 and w29819;
w29823 <= not w29820 and not w29822;
w29824 <= pi1153 and not w29823;
w29825 <= not pi1153 and not w29818;
w29826 <= not w29822 and w29825;
w29827 <= pi0778 and not w29826;
w29828 <= not w29824 and w29827;
w29829 <= not w29821 and not w29828;
w29830 <= not w15408 and not w29829;
w29831 <= not w15410 and w29830;
w29832 <= not w15412 and w29831;
w29833 <= not w15414 and w29832;
w29834 <= not w15420 and w29833;
w29835 <= not pi0647 and w29834;
w29836 <= pi0647 and w29818;
w29837 <= not pi1157 and not w29836;
w29838 <= not w29835 and w29837;
w29839 <= pi0630 and w29838;
w29840 <= pi0739 and w14807;
w29841 <= not w29818 and not w29840;
w29842 <= not w15437 and not w29841;
w29843 <= not pi0785 and not w29842;
w29844 <= w14859 and w29840;
w29845 <= w29842 and not w29844;
w29846 <= pi1155 and not w29845;
w29847 <= not pi1155 and not w29818;
w29848 <= not w29844 and w29847;
w29849 <= not w29846 and not w29848;
w29850 <= pi0785 and not w29849;
w29851 <= not w29843 and not w29850;
w29852 <= not pi0781 and not w29851;
w29853 <= not w15452 and w29851;
w29854 <= pi1154 and not w29853;
w29855 <= not w15455 and w29851;
w29856 <= not pi1154 and not w29855;
w29857 <= not w29854 and not w29856;
w29858 <= pi0781 and not w29857;
w29859 <= not w29852 and not w29858;
w29860 <= not pi0789 and not w29859;
w29861 <= not w20641 and w29859;
w29862 <= pi1159 and not w29861;
w29863 <= not w20644 and w29859;
w29864 <= not pi1159 and not w29863;
w29865 <= not w29862 and not w29864;
w29866 <= pi0789 and not w29865;
w29867 <= not w29860 and not w29866;
w29868 <= not w15532 and w29867;
w29869 <= w15532 and w29818;
w29870 <= not w29868 and not w29869;
w29871 <= not w15342 and not w29870;
w29872 <= w15342 and w29818;
w29873 <= not w29871 and not w29872;
w29874 <= not w18122 and w29873;
w29875 <= pi0647 and not w29834;
w29876 <= not pi0647 and not w29818;
w29877 <= not w29875 and not w29876;
w29878 <= w15364 and not w29877;
w29879 <= not w29839 and not w29878;
w29880 <= not w29874 and w29879;
w29881 <= pi0787 and not w29880;
w29882 <= w15434 and w29832;
w29883 <= not pi0626 and not w29867;
w29884 <= pi0626 and not w29818;
w29885 <= w14192 and not w29884;
w29886 <= not w29883 and w29885;
w29887 <= pi0626 and not w29867;
w29888 <= not pi0626 and not w29818;
w29889 <= w14191 and not w29888;
w29890 <= not w29887 and w29889;
w29891 <= not w29882 and not w29886;
w29892 <= not w29890 and w29891;
w29893 <= pi0788 and not w29892;
w29894 <= pi0618 and w29830;
w29895 <= not w14731 and not w29820;
w29896 <= pi0625 and w29895;
w29897 <= w29841 and not w29895;
w29898 <= not w29896 and not w29897;
w29899 <= w29825 and not w29898;
w29900 <= not pi0608 and not w29824;
w29901 <= not w29899 and w29900;
w29902 <= pi1153 and w29841;
w29903 <= not w29896 and w29902;
w29904 <= pi0608 and not w29826;
w29905 <= not w29903 and w29904;
w29906 <= not w29901 and not w29905;
w29907 <= pi0778 and not w29906;
w29908 <= not pi0778 and not w29897;
w29909 <= not w29907 and not w29908;
w29910 <= not pi0609 and not w29909;
w29911 <= pi0609 and not w29829;
w29912 <= not pi1155 and not w29911;
w29913 <= not w29910 and w29912;
w29914 <= not pi0660 and not w29846;
w29915 <= not w29913 and w29914;
w29916 <= pi0609 and not w29909;
w29917 <= not pi0609 and not w29829;
w29918 <= pi1155 and not w29917;
w29919 <= not w29916 and w29918;
w29920 <= pi0660 and not w29848;
w29921 <= not w29919 and w29920;
w29922 <= not w29915 and not w29921;
w29923 <= pi0785 and not w29922;
w29924 <= not pi0785 and not w29909;
w29925 <= not w29923 and not w29924;
w29926 <= not pi0618 and not w29925;
w29927 <= not pi1154 and not w29894;
w29928 <= not w29926 and w29927;
w29929 <= not pi0627 and not w29854;
w29930 <= not w29928 and w29929;
w29931 <= not pi0618 and w29830;
w29932 <= pi0618 and not w29925;
w29933 <= pi1154 and not w29931;
w29934 <= not w29932 and w29933;
w29935 <= pi0627 and not w29856;
w29936 <= not w29934 and w29935;
w29937 <= not w29930 and not w29936;
w29938 <= pi0781 and not w29937;
w29939 <= not pi0781 and not w29925;
w29940 <= not w29938 and not w29939;
w29941 <= not pi0789 and w29940;
w29942 <= not pi0619 and not w29940;
w29943 <= pi0619 and w29831;
w29944 <= not pi1159 and not w29943;
w29945 <= not w29942 and w29944;
w29946 <= not pi0648 and not w29862;
w29947 <= not w29945 and w29946;
w29948 <= pi0619 and not w29940;
w29949 <= not pi0619 and w29831;
w29950 <= pi1159 and not w29949;
w29951 <= not w29948 and w29950;
w29952 <= pi0648 and not w29864;
w29953 <= not w29951 and w29952;
w29954 <= pi0789 and not w29947;
w29955 <= not w29953 and w29954;
w29956 <= w15533 and not w29941;
w29957 <= not w29955 and w29956;
w29958 <= not w29893 and not w29957;
w29959 <= not w17927 and not w29958;
w29960 <= w15417 and not w29870;
w29961 <= w18414 and w29833;
w29962 <= not w29960 and not w29961;
w29963 <= not pi0629 and not w29962;
w29964 <= w18418 and w29833;
w29965 <= w15416 and not w29870;
w29966 <= not w29964 and not w29965;
w29967 <= pi0629 and not w29966;
w29968 <= not w29963 and not w29967;
w29969 <= pi0792 and not w29968;
w29970 <= not w17769 and not w29969;
w29971 <= not w29959 and w29970;
w29972 <= not w29881 and not w29971;
w29973 <= not pi0790 and w29972;
w29974 <= not pi0787 and not w29834;
w29975 <= pi1157 and not w29877;
w29976 <= not w29838 and not w29975;
w29977 <= pi0787 and not w29976;
w29978 <= not w29974 and not w29977;
w29979 <= not pi0644 and w29978;
w29980 <= pi0644 and w29972;
w29981 <= pi0715 and not w29979;
w29982 <= not w29980 and w29981;
w29983 <= not w15367 and not w29873;
w29984 <= w15367 and w29818;
w29985 <= not w29983 and not w29984;
w29986 <= pi0644 and not w29985;
w29987 <= not pi0644 and w29818;
w29988 <= not pi0715 and not w29987;
w29989 <= not w29986 and w29988;
w29990 <= pi1160 and not w29989;
w29991 <= not w29982 and w29990;
w29992 <= not pi0644 and not w29985;
w29993 <= pi0644 and w29818;
w29994 <= pi0715 and not w29993;
w29995 <= not w29992 and w29994;
w29996 <= pi0644 and w29978;
w29997 <= not pi0644 and w29972;
w29998 <= not pi0715 and not w29996;
w29999 <= not w29997 and w29998;
w30000 <= not pi1160 and not w29995;
w30001 <= not w29999 and w30000;
w30002 <= not w29991 and not w30001;
w30003 <= pi0790 and not w30002;
w30004 <= pi0832 and not w29973;
w30005 <= not w30003 and w30004;
w30006 <= not pi0193 and not w4989;
w30007 <= not pi0193 and not w14622;
w30008 <= w14198 and not w30007;
w30009 <= pi0690 and w134;
w30010 <= w30007 and not w30009;
w30011 <= not pi0193 and not w14204;
w30012 <= w14210 and not w30011;
w30013 <= pi0193 and not w15639;
w30014 <= not pi0038 and not w30013;
w30015 <= w134 and not w30014;
w30016 <= not pi0193 and w15635;
w30017 <= not w30015 and not w30016;
w30018 <= pi0690 and not w30012;
w30019 <= not w30017 and w30018;
w30020 <= not w30010 and not w30019;
w30021 <= not pi0778 and w30020;
w30022 <= not pi0625 and w30007;
w30023 <= pi0625 and not w30020;
w30024 <= pi1153 and not w30022;
w30025 <= not w30023 and w30024;
w30026 <= pi0625 and w30007;
w30027 <= not pi0625 and not w30020;
w30028 <= not pi1153 and not w30026;
w30029 <= not w30027 and w30028;
w30030 <= not w30025 and not w30029;
w30031 <= pi0778 and not w30030;
w30032 <= not w30021 and not w30031;
w30033 <= not w14638 and not w30032;
w30034 <= w14638 and not w30007;
w30035 <= not w30033 and not w30034;
w30036 <= not w14202 and w30035;
w30037 <= w14202 and w30007;
w30038 <= not w30036 and not w30037;
w30039 <= not w14198 and w30038;
w30040 <= not w30008 and not w30039;
w30041 <= not w14194 and w30040;
w30042 <= w14194 and w30007;
w30043 <= not w30041 and not w30042;
w30044 <= not pi0792 and w30043;
w30045 <= pi0628 and not w30043;
w30046 <= not pi0628 and w30007;
w30047 <= pi1156 and not w30046;
w30048 <= not w30045 and w30047;
w30049 <= pi0628 and w30007;
w30050 <= not pi0628 and not w30043;
w30051 <= not pi1156 and not w30049;
w30052 <= not w30050 and w30051;
w30053 <= not w30048 and not w30052;
w30054 <= pi0792 and not w30053;
w30055 <= not w30044 and not w30054;
w30056 <= not pi0647 and not w30055;
w30057 <= pi0647 and not w30007;
w30058 <= not w30056 and not w30057;
w30059 <= not pi1157 and w30058;
w30060 <= pi0647 and not w30055;
w30061 <= not pi0647 and not w30007;
w30062 <= not w30060 and not w30061;
w30063 <= pi1157 and w30062;
w30064 <= not w30059 and not w30063;
w30065 <= pi0787 and not w30064;
w30066 <= not pi0787 and w30055;
w30067 <= not w30065 and not w30066;
w30068 <= not pi0644 and not w30067;
w30069 <= pi0715 and not w30068;
w30070 <= pi0193 and not w134;
w30071 <= pi0739 and w14843;
w30072 <= not w30011 and not w30071;
w30073 <= pi0038 and not w30072;
w30074 <= not pi0193 and w14784;
w30075 <= pi0193 and not w14838;
w30076 <= pi0739 and not w30075;
w30077 <= not w30074 and w30076;
w30078 <= not pi0193 and not pi0739;
w30079 <= not w14611 and w30078;
w30080 <= not w30077 and not w30079;
w30081 <= not pi0038 and not w30080;
w30082 <= not w30073 and not w30081;
w30083 <= w134 and w30082;
w30084 <= not w30070 and not w30083;
w30085 <= not w14680 and not w30084;
w30086 <= w14680 and not w30007;
w30087 <= not w30085 and not w30086;
w30088 <= not pi0785 and not w30087;
w30089 <= not w14854 and not w30007;
w30090 <= pi0609 and w30085;
w30091 <= not w30089 and not w30090;
w30092 <= pi1155 and not w30091;
w30093 <= not w14859 and not w30007;
w30094 <= not pi0609 and w30085;
w30095 <= not w30093 and not w30094;
w30096 <= not pi1155 and not w30095;
w30097 <= not w30092 and not w30096;
w30098 <= pi0785 and not w30097;
w30099 <= not w30088 and not w30098;
w30100 <= not pi0781 and not w30099;
w30101 <= not pi0618 and w30007;
w30102 <= pi0618 and w30099;
w30103 <= pi1154 and not w30101;
w30104 <= not w30102 and w30103;
w30105 <= not pi0618 and w30099;
w30106 <= pi0618 and w30007;
w30107 <= not pi1154 and not w30106;
w30108 <= not w30105 and w30107;
w30109 <= not w30104 and not w30108;
w30110 <= pi0781 and not w30109;
w30111 <= not w30100 and not w30110;
w30112 <= not pi0789 and not w30111;
w30113 <= not pi0619 and w30007;
w30114 <= pi0619 and w30111;
w30115 <= pi1159 and not w30113;
w30116 <= not w30114 and w30115;
w30117 <= not pi0619 and w30111;
w30118 <= pi0619 and w30007;
w30119 <= not pi1159 and not w30118;
w30120 <= not w30117 and w30119;
w30121 <= not w30116 and not w30120;
w30122 <= pi0789 and not w30121;
w30123 <= not w30112 and not w30122;
w30124 <= not w15532 and w30123;
w30125 <= w15532 and w30007;
w30126 <= not w30124 and not w30125;
w30127 <= not w15342 and not w30126;
w30128 <= w15342 and w30007;
w30129 <= not w30127 and not w30128;
w30130 <= not w15367 and not w30129;
w30131 <= w15367 and w30007;
w30132 <= not w30130 and not w30131;
w30133 <= pi0644 and not w30132;
w30134 <= not pi0644 and w30007;
w30135 <= not pi0715 and not w30134;
w30136 <= not w30133 and w30135;
w30137 <= pi1160 and not w30136;
w30138 <= not w30069 and w30137;
w30139 <= pi0644 and not w30067;
w30140 <= not pi0715 and not w30139;
w30141 <= not pi0644 and not w30132;
w30142 <= pi0644 and w30007;
w30143 <= pi0715 and not w30142;
w30144 <= not w30141 and w30143;
w30145 <= not pi1160 and not w30144;
w30146 <= not w30140 and w30145;
w30147 <= not w30138 and not w30146;
w30148 <= pi0790 and not w30147;
w30149 <= not pi0629 and w30048;
w30150 <= not w18133 and w30126;
w30151 <= pi0629 and w30052;
w30152 <= not w30149 and not w30151;
w30153 <= not w30150 and w30152;
w30154 <= pi0792 and not w30153;
w30155 <= pi0609 and w30032;
w30156 <= not pi0690 and not w30082;
w30157 <= not pi0193 and w15192;
w30158 <= pi0193 and w15194;
w30159 <= pi0739 and not w30158;
w30160 <= not w30157 and w30159;
w30161 <= pi0193 and not w15188;
w30162 <= not pi0193 and not w15175;
w30163 <= not pi0739 and not w30161;
w30164 <= not w30162 and w30163;
w30165 <= not w30160 and not w30164;
w30166 <= not pi0039 and not w30165;
w30167 <= pi0193 and w15168;
w30168 <= not pi0193 and not w15109;
w30169 <= pi0739 and not w30168;
w30170 <= not w30167 and w30169;
w30171 <= not pi0193 and w14967;
w30172 <= pi0193 and w15048;
w30173 <= not pi0739 and not w30172;
w30174 <= not w30171 and w30173;
w30175 <= pi0039 and not w30170;
w30176 <= not w30174 and w30175;
w30177 <= not pi0038 and not w30166;
w30178 <= not w30176 and w30177;
w30179 <= not pi0739 and w21618;
w30180 <= not w15053 and not w30179;
w30181 <= not pi0039 and not w30180;
w30182 <= not pi0193 and not w30181;
w30183 <= not w15032 and not w29840;
w30184 <= pi0193 and not w30183;
w30185 <= w3847 and w30184;
w30186 <= pi0038 and not w30185;
w30187 <= not w30182 and w30186;
w30188 <= pi0690 and not w30187;
w30189 <= not w30178 and w30188;
w30190 <= w134 and not w30189;
w30191 <= not w30156 and w30190;
w30192 <= not w30070 and not w30191;
w30193 <= not pi0625 and w30192;
w30194 <= pi0625 and w30084;
w30195 <= not pi1153 and not w30194;
w30196 <= not w30193 and w30195;
w30197 <= not pi0608 and not w30025;
w30198 <= not w30196 and w30197;
w30199 <= not pi0625 and w30084;
w30200 <= pi0625 and w30192;
w30201 <= pi1153 and not w30199;
w30202 <= not w30200 and w30201;
w30203 <= pi0608 and not w30029;
w30204 <= not w30202 and w30203;
w30205 <= not w30198 and not w30204;
w30206 <= pi0778 and not w30205;
w30207 <= not pi0778 and w30192;
w30208 <= not w30206 and not w30207;
w30209 <= not pi0609 and not w30208;
w30210 <= not pi1155 and not w30155;
w30211 <= not w30209 and w30210;
w30212 <= not pi0660 and not w30092;
w30213 <= not w30211 and w30212;
w30214 <= not pi0609 and w30032;
w30215 <= pi0609 and not w30208;
w30216 <= pi1155 and not w30214;
w30217 <= not w30215 and w30216;
w30218 <= pi0660 and not w30096;
w30219 <= not w30217 and w30218;
w30220 <= not w30213 and not w30219;
w30221 <= pi0785 and not w30220;
w30222 <= not pi0785 and not w30208;
w30223 <= not w30221 and not w30222;
w30224 <= not pi0618 and not w30223;
w30225 <= pi0618 and w30035;
w30226 <= not pi1154 and not w30225;
w30227 <= not w30224 and w30226;
w30228 <= not pi0627 and not w30104;
w30229 <= not w30227 and w30228;
w30230 <= not pi0618 and w30035;
w30231 <= pi0618 and not w30223;
w30232 <= pi1154 and not w30230;
w30233 <= not w30231 and w30232;
w30234 <= pi0627 and not w30108;
w30235 <= not w30233 and w30234;
w30236 <= not w30229 and not w30235;
w30237 <= pi0781 and not w30236;
w30238 <= not pi0781 and not w30223;
w30239 <= not w30237 and not w30238;
w30240 <= not pi0789 and w30239;
w30241 <= pi0619 and not w30038;
w30242 <= not pi0619 and not w30239;
w30243 <= not pi1159 and not w30241;
w30244 <= not w30242 and w30243;
w30245 <= not pi0648 and not w30116;
w30246 <= not w30244 and w30245;
w30247 <= not pi0619 and not w30038;
w30248 <= pi0619 and not w30239;
w30249 <= pi1159 and not w30247;
w30250 <= not w30248 and w30249;
w30251 <= pi0648 and not w30120;
w30252 <= not w30250 and w30251;
w30253 <= pi0789 and not w30246;
w30254 <= not w30252 and w30253;
w30255 <= w15533 and not w30240;
w30256 <= not w30254 and w30255;
w30257 <= w15434 and w30040;
w30258 <= not pi0626 and not w30123;
w30259 <= pi0626 and not w30007;
w30260 <= w14192 and not w30259;
w30261 <= not w30258 and w30260;
w30262 <= pi0626 and not w30123;
w30263 <= not pi0626 and not w30007;
w30264 <= w14191 and not w30263;
w30265 <= not w30262 and w30264;
w30266 <= not w30257 and not w30261;
w30267 <= not w30265 and w30266;
w30268 <= pi0788 and not w30267;
w30269 <= not w17927 and not w30268;
w30270 <= not w30256 and w30269;
w30271 <= not w30154 and not w30270;
w30272 <= not w17769 and not w30271;
w30273 <= w15365 and not w30058;
w30274 <= not w18122 and w30129;
w30275 <= w15364 and not w30062;
w30276 <= not w30273 and not w30275;
w30277 <= not w30274 and w30276;
w30278 <= pi0787 and not w30277;
w30279 <= not pi0644 and w30145;
w30280 <= pi0644 and w30137;
w30281 <= pi0790 and not w30279;
w30282 <= not w30280 and w30281;
w30283 <= not w30272 and not w30278;
w30284 <= not w30282 and w30283;
w30285 <= not w30148 and not w30284;
w30286 <= w4989 and not w30285;
w30287 <= not pi0832 and not w30006;
w30288 <= not w30286 and w30287;
w30289 <= not w30005 and not w30288;
w30290 <= not pi0194 and not w14622;
w30291 <= w14198 and not w30290;
w30292 <= pi0194 and not w21948;
w30293 <= not pi0194 and w21951;
w30294 <= pi0730 and not w30293;
w30295 <= not pi0194 and not w14615;
w30296 <= not pi0730 and w30295;
w30297 <= w134 and not w30296;
w30298 <= not w30294 and w30297;
w30299 <= not w30292 and not w30298;
w30300 <= not pi0778 and not w30299;
w30301 <= not pi0625 and w30290;
w30302 <= pi0625 and w30299;
w30303 <= pi1153 and not w30301;
w30304 <= not w30302 and w30303;
w30305 <= not pi0625 and w30299;
w30306 <= pi0625 and w30290;
w30307 <= not pi1153 and not w30306;
w30308 <= not w30305 and w30307;
w30309 <= not w30304 and not w30308;
w30310 <= pi0778 and not w30309;
w30311 <= not w30300 and not w30310;
w30312 <= not w14638 and not w30311;
w30313 <= w14638 and not w30290;
w30314 <= not w30312 and not w30313;
w30315 <= not w14202 and w30314;
w30316 <= w14202 and w30290;
w30317 <= not w30315 and not w30316;
w30318 <= not w14198 and w30317;
w30319 <= not w30291 and not w30318;
w30320 <= not w14194 and w30319;
w30321 <= w14194 and w30290;
w30322 <= not w30320 and not w30321;
w30323 <= not pi0792 and w30322;
w30324 <= not pi0628 and w30290;
w30325 <= pi0628 and not w30322;
w30326 <= pi1156 and not w30324;
w30327 <= not w30325 and w30326;
w30328 <= pi0628 and w30290;
w30329 <= not pi0628 and not w30322;
w30330 <= not pi1156 and not w30328;
w30331 <= not w30329 and w30330;
w30332 <= not w30327 and not w30331;
w30333 <= pi0792 and not w30332;
w30334 <= not w30323 and not w30333;
w30335 <= not pi0787 and not w30334;
w30336 <= not pi0647 and w30290;
w30337 <= pi0647 and w30334;
w30338 <= pi1157 and not w30336;
w30339 <= not w30337 and w30338;
w30340 <= not pi0647 and w30334;
w30341 <= pi0647 and w30290;
w30342 <= not pi1157 and not w30341;
w30343 <= not w30340 and w30342;
w30344 <= not w30339 and not w30343;
w30345 <= pi0787 and not w30344;
w30346 <= not w30335 and not w30345;
w30347 <= not pi0644 and w30346;
w30348 <= not pi0618 and w30290;
w30349 <= pi0194 and not w134;
w30350 <= not pi0194 and w17002;
w30351 <= pi0194 and w22010;
w30352 <= not w30350 and not w30351;
w30353 <= pi0748 and not w30352;
w30354 <= not pi0748 and not w30295;
w30355 <= not w30353 and not w30354;
w30356 <= w134 and not w30355;
w30357 <= not w30349 and not w30356;
w30358 <= not w14680 and not w30357;
w30359 <= w14680 and not w30290;
w30360 <= not w30358 and not w30359;
w30361 <= not pi0785 and not w30360;
w30362 <= not w14854 and not w30290;
w30363 <= pi0609 and w30358;
w30364 <= not w30362 and not w30363;
w30365 <= pi1155 and not w30364;
w30366 <= not w14859 and not w30290;
w30367 <= not pi0609 and w30358;
w30368 <= not w30366 and not w30367;
w30369 <= not pi1155 and not w30368;
w30370 <= not w30365 and not w30369;
w30371 <= pi0785 and not w30370;
w30372 <= not w30361 and not w30371;
w30373 <= pi0618 and w30372;
w30374 <= pi1154 and not w30348;
w30375 <= not w30373 and w30374;
w30376 <= not pi0730 and w30355;
w30377 <= pi0194 and w17059;
w30378 <= not pi0194 and not w17051;
w30379 <= pi0748 and not w30378;
w30380 <= not w30377 and w30379;
w30381 <= pi0194 and not w22112;
w30382 <= not pi0194 and w17040;
w30383 <= not pi0748 and not w30381;
w30384 <= not w30382 and w30383;
w30385 <= pi0730 and not w30380;
w30386 <= not w30384 and w30385;
w30387 <= w134 and not w30376;
w30388 <= not w30386 and w30387;
w30389 <= not w30349 and not w30388;
w30390 <= not pi0625 and w30389;
w30391 <= pi0625 and w30357;
w30392 <= not pi1153 and not w30391;
w30393 <= not w30390 and w30392;
w30394 <= not pi0608 and not w30304;
w30395 <= not w30393 and w30394;
w30396 <= not pi0625 and w30357;
w30397 <= pi0625 and w30389;
w30398 <= pi1153 and not w30396;
w30399 <= not w30397 and w30398;
w30400 <= pi0608 and not w30308;
w30401 <= not w30399 and w30400;
w30402 <= not w30395 and not w30401;
w30403 <= pi0778 and not w30402;
w30404 <= not pi0778 and w30389;
w30405 <= not w30403 and not w30404;
w30406 <= not pi0609 and not w30405;
w30407 <= pi0609 and w30311;
w30408 <= not pi1155 and not w30407;
w30409 <= not w30406 and w30408;
w30410 <= not pi0660 and not w30365;
w30411 <= not w30409 and w30410;
w30412 <= not pi0609 and w30311;
w30413 <= pi0609 and not w30405;
w30414 <= pi1155 and not w30412;
w30415 <= not w30413 and w30414;
w30416 <= pi0660 and not w30369;
w30417 <= not w30415 and w30416;
w30418 <= not w30411 and not w30417;
w30419 <= pi0785 and not w30418;
w30420 <= not pi0785 and not w30405;
w30421 <= not w30419 and not w30420;
w30422 <= not pi0618 and not w30421;
w30423 <= pi0618 and w30314;
w30424 <= not pi1154 and not w30423;
w30425 <= not w30422 and w30424;
w30426 <= not pi0627 and not w30375;
w30427 <= not w30425 and w30426;
w30428 <= not pi0618 and w30372;
w30429 <= pi0618 and w30290;
w30430 <= not pi1154 and not w30429;
w30431 <= not w30428 and w30430;
w30432 <= not pi0618 and w30314;
w30433 <= pi0618 and not w30421;
w30434 <= pi1154 and not w30432;
w30435 <= not w30433 and w30434;
w30436 <= pi0627 and not w30431;
w30437 <= not w30435 and w30436;
w30438 <= not w30427 and not w30437;
w30439 <= pi0781 and not w30438;
w30440 <= not pi0781 and not w30421;
w30441 <= not w30439 and not w30440;
w30442 <= not pi0619 and not w30441;
w30443 <= pi0619 and not w30317;
w30444 <= not pi1159 and not w30443;
w30445 <= not w30442 and w30444;
w30446 <= not pi0619 and w30290;
w30447 <= not pi0781 and not w30372;
w30448 <= not w30375 and not w30431;
w30449 <= pi0781 and not w30448;
w30450 <= not w30447 and not w30449;
w30451 <= pi0619 and w30450;
w30452 <= pi1159 and not w30446;
w30453 <= not w30451 and w30452;
w30454 <= not pi0648 and not w30453;
w30455 <= not w30445 and w30454;
w30456 <= pi0619 and not w30441;
w30457 <= not pi0619 and not w30317;
w30458 <= pi1159 and not w30457;
w30459 <= not w30456 and w30458;
w30460 <= not pi0619 and w30450;
w30461 <= pi0619 and w30290;
w30462 <= not pi1159 and not w30461;
w30463 <= not w30460 and w30462;
w30464 <= pi0648 and not w30463;
w30465 <= not w30459 and w30464;
w30466 <= not w30455 and not w30465;
w30467 <= pi0789 and not w30466;
w30468 <= not pi0789 and not w30441;
w30469 <= not w30467 and not w30468;
w30470 <= not pi0788 and w30469;
w30471 <= not pi0626 and w30469;
w30472 <= pi0626 and not w30319;
w30473 <= not pi0641 and not w30472;
w30474 <= not w30471 and w30473;
w30475 <= not pi0789 and not w30450;
w30476 <= not w30453 and not w30463;
w30477 <= pi0789 and not w30476;
w30478 <= not w30475 and not w30477;
w30479 <= not pi0626 and not w30478;
w30480 <= pi0626 and not w30290;
w30481 <= pi0641 and not w30480;
w30482 <= not w30479 and w30481;
w30483 <= not pi1158 and not w30482;
w30484 <= not w30474 and w30483;
w30485 <= pi0626 and w30469;
w30486 <= not pi0626 and not w30319;
w30487 <= pi0641 and not w30486;
w30488 <= not w30485 and w30487;
w30489 <= pi0626 and not w30478;
w30490 <= not pi0626 and not w30290;
w30491 <= not pi0641 and not w30490;
w30492 <= not w30489 and w30491;
w30493 <= pi1158 and not w30492;
w30494 <= not w30488 and w30493;
w30495 <= not w30484 and not w30494;
w30496 <= pi0788 and not w30495;
w30497 <= not w30470 and not w30496;
w30498 <= not pi0628 and w30497;
w30499 <= not w15532 and w30478;
w30500 <= w15532 and w30290;
w30501 <= not w30499 and not w30500;
w30502 <= pi0628 and not w30501;
w30503 <= not pi1156 and not w30502;
w30504 <= not w30498 and w30503;
w30505 <= not pi0629 and not w30327;
w30506 <= not w30504 and w30505;
w30507 <= pi0628 and w30497;
w30508 <= not pi0628 and not w30501;
w30509 <= pi1156 and not w30508;
w30510 <= not w30507 and w30509;
w30511 <= pi0629 and not w30331;
w30512 <= not w30510 and w30511;
w30513 <= not w30506 and not w30512;
w30514 <= pi0792 and not w30513;
w30515 <= not pi0792 and w30497;
w30516 <= not w30514 and not w30515;
w30517 <= not pi0647 and not w30516;
w30518 <= not w15342 and not w30501;
w30519 <= w15342 and w30290;
w30520 <= not w30518 and not w30519;
w30521 <= pi0647 and not w30520;
w30522 <= not pi1157 and not w30521;
w30523 <= not w30517 and w30522;
w30524 <= not pi0630 and not w30339;
w30525 <= not w30523 and w30524;
w30526 <= pi0647 and not w30516;
w30527 <= not pi0647 and not w30520;
w30528 <= pi1157 and not w30527;
w30529 <= not w30526 and w30528;
w30530 <= pi0630 and not w30343;
w30531 <= not w30529 and w30530;
w30532 <= not w30525 and not w30531;
w30533 <= pi0787 and not w30532;
w30534 <= not pi0787 and not w30516;
w30535 <= not w30533 and not w30534;
w30536 <= pi0644 and not w30535;
w30537 <= pi0715 and not w30347;
w30538 <= not w30536 and w30537;
w30539 <= w15367 and not w30290;
w30540 <= not w15367 and w30520;
w30541 <= not w30539 and not w30540;
w30542 <= pi0644 and w30541;
w30543 <= not pi0644 and w30290;
w30544 <= not pi0715 and not w30543;
w30545 <= not w30542 and w30544;
w30546 <= pi1160 and not w30545;
w30547 <= not w30538 and w30546;
w30548 <= not pi0644 and not w30535;
w30549 <= pi0644 and w30346;
w30550 <= not pi0715 and not w30549;
w30551 <= not w30548 and w30550;
w30552 <= not pi0644 and w30541;
w30553 <= pi0644 and w30290;
w30554 <= pi0715 and not w30553;
w30555 <= not w30552 and w30554;
w30556 <= not pi1160 and not w30555;
w30557 <= not w30551 and w30556;
w30558 <= pi0790 and not w30547;
w30559 <= not w30557 and w30558;
w30560 <= not pi0790 and w30535;
w30561 <= w4989 and not w30560;
w30562 <= not w30559 and w30561;
w30563 <= not pi0194 and not w4989;
w30564 <= not pi0832 and not w30563;
w30565 <= not w30562 and w30564;
w30566 <= not pi0194 and not w489;
w30567 <= pi0730 and w14208;
w30568 <= not w30566 and not w30567;
w30569 <= not pi0778 and w30568;
w30570 <= not pi0625 and w30567;
w30571 <= not w30568 and not w30570;
w30572 <= pi1153 and not w30571;
w30573 <= not pi1153 and not w30566;
w30574 <= not w30570 and w30573;
w30575 <= not w30572 and not w30574;
w30576 <= pi0778 and not w30575;
w30577 <= not w30569 and not w30576;
w30578 <= not w15408 and w30577;
w30579 <= not w15410 and w30578;
w30580 <= not w15412 and w30579;
w30581 <= not w15414 and w30580;
w30582 <= not w15420 and w30581;
w30583 <= not pi0647 and w30582;
w30584 <= pi0647 and w30566;
w30585 <= not pi1157 and not w30584;
w30586 <= not w30583 and w30585;
w30587 <= pi0630 and w30586;
w30588 <= pi0748 and w14807;
w30589 <= not w30566 and not w30588;
w30590 <= not w15437 and not w30589;
w30591 <= not pi0785 and not w30590;
w30592 <= not w15442 and not w30589;
w30593 <= pi1155 and not w30592;
w30594 <= not w15445 and w30590;
w30595 <= not pi1155 and not w30594;
w30596 <= not w30593 and not w30595;
w30597 <= pi0785 and not w30596;
w30598 <= not w30591 and not w30597;
w30599 <= not pi0781 and not w30598;
w30600 <= not w15452 and w30598;
w30601 <= pi1154 and not w30600;
w30602 <= not w15455 and w30598;
w30603 <= not pi1154 and not w30602;
w30604 <= not w30601 and not w30603;
w30605 <= pi0781 and not w30604;
w30606 <= not w30599 and not w30605;
w30607 <= not pi0789 and not w30606;
w30608 <= not pi0619 and w30566;
w30609 <= pi0619 and w30606;
w30610 <= pi1159 and not w30608;
w30611 <= not w30609 and w30610;
w30612 <= not pi0619 and w30606;
w30613 <= pi0619 and w30566;
w30614 <= not pi1159 and not w30613;
w30615 <= not w30612 and w30614;
w30616 <= not w30611 and not w30615;
w30617 <= pi0789 and not w30616;
w30618 <= not w30607 and not w30617;
w30619 <= not w15532 and w30618;
w30620 <= w15532 and w30566;
w30621 <= not w30619 and not w30620;
w30622 <= not w15342 and not w30621;
w30623 <= w15342 and w30566;
w30624 <= not w30622 and not w30623;
w30625 <= not w18122 and w30624;
w30626 <= pi0647 and not w30582;
w30627 <= not pi0647 and not w30566;
w30628 <= not w30626 and not w30627;
w30629 <= w15364 and not w30628;
w30630 <= not w30587 and not w30629;
w30631 <= not w30625 and w30630;
w30632 <= pi0787 and not w30631;
w30633 <= w15434 and w30580;
w30634 <= not pi0626 and not w30618;
w30635 <= pi0626 and not w30566;
w30636 <= w14192 and not w30635;
w30637 <= not w30634 and w30636;
w30638 <= pi0626 and not w30618;
w30639 <= not pi0626 and not w30566;
w30640 <= w14191 and not w30639;
w30641 <= not w30638 and w30640;
w30642 <= not w30633 and not w30637;
w30643 <= not w30641 and w30642;
w30644 <= pi0788 and not w30643;
w30645 <= pi0618 and w30578;
w30646 <= pi0609 and w30577;
w30647 <= not w14731 and not w30568;
w30648 <= pi0625 and w30647;
w30649 <= w30589 and not w30647;
w30650 <= not w30648 and not w30649;
w30651 <= w30573 and not w30650;
w30652 <= not pi0608 and not w30572;
w30653 <= not w30651 and w30652;
w30654 <= pi1153 and w30589;
w30655 <= not w30648 and w30654;
w30656 <= pi0608 and not w30574;
w30657 <= not w30655 and w30656;
w30658 <= not w30653 and not w30657;
w30659 <= pi0778 and not w30658;
w30660 <= not pi0778 and not w30649;
w30661 <= not w30659 and not w30660;
w30662 <= not pi0609 and not w30661;
w30663 <= not pi1155 and not w30646;
w30664 <= not w30662 and w30663;
w30665 <= not pi0660 and not w30593;
w30666 <= not w30664 and w30665;
w30667 <= not pi0609 and w30577;
w30668 <= pi0609 and not w30661;
w30669 <= pi1155 and not w30667;
w30670 <= not w30668 and w30669;
w30671 <= pi0660 and not w30595;
w30672 <= not w30670 and w30671;
w30673 <= not w30666 and not w30672;
w30674 <= pi0785 and not w30673;
w30675 <= not pi0785 and not w30661;
w30676 <= not w30674 and not w30675;
w30677 <= not pi0618 and not w30676;
w30678 <= not pi1154 and not w30645;
w30679 <= not w30677 and w30678;
w30680 <= not pi0627 and not w30601;
w30681 <= not w30679 and w30680;
w30682 <= not pi0618 and w30578;
w30683 <= pi0618 and not w30676;
w30684 <= pi1154 and not w30682;
w30685 <= not w30683 and w30684;
w30686 <= pi0627 and not w30603;
w30687 <= not w30685 and w30686;
w30688 <= not w30681 and not w30687;
w30689 <= pi0781 and not w30688;
w30690 <= not pi0781 and not w30676;
w30691 <= not w30689 and not w30690;
w30692 <= not pi0789 and w30691;
w30693 <= not pi0619 and not w30691;
w30694 <= pi0619 and w30579;
w30695 <= not pi1159 and not w30694;
w30696 <= not w30693 and w30695;
w30697 <= not pi0648 and not w30611;
w30698 <= not w30696 and w30697;
w30699 <= pi0619 and not w30691;
w30700 <= not pi0619 and w30579;
w30701 <= pi1159 and not w30700;
w30702 <= not w30699 and w30701;
w30703 <= pi0648 and not w30615;
w30704 <= not w30702 and w30703;
w30705 <= pi0789 and not w30698;
w30706 <= not w30704 and w30705;
w30707 <= w15533 and not w30692;
w30708 <= not w30706 and w30707;
w30709 <= not w30644 and not w30708;
w30710 <= not w17927 and not w30709;
w30711 <= w15417 and not w30621;
w30712 <= w18414 and w30581;
w30713 <= not w30711 and not w30712;
w30714 <= not pi0629 and not w30713;
w30715 <= w18418 and w30581;
w30716 <= w15416 and not w30621;
w30717 <= not w30715 and not w30716;
w30718 <= pi0629 and not w30717;
w30719 <= not w30714 and not w30718;
w30720 <= pi0792 and not w30719;
w30721 <= not w17769 and not w30720;
w30722 <= not w30710 and w30721;
w30723 <= not w30632 and not w30722;
w30724 <= not pi0790 and w30723;
w30725 <= not pi0787 and not w30582;
w30726 <= pi1157 and not w30628;
w30727 <= not w30586 and not w30726;
w30728 <= pi0787 and not w30727;
w30729 <= not w30725 and not w30728;
w30730 <= not pi0644 and w30729;
w30731 <= pi0644 and w30723;
w30732 <= pi0715 and not w30730;
w30733 <= not w30731 and w30732;
w30734 <= not w15367 and not w30624;
w30735 <= w15367 and w30566;
w30736 <= not w30734 and not w30735;
w30737 <= pi0644 and not w30736;
w30738 <= not pi0644 and w30566;
w30739 <= not pi0715 and not w30738;
w30740 <= not w30737 and w30739;
w30741 <= pi1160 and not w30740;
w30742 <= not w30733 and w30741;
w30743 <= not pi0644 and not w30736;
w30744 <= pi0644 and w30566;
w30745 <= pi0715 and not w30744;
w30746 <= not w30743 and w30745;
w30747 <= pi0644 and w30729;
w30748 <= not pi0644 and w30723;
w30749 <= not pi0715 and not w30747;
w30750 <= not w30748 and w30749;
w30751 <= not pi1160 and not w30746;
w30752 <= not w30750 and w30751;
w30753 <= not w30742 and not w30752;
w30754 <= pi0790 and not w30753;
w30755 <= pi0832 and not w30724;
w30756 <= not w30754 and w30755;
w30757 <= not w30565 and not w30756;
w30758 <= not pi0138 and w14128;
w30759 <= not pi0196 and w30758;
w30760 <= pi0195 and not w30759;
w30761 <= not w9040 and w13756;
w30762 <= not w3761 and w13731;
w30763 <= w13730 and not w14056;
w30764 <= not w9043 and not w30762;
w30765 <= not w30761 and not w30763;
w30766 <= w30764 and w30765;
w30767 <= pi0232 and not w30766;
w30768 <= not w14054 and not w30767;
w30769 <= pi0039 and not w30768;
w30770 <= w11473 and not w13733;
w30771 <= not pi0039 and not w30770;
w30772 <= w7763 and not w30760;
w30773 <= not w30771 and w30772;
w30774 <= not w30769 and w30773;
w30775 <= not pi0171 and w6889;
w30776 <= not w14085 and not w30775;
w30777 <= w6599 and not w30776;
w30778 <= w6854 and not w30777;
w30779 <= not pi0192 and w14074;
w30780 <= pi0192 and w14083;
w30781 <= not w30778 and not w30779;
w30782 <= not w30780 and w30781;
w30783 <= pi0232 and not w30782;
w30784 <= not w14080 and not w30783;
w30785 <= pi0039 and not w30784;
w30786 <= pi0192 and w14102;
w30787 <= not w7168 and not w13725;
w30788 <= pi0171 and w11300;
w30789 <= not w30787 and not w30788;
w30790 <= pi0299 and not w30789;
w30791 <= not pi0192 and w14096;
w30792 <= pi0232 and not w30791;
w30793 <= not w30786 and w30792;
w30794 <= not w30790 and w30793;
w30795 <= w14099 and not w30794;
w30796 <= w171 and not w30785;
w30797 <= not w30795 and w30796;
w30798 <= not pi0087 and not w30797;
w30799 <= w14071 and not w30798;
w30800 <= not pi0092 and not w30799;
w30801 <= w14070 and not w30800;
w30802 <= not pi0055 and not w30801;
w30803 <= not w14122 and not w30802;
w30804 <= w92 and not w30803;
w30805 <= w7446 and w30760;
w30806 <= not w30804 and w30805;
w30807 <= not w30774 and not w30806;
w30808 <= w10695 and w14055;
w30809 <= not pi0170 and w6602;
w30810 <= not w14055 and not w30809;
w30811 <= w10693 and not w30810;
w30812 <= pi0232 and not w30808;
w30813 <= not w30811 and w30812;
w30814 <= not w14054 and not w30813;
w30815 <= pi0039 and not w30814;
w30816 <= w11473 and w13850;
w30817 <= not pi0039 and not w30816;
w30818 <= not pi0038 and not w30817;
w30819 <= not w30815 and w30818;
w30820 <= pi0194 and not w30819;
w30821 <= pi0299 and not w30814;
w30822 <= not w9041 and not w30821;
w30823 <= pi0039 and not w30822;
w30824 <= w11473 and not w13838;
w30825 <= not pi0039 and not w30824;
w30826 <= not pi0038 and not w30825;
w30827 <= not w30823 and w30826;
w30828 <= not pi0194 and not w30827;
w30829 <= w7760 and not w30820;
w30830 <= not w30828 and w30829;
w30831 <= not pi0196 and not w30830;
w30832 <= not pi0170 and w6889;
w30833 <= not w14085 and not w30832;
w30834 <= w6599 and not w30833;
w30835 <= w6854 and not w30834;
w30836 <= not w14074 and not w30835;
w30837 <= pi0232 and not w30836;
w30838 <= not w14080 and not w30837;
w30839 <= pi0232 and w14083;
w30840 <= w30838 and not w30839;
w30841 <= pi0039 and not w30840;
w30842 <= not pi0038 and pi0194;
w30843 <= not w30841 and w30842;
w30844 <= pi0039 and not w30838;
w30845 <= not pi0038 and not pi0194;
w30846 <= not w30844 and w30845;
w30847 <= not w30843 and not w30846;
w30848 <= not w14099 and not w30847;
w30849 <= not w7168 and not w13837;
w30850 <= pi0170 and w11300;
w30851 <= not w30849 and not w30850;
w30852 <= pi0299 and not w30851;
w30853 <= not w14102 and w30843;
w30854 <= not w14096 and w30846;
w30855 <= not w30853 and not w30854;
w30856 <= pi0232 and not w30852;
w30857 <= not w30855 and w30856;
w30858 <= not w30848 and not w30857;
w30859 <= not pi0100 and not w30858;
w30860 <= not pi0087 and not w30859;
w30861 <= w14071 and not w30860;
w30862 <= not pi0092 and not w30861;
w30863 <= w14070 and not w30862;
w30864 <= not pi0055 and not w30863;
w30865 <= not w14122 and not w30864;
w30866 <= w92 and not w30865;
w30867 <= w7446 and not w30866;
w30868 <= pi0196 and not w30867;
w30869 <= not w30758 and not w30831;
w30870 <= not w30868 and w30869;
w30871 <= pi0195 and not pi0196;
w30872 <= not w30830 and not w30871;
w30873 <= not w30867 and w30871;
w30874 <= w30758 and not w30872;
w30875 <= not w30873 and w30874;
w30876 <= not w30870 and not w30875;
w30877 <= not pi0197 and not w489;
w30878 <= not pi0767 and pi0947;
w30879 <= not pi0698 and w18465;
w30880 <= not w30878 and not w30879;
w30881 <= w489 and not w30880;
w30882 <= pi0832 and not w30877;
w30883 <= not w30881 and w30882;
w30884 <= not pi0197 and not w7760;
w30885 <= w14204 and not w30878;
w30886 <= pi0197 and not w14613;
w30887 <= pi0038 and not w30885;
w30888 <= not w30886 and w30887;
w30889 <= not pi0197 and not w14521;
w30890 <= w14521 and w30878;
w30891 <= not pi0039 and not w30889;
w30892 <= not w30890 and w30891;
w30893 <= not pi0197 and not w18564;
w30894 <= pi0197 and not w18725;
w30895 <= pi0299 and not w30894;
w30896 <= not w30893 and w30895;
w30897 <= not pi0197 and not w14587;
w30898 <= w18582 and not w30897;
w30899 <= not pi0767 and not w30898;
w30900 <= not w30896 and w30899;
w30901 <= not pi0197 and pi0767;
w30902 <= not w14609 and w30901;
w30903 <= pi0039 and not w30902;
w30904 <= not w30900 and w30903;
w30905 <= not pi0038 and not w30892;
w30906 <= not w30904 and w30905;
w30907 <= not w30888 and not w30906;
w30908 <= pi0698 and not w30907;
w30909 <= not w18677 and w30892;
w30910 <= w18674 and not w30897;
w30911 <= pi0197 and w18671;
w30912 <= not pi0197 and w18655;
w30913 <= pi0299 and not w30911;
w30914 <= not w30912 and w30913;
w30915 <= pi0767 and not w30910;
w30916 <= not w30914 and w30915;
w30917 <= not pi0197 and w18627;
w30918 <= pi0197 and w18643;
w30919 <= not pi0767 and not w30918;
w30920 <= not w30917 and w30919;
w30921 <= pi0039 and not w30916;
w30922 <= not w30920 and w30921;
w30923 <= not w30909 and not w30922;
w30924 <= not pi0038 and not w30923;
w30925 <= not pi0197 and not w14204;
w30926 <= pi0767 and pi0947;
w30927 <= not pi0039 and not w30926;
w30928 <= w18802 and w30927;
w30929 <= pi0038 and not w30925;
w30930 <= not w30928 and w30929;
w30931 <= not pi0698 and not w30930;
w30932 <= not w30924 and w30931;
w30933 <= not w30908 and not w30932;
w30934 <= w7760 and not w30933;
w30935 <= not pi0832 and not w30884;
w30936 <= not w30934 and w30935;
w30937 <= not w30883 and not w30936;
w30938 <= w93 and not w14521;
w30939 <= w16154 and not w30938;
w30940 <= pi0198 and not w30939;
w30941 <= pi0198 and not w14360;
w30942 <= pi0198 and not w14216;
w30943 <= w3759 and not w30942;
w30944 <= w30941 and not w30943;
w30945 <= w3755 and not w14284;
w30946 <= not w3755 and not w14286;
w30947 <= pi0198 and not w30945;
w30948 <= not w30946 and w30947;
w30949 <= not w3805 and w30948;
w30950 <= not w30944 and not w30949;
w30951 <= pi0215 and not w30950;
w30952 <= w1011 and not w30942;
w30953 <= pi0198 and not w14247;
w30954 <= not w3759 and not w30953;
w30955 <= not w30943 and not w30954;
w30956 <= w3805 and w30955;
w30957 <= pi0198 and not w14706;
w30958 <= not w3805 and w30957;
w30959 <= not w1011 and not w30956;
w30960 <= not w30958 and w30959;
w30961 <= not pi0215 and not w30952;
w30962 <= not w30960 and w30961;
w30963 <= pi0299 and not w30951;
w30964 <= not w30962 and w30963;
w30965 <= not w3768 and w30948;
w30966 <= not w30944 and not w30965;
w30967 <= pi0223 and not w30966;
w30968 <= w166 and not w30942;
w30969 <= not w3768 and w30957;
w30970 <= w3768 and w30955;
w30971 <= not w166 and not w30970;
w30972 <= not w30969 and w30971;
w30973 <= not pi0223 and not w30968;
w30974 <= not w30972 and w30973;
w30975 <= not pi0299 and not w30967;
w30976 <= not w30974 and w30975;
w30977 <= w134 and w8545;
w30978 <= not w30964 and w30977;
w30979 <= not w30976 and w30978;
w30980 <= not w30940 and not w30979;
w30981 <= not w16712 and w30980;
w30982 <= w14202 and not w30980;
w30983 <= pi0198 and not w134;
w30984 <= pi0039 and pi0198;
w30985 <= pi0038 and not w30984;
w30986 <= pi0198 and not w14230;
w30987 <= pi0634 and w14207;
w30988 <= w14230 and w30987;
w30989 <= not w30986 and not w30988;
w30990 <= not pi0039 and not w30989;
w30991 <= w30985 and not w30990;
w30992 <= pi0198 and w14284;
w30993 <= pi0634 and not w14284;
w30994 <= w14221 and w30993;
w30995 <= not w30992 and not w30994;
w30996 <= w3758 and not w30995;
w30997 <= not pi0680 and w30948;
w30998 <= w3755 and w30995;
w30999 <= not w14221 and not w30942;
w31000 <= pi0634 and not w30999;
w31001 <= not w30942 and not w31000;
w31002 <= not w3760 and w31001;
w31003 <= w3760 and w30995;
w31004 <= not w31002 and not w31003;
w31005 <= not w3755 and not w31004;
w31006 <= w14886 and not w30998;
w31007 <= not w31005 and w31006;
w31008 <= not w30996 and not w30997;
w31009 <= not w31007 and w31008;
w31010 <= not w3768 and w31009;
w31011 <= w30941 and w30997;
w31012 <= w3760 and not w31001;
w31013 <= not w3760 and not w30995;
w31014 <= not w31012 and not w31013;
w31015 <= w3755 and w31014;
w31016 <= not w3755 and w31001;
w31017 <= w14886 and not w31016;
w31018 <= not w31015 and w31017;
w31019 <= w3758 and not w31014;
w31020 <= not w31011 and not w31019;
w31021 <= not w31018 and w31020;
w31022 <= w3768 and w31021;
w31023 <= pi0223 and not w31010;
w31024 <= not w31022 and w31023;
w31025 <= pi0680 and w31000;
w31026 <= not w30942 and not w31025;
w31027 <= w166 and w31026;
w31028 <= pi0198 and w14244;
w31029 <= pi0634 and w14249;
w31030 <= not w31028 and not w31029;
w31031 <= not w3760 and not w31030;
w31032 <= not w31012 and not w31031;
w31033 <= w3758 and not w31032;
w31034 <= w3755 and w31032;
w31035 <= w31017 and not w31034;
w31036 <= not w3755 and not w30942;
w31037 <= w3755 and not w30953;
w31038 <= not pi0680 and not w31036;
w31039 <= not w31037 and w31038;
w31040 <= not w31033 and not w31039;
w31041 <= not w31035 and w31040;
w31042 <= w3768 and not w31041;
w31043 <= pi0198 and w14316;
w31044 <= w3758 and not w31030;
w31045 <= w3755 and w31030;
w31046 <= w3760 and w31030;
w31047 <= not w31002 and not w31046;
w31048 <= not w3755 and not w31047;
w31049 <= w14886 and not w31045;
w31050 <= not w31048 and w31049;
w31051 <= not w31043 and not w31044;
w31052 <= not w31050 and w31051;
w31053 <= not w3768 and not w31052;
w31054 <= not w166 and not w31042;
w31055 <= not w31053 and w31054;
w31056 <= not pi0223 and not w31027;
w31057 <= not w31055 and w31056;
w31058 <= not pi0299 and not w31024;
w31059 <= not w31057 and w31058;
w31060 <= not w3805 and w31009;
w31061 <= w3805 and w31021;
w31062 <= pi0215 and not w31060;
w31063 <= not w31061 and w31062;
w31064 <= w1011 and w31026;
w31065 <= not w3805 and not w31052;
w31066 <= w3805 and not w31041;
w31067 <= not w1011 and not w31065;
w31068 <= not w31066 and w31067;
w31069 <= not pi0215 and not w31064;
w31070 <= not w31068 and w31069;
w31071 <= pi0299 and not w31063;
w31072 <= not w31070 and w31071;
w31073 <= not w31059 and not w31072;
w31074 <= pi0039 and not w31073;
w31075 <= pi0634 and pi0680;
w31076 <= pi0198 and w14494;
w31077 <= not w14459 and w31075;
w31078 <= not w31076 and w31077;
w31079 <= not w14492 and not w31078;
w31080 <= not pi0299 and not w31079;
w31081 <= not pi0198 and w14486;
w31082 <= pi0198 and not w14507;
w31083 <= not w31081 and not w31082;
w31084 <= w31075 and not w31083;
w31085 <= pi0198 and not w14504;
w31086 <= not w31075 and w31085;
w31087 <= not w31084 and not w31086;
w31088 <= pi0299 and not w31087;
w31089 <= not pi0039 and not w31080;
w31090 <= not w31088 and w31089;
w31091 <= not w31074 and not w31090;
w31092 <= not pi0038 and not w31091;
w31093 <= w134 and not w30991;
w31094 <= not w31092 and w31093;
w31095 <= not w30983 and not w31094;
w31096 <= not pi0778 and not w31095;
w31097 <= not pi0625 and w30980;
w31098 <= pi0625 and w31095;
w31099 <= pi1153 and not w31097;
w31100 <= not w31098 and w31099;
w31101 <= not pi0625 and w31095;
w31102 <= pi0625 and w30980;
w31103 <= not pi1153 and not w31102;
w31104 <= not w31101 and w31103;
w31105 <= not w31100 and not w31104;
w31106 <= pi0778 and not w31105;
w31107 <= not w31096 and not w31106;
w31108 <= not w14638 and w31107;
w31109 <= w14638 and w30980;
w31110 <= not w31108 and not w31109;
w31111 <= not w14202 and w31110;
w31112 <= not w30982 and not w31111;
w31113 <= not w14198 and w31112;
w31114 <= not w14194 and w31113;
w31115 <= not w30981 and not w31114;
w31116 <= not pi0792 and w31115;
w31117 <= pi0628 and not w31115;
w31118 <= not pi0628 and w30980;
w31119 <= not w31117 and not w31118;
w31120 <= pi1156 and w31119;
w31121 <= pi0628 and w30980;
w31122 <= not pi0628 and not w31115;
w31123 <= not pi1156 and not w31121;
w31124 <= not w31122 and w31123;
w31125 <= not w31120 and not w31124;
w31126 <= pi0792 and not w31125;
w31127 <= not w31116 and not w31126;
w31128 <= not pi0647 and w31127;
w31129 <= pi0647 and w30980;
w31130 <= not pi1157 and not w31129;
w31131 <= not w31128 and w31130;
w31132 <= pi0630 and w31131;
w31133 <= w15342 and not w30980;
w31134 <= not w14690 and not w14694;
w31135 <= pi0633 and not w31134;
w31136 <= not w14492 and not w31135;
w31137 <= not w14699 and not w31136;
w31138 <= not pi0299 and w31137;
w31139 <= pi0603 and pi0633;
w31140 <= not w31085 and not w31139;
w31141 <= pi0198 and not w14685;
w31142 <= not pi0198 and w14793;
w31143 <= not w31141 and not w31142;
w31144 <= w31139 and w31143;
w31145 <= not w31140 and not w31144;
w31146 <= pi0299 and w31145;
w31147 <= not pi0039 and not w31138;
w31148 <= not w31146 and w31147;
w31149 <= pi0633 and w14802;
w31150 <= not w30948 and not w31149;
w31151 <= not w3758 and not w31150;
w31152 <= pi0633 and w14216;
w31153 <= not w14707 and w31152;
w31154 <= not w14284 and w31153;
w31155 <= not w30992 and not w31154;
w31156 <= w14751 and not w31155;
w31157 <= not w31151 and not w31156;
w31158 <= not w3768 and w31157;
w31159 <= not w30942 and not w31153;
w31160 <= pi0603 and not w31159;
w31161 <= not pi0603 and w30942;
w31162 <= not w31160 and not w31161;
w31163 <= not w14730 and w31162;
w31164 <= w3760 and not w31159;
w31165 <= not w30941 and not w31154;
w31166 <= not w31164 and w31165;
w31167 <= pi0603 and not w31166;
w31168 <= w14730 and not w31161;
w31169 <= not w31167 and w31168;
w31170 <= not w31163 and not w31169;
w31171 <= not w3758 and w31170;
w31172 <= not w30941 and not w31167;
w31173 <= w3758 and not w31172;
w31174 <= not w31171 and not w31173;
w31175 <= w3768 and w31174;
w31176 <= pi0223 and not w31158;
w31177 <= not w31175 and w31176;
w31178 <= w166 and w31162;
w31179 <= pi0642 and not w31160;
w31180 <= pi0633 and w14710;
w31181 <= not w31028 and not w31180;
w31182 <= not w3760 and not w31181;
w31183 <= not w31164 and not w31182;
w31184 <= pi0603 and not w31183;
w31185 <= not pi0642 and not w31184;
w31186 <= w3754 and not w31179;
w31187 <= not w31185 and w31186;
w31188 <= not w3754 and w31160;
w31189 <= not w31161 and not w31188;
w31190 <= not w31187 and w31189;
w31191 <= not w3758 and w31190;
w31192 <= not pi0603 and w30953;
w31193 <= w3758 and not w31192;
w31194 <= not w31184 and w31193;
w31195 <= not w31191 and not w31194;
w31196 <= w3768 and w31195;
w31197 <= pi0603 and not w31181;
w31198 <= w14730 and w31197;
w31199 <= pi0198 and w14712;
w31200 <= w3760 and w31181;
w31201 <= not w3760 and w31159;
w31202 <= pi0603 and not w14730;
w31203 <= not w31201 and w31202;
w31204 <= not w31200 and w31203;
w31205 <= not w31198 and not w31199;
w31206 <= not w31204 and w31205;
w31207 <= not w3758 and w31206;
w31208 <= w3758 and not w31028;
w31209 <= not w31197 and w31208;
w31210 <= not w31207 and not w31209;
w31211 <= not w3768 and w31210;
w31212 <= not w166 and not w31211;
w31213 <= not w31196 and w31212;
w31214 <= not pi0223 and not w31178;
w31215 <= not w31213 and w31214;
w31216 <= not w31177 and not w31215;
w31217 <= not pi0299 and not w31216;
w31218 <= not w3805 and w31157;
w31219 <= w3805 and w31174;
w31220 <= pi0215 and not w31218;
w31221 <= not w31219 and w31220;
w31222 <= w1011 and w31162;
w31223 <= not w3805 and w31210;
w31224 <= w3805 and w31195;
w31225 <= not w1011 and not w31223;
w31226 <= not w31224 and w31225;
w31227 <= not pi0215 and not w31222;
w31228 <= not w31226 and w31227;
w31229 <= not w31221 and not w31228;
w31230 <= pi0299 and not w31229;
w31231 <= pi0039 and not w31217;
w31232 <= not w31230 and w31231;
w31233 <= not w31148 and not w31232;
w31234 <= not pi0038 and not w31233;
w31235 <= pi0633 and w14731;
w31236 <= w14230 and w31235;
w31237 <= not w30986 and not w31236;
w31238 <= not pi0039 and not w31237;
w31239 <= w30985 and not w31238;
w31240 <= w134 and not w31239;
w31241 <= not w31234 and w31240;
w31242 <= not w30983 and not w31241;
w31243 <= not w14680 and not w31242;
w31244 <= w14680 and not w30980;
w31245 <= not w31243 and not w31244;
w31246 <= not pi0785 and not w31245;
w31247 <= not w14854 and not w30980;
w31248 <= pi0609 and w31243;
w31249 <= not w31247 and not w31248;
w31250 <= pi1155 and not w31249;
w31251 <= not w14859 and not w30980;
w31252 <= not pi0609 and w31243;
w31253 <= not w31251 and not w31252;
w31254 <= not pi1155 and not w31253;
w31255 <= not w31250 and not w31254;
w31256 <= pi0785 and not w31255;
w31257 <= not w31246 and not w31256;
w31258 <= not pi0781 and not w31257;
w31259 <= not pi0618 and w30980;
w31260 <= pi0618 and w31257;
w31261 <= pi1154 and not w31259;
w31262 <= not w31260 and w31261;
w31263 <= not pi0618 and w31257;
w31264 <= pi0618 and w30980;
w31265 <= not pi1154 and not w31264;
w31266 <= not w31263 and w31265;
w31267 <= not w31262 and not w31266;
w31268 <= pi0781 and not w31267;
w31269 <= not w31258 and not w31268;
w31270 <= not pi0789 and not w31269;
w31271 <= not pi0619 and w30980;
w31272 <= pi0619 and w31269;
w31273 <= pi1159 and not w31271;
w31274 <= not w31272 and w31273;
w31275 <= not pi0619 and w31269;
w31276 <= pi0619 and w30980;
w31277 <= not pi1159 and not w31276;
w31278 <= not w31275 and w31277;
w31279 <= not w31274 and not w31278;
w31280 <= pi0789 and not w31279;
w31281 <= not w31270 and not w31280;
w31282 <= not w15532 and w31281;
w31283 <= w15532 and w30980;
w31284 <= not w31282 and not w31283;
w31285 <= not w15342 and w31284;
w31286 <= not w31133 and not w31285;
w31287 <= not w18122 and not w31286;
w31288 <= pi0647 and not w31127;
w31289 <= not pi0647 and not w30980;
w31290 <= not w31288 and not w31289;
w31291 <= w15364 and not w31290;
w31292 <= not w31132 and not w31291;
w31293 <= not w31287 and w31292;
w31294 <= pi0787 and not w31293;
w31295 <= pi0629 and w31124;
w31296 <= not w18133 and w31284;
w31297 <= w15339 and w31119;
w31298 <= not w31295 and not w31297;
w31299 <= not w31296 and w31298;
w31300 <= pi0792 and not w31299;
w31301 <= w14198 and w30980;
w31302 <= not w31113 and not w31301;
w31303 <= w15434 and not w31302;
w31304 <= not pi0626 and not w31281;
w31305 <= pi0626 and not w30980;
w31306 <= w14192 and not w31305;
w31307 <= not w31304 and w31306;
w31308 <= pi0626 and not w31281;
w31309 <= not pi0626 and not w30980;
w31310 <= w14191 and not w31309;
w31311 <= not w31308 and w31310;
w31312 <= not w31303 and not w31307;
w31313 <= not w31311 and w31312;
w31314 <= pi0788 and not w31313;
w31315 <= pi0609 and w31107;
w31316 <= pi0634 and w15208;
w31317 <= w31237 and not w31316;
w31318 <= not pi0039 and not w31317;
w31319 <= w30985 and not w31318;
w31320 <= not w31075 and w31145;
w31321 <= not pi0603 and not w31083;
w31322 <= not pi0198 and not pi0665;
w31323 <= w14685 and w31322;
w31324 <= not w14793 and w31082;
w31325 <= not pi0633 and not w31323;
w31326 <= not w31324 and w31325;
w31327 <= pi0198 and not pi0665;
w31328 <= pi0633 and not w31327;
w31329 <= not w31081 and w31328;
w31330 <= w31143 and w31329;
w31331 <= pi0603 and not w31326;
w31332 <= not w31330 and w31331;
w31333 <= not w31321 and not w31332;
w31334 <= w31075 and not w31333;
w31335 <= pi0299 and not w31320;
w31336 <= not w31334 and w31335;
w31337 <= not pi0680 and w31137;
w31338 <= not pi0603 and w31079;
w31339 <= pi0198 and not pi0633;
w31340 <= pi0634 and not pi0665;
w31341 <= not w31339 and w31340;
w31342 <= not w14689 and w31341;
w31343 <= not pi0634 and w14492;
w31344 <= pi0634 and w14495;
w31345 <= not w14696 and w31344;
w31346 <= not w31343 and not w31345;
w31347 <= not pi0633 and not w31346;
w31348 <= pi0603 and not w31342;
w31349 <= not w31135 and w31348;
w31350 <= not w31347 and w31349;
w31351 <= pi0680 and not w31338;
w31352 <= not w31350 and w31351;
w31353 <= not pi0299 and not w31337;
w31354 <= not w31352 and w31353;
w31355 <= not w31336 and not w31354;
w31356 <= not pi0039 and not w31355;
w31357 <= w14918 and w31000;
w31358 <= w31162 and not w31357;
w31359 <= w166 and w31358;
w31360 <= not pi0680 and w31190;
w31361 <= not pi0603 and not w31001;
w31362 <= w14722 and w31340;
w31363 <= w31159 and not w31362;
w31364 <= pi0603 and not w31363;
w31365 <= not w31361 and not w31364;
w31366 <= not w3754 and not w31365;
w31367 <= w3760 and not w31363;
w31368 <= pi0634 and w14987;
w31369 <= w31181 and not w31368;
w31370 <= not w3760 and not w31369;
w31371 <= not w31367 and not w31370;
w31372 <= pi0603 and not w31371;
w31373 <= not pi0642 and w31372;
w31374 <= pi0642 and w31364;
w31375 <= not w31361 and not w31374;
w31376 <= not w31373 and w31375;
w31377 <= w3754 and not w31376;
w31378 <= not w14220 and not w31366;
w31379 <= not w31377 and w31378;
w31380 <= not pi0603 and not w31032;
w31381 <= w14220 and not w31380;
w31382 <= not w31372 and w31381;
w31383 <= not w31379 and not w31382;
w31384 <= pi0680 and not w31383;
w31385 <= not w31360 and not w31384;
w31386 <= w3768 and w31385;
w31387 <= not pi0680 and not w31206;
w31388 <= not pi0603 and w31047;
w31389 <= not w14730 and w31364;
w31390 <= not w31203 and not w31389;
w31391 <= not w3755 and w31390;
w31392 <= not w3760 and not w31390;
w31393 <= w31369 and not w31392;
w31394 <= not w31391 and not w31393;
w31395 <= not w31388 and not w31394;
w31396 <= w14886 and not w31395;
w31397 <= not w14731 and not w31030;
w31398 <= not w31197 and not w31397;
w31399 <= w3758 and not w31398;
w31400 <= not w31387 and not w31399;
w31401 <= not w31396 and w31400;
w31402 <= not w3768 and not w31401;
w31403 <= not w166 and not w31402;
w31404 <= not w31386 and w31403;
w31405 <= not pi0223 and not w31359;
w31406 <= not w31404 and w31405;
w31407 <= not pi0680 and not w31150;
w31408 <= w14754 and w31322;
w31409 <= w14707 and w31327;
w31410 <= not w30992 and not w31409;
w31411 <= not w31408 and w31410;
w31412 <= pi0634 and not w31411;
w31413 <= not pi0634 and w30992;
w31414 <= not w31154 and not w31413;
w31415 <= not w31412 and w31414;
w31416 <= pi0603 and not w31415;
w31417 <= not pi0603 and not w30995;
w31418 <= not w31416 and not w31417;
w31419 <= w3758 and not w31418;
w31420 <= w14730 and w31416;
w31421 <= not pi0603 and w31004;
w31422 <= not w31390 and not w31415;
w31423 <= not w31392 and not w31421;
w31424 <= not w31420 and not w31422;
w31425 <= w31423 and w31424;
w31426 <= w14886 and not w31425;
w31427 <= not w31407 and not w31419;
w31428 <= not w31426 and w31427;
w31429 <= not w3768 and w31428;
w31430 <= not pi0680 and w31170;
w31431 <= not w3760 and not w31415;
w31432 <= not w31367 and not w31431;
w31433 <= pi0603 and not w31432;
w31434 <= not pi0603 and not w31014;
w31435 <= not w31433 and not w31434;
w31436 <= w3758 and not w31435;
w31437 <= not w14730 and w31365;
w31438 <= w14730 and not w31361;
w31439 <= not w31433 and w31438;
w31440 <= w14886 and not w31437;
w31441 <= not w31439 and w31440;
w31442 <= not w31430 and not w31436;
w31443 <= not w31441 and w31442;
w31444 <= w3768 and w31443;
w31445 <= pi0223 and not w31429;
w31446 <= not w31444 and w31445;
w31447 <= not w31406 and not w31446;
w31448 <= not pi0299 and not w31447;
w31449 <= w1011 and w31358;
w31450 <= w3805 and w31385;
w31451 <= not w3805 and not w31401;
w31452 <= not w1011 and not w31451;
w31453 <= not w31450 and w31452;
w31454 <= not pi0215 and not w31449;
w31455 <= not w31453 and w31454;
w31456 <= not w3805 and w31428;
w31457 <= w3805 and w31443;
w31458 <= pi0215 and not w31456;
w31459 <= not w31457 and w31458;
w31460 <= not w31455 and not w31459;
w31461 <= pi0299 and not w31460;
w31462 <= pi0039 and not w31448;
w31463 <= not w31461 and w31462;
w31464 <= not w31356 and not w31463;
w31465 <= not pi0038 and not w31464;
w31466 <= w134 and not w31319;
w31467 <= not w31465 and w31466;
w31468 <= not w30983 and not w31467;
w31469 <= not pi0625 and w31468;
w31470 <= pi0625 and w31242;
w31471 <= not pi1153 and not w31470;
w31472 <= not w31469 and w31471;
w31473 <= not pi0608 and not w31100;
w31474 <= not w31472 and w31473;
w31475 <= not pi0625 and w31242;
w31476 <= pi0625 and w31468;
w31477 <= pi1153 and not w31475;
w31478 <= not w31476 and w31477;
w31479 <= pi0608 and not w31104;
w31480 <= not w31478 and w31479;
w31481 <= not w31474 and not w31480;
w31482 <= pi0778 and not w31481;
w31483 <= not pi0778 and w31468;
w31484 <= not w31482 and not w31483;
w31485 <= not pi0609 and not w31484;
w31486 <= not pi1155 and not w31315;
w31487 <= not w31485 and w31486;
w31488 <= not pi0660 and not w31250;
w31489 <= not w31487 and w31488;
w31490 <= not pi0609 and w31107;
w31491 <= pi0609 and not w31484;
w31492 <= pi1155 and not w31490;
w31493 <= not w31491 and w31492;
w31494 <= pi0660 and not w31254;
w31495 <= not w31493 and w31494;
w31496 <= not w31489 and not w31495;
w31497 <= pi0785 and not w31496;
w31498 <= not pi0785 and not w31484;
w31499 <= not w31497 and not w31498;
w31500 <= not pi0618 and not w31499;
w31501 <= pi0618 and not w31110;
w31502 <= not pi1154 and not w31501;
w31503 <= not w31500 and w31502;
w31504 <= not pi0627 and not w31262;
w31505 <= not w31503 and w31504;
w31506 <= pi0618 and not w31499;
w31507 <= not pi0618 and not w31110;
w31508 <= pi1154 and not w31507;
w31509 <= not w31506 and w31508;
w31510 <= pi0627 and not w31266;
w31511 <= not w31509 and w31510;
w31512 <= not w31505 and not w31511;
w31513 <= pi0781 and not w31512;
w31514 <= not pi0781 and not w31499;
w31515 <= not w31513 and not w31514;
w31516 <= not pi0789 and w31515;
w31517 <= not pi0619 and not w31515;
w31518 <= pi0619 and w31112;
w31519 <= not pi1159 and not w31518;
w31520 <= not w31517 and w31519;
w31521 <= not pi0648 and not w31274;
w31522 <= not w31520 and w31521;
w31523 <= not pi0619 and w31112;
w31524 <= pi0619 and not w31515;
w31525 <= pi1159 and not w31523;
w31526 <= not w31524 and w31525;
w31527 <= pi0648 and not w31278;
w31528 <= not w31526 and w31527;
w31529 <= pi0789 and not w31522;
w31530 <= not w31528 and w31529;
w31531 <= w15533 and not w31516;
w31532 <= not w31530 and w31531;
w31533 <= not w31314 and not w31532;
w31534 <= not w31300 and not w31533;
w31535 <= w17927 and w31299;
w31536 <= not w17769 and not w31535;
w31537 <= not w31534 and w31536;
w31538 <= not w31294 and not w31537;
w31539 <= not pi0790 and not w31538;
w31540 <= not pi0787 and not w31127;
w31541 <= pi1157 and not w31290;
w31542 <= not w31131 and not w31541;
w31543 <= pi0787 and not w31542;
w31544 <= not w31540 and not w31543;
w31545 <= not pi0644 and w31544;
w31546 <= pi0644 and w31538;
w31547 <= pi0715 and not w31545;
w31548 <= not w31546 and w31547;
w31549 <= not w15367 and w31286;
w31550 <= w15367 and w30980;
w31551 <= not w31549 and not w31550;
w31552 <= pi0644 and not w31551;
w31553 <= not pi0644 and w30980;
w31554 <= not pi0715 and not w31553;
w31555 <= not w31552 and w31554;
w31556 <= pi1160 and not w31555;
w31557 <= not w31548 and w31556;
w31558 <= not pi0644 and not w31551;
w31559 <= pi0644 and w30980;
w31560 <= pi0715 and not w31559;
w31561 <= not w31558 and w31560;
w31562 <= pi0644 and w31544;
w31563 <= not pi0644 and w31538;
w31564 <= not pi0715 and not w31562;
w31565 <= not w31563 and w31564;
w31566 <= not pi1160 and not w31561;
w31567 <= not w31565 and w31566;
w31568 <= pi0790 and not w31557;
w31569 <= not w31567 and w31568;
w31570 <= not w31539 and not w31569;
w31571 <= w4989 and not w31570;
w31572 <= pi0198 and not w4989;
w31573 <= not w31571 and not w31572;
w31574 <= pi0199 and not w14622;
w31575 <= not pi0619 and not w31574;
w31576 <= not pi0617 and not w31574;
w31577 <= not pi0199 and not w16995;
w31578 <= w17001 and not w31577;
w31579 <= not pi0199 and not w14838;
w31580 <= pi0199 and w14784;
w31581 <= not pi0038 and not w31579;
w31582 <= not w31580 and w31581;
w31583 <= not w31578 and not w31582;
w31584 <= w134 and not w31583;
w31585 <= pi0199 and not w134;
w31586 <= pi0617 and not w31585;
w31587 <= not w31584 and w31586;
w31588 <= not w31576 and not w31587;
w31589 <= not w14680 and not w31588;
w31590 <= w14680 and not w31574;
w31591 <= not w31589 and not w31590;
w31592 <= not pi0785 and w31591;
w31593 <= not pi0609 and not w31574;
w31594 <= pi0609 and not w31591;
w31595 <= pi1155 and not w31593;
w31596 <= not w31594 and w31595;
w31597 <= not pi0609 and not w31591;
w31598 <= pi0609 and not w31574;
w31599 <= not pi1155 and not w31598;
w31600 <= not w31597 and w31599;
w31601 <= not w31596 and not w31600;
w31602 <= pi0785 and not w31601;
w31603 <= not w31592 and not w31602;
w31604 <= not pi0781 and not w31603;
w31605 <= not pi0618 and not w31574;
w31606 <= pi0618 and w31603;
w31607 <= pi1154 and not w31605;
w31608 <= not w31606 and w31607;
w31609 <= pi0618 and not w31574;
w31610 <= not pi0618 and w31603;
w31611 <= not pi1154 and not w31609;
w31612 <= not w31610 and w31611;
w31613 <= not w31608 and not w31612;
w31614 <= pi0781 and not w31613;
w31615 <= not w31604 and not w31614;
w31616 <= pi0619 and w31615;
w31617 <= pi1159 and not w31575;
w31618 <= not w31616 and w31617;
w31619 <= not pi0625 and not w31574;
w31620 <= not pi0637 and not w31574;
w31621 <= not pi0199 and not w14204;
w31622 <= w17462 and not w31621;
w31623 <= pi0199 and not w14403;
w31624 <= not pi0199 and not w14312;
w31625 <= pi0039 and not w31624;
w31626 <= not w31623 and w31625;
w31627 <= pi0199 and not w14511;
w31628 <= not pi0199 and w14489;
w31629 <= not pi0039 and not w31627;
w31630 <= not w31628 and w31629;
w31631 <= not pi0038 and not w31630;
w31632 <= not w31626 and w31631;
w31633 <= not w31622 and not w31632;
w31634 <= w134 and not w31633;
w31635 <= pi0637 and not w31585;
w31636 <= not w31634 and w31635;
w31637 <= not w31620 and not w31636;
w31638 <= pi0625 and not w31637;
w31639 <= pi1153 and not w31619;
w31640 <= not w31638 and w31639;
w31641 <= not pi0637 and w31588;
w31642 <= pi0199 and w17039;
w31643 <= w134 and not w22112;
w31644 <= not pi0199 and not w31643;
w31645 <= not pi0617 and not w17035;
w31646 <= not w31644 and w31645;
w31647 <= not w31642 and w31646;
w31648 <= w134 and w17059;
w31649 <= not pi0199 and not w31648;
w31650 <= pi0199 and w17051;
w31651 <= pi0617 and not w31650;
w31652 <= not w31649 and w31651;
w31653 <= not w31585 and not w31652;
w31654 <= not w31647 and w31653;
w31655 <= pi0637 and not w31654;
w31656 <= not w31641 and not w31655;
w31657 <= not pi0625 and w31656;
w31658 <= pi0625 and not w31588;
w31659 <= not pi1153 and not w31658;
w31660 <= not w31657 and w31659;
w31661 <= not pi0608 and not w31640;
w31662 <= not w31660 and w31661;
w31663 <= not pi0625 and not w31637;
w31664 <= pi0625 and not w31574;
w31665 <= not pi1153 and not w31664;
w31666 <= not w31663 and w31665;
w31667 <= pi0625 and w31656;
w31668 <= not pi0625 and not w31588;
w31669 <= pi1153 and not w31668;
w31670 <= not w31667 and w31669;
w31671 <= pi0608 and not w31666;
w31672 <= not w31670 and w31671;
w31673 <= not w31662 and not w31672;
w31674 <= pi0778 and not w31673;
w31675 <= not pi0778 and w31656;
w31676 <= not w31674 and not w31675;
w31677 <= not pi0609 and not w31676;
w31678 <= not pi0778 and w31637;
w31679 <= not w31640 and not w31666;
w31680 <= pi0778 and not w31679;
w31681 <= not w31678 and not w31680;
w31682 <= pi0609 and w31681;
w31683 <= not pi1155 and not w31682;
w31684 <= not w31677 and w31683;
w31685 <= not pi0660 and not w31596;
w31686 <= not w31684 and w31685;
w31687 <= not pi0609 and w31681;
w31688 <= pi0609 and not w31676;
w31689 <= pi1155 and not w31687;
w31690 <= not w31688 and w31689;
w31691 <= pi0660 and not w31600;
w31692 <= not w31690 and w31691;
w31693 <= not w31686 and not w31692;
w31694 <= pi0785 and not w31693;
w31695 <= not pi0785 and not w31676;
w31696 <= not w31694 and not w31695;
w31697 <= not pi0618 and not w31696;
w31698 <= w14638 and not w31574;
w31699 <= not w14638 and w31681;
w31700 <= not w31698 and not w31699;
w31701 <= pi0618 and not w31700;
w31702 <= not pi1154 and not w31701;
w31703 <= not w31697 and w31702;
w31704 <= not pi0627 and not w31608;
w31705 <= not w31703 and w31704;
w31706 <= pi0618 and not w31696;
w31707 <= not pi0618 and not w31700;
w31708 <= pi1154 and not w31707;
w31709 <= not w31706 and w31708;
w31710 <= pi0627 and not w31612;
w31711 <= not w31709 and w31710;
w31712 <= not w31705 and not w31711;
w31713 <= pi0781 and not w31712;
w31714 <= not pi0781 and not w31696;
w31715 <= not w31713 and not w31714;
w31716 <= not pi0619 and not w31715;
w31717 <= not w14202 and w31700;
w31718 <= w14202 and w31574;
w31719 <= not w31717 and not w31718;
w31720 <= pi0619 and w31719;
w31721 <= not pi1159 and not w31720;
w31722 <= not w31716 and w31721;
w31723 <= not pi0648 and not w31618;
w31724 <= not w31722 and w31723;
w31725 <= pi0619 and not w31574;
w31726 <= not pi0619 and w31615;
w31727 <= not pi1159 and not w31725;
w31728 <= not w31726 and w31727;
w31729 <= not pi0619 and w31719;
w31730 <= pi0619 and not w31715;
w31731 <= pi1159 and not w31729;
w31732 <= not w31730 and w31731;
w31733 <= pi0648 and not w31728;
w31734 <= not w31732 and w31733;
w31735 <= not w31724 and not w31734;
w31736 <= pi0789 and not w31735;
w31737 <= not pi0789 and not w31715;
w31738 <= not w31736 and not w31737;
w31739 <= not pi0788 and w31738;
w31740 <= not pi0626 and w31738;
w31741 <= w14198 and not w31574;
w31742 <= not w14198 and w31719;
w31743 <= not w31741 and not w31742;
w31744 <= pi0626 and w31743;
w31745 <= not pi0641 and not w31744;
w31746 <= not w31740 and w31745;
w31747 <= not pi0789 and not w31615;
w31748 <= not w31618 and not w31728;
w31749 <= pi0789 and not w31748;
w31750 <= not w31747 and not w31749;
w31751 <= not pi0626 and not w31750;
w31752 <= pi0626 and w31574;
w31753 <= pi0641 and not w31752;
w31754 <= not w31751 and w31753;
w31755 <= not pi1158 and not w31754;
w31756 <= not w31746 and w31755;
w31757 <= not pi0626 and w31743;
w31758 <= pi0626 and w31738;
w31759 <= pi0641 and not w31757;
w31760 <= not w31758 and w31759;
w31761 <= pi0626 and not w31750;
w31762 <= not pi0626 and w31574;
w31763 <= not pi0641 and not w31762;
w31764 <= not w31761 and w31763;
w31765 <= pi1158 and not w31764;
w31766 <= not w31760 and w31765;
w31767 <= not w31756 and not w31766;
w31768 <= pi0788 and not w31767;
w31769 <= not w31739 and not w31768;
w31770 <= not pi0628 and w31769;
w31771 <= not w15532 and not w31750;
w31772 <= w15532 and w31574;
w31773 <= not w31771 and not w31772;
w31774 <= pi0628 and w31773;
w31775 <= not pi1156 and not w31774;
w31776 <= not w31770 and w31775;
w31777 <= not pi0628 and not w31574;
w31778 <= not w14194 and w31743;
w31779 <= w14194 and w31574;
w31780 <= not w31778 and not w31779;
w31781 <= pi0628 and w31780;
w31782 <= pi1156 and not w31777;
w31783 <= not w31781 and w31782;
w31784 <= not pi0629 and not w31783;
w31785 <= not w31776 and w31784;
w31786 <= pi0628 and w31769;
w31787 <= not pi0628 and w31773;
w31788 <= pi1156 and not w31787;
w31789 <= not w31786 and w31788;
w31790 <= pi0628 and not w31574;
w31791 <= not pi0628 and w31780;
w31792 <= not pi1156 and not w31790;
w31793 <= not w31791 and w31792;
w31794 <= pi0629 and not w31793;
w31795 <= not w31789 and w31794;
w31796 <= not w31785 and not w31795;
w31797 <= pi0792 and not w31796;
w31798 <= not pi0792 and w31769;
w31799 <= not w31797 and not w31798;
w31800 <= not pi0647 and not w31799;
w31801 <= not w15342 and not w31773;
w31802 <= w15342 and w31574;
w31803 <= not w31801 and not w31802;
w31804 <= pi0647 and w31803;
w31805 <= not pi1157 and not w31804;
w31806 <= not w31800 and w31805;
w31807 <= not pi0647 and not w31574;
w31808 <= not pi0792 and not w31780;
w31809 <= not w31783 and not w31793;
w31810 <= pi0792 and not w31809;
w31811 <= not w31808 and not w31810;
w31812 <= pi0647 and w31811;
w31813 <= pi1157 and not w31807;
w31814 <= not w31812 and w31813;
w31815 <= not pi0630 and not w31814;
w31816 <= not w31806 and w31815;
w31817 <= pi0647 and not w31799;
w31818 <= not pi0647 and w31803;
w31819 <= pi1157 and not w31818;
w31820 <= not w31817 and w31819;
w31821 <= pi0647 and not w31574;
w31822 <= not pi0647 and w31811;
w31823 <= not pi1157 and not w31821;
w31824 <= not w31822 and w31823;
w31825 <= pi0630 and not w31824;
w31826 <= not w31820 and w31825;
w31827 <= not w31816 and not w31826;
w31828 <= pi0787 and not w31827;
w31829 <= not pi0787 and not w31799;
w31830 <= not w31828 and not w31829;
w31831 <= not pi0790 and w31830;
w31832 <= not pi0787 and not w31811;
w31833 <= not w31814 and not w31824;
w31834 <= pi0787 and not w31833;
w31835 <= not w31832 and not w31834;
w31836 <= not pi0644 and w31835;
w31837 <= pi0644 and not w31830;
w31838 <= pi0715 and not w31836;
w31839 <= not w31837 and w31838;
w31840 <= w15367 and not w31574;
w31841 <= not w15367 and w31803;
w31842 <= not w31840 and not w31841;
w31843 <= pi0644 and not w31842;
w31844 <= not pi0644 and not w31574;
w31845 <= not pi0715 and not w31844;
w31846 <= not w31843 and w31845;
w31847 <= pi1160 and not w31846;
w31848 <= not w31839 and w31847;
w31849 <= not pi0644 and not w31830;
w31850 <= pi0644 and w31835;
w31851 <= not pi0715 and not w31850;
w31852 <= not w31849 and w31851;
w31853 <= not pi0644 and not w31842;
w31854 <= pi0644 and not w31574;
w31855 <= pi0715 and not w31854;
w31856 <= not w31853 and w31855;
w31857 <= not pi1160 and not w31856;
w31858 <= not w31852 and w31857;
w31859 <= pi0790 and not w31848;
w31860 <= not w31858 and w31859;
w31861 <= not w31831 and not w31860;
w31862 <= w4989 and not w31861;
w31863 <= pi0199 and not w4989;
w31864 <= not w31862 and not w31863;
w31865 <= pi0200 and not w14622;
w31866 <= not pi0606 and not w31865;
w31867 <= pi0200 and not w134;
w31868 <= not pi0200 and not w16995;
w31869 <= w17001 and not w31868;
w31870 <= not pi0200 and not w14838;
w31871 <= pi0200 and w14784;
w31872 <= not pi0038 and not w31870;
w31873 <= not w31871 and w31872;
w31874 <= not w31869 and not w31873;
w31875 <= w134 and not w31874;
w31876 <= pi0606 and not w31867;
w31877 <= not w31875 and w31876;
w31878 <= not w31866 and not w31877;
w31879 <= not w14680 and not w31878;
w31880 <= w14680 and not w31865;
w31881 <= not w31879 and not w31880;
w31882 <= not pi0785 and w31881;
w31883 <= not pi0609 and not w31865;
w31884 <= pi0609 and not w31881;
w31885 <= pi1155 and not w31883;
w31886 <= not w31884 and w31885;
w31887 <= not pi0609 and not w31881;
w31888 <= pi0609 and not w31865;
w31889 <= not pi1155 and not w31888;
w31890 <= not w31887 and w31889;
w31891 <= not w31886 and not w31890;
w31892 <= pi0785 and not w31891;
w31893 <= not w31882 and not w31892;
w31894 <= not pi0781 and not w31893;
w31895 <= not pi0618 and not w31865;
w31896 <= pi0618 and w31893;
w31897 <= pi1154 and not w31895;
w31898 <= not w31896 and w31897;
w31899 <= pi0618 and not w31865;
w31900 <= not pi0618 and w31893;
w31901 <= not pi1154 and not w31899;
w31902 <= not w31900 and w31901;
w31903 <= not w31898 and not w31902;
w31904 <= pi0781 and not w31903;
w31905 <= not w31894 and not w31904;
w31906 <= not pi0789 and not w31905;
w31907 <= not pi0619 and not w31865;
w31908 <= pi0619 and w31905;
w31909 <= pi1159 and not w31907;
w31910 <= not w31908 and w31909;
w31911 <= pi0619 and not w31865;
w31912 <= not pi0619 and w31905;
w31913 <= not pi1159 and not w31911;
w31914 <= not w31912 and w31913;
w31915 <= not w31910 and not w31914;
w31916 <= pi0789 and not w31915;
w31917 <= not w31906 and not w31916;
w31918 <= not w15532 and not w31917;
w31919 <= w15532 and w31865;
w31920 <= not w31918 and not w31919;
w31921 <= not w15342 and not w31920;
w31922 <= w15342 and w31865;
w31923 <= not w31921 and not w31922;
w31924 <= not w15367 and not w31923;
w31925 <= w15367 and w31865;
w31926 <= not w31924 and not w31925;
w31927 <= not pi0644 and w31926;
w31928 <= pi0644 and not w31865;
w31929 <= pi0715 and not w31928;
w31930 <= not w31927 and w31929;
w31931 <= w14198 and not w31865;
w31932 <= w14638 and not w31865;
w31933 <= not pi0643 and not w31865;
w31934 <= not pi0200 and not w14204;
w31935 <= w17462 and not w31934;
w31936 <= not pi0200 and w14296;
w31937 <= pi0200 and w14386;
w31938 <= not pi0299 and not w31936;
w31939 <= not w31937 and w31938;
w31940 <= not pi0200 and w14310;
w31941 <= pi0200 and w14401;
w31942 <= pi0299 and not w31940;
w31943 <= not w31941 and w31942;
w31944 <= not w31939 and not w31943;
w31945 <= pi0039 and not w31944;
w31946 <= not pi0200 and not w14489;
w31947 <= pi0200 and w14511;
w31948 <= not pi0039 and not w31946;
w31949 <= not w31947 and w31948;
w31950 <= not w31945 and not w31949;
w31951 <= not pi0038 and not w31950;
w31952 <= not w31935 and not w31951;
w31953 <= w134 and not w31952;
w31954 <= pi0643 and not w31867;
w31955 <= not w31953 and w31954;
w31956 <= not w31933 and not w31955;
w31957 <= not pi0778 and w31956;
w31958 <= not pi0625 and not w31865;
w31959 <= pi0625 and not w31956;
w31960 <= pi1153 and not w31958;
w31961 <= not w31959 and w31960;
w31962 <= not pi0625 and not w31956;
w31963 <= pi0625 and not w31865;
w31964 <= not pi1153 and not w31963;
w31965 <= not w31962 and w31964;
w31966 <= not w31961 and not w31965;
w31967 <= pi0778 and not w31966;
w31968 <= not w31957 and not w31967;
w31969 <= not w14638 and w31968;
w31970 <= not w31932 and not w31969;
w31971 <= not w14202 and w31970;
w31972 <= w14202 and w31865;
w31973 <= not w31971 and not w31972;
w31974 <= not w14198 and w31973;
w31975 <= not w31931 and not w31974;
w31976 <= not w14194 and w31975;
w31977 <= w14194 and w31865;
w31978 <= not w31976 and not w31977;
w31979 <= not pi0792 and not w31978;
w31980 <= pi0628 and not w31865;
w31981 <= not pi0628 and w31978;
w31982 <= not pi1156 and not w31980;
w31983 <= not w31981 and w31982;
w31984 <= not pi0628 and not w31865;
w31985 <= pi0628 and w31978;
w31986 <= pi1156 and not w31984;
w31987 <= not w31985 and w31986;
w31988 <= not w31983 and not w31987;
w31989 <= pi0792 and not w31988;
w31990 <= not w31979 and not w31989;
w31991 <= not pi0787 and not w31990;
w31992 <= pi0647 and not w31990;
w31993 <= not pi0647 and w31865;
w31994 <= not w31992 and not w31993;
w31995 <= pi1157 and not w31994;
w31996 <= pi0647 and not w31865;
w31997 <= not pi0647 and w31990;
w31998 <= not pi1157 and not w31996;
w31999 <= not w31997 and w31998;
w32000 <= not w31995 and not w31999;
w32001 <= pi0787 and not w32000;
w32002 <= not w31991 and not w32001;
w32003 <= pi0644 and w32002;
w32004 <= not pi0629 and w31987;
w32005 <= not w18133 and not w31920;
w32006 <= pi0629 and w31983;
w32007 <= not w32004 and not w32006;
w32008 <= not w32005 and w32007;
w32009 <= pi0792 and not w32008;
w32010 <= pi0609 and w31968;
w32011 <= not pi0643 and w31878;
w32012 <= not w17054 and not w17055;
w32013 <= not pi0200 and not w32012;
w32014 <= pi0038 and pi0200;
w32015 <= w17048 and w32014;
w32016 <= not pi0200 and not w17056;
w32017 <= pi0200 and not w22317;
w32018 <= not pi0038 and not w32016;
w32019 <= not w32017 and w32018;
w32020 <= pi0606 and w134;
w32021 <= not w32015 and w32020;
w32022 <= not w32013 and w32021;
w32023 <= not w32019 and w32022;
w32024 <= not w14210 and not w14918;
w32025 <= w31935 and not w32024;
w32026 <= not pi0200 and not w17030;
w32027 <= pi0200 and not w17038;
w32028 <= not pi0038 and not w32026;
w32029 <= not w32027 and w32028;
w32030 <= not w32025 and not w32029;
w32031 <= not pi0606 and w134;
w32032 <= not w32030 and w32031;
w32033 <= not w31867 and not w32023;
w32034 <= not w32032 and w32033;
w32035 <= pi0643 and not w32034;
w32036 <= not w32011 and not w32035;
w32037 <= not pi0625 and w32036;
w32038 <= pi0625 and not w31878;
w32039 <= not pi1153 and not w32038;
w32040 <= not w32037 and w32039;
w32041 <= not pi0608 and not w31961;
w32042 <= not w32040 and w32041;
w32043 <= pi0625 and w32036;
w32044 <= not pi0625 and not w31878;
w32045 <= pi1153 and not w32044;
w32046 <= not w32043 and w32045;
w32047 <= pi0608 and not w31965;
w32048 <= not w32046 and w32047;
w32049 <= not w32042 and not w32048;
w32050 <= pi0778 and not w32049;
w32051 <= not pi0778 and w32036;
w32052 <= not w32050 and not w32051;
w32053 <= not pi0609 and not w32052;
w32054 <= not pi1155 and not w32010;
w32055 <= not w32053 and w32054;
w32056 <= not pi0660 and not w31886;
w32057 <= not w32055 and w32056;
w32058 <= not pi0609 and w31968;
w32059 <= pi0609 and not w32052;
w32060 <= pi1155 and not w32058;
w32061 <= not w32059 and w32060;
w32062 <= pi0660 and not w31890;
w32063 <= not w32061 and w32062;
w32064 <= not w32057 and not w32063;
w32065 <= pi0785 and not w32064;
w32066 <= not pi0785 and not w32052;
w32067 <= not w32065 and not w32066;
w32068 <= not pi0618 and not w32067;
w32069 <= pi0618 and not w31970;
w32070 <= not pi1154 and not w32069;
w32071 <= not w32068 and w32070;
w32072 <= not pi0627 and not w31898;
w32073 <= not w32071 and w32072;
w32074 <= pi0618 and not w32067;
w32075 <= not pi0618 and not w31970;
w32076 <= pi1154 and not w32075;
w32077 <= not w32074 and w32076;
w32078 <= pi0627 and not w31902;
w32079 <= not w32077 and w32078;
w32080 <= not w32073 and not w32079;
w32081 <= pi0781 and not w32080;
w32082 <= not pi0781 and not w32067;
w32083 <= not w32081 and not w32082;
w32084 <= not pi0789 and w32083;
w32085 <= not pi0619 and not w32083;
w32086 <= pi0619 and w31973;
w32087 <= not pi1159 and not w32086;
w32088 <= not w32085 and w32087;
w32089 <= not pi0648 and not w31910;
w32090 <= not w32088 and w32089;
w32091 <= pi0619 and not w32083;
w32092 <= not pi0619 and w31973;
w32093 <= pi1159 and not w32092;
w32094 <= not w32091 and w32093;
w32095 <= pi0648 and not w31914;
w32096 <= not w32094 and w32095;
w32097 <= pi0789 and not w32090;
w32098 <= not w32096 and w32097;
w32099 <= w15533 and not w32084;
w32100 <= not w32098 and w32099;
w32101 <= w15434 and not w31975;
w32102 <= pi0626 and w31865;
w32103 <= not pi0626 and not w31917;
w32104 <= w14192 and not w32102;
w32105 <= not w32103 and w32104;
w32106 <= not pi0626 and w31865;
w32107 <= pi0626 and not w31917;
w32108 <= w14191 and not w32106;
w32109 <= not w32107 and w32108;
w32110 <= not w32101 and not w32105;
w32111 <= not w32109 and w32110;
w32112 <= pi0788 and not w32111;
w32113 <= not w17927 and not w32112;
w32114 <= not w32100 and w32113;
w32115 <= not w32009 and not w32114;
w32116 <= not w17769 and not w32115;
w32117 <= pi0630 and w31999;
w32118 <= not w18122 and not w31923;
w32119 <= w15364 and not w31994;
w32120 <= not w32117 and not w32118;
w32121 <= not w32119 and w32120;
w32122 <= pi0787 and not w32121;
w32123 <= not w32116 and not w32122;
w32124 <= not pi0644 and w32123;
w32125 <= not pi0715 and not w32003;
w32126 <= not w32124 and w32125;
w32127 <= not pi1160 and not w31930;
w32128 <= not w32126 and w32127;
w32129 <= not pi0644 and w32002;
w32130 <= pi0644 and w32123;
w32131 <= pi0715 and not w32129;
w32132 <= not w32130 and w32131;
w32133 <= pi0644 and w31926;
w32134 <= not pi0644 and not w31865;
w32135 <= not pi0715 and not w32134;
w32136 <= not w32133 and w32135;
w32137 <= pi1160 and not w32136;
w32138 <= not w32132 and w32137;
w32139 <= not w32128 and not w32138;
w32140 <= pi0790 and not w32139;
w32141 <= not pi0790 and w32123;
w32142 <= not w32140 and not w32141;
w32143 <= w4989 and not w32142;
w32144 <= not pi0200 and not w4989;
w32145 <= not w32143 and not w32144;
w32146 <= pi0233 and pi0237;
w32147 <= pi0057 and pi0332;
w32148 <= w135 and w4136;
w32149 <= w84 and w32148;
w32150 <= not pi0332 and not w32149;
w32151 <= w3867 and not w32150;
w32152 <= pi0332 and not w3867;
w32153 <= pi0059 and not w32152;
w32154 <= not w32151 and w32153;
w32155 <= pi0332 and not w92;
w32156 <= not pi0059 and not w32155;
w32157 <= pi0055 and w32150;
w32158 <= pi0074 and pi0332;
w32159 <= not pi0055 and not w32158;
w32160 <= w289 and w8649;
w32161 <= pi0468 and w3755;
w32162 <= not pi0299 and pi0587;
w32163 <= not w18607 and not w32162;
w32164 <= not pi0468 and not w32163;
w32165 <= not w32161 and not w32164;
w32166 <= w32160 and not w32165;
w32167 <= not pi0332 and not w32166;
w32168 <= w4926 and not w32167;
w32169 <= w84 and w4148;
w32170 <= not pi0332 and not w32169;
w32171 <= w13188 and not w32170;
w32172 <= pi0332 and not w174;
w32173 <= not w32171 and not w32172;
w32174 <= not w32168 and w32173;
w32175 <= not pi0074 and not w32174;
w32176 <= w32159 and not w32175;
w32177 <= w92 and not w32157;
w32178 <= not w32176 and w32177;
w32179 <= w32156 and not w32178;
w32180 <= not pi0057 and not w32154;
w32181 <= not w32179 and w32180;
w32182 <= not w32147 and not w32181;
w32183 <= not w32146 and not w32182;
w32184 <= not pi0332 and not w3755;
w32185 <= not pi0947 and not w32184;
w32186 <= pi0096 and pi0210;
w32187 <= pi0332 and w32186;
w32188 <= not pi0032 and pi0070;
w32189 <= not pi0070 and not pi0841;
w32190 <= pi0032 and w32189;
w32191 <= not w32188 and not w32190;
w32192 <= not pi0210 and not w32191;
w32193 <= not pi0032 and not pi0096;
w32194 <= pi0070 and w32193;
w32195 <= not pi0332 and not w32194;
w32196 <= not w32192 and w32195;
w32197 <= not w32187 and not w32196;
w32198 <= not w3760 and w32197;
w32199 <= w3755 and not w32198;
w32200 <= w32185 and not w32199;
w32201 <= w3755 and not w32197;
w32202 <= pi0332 and pi0468;
w32203 <= not pi0468 and not w32196;
w32204 <= not w32202 and not w32203;
w32205 <= not w3755 and w32204;
w32206 <= pi0947 and not w32201;
w32207 <= not w32205 and w32206;
w32208 <= not w32200 and not w32207;
w32209 <= pi0057 and not w32208;
w32210 <= not w3867 and w32208;
w32211 <= not w135 and w32208;
w32212 <= pi0032 and not w32189;
w32213 <= not pi0095 and w299;
w32214 <= not w32212 and w32213;
w32215 <= w269 and w32214;
w32216 <= w291 and w32215;
w32217 <= w32191 and not w32216;
w32218 <= not pi0210 and not w32217;
w32219 <= not pi0095 and w538;
w32220 <= not pi0070 and not w32219;
w32221 <= w32193 and not w32220;
w32222 <= pi0210 and w32221;
w32223 <= not pi0332 and not w32218;
w32224 <= not w32222 and w32223;
w32225 <= not w32187 and not w32224;
w32226 <= not w3760 and w32225;
w32227 <= w3755 and not w32226;
w32228 <= w32185 and not w32227;
w32229 <= w3755 and not w32225;
w32230 <= not pi0468 and not w32224;
w32231 <= not w32202 and not w32230;
w32232 <= not w3755 and w32231;
w32233 <= pi0947 and not w32229;
w32234 <= not w32232 and w32233;
w32235 <= not w32228 and not w32234;
w32236 <= w135 and w32235;
w32237 <= not w32211 and not w32236;
w32238 <= w3867 and not w32237;
w32239 <= pi0059 and not w32210;
w32240 <= not w32238 and w32239;
w32241 <= not w92 and w32208;
w32242 <= pi0055 and w32237;
w32243 <= not pi0074 and w174;
w32244 <= pi0299 and not w32208;
w32245 <= pi0096 and pi0198;
w32246 <= pi0332 and w32245;
w32247 <= not pi0198 and not w32191;
w32248 <= w32195 and not w32247;
w32249 <= not w32246 and not w32248;
w32250 <= w3755 and not w32249;
w32251 <= w4146 and not w32248;
w32252 <= w32184 and not w32251;
w32253 <= not pi0299 and not w4145;
w32254 <= not w32250 and w32253;
w32255 <= not w32252 and w32254;
w32256 <= not w32243 and not w32255;
w32257 <= not w32244 and w32256;
w32258 <= w289 and w525;
w32259 <= w32214 and w32258;
w32260 <= w32191 and not w32259;
w32261 <= not pi0210 and not w32260;
w32262 <= not pi0095 and w80;
w32263 <= w32258 and w32262;
w32264 <= not pi0070 and not w32263;
w32265 <= w32193 and not w32264;
w32266 <= pi0210 and w32265;
w32267 <= not pi0332 and not w32261;
w32268 <= not w32266 and w32267;
w32269 <= not w32187 and not w32268;
w32270 <= not w3760 and w32269;
w32271 <= w3755 and not w32270;
w32272 <= w32185 and not w32271;
w32273 <= w3755 and not w32269;
w32274 <= not pi0468 and not w32268;
w32275 <= not w32202 and not w32274;
w32276 <= not w3755 and w32275;
w32277 <= pi0947 and not w32273;
w32278 <= not w32276 and w32277;
w32279 <= pi0299 and not w32272;
w32280 <= not w32278 and w32279;
w32281 <= not pi0587 and not w32184;
w32282 <= not pi0198 and not w32260;
w32283 <= pi0198 and w32265;
w32284 <= not pi0332 and not w32282;
w32285 <= not w32283 and w32284;
w32286 <= not w32246 and not w32285;
w32287 <= not w3760 and w32286;
w32288 <= w3755 and not w32287;
w32289 <= w32281 and not w32288;
w32290 <= w3755 and not w32286;
w32291 <= not pi0468 and not w32285;
w32292 <= not w3755 and not w32202;
w32293 <= not w32291 and w32292;
w32294 <= pi0587 and not w32290;
w32295 <= not w32293 and w32294;
w32296 <= not pi0299 and not w32289;
w32297 <= not w32295 and w32296;
w32298 <= not w32280 and not w32297;
w32299 <= w4926 and not w32298;
w32300 <= pi0299 and not w32235;
w32301 <= not pi0198 and not w32217;
w32302 <= pi0198 and w32221;
w32303 <= not pi0332 and not w32301;
w32304 <= not w32302 and w32303;
w32305 <= not w32246 and not w32304;
w32306 <= not w3760 and w32305;
w32307 <= w3755 and not w32306;
w32308 <= w32281 and not w32307;
w32309 <= w3755 and not w32305;
w32310 <= not pi0468 and not w32304;
w32311 <= w32292 and not w32310;
w32312 <= pi0587 and not w32309;
w32313 <= not w32311 and w32312;
w32314 <= not w32308 and not w32313;
w32315 <= not pi0299 and not w32314;
w32316 <= w13188 and not w32300;
w32317 <= not w32315 and w32316;
w32318 <= not w32299 and not w32317;
w32319 <= not pi0074 and not w32318;
w32320 <= not pi0055 and not w32257;
w32321 <= not w32319 and w32320;
w32322 <= w92 and not w32242;
w32323 <= not w32321 and w32322;
w32324 <= not pi0059 and not w32241;
w32325 <= not w32323 and w32324;
w32326 <= not w32240 and not w32325;
w32327 <= not pi0057 and not w32326;
w32328 <= not w32209 and not w32327;
w32329 <= w32146 and not w32328;
w32330 <= not w32183 and not w32329;
w32331 <= not pi0201 and not w32330;
w32332 <= not w4136 and not w14042;
w32333 <= w4146 and w32245;
w32334 <= w14042 and not w32333;
w32335 <= not w14042 and not w32186;
w32336 <= not w32332 and not w32334;
w32337 <= not w32335 and w32336;
w32338 <= w32146 and w32337;
w32339 <= pi0201 and not w32338;
w32340 <= not w32331 and not w32339;
w32341 <= not pi0233 and pi0237;
w32342 <= not w32182 and not w32341;
w32343 <= not w32328 and w32341;
w32344 <= not w32342 and not w32343;
w32345 <= not pi0202 and not w32344;
w32346 <= w32337 and w32341;
w32347 <= pi0202 and not w32346;
w32348 <= not w32345 and not w32347;
w32349 <= not pi0233 and not pi0237;
w32350 <= not w32182 and not w32349;
w32351 <= not w32328 and w32349;
w32352 <= not w32350 and not w32351;
w32353 <= not pi0203 and not w32352;
w32354 <= w32337 and w32349;
w32355 <= pi0203 and not w32354;
w32356 <= not w32353 and not w32355;
w32357 <= w135 and w3873;
w32358 <= w84 and w32357;
w32359 <= not pi0332 and not w32358;
w32360 <= w3867 and not w32359;
w32361 <= w32153 and not w32360;
w32362 <= pi0055 and w32359;
w32363 <= not pi0468 and pi0602;
w32364 <= pi0468 and w3758;
w32365 <= not w32363 and not w32364;
w32366 <= not pi0299 and not w32365;
w32367 <= not w3887 and not w32366;
w32368 <= w84 and not w32367;
w32369 <= not pi0332 and not w32368;
w32370 <= w13188 and not w32369;
w32371 <= not pi0299 and not pi0602;
w32372 <= pi0299 and not pi0907;
w32373 <= not pi0468 and not w32371;
w32374 <= not w32372 and w32373;
w32375 <= not w32364 and not w32374;
w32376 <= w32160 and not w32375;
w32377 <= not pi0332 and not w32376;
w32378 <= w4926 and not w32377;
w32379 <= not w32370 and not w32378;
w32380 <= not pi0074 and not w32379;
w32381 <= w32159 and not w32172;
w32382 <= not w32380 and w32381;
w32383 <= w92 and not w32362;
w32384 <= not w32382 and w32383;
w32385 <= w32156 and not w32384;
w32386 <= not pi0057 and not w32361;
w32387 <= not w32385 and w32386;
w32388 <= not w32147 and not w32387;
w32389 <= not w32146 and not w32388;
w32390 <= not pi0332 and not w3758;
w32391 <= not pi0907 and not w32390;
w32392 <= w3758 and not w32198;
w32393 <= w32391 and not w32392;
w32394 <= w3758 and not w32197;
w32395 <= not w3758 and w32204;
w32396 <= pi0907 and not w32394;
w32397 <= not w32395 and w32396;
w32398 <= not w32393 and not w32397;
w32399 <= pi0057 and not w32398;
w32400 <= not w3867 and w32398;
w32401 <= not w135 and w32398;
w32402 <= w3758 and not w32225;
w32403 <= not w3758 and w32231;
w32404 <= pi0907 and not w32402;
w32405 <= not w32403 and w32404;
w32406 <= pi0332 and not w14220;
w32407 <= pi0680 and not w32406;
w32408 <= not w32226 and w32407;
w32409 <= w32391 and not w32408;
w32410 <= not w32405 and not w32409;
w32411 <= w135 and w32410;
w32412 <= not w32401 and not w32411;
w32413 <= w3867 and not w32412;
w32414 <= pi0059 and not w32400;
w32415 <= not w32413 and w32414;
w32416 <= not w92 and w32398;
w32417 <= pi0055 and w32412;
w32418 <= pi0299 and w32410;
w32419 <= w3758 and w32245;
w32420 <= pi0332 and not w32419;
w32421 <= not pi0299 and not w32420;
w32422 <= w3889 and w32305;
w32423 <= w32421 and not w32422;
w32424 <= not w32418 and not w32423;
w32425 <= w13188 and not w32424;
w32426 <= w3889 and w32286;
w32427 <= w32421 and not w32426;
w32428 <= w3758 and not w32270;
w32429 <= w32391 and not w32428;
w32430 <= w3758 and not w32269;
w32431 <= not w3758 and w32275;
w32432 <= pi0907 and not w32430;
w32433 <= not w32431 and w32432;
w32434 <= pi0299 and not w32429;
w32435 <= not w32433 and w32434;
w32436 <= not w32427 and not w32435;
w32437 <= w4926 and not w32436;
w32438 <= not w32425 and not w32437;
w32439 <= not pi0074 and not w32438;
w32440 <= pi0299 and not w32398;
w32441 <= w32249 and not w32365;
w32442 <= not w32420 and not w32441;
w32443 <= not pi0299 and not w32442;
w32444 <= not w32243 and not w32443;
w32445 <= not w32440 and w32444;
w32446 <= not pi0055 and not w32445;
w32447 <= not w32439 and w32446;
w32448 <= w92 and not w32417;
w32449 <= not w32447 and w32448;
w32450 <= not pi0059 and not w32416;
w32451 <= not w32449 and w32450;
w32452 <= not w32415 and not w32451;
w32453 <= not pi0057 and not w32452;
w32454 <= not w32399 and not w32453;
w32455 <= w32146 and not w32454;
w32456 <= not w32389 and not w32455;
w32457 <= not pi0204 and not w32456;
w32458 <= not w3873 and not w14042;
w32459 <= w3889 and w32245;
w32460 <= w14042 and not w32459;
w32461 <= not w32335 and not w32458;
w32462 <= not w32460 and w32461;
w32463 <= w32146 and w32462;
w32464 <= pi0204 and not w32463;
w32465 <= not w32457 and not w32464;
w32466 <= not w32341 and not w32388;
w32467 <= w32341 and not w32454;
w32468 <= not w32466 and not w32467;
w32469 <= not pi0205 and not w32468;
w32470 <= w32341 and w32462;
w32471 <= pi0205 and not w32470;
w32472 <= not w32469 and not w32471;
w32473 <= pi0233 and not pi0237;
w32474 <= not w32388 and not w32473;
w32475 <= not w32454 and w32473;
w32476 <= not w32474 and not w32475;
w32477 <= not pi0206 and not w32476;
w32478 <= w32462 and w32473;
w32479 <= pi0206 and not w32478;
w32480 <= not w32477 and not w32479;
w32481 <= not w16709 and w21948;
w32482 <= w16714 and w32481;
w32483 <= not w16705 and w32482;
w32484 <= pi0207 and not w32483;
w32485 <= w14198 and not w14622;
w32486 <= w134 and w21951;
w32487 <= not pi0778 and not w32486;
w32488 <= not pi0625 and not w14622;
w32489 <= pi0625 and not w32486;
w32490 <= not w32488 and not w32489;
w32491 <= pi1153 and not w32490;
w32492 <= pi0625 and not w14622;
w32493 <= not pi0625 and not w32486;
w32494 <= not w32492 and not w32493;
w32495 <= not pi1153 and not w32494;
w32496 <= not w32491 and not w32495;
w32497 <= pi0778 and not w32496;
w32498 <= not w32487 and not w32497;
w32499 <= not w14638 and not w32498;
w32500 <= not w14622 and w14638;
w32501 <= not w32499 and not w32500;
w32502 <= not w14202 and w32501;
w32503 <= w14202 and w14622;
w32504 <= not w32502 and not w32503;
w32505 <= not w14198 and w32504;
w32506 <= not w32485 and not w32505;
w32507 <= not w14194 and w32506;
w32508 <= w14194 and w14622;
w32509 <= not w32507 and not w32508;
w32510 <= not w16705 and not w32509;
w32511 <= w14622 and w15419;
w32512 <= not w32510 and not w32511;
w32513 <= not pi0207 and not w32512;
w32514 <= not w32484 and not w32513;
w32515 <= pi0710 and not w32514;
w32516 <= not pi0207 and not w14622;
w32517 <= not pi0710 and not w32516;
w32518 <= not w32515 and not w32517;
w32519 <= not pi0787 and not w32518;
w32520 <= not pi0647 and w32518;
w32521 <= pi0647 and w32516;
w32522 <= not pi1157 and not w32521;
w32523 <= not w32520 and w32522;
w32524 <= not pi0647 and w32516;
w32525 <= pi0647 and w32518;
w32526 <= pi1157 and not w32524;
w32527 <= not w32525 and w32526;
w32528 <= not w32523 and not w32527;
w32529 <= pi0787 and not w32528;
w32530 <= not w32519 and not w32529;
w32531 <= not pi0644 and w32530;
w32532 <= not pi0630 and w32527;
w32533 <= not w14622 and w14680;
w32534 <= w134 and w17002;
w32535 <= not w14680 and not w32534;
w32536 <= not w32533 and not w32535;
w32537 <= not pi0785 and not w32536;
w32538 <= not w14622 and not w14859;
w32539 <= not pi0609 and w32535;
w32540 <= not w32538 and not w32539;
w32541 <= not pi1155 and not w32540;
w32542 <= not w14622 and not w14854;
w32543 <= pi0609 and w32535;
w32544 <= not w32542 and not w32543;
w32545 <= pi1155 and not w32544;
w32546 <= not w32541 and not w32545;
w32547 <= pi0785 and not w32546;
w32548 <= not w32537 and not w32547;
w32549 <= not pi0781 and not w32548;
w32550 <= not pi0618 and w32548;
w32551 <= pi0618 and w14622;
w32552 <= not pi1154 and not w32551;
w32553 <= not w32550 and w32552;
w32554 <= not pi0618 and w14622;
w32555 <= pi0618 and w32548;
w32556 <= pi1154 and not w32554;
w32557 <= not w32555 and w32556;
w32558 <= not w32553 and not w32557;
w32559 <= pi0781 and not w32558;
w32560 <= not w32549 and not w32559;
w32561 <= not pi0789 and not w32560;
w32562 <= not pi0619 and w32560;
w32563 <= pi0619 and w14622;
w32564 <= not pi1159 and not w32563;
w32565 <= not w32562 and w32564;
w32566 <= not pi0619 and w14622;
w32567 <= pi0619 and w32560;
w32568 <= pi1159 and not w32566;
w32569 <= not w32567 and w32568;
w32570 <= not w32565 and not w32569;
w32571 <= pi0789 and not w32570;
w32572 <= not w32561 and not w32571;
w32573 <= not w15532 and w32572;
w32574 <= w14622 and w15532;
w32575 <= not w32573 and not w32574;
w32576 <= not w15342 and not w32575;
w32577 <= w14622 and w15342;
w32578 <= not w32576 and not w32577;
w32579 <= not pi0207 and not w32578;
w32580 <= w134 and not w22010;
w32581 <= not w14680 and w32580;
w32582 <= not w17788 and w32581;
w32583 <= not w17798 and w32582;
w32584 <= not w17794 and w32583;
w32585 <= not w15532 and w32584;
w32586 <= not w15342 and w32585;
w32587 <= pi0207 and not w32586;
w32588 <= pi0623 and not w32587;
w32589 <= not w32579 and w32588;
w32590 <= not pi0623 and w32516;
w32591 <= not w32589 and not w32590;
w32592 <= not w18122 and w32591;
w32593 <= pi0630 and w32523;
w32594 <= not w32532 and not w32592;
w32595 <= not w32593 and w32594;
w32596 <= pi0787 and not w32595;
w32597 <= not pi0710 and not w32591;
w32598 <= not pi0628 and not w14622;
w32599 <= pi0628 and w32509;
w32600 <= not w32598 and not w32599;
w32601 <= not pi0629 and not w32600;
w32602 <= not w32598 and not w32601;
w32603 <= pi1156 and not w32602;
w32604 <= pi0628 and not w14622;
w32605 <= not pi1156 and w32604;
w32606 <= not pi0628 and w32509;
w32607 <= not w32604 and not w32606;
w32608 <= w15340 and not w32607;
w32609 <= not w32605 and not w32608;
w32610 <= not w32603 and w32609;
w32611 <= pi0792 and not w32610;
w32612 <= pi1159 and not w14622;
w32613 <= pi0619 and w32504;
w32614 <= pi1154 and not w14622;
w32615 <= pi0618 and not w32501;
w32616 <= pi1155 and not w14622;
w32617 <= pi0609 and not w32498;
w32618 <= w134 and not w17040;
w32619 <= not pi0778 and not w32618;
w32620 <= not pi0625 and not w32618;
w32621 <= not w32492 and not w32620;
w32622 <= not pi1153 and not w32621;
w32623 <= not pi0608 and not w32491;
w32624 <= not w32622 and w32623;
w32625 <= pi0625 and not w32618;
w32626 <= not w32488 and not w32625;
w32627 <= pi1153 and not w32626;
w32628 <= pi0608 and not w32495;
w32629 <= not w32627 and w32628;
w32630 <= pi0778 and not w32624;
w32631 <= not w32629 and w32630;
w32632 <= not w32619 and not w32631;
w32633 <= not pi0609 and not w32632;
w32634 <= not w32617 and not w32633;
w32635 <= not pi1155 and not w32634;
w32636 <= not pi0660 and not w32616;
w32637 <= not w32635 and w32636;
w32638 <= not pi1155 and not w14622;
w32639 <= not pi0609 and not w32498;
w32640 <= pi0609 and not w32632;
w32641 <= not w32639 and not w32640;
w32642 <= pi1155 and not w32641;
w32643 <= pi0660 and not w32638;
w32644 <= not w32642 and w32643;
w32645 <= not w32637 and not w32644;
w32646 <= pi0785 and not w32645;
w32647 <= not pi0785 and w32632;
w32648 <= not w32646 and not w32647;
w32649 <= not pi0618 and w32648;
w32650 <= not w32615 and not w32649;
w32651 <= not pi1154 and not w32650;
w32652 <= not pi0627 and not w32614;
w32653 <= not w32651 and w32652;
w32654 <= not pi1154 and not w14622;
w32655 <= not pi0618 and not w32501;
w32656 <= pi0618 and w32648;
w32657 <= not w32655 and not w32656;
w32658 <= pi1154 and not w32657;
w32659 <= pi0627 and not w32654;
w32660 <= not w32658 and w32659;
w32661 <= not w32653 and not w32660;
w32662 <= pi0781 and not w32661;
w32663 <= not pi0781 and not w32648;
w32664 <= not w32662 and not w32663;
w32665 <= not pi0619 and w32664;
w32666 <= not w32613 and not w32665;
w32667 <= not pi1159 and not w32666;
w32668 <= not pi0648 and not w32612;
w32669 <= not w32667 and w32668;
w32670 <= not pi1159 and not w14622;
w32671 <= not pi0619 and w32504;
w32672 <= pi0619 and w32664;
w32673 <= not w32671 and not w32672;
w32674 <= pi1159 and not w32673;
w32675 <= pi0648 and not w32670;
w32676 <= not w32674 and w32675;
w32677 <= not w32669 and not w32676;
w32678 <= pi0789 and not w32677;
w32679 <= not pi0789 and not w32664;
w32680 <= not w32678 and not w32679;
w32681 <= not pi0788 and not w32680;
w32682 <= pi0641 and not w14622;
w32683 <= pi0626 and w32506;
w32684 <= not pi0626 and not w32680;
w32685 <= not pi0641 and not w32683;
w32686 <= not w32684 and w32685;
w32687 <= not pi1158 and not w32682;
w32688 <= not w32686 and w32687;
w32689 <= not pi0641 and not w14622;
w32690 <= not pi0626 and w32506;
w32691 <= pi0626 and not w32680;
w32692 <= pi0641 and not w32690;
w32693 <= not w32691 and w32692;
w32694 <= pi1158 and not w32689;
w32695 <= not w32693 and w32694;
w32696 <= not w32688 and not w32695;
w32697 <= pi0788 and not w32696;
w32698 <= not w17927 and not w32681;
w32699 <= not w32697 and w32698;
w32700 <= not w32611 and not w32699;
w32701 <= not pi0207 and not w32700;
w32702 <= pi0609 and not w32481;
w32703 <= not pi0778 and not w31643;
w32704 <= not pi0625 and w31643;
w32705 <= not pi1153 and not w32704;
w32706 <= pi0625 and w21948;
w32707 <= pi1153 and not w32706;
w32708 <= not pi0608 and not w32707;
w32709 <= not w32705 and w32708;
w32710 <= pi0625 and w31643;
w32711 <= pi1153 and not w32710;
w32712 <= not pi0625 and w21948;
w32713 <= not pi1153 and not w32712;
w32714 <= pi0608 and not w32713;
w32715 <= not w32711 and w32714;
w32716 <= pi0778 and not w32709;
w32717 <= not w32715 and w32716;
w32718 <= not w32703 and not w32717;
w32719 <= not pi0609 and not w32718;
w32720 <= w14636 and not w32702;
w32721 <= not w32719 and w32720;
w32722 <= pi0609 and not w32718;
w32723 <= not pi0609 and not w32481;
w32724 <= w14635 and not w32723;
w32725 <= not w32722 and w32724;
w32726 <= not w32721 and not w32725;
w32727 <= pi0785 and not w32726;
w32728 <= not pi0785 and w32718;
w32729 <= not w32727 and not w32728;
w32730 <= not pi0781 and w32729;
w32731 <= not pi0618 and w32729;
w32732 <= not w14638 and w32481;
w32733 <= pi0618 and not w32732;
w32734 <= w14200 and not w32733;
w32735 <= not w32731 and w32734;
w32736 <= not pi0618 and not w32732;
w32737 <= pi0618 and w32729;
w32738 <= w14199 and not w32736;
w32739 <= not w32737 and w32738;
w32740 <= pi0781 and not w32735;
w32741 <= not w32739 and w32740;
w32742 <= not w21178 and not w32730;
w32743 <= not w32741 and w32742;
w32744 <= w16713 and w32481;
w32745 <= w14197 and w17794;
w32746 <= w32744 and w32745;
w32747 <= not w32743 and not w32746;
w32748 <= not pi0788 and w32747;
w32749 <= not w14198 and w32744;
w32750 <= pi0626 and not w32749;
w32751 <= not pi0641 and not w32750;
w32752 <= not pi0626 and w32747;
w32753 <= not pi1158 and w32751;
w32754 <= not w32752 and w32753;
w32755 <= pi0626 and w32747;
w32756 <= not pi0626 and not w32749;
w32757 <= pi0641 and not w32756;
w32758 <= pi1158 and w32757;
w32759 <= not w32755 and w32758;
w32760 <= pi0788 and not w32754;
w32761 <= not w32759 and w32760;
w32762 <= not w17927 and not w32748;
w32763 <= not w32761 and w32762;
w32764 <= w15342 and w15418;
w32765 <= w32482 and w32764;
w32766 <= not w32763 and not w32765;
w32767 <= pi0207 and not w32766;
w32768 <= not pi0623 and not w32767;
w32769 <= not w32701 and w32768;
w32770 <= not pi1156 and not w32482;
w32771 <= pi1156 and not w32585;
w32772 <= w18129 and not w32770;
w32773 <= not w32771 and w32772;
w32774 <= pi1156 and not w32482;
w32775 <= not pi1156 and not w32585;
w32776 <= w18131 and not w32774;
w32777 <= not w32775 and w32776;
w32778 <= not w32773 and not w32777;
w32779 <= pi0792 and not w32778;
w32780 <= w15431 and w32584;
w32781 <= not pi1159 and not w32583;
w32782 <= pi1159 and not w32744;
w32783 <= not pi0619 and pi0648;
w32784 <= not w32781 and w32783;
w32785 <= not w32782 and w32784;
w32786 <= pi1159 and not w32583;
w32787 <= not pi1159 and not w32744;
w32788 <= pi0619 and not pi0648;
w32789 <= not w32786 and w32788;
w32790 <= not w32787 and w32789;
w32791 <= pi0789 and not w32785;
w32792 <= not w32790 and w32791;
w32793 <= pi0789 and not w32792;
w32794 <= not pi1154 and not w32733;
w32795 <= w17796 and w32582;
w32796 <= not pi0627 and not w32795;
w32797 <= not w32794 and w32796;
w32798 <= w17795 and w32582;
w32799 <= not pi0778 and not w31648;
w32800 <= not pi0625 and w31648;
w32801 <= pi0625 and w32580;
w32802 <= not pi1153 and not w32801;
w32803 <= not w32800 and w32802;
w32804 <= w32708 and not w32803;
w32805 <= not pi0625 and w32580;
w32806 <= pi0625 and w31648;
w32807 <= pi1153 and not w32805;
w32808 <= not w32806 and w32807;
w32809 <= w32714 and not w32808;
w32810 <= pi0778 and not w32804;
w32811 <= not w32809 and w32810;
w32812 <= not w32799 and not w32811;
w32813 <= not pi0785 and not w32812;
w32814 <= w17786 and w32581;
w32815 <= not pi0609 and not w32812;
w32816 <= not pi1155 and not w32702;
w32817 <= not w32815 and w32816;
w32818 <= not pi0660 and not w32814;
w32819 <= not w32817 and w32818;
w32820 <= w17785 and w32581;
w32821 <= pi0609 and not w32812;
w32822 <= pi1155 and not w32723;
w32823 <= not w32821 and w32822;
w32824 <= pi0660 and not w32820;
w32825 <= not w32823 and w32824;
w32826 <= not w32819 and not w32825;
w32827 <= pi0785 and not w32826;
w32828 <= not w32813 and not w32827;
w32829 <= pi0618 and not w32828;
w32830 <= pi1154 and not w32736;
w32831 <= not w32829 and w32830;
w32832 <= pi0627 and not w32798;
w32833 <= not w32831 and w32832;
w32834 <= not w32797 and not w32833;
w32835 <= pi0781 and not w32834;
w32836 <= not pi0618 and not pi0627;
w32837 <= pi0781 and not w32836;
w32838 <= not w32828 and not w32837;
w32839 <= not w21177 and w32792;
w32840 <= not w32838 and not w32839;
w32841 <= not w32835 and w32840;
w32842 <= not w32793 and not w32841;
w32843 <= not pi0626 and w32842;
w32844 <= w32751 and not w32843;
w32845 <= not pi1158 and not w32780;
w32846 <= not w32844 and w32845;
w32847 <= w15432 and w32584;
w32848 <= pi0626 and w32842;
w32849 <= w32757 and not w32848;
w32850 <= pi1158 and not w32847;
w32851 <= not w32849 and w32850;
w32852 <= not w32846 and not w32851;
w32853 <= pi0788 and not w32852;
w32854 <= not pi0788 and w32842;
w32855 <= not w17927 and not w32854;
w32856 <= not w32853 and w32855;
w32857 <= not w32779 and not w32856;
w32858 <= pi0207 and not w32857;
w32859 <= w134 and w17051;
w32860 <= not pi0778 and not w32859;
w32861 <= not pi0625 and w32534;
w32862 <= pi0625 and w32859;
w32863 <= pi1153 and not w32862;
w32864 <= not w32861 and w32863;
w32865 <= w32628 and not w32864;
w32866 <= not pi0625 and w32859;
w32867 <= pi0625 and w32534;
w32868 <= not pi1153 and not w32866;
w32869 <= not w32867 and w32868;
w32870 <= w32623 and not w32869;
w32871 <= pi0778 and not w32865;
w32872 <= not w32870 and w32871;
w32873 <= not w32860 and not w32872;
w32874 <= not pi0609 and not w32873;
w32875 <= not w32617 and not w32874;
w32876 <= not pi1155 and not w32875;
w32877 <= not pi0660 and not w32545;
w32878 <= not w32876 and w32877;
w32879 <= pi0609 and not w32873;
w32880 <= not w32639 and not w32879;
w32881 <= pi1155 and not w32880;
w32882 <= pi0660 and not w32541;
w32883 <= not w32881 and w32882;
w32884 <= not w32878 and not w32883;
w32885 <= pi0785 and not w32884;
w32886 <= not pi0785 and w32873;
w32887 <= not w32885 and not w32886;
w32888 <= not pi0618 and w32887;
w32889 <= not w32615 and not w32888;
w32890 <= not pi1154 and not w32889;
w32891 <= not pi0627 and not w32557;
w32892 <= not w32890 and w32891;
w32893 <= pi0618 and w32887;
w32894 <= not w32655 and not w32893;
w32895 <= pi1154 and not w32894;
w32896 <= pi0627 and not w32553;
w32897 <= not w32895 and w32896;
w32898 <= not w32892 and not w32897;
w32899 <= pi0781 and not w32898;
w32900 <= not pi0781 and not w32887;
w32901 <= not w32899 and not w32900;
w32902 <= not pi0789 and w32901;
w32903 <= not pi0619 and w32901;
w32904 <= not w32613 and not w32903;
w32905 <= not pi1159 and not w32904;
w32906 <= not pi0648 and not w32569;
w32907 <= not w32905 and w32906;
w32908 <= pi0619 and w32901;
w32909 <= not w32671 and not w32908;
w32910 <= pi1159 and not w32909;
w32911 <= pi0648 and not w32565;
w32912 <= not w32910 and w32911;
w32913 <= pi0789 and not w32907;
w32914 <= not w32912 and w32913;
w32915 <= w15533 and not w32902;
w32916 <= not w32914 and w32915;
w32917 <= pi0641 and not w32506;
w32918 <= w15428 and not w32689;
w32919 <= not w32917 and w32918;
w32920 <= not w14193 and not w15433;
w32921 <= w32572 and w32920;
w32922 <= not pi0641 and not w32506;
w32923 <= w15429 and not w32682;
w32924 <= not w32922 and w32923;
w32925 <= not w32919 and not w32924;
w32926 <= not w32921 and w32925;
w32927 <= pi0788 and not w32926;
w32928 <= not w17927 and not w32927;
w32929 <= not w32916 and w32928;
w32930 <= not w18133 and w32575;
w32931 <= pi1156 and w32601;
w32932 <= not w32608 and not w32930;
w32933 <= not w32931 and w32932;
w32934 <= pi0792 and not w32933;
w32935 <= not w32929 and not w32934;
w32936 <= not pi0207 and not w32935;
w32937 <= pi0623 and not w32858;
w32938 <= not w32936 and w32937;
w32939 <= pi0710 and not w32938;
w32940 <= not w32769 and w32939;
w32941 <= not w17769 and not w32597;
w32942 <= not w32940 and w32941;
w32943 <= not w32596 and not w32942;
w32944 <= pi0644 and w32943;
w32945 <= pi0715 and not w32531;
w32946 <= not w32944 and w32945;
w32947 <= w15367 and not w32516;
w32948 <= not w15367 and w32591;
w32949 <= not w32947 and not w32948;
w32950 <= pi0644 and w32949;
w32951 <= not pi0644 and w32516;
w32952 <= not pi0715 and not w32951;
w32953 <= not w32950 and w32952;
w32954 <= pi1160 and not w32953;
w32955 <= not w32946 and w32954;
w32956 <= pi0644 and w32530;
w32957 <= not pi0644 and w32943;
w32958 <= not pi0715 and not w32956;
w32959 <= not w32957 and w32958;
w32960 <= not pi0644 and w32949;
w32961 <= pi0644 and w32516;
w32962 <= pi0715 and not w32961;
w32963 <= not w32960 and w32962;
w32964 <= not pi1160 and not w32963;
w32965 <= not w32959 and w32964;
w32966 <= not w32955 and not w32965;
w32967 <= pi0790 and not w32966;
w32968 <= not pi0790 and w32943;
w32969 <= not w32967 and not w32968;
w32970 <= w4989 and not w32969;
w32971 <= not pi0207 and not w4989;
w32972 <= not w32970 and not w32971;
w32973 <= pi0208 and not w32483;
w32974 <= not pi0208 and not w32512;
w32975 <= not w32973 and not w32974;
w32976 <= pi0638 and not w32975;
w32977 <= not pi0208 and not w14622;
w32978 <= not pi0638 and not w32977;
w32979 <= not w32976 and not w32978;
w32980 <= not pi0787 and not w32979;
w32981 <= not pi0647 and w32979;
w32982 <= pi0647 and w32977;
w32983 <= not pi1157 and not w32982;
w32984 <= not w32981 and w32983;
w32985 <= not pi0647 and w32977;
w32986 <= pi0647 and w32979;
w32987 <= pi1157 and not w32985;
w32988 <= not w32986 and w32987;
w32989 <= not w32984 and not w32988;
w32990 <= pi0787 and not w32989;
w32991 <= not w32980 and not w32990;
w32992 <= not pi0644 and w32991;
w32993 <= not pi0630 and w32988;
w32994 <= not pi0208 and not w32578;
w32995 <= pi0208 and not w32586;
w32996 <= pi0607 and not w32995;
w32997 <= not w32994 and w32996;
w32998 <= not pi0607 and w32977;
w32999 <= not w32997 and not w32998;
w33000 <= not w18122 and w32999;
w33001 <= pi0630 and w32984;
w33002 <= not w32993 and not w33000;
w33003 <= not w33001 and w33002;
w33004 <= pi0787 and not w33003;
w33005 <= not pi0638 and not w32999;
w33006 <= not pi0208 and not w32700;
w33007 <= pi0208 and not w32766;
w33008 <= not pi0607 and not w33007;
w33009 <= not w33006 and w33008;
w33010 <= pi0208 and not w32857;
w33011 <= not pi0208 and not w32935;
w33012 <= pi0607 and not w33010;
w33013 <= not w33011 and w33012;
w33014 <= pi0638 and not w33013;
w33015 <= not w33009 and w33014;
w33016 <= not w17769 and not w33005;
w33017 <= not w33015 and w33016;
w33018 <= not w33004 and not w33017;
w33019 <= pi0644 and w33018;
w33020 <= pi0715 and not w32992;
w33021 <= not w33019 and w33020;
w33022 <= w15367 and not w32977;
w33023 <= not w15367 and w32999;
w33024 <= not w33022 and not w33023;
w33025 <= pi0644 and w33024;
w33026 <= not pi0644 and w32977;
w33027 <= not pi0715 and not w33026;
w33028 <= not w33025 and w33027;
w33029 <= pi1160 and not w33028;
w33030 <= not w33021 and w33029;
w33031 <= pi0644 and w32991;
w33032 <= not pi0644 and w33018;
w33033 <= not pi0715 and not w33031;
w33034 <= not w33032 and w33033;
w33035 <= not pi0644 and w33024;
w33036 <= pi0644 and w32977;
w33037 <= pi0715 and not w33036;
w33038 <= not w33035 and w33037;
w33039 <= not pi1160 and not w33038;
w33040 <= not w33034 and w33039;
w33041 <= not w33030 and not w33040;
w33042 <= pi0790 and not w33041;
w33043 <= not pi0790 and w33018;
w33044 <= not w33042 and not w33043;
w33045 <= w4989 and not w33044;
w33046 <= not pi0208 and not w4989;
w33047 <= not w33045 and not w33046;
w33048 <= w7760 and w14615;
w33049 <= not pi0639 and w33048;
w33050 <= pi0715 and w14622;
w33051 <= not w17769 and not w32700;
w33052 <= not pi0647 and not w14622;
w33053 <= pi0647 and w32512;
w33054 <= not w33052 and not w33053;
w33055 <= not pi0630 and not w33054;
w33056 <= not w33052 and not w33055;
w33057 <= pi1157 and not w33056;
w33058 <= pi0647 and not w14622;
w33059 <= not pi1157 and w33058;
w33060 <= not pi0647 and w32512;
w33061 <= not w33058 and not w33060;
w33062 <= w15365 and not w33061;
w33063 <= not w33059 and not w33062;
w33064 <= not w33057 and w33063;
w33065 <= pi0787 and not w33064;
w33066 <= not w33051 and not w33065;
w33067 <= not pi0644 and not w33066;
w33068 <= not w16905 and w32512;
w33069 <= not w14622 and w16905;
w33070 <= not w33068 and not w33069;
w33071 <= pi0644 and not w33070;
w33072 <= not pi0715 and not w33071;
w33073 <= not w33067 and w33072;
w33074 <= not pi1160 and not w33050;
w33075 <= not w33073 and w33074;
w33076 <= not pi0715 and w14622;
w33077 <= pi0644 and not w33066;
w33078 <= not pi0644 and not w33070;
w33079 <= pi0715 and not w33078;
w33080 <= not w33077 and w33079;
w33081 <= pi1160 and not w33076;
w33082 <= not w33080 and w33081;
w33083 <= not w33075 and not w33082;
w33084 <= pi0790 and not w33083;
w33085 <= not pi0790 and not w33066;
w33086 <= w4989 and not w33085;
w33087 <= not w33084 and w33086;
w33088 <= pi0639 and w33087;
w33089 <= not pi0622 and not w33049;
w33090 <= not w33088 and w33089;
w33091 <= not w14622 and w15367;
w33092 <= not w15367 and w32578;
w33093 <= not w33091 and not w33092;
w33094 <= not pi0790 and not w33093;
w33095 <= pi0644 and not w33093;
w33096 <= not pi0644 and not w14622;
w33097 <= not w33095 and not w33096;
w33098 <= pi1160 and w33097;
w33099 <= not pi0644 and not w33093;
w33100 <= pi0644 and not w14622;
w33101 <= not w33099 and not w33100;
w33102 <= not pi1160 and w33101;
w33103 <= pi0790 and not w33098;
w33104 <= not w33102 and w33103;
w33105 <= w4989 and not w33094;
w33106 <= not w33104 and w33105;
w33107 <= not pi0639 and w33106;
w33108 <= pi0715 and w33101;
w33109 <= not w17769 and not w32935;
w33110 <= not w18122 and w32578;
w33111 <= pi1157 and w33055;
w33112 <= not w33062 and not w33110;
w33113 <= not w33111 and w33112;
w33114 <= pi0787 and not w33113;
w33115 <= not w33109 and not w33114;
w33116 <= not pi0644 and not w33115;
w33117 <= w33072 and not w33116;
w33118 <= not pi1160 and not w33108;
w33119 <= not w33117 and w33118;
w33120 <= not pi0715 and w33097;
w33121 <= pi0644 and not w33115;
w33122 <= w33079 and not w33121;
w33123 <= pi1160 and not w33120;
w33124 <= not w33122 and w33123;
w33125 <= not w33119 and not w33124;
w33126 <= pi0790 and not w33125;
w33127 <= not pi0790 and not w33115;
w33128 <= w4989 and not w33127;
w33129 <= not w33126 and w33128;
w33130 <= pi0639 and w33129;
w33131 <= pi0622 and not w33107;
w33132 <= not w33130 and w33131;
w33133 <= not w33090 and not w33132;
w33134 <= not pi0209 and not w33133;
w33135 <= not pi0644 and pi1160;
w33136 <= pi0644 and not pi1160;
w33137 <= not w33135 and not w33136;
w33138 <= pi0790 and not w33137;
w33139 <= w21247 and w32585;
w33140 <= w4989 and not w33138;
w33141 <= w33139 and w33140;
w33142 <= pi0622 and w33141;
w33143 <= not pi0639 and not w33142;
w33144 <= not w17769 and not w32766;
w33145 <= w15367 and w16904;
w33146 <= w32483 and w33145;
w33147 <= not w33144 and not w33146;
w33148 <= not pi0790 and w33147;
w33149 <= not w16905 and w32483;
w33150 <= not pi0644 and not w33149;
w33151 <= pi0715 and not w33150;
w33152 <= pi0644 and w33147;
w33153 <= pi1160 and w33151;
w33154 <= not w33152 and w33153;
w33155 <= pi0644 and not w33149;
w33156 <= not pi0715 and not w33155;
w33157 <= not pi0644 and w33147;
w33158 <= not pi1160 and w33156;
w33159 <= not w33157 and w33158;
w33160 <= pi0790 and not w33154;
w33161 <= not w33159 and w33160;
w33162 <= w4989 and not w33148;
w33163 <= not w33161 and w33162;
w33164 <= not pi0622 and not w33163;
w33165 <= not pi0644 and pi0715;
w33166 <= w33139 and w33165;
w33167 <= pi0647 and w32483;
w33168 <= pi1157 and not w33167;
w33169 <= pi0647 and w32586;
w33170 <= not pi0647 and not w32857;
w33171 <= not pi1157 and not w33169;
w33172 <= not w33170 and w33171;
w33173 <= not pi0630 and not w33168;
w33174 <= not w33172 and w33173;
w33175 <= not pi0647 and w32483;
w33176 <= not pi1157 and not w33175;
w33177 <= not pi0647 and w32586;
w33178 <= pi0647 and not w32857;
w33179 <= pi1157 and not w33177;
w33180 <= not w33178 and w33179;
w33181 <= pi0630 and not w33176;
w33182 <= not w33180 and w33181;
w33183 <= not w33174 and not w33182;
w33184 <= pi0787 and not w33183;
w33185 <= not pi0787 and not w32857;
w33186 <= not w33184 and not w33185;
w33187 <= not pi0644 and w33186;
w33188 <= w33156 and not w33187;
w33189 <= not pi1160 and not w33166;
w33190 <= not w33188 and w33189;
w33191 <= pi0644 and not pi0715;
w33192 <= w33139 and w33191;
w33193 <= pi0644 and w33186;
w33194 <= w33151 and not w33193;
w33195 <= pi1160 and not w33192;
w33196 <= not w33194 and w33195;
w33197 <= not w33190 and not w33196;
w33198 <= pi0790 and not w33197;
w33199 <= not pi0790 and w33186;
w33200 <= w4989 and not w33199;
w33201 <= not w33198 and w33200;
w33202 <= pi0622 and pi0639;
w33203 <= not w33201 and w33202;
w33204 <= pi0209 and not w33143;
w33205 <= not w33164 and w33204;
w33206 <= not w33203 and w33205;
w33207 <= not w33134 and not w33206;
w33208 <= pi0210 and not w14204;
w33209 <= pi0634 and w18465;
w33210 <= pi0633 and pi0947;
w33211 <= not w33209 and not w33210;
w33212 <= w14204 and not w33211;
w33213 <= pi0038 and not w33208;
w33214 <= not w33212 and w33213;
w33215 <= not w14502 and not w33211;
w33216 <= pi0299 and not w33215;
w33217 <= not w14503 and w33216;
w33218 <= pi0210 and not w14493;
w33219 <= w14493 and not w33211;
w33220 <= not pi0299 and not w33218;
w33221 <= not w33219 and w33220;
w33222 <= not pi0039 and not w33217;
w33223 <= not w33221 and w33222;
w33224 <= pi0210 and not w14216;
w33225 <= not w31152 and not w33224;
w33226 <= w3790 and w33225;
w33227 <= pi0947 and not w33226;
w33228 <= pi0210 and w14284;
w33229 <= pi0633 and not w14284;
w33230 <= not w33228 and not w33229;
w33231 <= not w3790 and w33230;
w33232 <= w33227 and not w33231;
w33233 <= pi0634 and w14216;
w33234 <= not w33224 and not w33233;
w33235 <= w3790 and w33234;
w33236 <= pi0907 and not w33235;
w33237 <= not w30993 and not w33228;
w33238 <= not w3790 and w33237;
w33239 <= w33236 and not w33238;
w33240 <= w3790 and w14215;
w33241 <= w489 and w33240;
w33242 <= w33228 and not w33241;
w33243 <= not w33239 and not w33242;
w33244 <= not pi0947 and not w33243;
w33245 <= not w3768 and not w33232;
w33246 <= not w33244 and w33245;
w33247 <= w3759 and w33225;
w33248 <= pi0947 and not w33247;
w33249 <= not w3760 and not w33230;
w33250 <= not w3759 and w33225;
w33251 <= not w3761 and not w33250;
w33252 <= not w33249 and not w33251;
w33253 <= w33248 and not w33252;
w33254 <= not w3761 and not w33234;
w33255 <= pi0907 and not w33254;
w33256 <= w3761 and not w33237;
w33257 <= w33255 and not w33256;
w33258 <= w3759 and w33224;
w33259 <= pi0210 and not w3759;
w33260 <= not w14360 and w33259;
w33261 <= not w33258 and not w33260;
w33262 <= not pi0907 and w33261;
w33263 <= not pi0947 and not w33257;
w33264 <= not w33262 and w33263;
w33265 <= w3768 and not w33253;
w33266 <= not w33264 and w33265;
w33267 <= pi0223 and not w33246;
w33268 <= not w33266 and w33267;
w33269 <= w14216 and not w33211;
w33270 <= not w33224 and not w33269;
w33271 <= w166 and w33270;
w33272 <= pi0210 and w14244;
w33273 <= pi0633 and not w14244;
w33274 <= not w33272 and not w33273;
w33275 <= not w3760 and not w33274;
w33276 <= not w33251 and not w33275;
w33277 <= w33248 and not w33276;
w33278 <= pi0634 and not w14244;
w33279 <= not w33272 and not w33278;
w33280 <= w3761 and not w33279;
w33281 <= w33255 and not w33280;
w33282 <= not w14247 and w33259;
w33283 <= not w33258 and not w33282;
w33284 <= not pi0907 and w33283;
w33285 <= not pi0947 and not w33281;
w33286 <= not w33284 and w33285;
w33287 <= w3768 and not w33277;
w33288 <= not w33286 and w33287;
w33289 <= not w3790 and w33279;
w33290 <= w33236 and not w33289;
w33291 <= pi0210 and not w14706;
w33292 <= not pi0907 and w33291;
w33293 <= not w33290 and not w33292;
w33294 <= not pi0947 and not w33293;
w33295 <= not w3790 and w33274;
w33296 <= w33227 and not w33295;
w33297 <= not w3768 and not w33296;
w33298 <= not w33294 and w33297;
w33299 <= not w33288 and not w33298;
w33300 <= not w166 and not w33299;
w33301 <= not pi0223 and not w33271;
w33302 <= not w33300 and w33301;
w33303 <= not pi0299 and not w33268;
w33304 <= not w33302 and w33303;
w33305 <= not w3804 and not w33242;
w33306 <= w3804 and w33261;
w33307 <= not pi0907 and not w33305;
w33308 <= not w33306 and w33307;
w33309 <= not w33239 and not w33308;
w33310 <= not pi0947 and not w33309;
w33311 <= not w33232 and not w33310;
w33312 <= pi0215 and not w33311;
w33313 <= w1011 and w33270;
w33314 <= not w3804 and not w33291;
w33315 <= w3804 and w33283;
w33316 <= not pi0907 and not w33315;
w33317 <= not w33314 and w33316;
w33318 <= not w33290 and not w33317;
w33319 <= not pi0947 and not w33318;
w33320 <= not w1011 and not w33296;
w33321 <= not w33319 and w33320;
w33322 <= not pi0215 and not w33313;
w33323 <= not w33321 and w33322;
w33324 <= pi0299 and not w33312;
w33325 <= not w33323 and w33324;
w33326 <= pi0039 and not w33325;
w33327 <= not w33304 and w33326;
w33328 <= not pi0038 and not w33223;
w33329 <= not w33327 and w33328;
w33330 <= not w33214 and not w33329;
w33331 <= w7760 and not w33330;
w33332 <= not pi0210 and not w7760;
w33333 <= not w33331 and not w33332;
w33334 <= w134 and not w19204;
w33335 <= not pi0606 and w33334;
w33336 <= w134 and not w19200;
w33337 <= pi0606 and w33336;
w33338 <= pi0643 and not w33335;
w33339 <= not w33337 and w33338;
w33340 <= not pi0606 and w14622;
w33341 <= w134 and not w18573;
w33342 <= pi0606 and w33341;
w33343 <= not pi0643 and not w33340;
w33344 <= not w33342 and w33343;
w33345 <= w4989 and not w33344;
w33346 <= not w33339 and w33345;
w33347 <= pi0211 and not w33346;
w33348 <= w134 and w19191;
w33349 <= not pi0606 and not w33348;
w33350 <= w134 and w19188;
w33351 <= pi0606 and not w33350;
w33352 <= pi0643 and not w33349;
w33353 <= not w33351 and w33352;
w33354 <= w134 and w18597;
w33355 <= pi0606 and not pi0643;
w33356 <= w33354 and w33355;
w33357 <= not w33353 and not w33356;
w33358 <= not pi0211 and w4989;
w33359 <= not w33357 and w33358;
w33360 <= not w33347 and not w33359;
w33361 <= not pi0607 and w33334;
w33362 <= pi0607 and w33336;
w33363 <= pi0638 and not w33361;
w33364 <= not w33362 and w33363;
w33365 <= not pi0607 and w14622;
w33366 <= pi0607 and w33341;
w33367 <= not pi0638 and not w33365;
w33368 <= not w33366 and w33367;
w33369 <= w4989 and not w33368;
w33370 <= not w33364 and w33369;
w33371 <= not pi0212 and not w33370;
w33372 <= pi0607 and not w33350;
w33373 <= not pi0607 and not w33348;
w33374 <= pi0638 and not w33372;
w33375 <= not w33373 and w33374;
w33376 <= pi0607 and not pi0638;
w33377 <= w33354 and w33376;
w33378 <= not w33375 and not w33377;
w33379 <= pi0212 and w4989;
w33380 <= not w33378 and w33379;
w33381 <= not w33371 and not w33380;
w33382 <= pi0213 and w4989;
w33383 <= pi0622 and not w33350;
w33384 <= not pi0622 and not w33348;
w33385 <= pi0639 and not w33383;
w33386 <= not w33384 and w33385;
w33387 <= pi0622 and not pi0639;
w33388 <= w33354 and w33387;
w33389 <= not w33386 and not w33388;
w33390 <= w33382 and not w33389;
w33391 <= not pi0639 and w33341;
w33392 <= pi0639 and w33336;
w33393 <= pi0622 and not w33391;
w33394 <= not w33392 and w33393;
w33395 <= not pi0639 and w14622;
w33396 <= pi0639 and w33334;
w33397 <= not pi0622 and not w33395;
w33398 <= not w33396 and w33397;
w33399 <= w4989 and not w33398;
w33400 <= not w33394 and w33399;
w33401 <= not pi0213 and not w33400;
w33402 <= not w33390 and not w33401;
w33403 <= not pi0623 and w33334;
w33404 <= pi0623 and w33336;
w33405 <= pi0710 and not w33403;
w33406 <= not w33404 and w33405;
w33407 <= not pi0623 and w14622;
w33408 <= pi0623 and w33341;
w33409 <= not pi0710 and not w33407;
w33410 <= not w33408 and w33409;
w33411 <= w4989 and not w33410;
w33412 <= not w33406 and w33411;
w33413 <= not pi0214 and not w33412;
w33414 <= pi0623 and not w33350;
w33415 <= not pi0623 and not w33348;
w33416 <= pi0710 and not w33414;
w33417 <= not w33415 and w33416;
w33418 <= pi0623 and not pi0710;
w33419 <= w33354 and w33418;
w33420 <= not w33417 and not w33419;
w33421 <= pi0214 and w4989;
w33422 <= not w33420 and w33421;
w33423 <= not w33413 and not w33422;
w33424 <= pi0215 and not w7760;
w33425 <= pi0681 and pi0907;
w33426 <= not pi0947 and w33425;
w33427 <= pi0642 and pi0947;
w33428 <= not w33426 and not w33427;
w33429 <= w14204 and not w33428;
w33430 <= pi0215 and not w14204;
w33431 <= pi0038 and not w33429;
w33432 <= not w33430 and w33431;
w33433 <= pi0215 and not w14504;
w33434 <= w14504 and not w33428;
w33435 <= pi0299 and not w33433;
w33436 <= not w33434 and w33435;
w33437 <= w14493 and not w33428;
w33438 <= pi0215 and not w14493;
w33439 <= not pi0299 and not w33437;
w33440 <= not w33438 and w33439;
w33441 <= not pi0039 and not w33436;
w33442 <= not w33440 and w33441;
w33443 <= not pi0947 and w18889;
w33444 <= w14219 and w14526;
w33445 <= not w3758 and not w14377;
w33446 <= not pi0642 and not w33444;
w33447 <= not w33445 and w33446;
w33448 <= pi0947 and not w33447;
w33449 <= not w33426 and not w33448;
w33450 <= not w33443 and w33449;
w33451 <= pi0299 and not w33450;
w33452 <= w166 and not w33428;
w33453 <= w166 and not w14216;
w33454 <= w18994 and not w33425;
w33455 <= not pi0642 and w14706;
w33456 <= not w3768 and not w33455;
w33457 <= not pi0642 and w14247;
w33458 <= w3758 and not w33457;
w33459 <= w14332 and w14730;
w33460 <= not w3754 and w14216;
w33461 <= not pi0642 and w33460;
w33462 <= not w3758 and not w33461;
w33463 <= not w33459 and w33462;
w33464 <= not w33458 and not w33463;
w33465 <= w3768 and not w33464;
w33466 <= pi0947 and not w33456;
w33467 <= not w33465 and w33466;
w33468 <= not w166 and not w33467;
w33469 <= not w33454 and w33468;
w33470 <= not pi0223 and not w33452;
w33471 <= not w33453 and w33470;
w33472 <= not w33469 and w33471;
w33473 <= not w3768 and not w33447;
w33474 <= w3758 and not w14360;
w33475 <= not w3758 and not w14366;
w33476 <= not pi0642 and not w33474;
w33477 <= not w33475 and w33476;
w33478 <= w3768 and not w33477;
w33479 <= pi0947 and not w33473;
w33480 <= not w33478 and w33479;
w33481 <= not w18615 and not w33480;
w33482 <= pi0223 and not w33426;
w33483 <= not w33481 and w33482;
w33484 <= not pi0299 and not w33483;
w33485 <= not w33472 and w33484;
w33486 <= not w33451 and not w33485;
w33487 <= pi0215 and not w33486;
w33488 <= w14216 and w33452;
w33489 <= w14265 and w33425;
w33490 <= not pi0947 and not w33489;
w33491 <= pi0642 and w14220;
w33492 <= not w3758 and w14262;
w33493 <= not w14705 and not w33492;
w33494 <= w33491 and w33493;
w33495 <= pi0642 and not w14220;
w33496 <= not w14262 and w33495;
w33497 <= pi0947 and not w33496;
w33498 <= not w33494 and w33497;
w33499 <= not w33490 and not w33498;
w33500 <= not w3768 and not w33499;
w33501 <= w14216 and w33495;
w33502 <= not w14537 and w33491;
w33503 <= not w14558 and w33502;
w33504 <= not w33501 and not w33503;
w33505 <= pi0947 and not w33504;
w33506 <= w14339 and w33426;
w33507 <= w3768 and not w33505;
w33508 <= not w33506 and w33507;
w33509 <= not w166 and not w33500;
w33510 <= not w33508 and w33509;
w33511 <= not pi0223 and not w33488;
w33512 <= not w33510 and w33511;
w33513 <= w3768 and not w14366;
w33514 <= w33425 and not w33513;
w33515 <= not pi0947 and not w33514;
w33516 <= pi0947 and not w14286;
w33517 <= not w14377 and not w33516;
w33518 <= not w3768 and w33517;
w33519 <= not w14536 and w33502;
w33520 <= pi0947 and not w33501;
w33521 <= not w33519 and w33520;
w33522 <= not w33518 and not w33521;
w33523 <= not w33515 and w33522;
w33524 <= pi0223 and not w33523;
w33525 <= not w33512 and not w33524;
w33526 <= not pi0299 and not w33525;
w33527 <= w14589 and not w33428;
w33528 <= not w1011 and w33499;
w33529 <= pi0299 and not w33527;
w33530 <= not w33528 and w33529;
w33531 <= not pi0215 and not w33530;
w33532 <= not w33526 and w33531;
w33533 <= not w33487 and not w33532;
w33534 <= pi0039 and not w33533;
w33535 <= not pi0038 and not w33442;
w33536 <= not w33534 and w33535;
w33537 <= w7760 and not w33432;
w33538 <= not w33536 and w33537;
w33539 <= not w33424 and not w33538;
w33540 <= pi0662 and pi0907;
w33541 <= not pi0947 and w33540;
w33542 <= pi0614 and pi0947;
w33543 <= not w33541 and not w33542;
w33544 <= w14204 and not w33543;
w33545 <= pi0216 and not w14204;
w33546 <= pi0038 and not w33544;
w33547 <= not w33545 and w33546;
w33548 <= pi0216 and not w14504;
w33549 <= w14504 and not w33543;
w33550 <= pi0299 and not w33548;
w33551 <= not w33549 and w33550;
w33552 <= w14493 and not w33543;
w33553 <= pi0216 and not w14493;
w33554 <= not pi0299 and not w33552;
w33555 <= not w33553 and w33554;
w33556 <= not pi0039 and not w33551;
w33557 <= not w33555 and w33556;
w33558 <= not w33513 and w33540;
w33559 <= not pi0947 and not w33558;
w33560 <= not w14536 and w14560;
w33561 <= pi0947 and not w14563;
w33562 <= not w33560 and w33561;
w33563 <= not w33518 and not w33562;
w33564 <= not w33559 and w33563;
w33565 <= pi0223 and not w33564;
w33566 <= w166 and not w33543;
w33567 <= w14216 and w33566;
w33568 <= w33493 and w33542;
w33569 <= w14265 and w33541;
w33570 <= not w33568 and not w33569;
w33571 <= not w3768 and w33570;
w33572 <= w14339 and w33541;
w33573 <= pi0947 and not w14564;
w33574 <= w3768 and not w33573;
w33575 <= not w33572 and w33574;
w33576 <= not w166 and not w33571;
w33577 <= not w33575 and w33576;
w33578 <= not pi0223 and not w33567;
w33579 <= not w33577 and w33578;
w33580 <= not pi0216 and not w33565;
w33581 <= not w33579 and w33580;
w33582 <= not pi0616 and w14362;
w33583 <= not w3758 and not w14541;
w33584 <= not w33582 and w33583;
w33585 <= not pi0614 and not w33474;
w33586 <= not w33584 and w33585;
w33587 <= w3768 and not w33586;
w33588 <= not w15015 and not w30945;
w33589 <= not w30946 and w33588;
w33590 <= w14565 and not w33589;
w33591 <= not pi0614 and not w14284;
w33592 <= w3758 and w33591;
w33593 <= not w33590 and not w33592;
w33594 <= not w3768 and w33593;
w33595 <= pi0947 and not w33594;
w33596 <= not w33587 and w33595;
w33597 <= not w18615 and not w33596;
w33598 <= pi0223 and not w33541;
w33599 <= not w33597 and w33598;
w33600 <= not pi0614 and w14706;
w33601 <= pi0947 and not w33600;
w33602 <= not pi0947 and not w14581;
w33603 <= not w3768 and not w33541;
w33604 <= not w33601 and w33603;
w33605 <= not w33602 and w33604;
w33606 <= pi0947 and not w14571;
w33607 <= not pi0947 and w14574;
w33608 <= not w33540 and w33607;
w33609 <= not w33606 and not w33608;
w33610 <= w3768 and not w33609;
w33611 <= not w166 and not w33605;
w33612 <= not w33610 and w33611;
w33613 <= not pi0223 and not w33566;
w33614 <= not w33453 and w33613;
w33615 <= not w33612 and w33614;
w33616 <= pi0216 and not w33599;
w33617 <= not w33615 and w33616;
w33618 <= not pi0299 and not w33581;
w33619 <= not w33617 and w33618;
w33620 <= w3340 and not w33570;
w33621 <= w14589 and not w33543;
w33622 <= not pi0947 and w18557;
w33623 <= not w33541 and not w33601;
w33624 <= not w33622 and w33623;
w33625 <= pi0216 and not w33624;
w33626 <= not w33620 and not w33621;
w33627 <= not w33625 and w33626;
w33628 <= not pi0215 and not w33627;
w33629 <= w14377 and w33540;
w33630 <= not pi0947 and not w33629;
w33631 <= pi0947 and w14286;
w33632 <= not w33562 and not w33631;
w33633 <= not w33630 and w33632;
w33634 <= not pi0216 and not w33633;
w33635 <= pi0947 and w33593;
w33636 <= pi0216 and not w33541;
w33637 <= not w33635 and w33636;
w33638 <= not w33443 and w33637;
w33639 <= pi0215 and not w33634;
w33640 <= not w33638 and w33639;
w33641 <= pi0299 and not w33640;
w33642 <= not w33628 and w33641;
w33643 <= pi0039 and not w33619;
w33644 <= not w33642 and w33643;
w33645 <= not pi0038 and not w33557;
w33646 <= not w33644 and w33645;
w33647 <= not w33547 and not w33646;
w33648 <= w7760 and not w33647;
w33649 <= not pi0216 and not w7760;
w33650 <= not w33648 and not w33649;
w33651 <= not pi0695 and w33163;
w33652 <= pi0217 and not w33651;
w33653 <= pi0695 and not w33048;
w33654 <= not pi0695 and not w33087;
w33655 <= not pi0217 and not w33653;
w33656 <= not w33654 and w33655;
w33657 <= not pi0612 and not w33652;
w33658 <= not w33656 and w33657;
w33659 <= not pi0695 and w33201;
w33660 <= pi0695 and w33141;
w33661 <= pi0217 and not w33660;
w33662 <= not w33659 and w33661;
w33663 <= pi0695 and not w33106;
w33664 <= not pi0695 and not w33129;
w33665 <= not pi0217 and not w33663;
w33666 <= not w33664 and w33665;
w33667 <= pi0612 and not w33662;
w33668 <= not w33666 and w33667;
w33669 <= not w33658 and not w33668;
w33670 <= not w32349 and not w32388;
w33671 <= w32349 and not w32454;
w33672 <= not w33670 and not w33671;
w33673 <= not pi0218 and not w33672;
w33674 <= w32349 and w32462;
w33675 <= pi0218 and not w33674;
w33676 <= not w33673 and not w33675;
w33677 <= not pi0219 and w4989;
w33678 <= pi0617 and not w33350;
w33679 <= not pi0617 and not w33348;
w33680 <= pi0637 and not w33678;
w33681 <= not w33679 and w33680;
w33682 <= pi0617 and not pi0637;
w33683 <= w33354 and w33682;
w33684 <= not w33681 and not w33683;
w33685 <= w33677 and not w33684;
w33686 <= not pi0617 and w33334;
w33687 <= pi0617 and w33336;
w33688 <= pi0637 and not w33686;
w33689 <= not w33687 and w33688;
w33690 <= not pi0617 and w14622;
w33691 <= pi0617 and w33341;
w33692 <= not pi0637 and not w33690;
w33693 <= not w33691 and w33692;
w33694 <= w4989 and not w33693;
w33695 <= not w33689 and w33694;
w33696 <= pi0219 and not w33695;
w33697 <= not w33685 and not w33696;
w33698 <= not w32182 and not w32473;
w33699 <= not w32328 and w32473;
w33700 <= not w33698 and not w33699;
w33701 <= not pi0220 and not w33700;
w33702 <= w32337 and w32473;
w33703 <= pi0220 and not w33702;
w33704 <= not w33701 and not w33703;
w33705 <= pi0661 and pi0907;
w33706 <= not pi0947 and w33705;
w33707 <= pi0616 and pi0947;
w33708 <= not w33706 and not w33707;
w33709 <= w14204 and not w33708;
w33710 <= pi0221 and not w14204;
w33711 <= pi0038 and not w33709;
w33712 <= not w33710 and w33711;
w33713 <= pi0221 and not w14504;
w33714 <= w14504 and not w33708;
w33715 <= pi0299 and not w33713;
w33716 <= not w33714 and w33715;
w33717 <= w14493 and not w33708;
w33718 <= pi0221 and not w14493;
w33719 <= not pi0299 and not w33717;
w33720 <= not w33718 and w33719;
w33721 <= not pi0039 and not w33716;
w33722 <= not w33720 and w33721;
w33723 <= pi0947 and not w14543;
w33724 <= not w33706 and not w33723;
w33725 <= w33513 and not w33723;
w33726 <= not w33518 and not w33724;
w33727 <= not w33725 and w33726;
w33728 <= pi0223 and not w33727;
w33729 <= w14216 and not w33708;
w33730 <= w166 and w33729;
w33731 <= not pi0223 and not w33730;
w33732 <= w14539 and not w14558;
w33733 <= not w14542 and not w33732;
w33734 <= pi0947 and not w33733;
w33735 <= w14339 and w33706;
w33736 <= w3768 and not w33734;
w33737 <= not w33735 and w33736;
w33738 <= w33493 and w33707;
w33739 <= w14265 and w33706;
w33740 <= not w33738 and not w33739;
w33741 <= not w3768 and w33740;
w33742 <= not w166 and not w33741;
w33743 <= not w33737 and w33742;
w33744 <= w33731 and not w33743;
w33745 <= not pi0221 and not w33728;
w33746 <= not w33744 and w33745;
w33747 <= not w33455 and not w33494;
w33748 <= w14547 and not w33747;
w33749 <= not w3760 and w14337;
w33750 <= not w14260 and not w33749;
w33751 <= w14544 and not w33750;
w33752 <= pi0947 and not w33748;
w33753 <= not w33751 and w33752;
w33754 <= not w33602 and not w33753;
w33755 <= not w3768 and not w33754;
w33756 <= w14337 and w14544;
w33757 <= not w14561 and w14571;
w33758 <= w14547 and not w33757;
w33759 <= not w33756 and not w33758;
w33760 <= pi0947 and not w33759;
w33761 <= w3768 and not w33607;
w33762 <= not w33760 and w33761;
w33763 <= not w33706 and not w33755;
w33764 <= not w33762 and w33763;
w33765 <= not w166 and not w33764;
w33766 <= not w33453 and w33731;
w33767 <= not w33765 and w33766;
w33768 <= not pi0947 and w14553;
w33769 <= pi0947 and not w14550;
w33770 <= w3768 and not w33769;
w33771 <= not w33768 and w33770;
w33772 <= not pi0947 and not w14533;
w33773 <= not w14286 and not w14363;
w33774 <= not w3758 and not w33773;
w33775 <= not pi0616 and not w33444;
w33776 <= not w33774 and w33775;
w33777 <= pi0947 and not w33776;
w33778 <= not w33772 and not w33777;
w33779 <= not w3768 and not w33778;
w33780 <= pi0223 and not w33706;
w33781 <= not w33771 and w33780;
w33782 <= not w33779 and w33781;
w33783 <= pi0221 and not w33782;
w33784 <= not w33767 and w33783;
w33785 <= not pi0299 and not w33746;
w33786 <= not w33784 and w33785;
w33787 <= not w18557 and not w33705;
w33788 <= not pi0947 and not w33787;
w33789 <= pi0221 and not w33753;
w33790 <= not w33788 and w33789;
w33791 <= pi0216 and not w33740;
w33792 <= not pi0216 and w33729;
w33793 <= not pi0221 and not w33792;
w33794 <= not w33791 and w33793;
w33795 <= not pi0215 and not w33794;
w33796 <= not w33790 and w33795;
w33797 <= pi0221 and not w33706;
w33798 <= not w33777 and w33797;
w33799 <= not w33443 and w33798;
w33800 <= not w33517 and not w33724;
w33801 <= not pi0221 and not w33800;
w33802 <= pi0215 and not w33801;
w33803 <= not w33799 and w33802;
w33804 <= pi0299 and not w33803;
w33805 <= not w33796 and w33804;
w33806 <= pi0039 and not w33786;
w33807 <= not w33805 and w33806;
w33808 <= not pi0038 and not w33722;
w33809 <= not w33807 and w33808;
w33810 <= not w33712 and not w33809;
w33811 <= w7760 and not w33810;
w33812 <= not pi0221 and not w7760;
w33813 <= not w33811 and not w33812;
w33814 <= not pi0223 and not w14583;
w33815 <= not w14556 and not w33814;
w33816 <= not pi0299 and not w33815;
w33817 <= pi0039 and not w33816;
w33818 <= not w14608 and w33817;
w33819 <= not pi0038 and not w15710;
w33820 <= not w33818 and w33819;
w33821 <= w16154 and not w33820;
w33822 <= pi0222 and not w33821;
w33823 <= not w16712 and not w33822;
w33824 <= pi0222 and not w134;
w33825 <= pi0222 and not w14204;
w33826 <= pi0038 and not w33825;
w33827 <= pi0661 and w14209;
w33828 <= w33826 and not w33827;
w33829 <= pi0661 and pi0680;
w33830 <= w14481 and not w33829;
w33831 <= not pi0222 and not w14481;
w33832 <= pi0222 and w14498;
w33833 <= not pi0299 and not w33832;
w33834 <= not w33830 and w33833;
w33835 <= not w33831 and w33834;
w33836 <= pi0222 and w14507;
w33837 <= w14486 and not w33829;
w33838 <= not pi0222 and not w14486;
w33839 <= pi0299 and not w33836;
w33840 <= not w33837 and w33839;
w33841 <= not w33838 and w33840;
w33842 <= not pi0039 and not w33835;
w33843 <= not w33841 and w33842;
w33844 <= not pi0661 and not w14581;
w33845 <= pi0680 and w14321;
w33846 <= not w14316 and not w33845;
w33847 <= pi0661 and not w33846;
w33848 <= not w33844 and not w33847;
w33849 <= not w3768 and w33848;
w33850 <= not pi0661 and w14557;
w33851 <= not w3756 and not w14339;
w33852 <= not pi0662 and w14558;
w33853 <= not w33851 and not w33852;
w33854 <= w14219 and not w33853;
w33855 <= pi0661 and not w14349;
w33856 <= not w33850 and not w33854;
w33857 <= not w33855 and w33856;
w33858 <= w3768 and w33857;
w33859 <= pi0222 and not w33849;
w33860 <= not w33858 and w33859;
w33861 <= not w14253 and w33829;
w33862 <= w3768 and w33861;
w33863 <= pi0661 and w14266;
w33864 <= not w3768 and w33863;
w33865 <= pi0224 and not w33862;
w33866 <= not w33864 and w33865;
w33867 <= pi0661 and w14302;
w33868 <= not pi0224 and not w33867;
w33869 <= not pi0222 and not w33868;
w33870 <= not w33866 and w33869;
w33871 <= not pi0223 and not w33870;
w33872 <= not w33860 and w33871;
w33873 <= not pi0222 and pi0661;
w33874 <= w14292 and w33873;
w33875 <= not pi0661 and w14523;
w33876 <= w14219 and w14529;
w33877 <= pi0661 and not w14381;
w33878 <= not w33875 and not w33877;
w33879 <= not w33876 and w33878;
w33880 <= not w3768 and w33879;
w33881 <= not pi0661 and not w14553;
w33882 <= not w14367 and not w14372;
w33883 <= pi0661 and not w33882;
w33884 <= not w33881 and not w33883;
w33885 <= w3768 and w33884;
w33886 <= pi0222 and not w33880;
w33887 <= not w33885 and w33886;
w33888 <= pi0223 and not w33874;
w33889 <= not w33887 and w33888;
w33890 <= not w33872 and not w33889;
w33891 <= not pi0299 and not w33890;
w33892 <= w14307 and w33873;
w33893 <= not w3805 and w33879;
w33894 <= w3805 and w33884;
w33895 <= pi0222 and not w33893;
w33896 <= not w33894 and w33895;
w33897 <= not w33892 and not w33896;
w33898 <= pi0215 and not w33897;
w33899 <= pi0222 and not w14216;
w33900 <= w1011 and not w33899;
w33901 <= not w33867 and w33900;
w33902 <= not w3805 and w33848;
w33903 <= w3805 and w33857;
w33904 <= pi0222 and not w33902;
w33905 <= not w33903 and w33904;
w33906 <= not w3805 and not w33863;
w33907 <= w3805 and not w33861;
w33908 <= not pi0222 and not w33906;
w33909 <= not w33907 and w33908;
w33910 <= not w1011 and not w33909;
w33911 <= not w33905 and w33910;
w33912 <= not pi0215 and not w33901;
w33913 <= not w33911 and w33912;
w33914 <= pi0299 and not w33898;
w33915 <= not w33913 and w33914;
w33916 <= not w33891 and not w33915;
w33917 <= pi0039 and not w33916;
w33918 <= not w33843 and not w33917;
w33919 <= not pi0038 and not w33918;
w33920 <= w134 and not w33828;
w33921 <= not w33919 and w33920;
w33922 <= not w33824 and not w33921;
w33923 <= not pi0778 and not w33922;
w33924 <= pi0625 and w33922;
w33925 <= not pi0625 and not w33822;
w33926 <= pi1153 and not w33925;
w33927 <= not w33924 and w33926;
w33928 <= not pi0625 and w33922;
w33929 <= pi0625 and not w33822;
w33930 <= not pi1153 and not w33929;
w33931 <= not w33928 and w33930;
w33932 <= not w33927 and not w33931;
w33933 <= pi0778 and not w33932;
w33934 <= not w33923 and not w33933;
w33935 <= not w14638 and not w33934;
w33936 <= w14638 and w33822;
w33937 <= not w33935 and not w33936;
w33938 <= not w14202 and not w33937;
w33939 <= w14202 and w33822;
w33940 <= not w33938 and not w33939;
w33941 <= not w14198 and w33940;
w33942 <= not w14194 and w33941;
w33943 <= not w33823 and not w33942;
w33944 <= not w16705 and not w33943;
w33945 <= w15419 and not w33822;
w33946 <= not w33944 and not w33945;
w33947 <= not pi0787 and w33946;
w33948 <= not pi0647 and not w33946;
w33949 <= pi0647 and not w33822;
w33950 <= not pi1157 and not w33949;
w33951 <= not w33948 and w33950;
w33952 <= pi0647 and not w33946;
w33953 <= not pi0647 and not w33822;
w33954 <= pi1157 and not w33953;
w33955 <= not w33952 and w33954;
w33956 <= not w33951 and not w33955;
w33957 <= pi0787 and not w33956;
w33958 <= not w33947 and not w33957;
w33959 <= not pi0644 and w33958;
w33960 <= pi0628 and not w33822;
w33961 <= not pi0628 and not w33943;
w33962 <= w15340 and not w33960;
w33963 <= not w33961 and w33962;
w33964 <= w15532 and not w33822;
w33965 <= pi0616 and w14843;
w33966 <= w33826 and not w33965;
w33967 <= not pi0616 and w14796;
w33968 <= not pi0222 and not w14796;
w33969 <= pi0222 and w14702;
w33970 <= not pi0039 and not w33967;
w33971 <= not w33968 and w33970;
w33972 <= not w33969 and w33971;
w33973 <= not w3758 and w14798;
w33974 <= not w14799 and not w33973;
w33975 <= pi0616 and not w33974;
w33976 <= not pi0222 and w33975;
w33977 <= not w14306 and w33976;
w33978 <= pi0616 and not w14745;
w33979 <= w14377 and not w33978;
w33980 <= not w14219 and not w33979;
w33981 <= not w3756 and not w14377;
w33982 <= not w14526 and not w33978;
w33983 <= not w33981 and w33982;
w33984 <= w14219 and not w33983;
w33985 <= not w33980 and not w33984;
w33986 <= not w3805 and w33985;
w33987 <= pi0616 and not w14732;
w33988 <= not w14365 and not w33987;
w33989 <= not w14219 and not w33988;
w33990 <= pi0616 and w14731;
w33991 <= w3756 and not w33990;
w33992 <= w14360 and w33991;
w33993 <= not w3756 and w33988;
w33994 <= w14219 and not w33992;
w33995 <= not w33993 and w33994;
w33996 <= not w33989 and not w33995;
w33997 <= w3805 and w33996;
w33998 <= pi0222 and not w33986;
w33999 <= not w33997 and w33998;
w34000 <= not w33977 and not w33999;
w34001 <= pi0215 and not w34000;
w34002 <= w14541 and w14731;
w34003 <= w33900 and not w34002;
w34004 <= not w14338 and not w33987;
w34005 <= not w14219 and not w34004;
w34006 <= w14247 and w33991;
w34007 <= not w3756 and w34004;
w34008 <= w14219 and not w34006;
w34009 <= not w34007 and w34008;
w34010 <= not w34005 and not w34009;
w34011 <= w3805 and w34010;
w34012 <= pi0616 and not w14717;
w34013 <= not pi0616 and w33750;
w34014 <= not w34012 and not w34013;
w34015 <= not w14219 and not w34014;
w34016 <= w14710 and not w33990;
w34017 <= not w14708 and not w34016;
w34018 <= w3756 and not w34017;
w34019 <= not w3756 and w34014;
w34020 <= w14219 and not w34018;
w34021 <= not w34019 and w34020;
w34022 <= not w34015 and not w34021;
w34023 <= not w3805 and w34022;
w34024 <= pi0222 and not w34011;
w34025 <= not w34023 and w34024;
w34026 <= not w14810 and not w33973;
w34027 <= pi0616 and not w34026;
w34028 <= w3805 and not w34027;
w34029 <= not w14262 and w33990;
w34030 <= not w14219 and not w34029;
w34031 <= pi0616 and w3756;
w34032 <= w14938 and w34031;
w34033 <= not w3756 and w34029;
w34034 <= w14219 and not w34032;
w34035 <= not w34033 and w34034;
w34036 <= not w34030 and not w34035;
w34037 <= not w3805 and not w34036;
w34038 <= not pi0222 and not w34028;
w34039 <= not w34037 and w34038;
w34040 <= not w1011 and not w34039;
w34041 <= not w34025 and w34040;
w34042 <= not pi0215 and not w34003;
w34043 <= not w34041 and w34042;
w34044 <= pi0299 and not w34001;
w34045 <= not w34043 and w34044;
w34046 <= w3768 and w34027;
w34047 <= not w3768 and w34036;
w34048 <= pi0224 and not w34046;
w34049 <= not w34047 and w34048;
w34050 <= not pi0224 and not w34002;
w34051 <= not pi0222 and not w34050;
w34052 <= not w34049 and w34051;
w34053 <= w3768 and w34010;
w34054 <= not w3768 and w34022;
w34055 <= pi0222 and not w34053;
w34056 <= not w34054 and w34055;
w34057 <= not pi0223 and not w34052;
w34058 <= not w34056 and w34057;
w34059 <= not w14287 and w33976;
w34060 <= not w3768 and w33985;
w34061 <= w3768 and w33996;
w34062 <= pi0222 and not w34060;
w34063 <= not w34061 and w34062;
w34064 <= pi0223 and not w34059;
w34065 <= not w34063 and w34064;
w34066 <= not w34058 and not w34065;
w34067 <= not pi0299 and not w34066;
w34068 <= pi0039 and not w34045;
w34069 <= not w34067 and w34068;
w34070 <= not pi0038 and not w33972;
w34071 <= not w34069 and w34070;
w34072 <= w134 and not w33966;
w34073 <= not w34071 and w34072;
w34074 <= not w33824 and not w34073;
w34075 <= not w14680 and not w34074;
w34076 <= w14680 and w33822;
w34077 <= not w34075 and not w34076;
w34078 <= not pi0785 and not w34077;
w34079 <= pi0609 and w34077;
w34080 <= not pi0609 and not w33822;
w34081 <= pi1155 and not w34080;
w34082 <= not w34079 and w34081;
w34083 <= not pi0609 and w34077;
w34084 <= pi0609 and not w33822;
w34085 <= not pi1155 and not w34084;
w34086 <= not w34083 and w34085;
w34087 <= not w34082 and not w34086;
w34088 <= pi0785 and not w34087;
w34089 <= not w34078 and not w34088;
w34090 <= not pi0781 and not w34089;
w34091 <= pi0618 and w34089;
w34092 <= not pi0618 and not w33822;
w34093 <= pi1154 and not w34092;
w34094 <= not w34091 and w34093;
w34095 <= not pi0618 and w34089;
w34096 <= pi0618 and not w33822;
w34097 <= not pi1154 and not w34096;
w34098 <= not w34095 and w34097;
w34099 <= not w34094 and not w34098;
w34100 <= pi0781 and not w34099;
w34101 <= not w34090 and not w34100;
w34102 <= not pi0789 and not w34101;
w34103 <= pi0619 and w34101;
w34104 <= not pi0619 and not w33822;
w34105 <= pi1159 and not w34104;
w34106 <= not w34103 and w34105;
w34107 <= not pi0619 and w34101;
w34108 <= pi0619 and not w33822;
w34109 <= not pi1159 and not w34108;
w34110 <= not w34107 and w34109;
w34111 <= not w34106 and not w34110;
w34112 <= pi0789 and not w34111;
w34113 <= not w34102 and not w34112;
w34114 <= not w15532 and w34113;
w34115 <= not w33964 and not w34114;
w34116 <= not w18133 and w34115;
w34117 <= not pi0628 and not w33822;
w34118 <= pi0628 and not w33943;
w34119 <= w15339 and not w34117;
w34120 <= not w34118 and w34119;
w34121 <= not w33963 and not w34120;
w34122 <= not w34116 and w34121;
w34123 <= pi0792 and not w34122;
w34124 <= pi0609 and w33934;
w34125 <= w14230 and w15056;
w34126 <= not pi0222 and not pi0616;
w34127 <= not pi0039 and pi0616;
w34128 <= w33829 and w34127;
w34129 <= not w34126 and not w34128;
w34130 <= w34125 and not w34129;
w34131 <= not w33829 and not w33990;
w34132 <= not pi0616 and not w14918;
w34133 <= not w34131 and not w34132;
w34134 <= w14204 and w34133;
w34135 <= not w33825 and not w34134;
w34136 <= not w34130 and not w34135;
w34137 <= pi0038 and not w34136;
w34138 <= not pi0661 and pi0681;
w34139 <= not w33988 and w34138;
w34140 <= not pi0680 and w33988;
w34141 <= pi0616 and not w15067;
w34142 <= pi0680 and not w34141;
w34143 <= not w14910 and w34142;
w34144 <= pi0661 and not w34140;
w34145 <= not w34143 and w34144;
w34146 <= not w33995 and not w34139;
w34147 <= not w34145 and w34146;
w34148 <= w3805 and not w34147;
w34149 <= not w33979 and w34138;
w34150 <= not pi0680 and w33979;
w34151 <= not w14887 and w15056;
w34152 <= pi0616 and not w34151;
w34153 <= pi0680 and not w34152;
w34154 <= w14893 and w34153;
w34155 <= pi0661 and not w34154;
w34156 <= not w34150 and w34155;
w34157 <= not w33984 and not w34149;
w34158 <= not w34156 and w34157;
w34159 <= not w3805 and not w34158;
w34160 <= pi0222 and not w34148;
w34161 <= not w34159 and w34160;
w34162 <= w15007 and w33829;
w34163 <= not w33975 and not w34162;
w34164 <= w3805 and not w34163;
w34165 <= pi0616 and w14800;
w34166 <= not pi0661 and not w34165;
w34167 <= not w14284 and w34002;
w34168 <= w3758 and not w34167;
w34169 <= not pi0680 and w34165;
w34170 <= not w14800 and not w15122;
w34171 <= pi0616 and w34170;
w34172 <= pi0680 and not w34171;
w34173 <= w15021 and w34172;
w34174 <= pi0661 and not w34169;
w34175 <= not w34173 and w34174;
w34176 <= not w34166 and not w34168;
w34177 <= not w34175 and w34176;
w34178 <= not w3805 and w34177;
w34179 <= not pi0222 and not w34164;
w34180 <= not w34178 and w34179;
w34181 <= pi0215 and not w34180;
w34182 <= not w34161 and w34181;
w34183 <= pi0616 and not w15111;
w34184 <= not pi0616 and not w14970;
w34185 <= not w34183 and not w34184;
w34186 <= not w34131 and w34185;
w34187 <= w33900 and not w34186;
w34188 <= not w34014 and w34138;
w34189 <= pi0603 and w14244;
w34190 <= w3760 and w14317;
w34191 <= not w14319 and not w34190;
w34192 <= not pi0603 and w34191;
w34193 <= not w14931 and not w34189;
w34194 <= not w34192 and w34193;
w34195 <= not pi0642 and w34194;
w34196 <= not w15140 and w34191;
w34197 <= pi0642 and not w34196;
w34198 <= w3754 and not w34195;
w34199 <= not w34197 and w34198;
w34200 <= w15015 and w34196;
w34201 <= w15056 and not w34191;
w34202 <= pi0616 and not w34201;
w34203 <= pi0680 and not w34202;
w34204 <= not w34200 and w34203;
w34205 <= not w34199 and w34204;
w34206 <= not pi0680 and w34014;
w34207 <= pi0661 and not w34205;
w34208 <= not w34206 and w34207;
w34209 <= not w34021 and not w34188;
w34210 <= not w34208 and w34209;
w34211 <= not w3805 and not w34210;
w34212 <= not w34004 and w34138;
w34213 <= not pi0680 and w34004;
w34214 <= not w14926 and w34142;
w34215 <= pi0661 and not w34213;
w34216 <= not w34214 and w34215;
w34217 <= not w34009 and not w34212;
w34218 <= not w34216 and w34217;
w34219 <= w3805 and not w34218;
w34220 <= pi0222 and not w34219;
w34221 <= not w34211 and w34220;
w34222 <= not w34029 and w34138;
w34223 <= not pi0680 and w34029;
w34224 <= pi0616 and w15141;
w34225 <= pi0680 and not w34224;
w34226 <= not w14996 and w34225;
w34227 <= pi0661 and not w34223;
w34228 <= not w34226 and w34227;
w34229 <= not w34035 and not w34222;
w34230 <= not w34228 and w34229;
w34231 <= not w3805 and w34230;
w34232 <= not w3756 and w34002;
w34233 <= w14809 and w34031;
w34234 <= w14219 and not w34232;
w34235 <= not w34233 and w34234;
w34236 <= not w34002 and w34138;
w34237 <= not pi0680 and w34002;
w34238 <= pi0680 and not w14980;
w34239 <= not w34183 and w34238;
w34240 <= pi0661 and not w34237;
w34241 <= not w34239 and w34240;
w34242 <= not w34235 and not w34236;
w34243 <= not w34241 and w34242;
w34244 <= w3805 and w34243;
w34245 <= not pi0222 and not w34244;
w34246 <= not w34231 and w34245;
w34247 <= not w34221 and not w34246;
w34248 <= not w1011 and not w34247;
w34249 <= not pi0215 and not w34187;
w34250 <= not w34248 and w34249;
w34251 <= pi0299 and not w34182;
w34252 <= not w34250 and w34251;
w34253 <= w33829 and not w34185;
w34254 <= not w33829 and not w34002;
w34255 <= not pi0222 and not w34254;
w34256 <= not w34253 and w34255;
w34257 <= not w914 and not w34256;
w34258 <= not w3768 and w34230;
w34259 <= w3768 and w34243;
w34260 <= pi0224 and not w34259;
w34261 <= not w34258 and w34260;
w34262 <= not w34257 and not w34261;
w34263 <= w3768 and w34218;
w34264 <= not w3768 and w34210;
w34265 <= pi0222 and not w34263;
w34266 <= not w34264 and w34265;
w34267 <= not w34262 and not w34266;
w34268 <= not pi0223 and not w34267;
w34269 <= w3768 and not w34147;
w34270 <= not w3768 and not w34158;
w34271 <= pi0222 and not w34269;
w34272 <= not w34270 and w34271;
w34273 <= w3768 and not w34163;
w34274 <= not w3768 and w34177;
w34275 <= not pi0222 and not w34273;
w34276 <= not w34274 and w34275;
w34277 <= pi0223 and not w34276;
w34278 <= not w34272 and w34277;
w34279 <= not pi0299 and not w34278;
w34280 <= not w34268 and w34279;
w34281 <= pi0039 and not w34280;
w34282 <= not w34252 and w34281;
w34283 <= pi0661 and w15181;
w34284 <= pi0616 and w14789;
w34285 <= not pi0222 and not w34284;
w34286 <= not w34283 and w34285;
w34287 <= not pi0616 and w14789;
w34288 <= w15180 and not w33829;
w34289 <= not pi0603 and not w14498;
w34290 <= not w14930 and not w15177;
w34291 <= not w34289 and w34290;
w34292 <= not w34287 and not w34291;
w34293 <= not w34288 and w34292;
w34294 <= pi0222 and not w34293;
w34295 <= not w34286 and not w34294;
w34296 <= not pi0299 and not w34295;
w34297 <= not pi0616 and w14794;
w34298 <= w15185 and not w33829;
w34299 <= not pi0603 and not w14507;
w34300 <= not w14686 and not w14930;
w34301 <= not w34299 and w34300;
w34302 <= not w34297 and not w34301;
w34303 <= not w34298 and w34302;
w34304 <= pi0222 and not w34303;
w34305 <= pi0661 and w15186;
w34306 <= pi0616 and w14794;
w34307 <= not pi0222 and not w34306;
w34308 <= not w34305 and w34307;
w34309 <= not w34304 and not w34308;
w34310 <= pi0299 and not w34309;
w34311 <= not pi0039 and not w34296;
w34312 <= not w34310 and w34311;
w34313 <= not pi0038 and not w34312;
w34314 <= not w34282 and w34313;
w34315 <= w134 and not w34137;
w34316 <= not w34314 and w34315;
w34317 <= not w33824 and not w34316;
w34318 <= not pi0625 and w34317;
w34319 <= pi0625 and w34074;
w34320 <= not pi1153 and not w34319;
w34321 <= not w34318 and w34320;
w34322 <= not pi0608 and not w33927;
w34323 <= not w34321 and w34322;
w34324 <= not pi0625 and w34074;
w34325 <= pi0625 and w34317;
w34326 <= pi1153 and not w34324;
w34327 <= not w34325 and w34326;
w34328 <= pi0608 and not w33931;
w34329 <= not w34327 and w34328;
w34330 <= not w34323 and not w34329;
w34331 <= pi0778 and not w34330;
w34332 <= not pi0778 and w34317;
w34333 <= not w34331 and not w34332;
w34334 <= not pi0609 and not w34333;
w34335 <= not pi1155 and not w34124;
w34336 <= not w34334 and w34335;
w34337 <= not pi0660 and not w34082;
w34338 <= not w34336 and w34337;
w34339 <= not pi0609 and w33934;
w34340 <= pi0609 and not w34333;
w34341 <= pi1155 and not w34339;
w34342 <= not w34340 and w34341;
w34343 <= pi0660 and not w34086;
w34344 <= not w34342 and w34343;
w34345 <= not w34338 and not w34344;
w34346 <= pi0785 and not w34345;
w34347 <= not pi0785 and not w34333;
w34348 <= not w34346 and not w34347;
w34349 <= not pi0618 and not w34348;
w34350 <= pi0618 and w33937;
w34351 <= not pi1154 and not w34350;
w34352 <= not w34349 and w34351;
w34353 <= not pi0627 and not w34094;
w34354 <= not w34352 and w34353;
w34355 <= not pi0618 and w33937;
w34356 <= pi0618 and not w34348;
w34357 <= pi1154 and not w34355;
w34358 <= not w34356 and w34357;
w34359 <= pi0627 and not w34098;
w34360 <= not w34358 and w34359;
w34361 <= not w34354 and not w34360;
w34362 <= pi0781 and not w34361;
w34363 <= not pi0781 and not w34348;
w34364 <= not w34362 and not w34363;
w34365 <= not pi0789 and w34364;
w34366 <= not pi0626 and w34113;
w34367 <= pi0626 and not w33822;
w34368 <= w14192 and not w34367;
w34369 <= not w34366 and w34368;
w34370 <= w14198 and not w33822;
w34371 <= w15434 and not w34370;
w34372 <= not w33941 and w34371;
w34373 <= pi0626 and w34113;
w34374 <= not pi0626 and not w33822;
w34375 <= w14191 and not w34374;
w34376 <= not w34373 and w34375;
w34377 <= not w34369 and not w34372;
w34378 <= not w34376 and w34377;
w34379 <= pi0788 and not w34378;
w34380 <= not pi0619 and not w34364;
w34381 <= pi0619 and w33940;
w34382 <= not pi1159 and not w34381;
w34383 <= not w34380 and w34382;
w34384 <= not pi0648 and not w34106;
w34385 <= not w34383 and w34384;
w34386 <= pi0619 and not w34364;
w34387 <= not pi0619 and w33940;
w34388 <= pi1159 and not w34387;
w34389 <= not w34386 and w34388;
w34390 <= pi0648 and not w34110;
w34391 <= not w34389 and w34390;
w34392 <= pi0789 and not w34385;
w34393 <= not w34391 and w34392;
w34394 <= not w34365 and not w34379;
w34395 <= not w34393 and w34394;
w34396 <= not w15533 and w34378;
w34397 <= not w17927 and not w34396;
w34398 <= not w34395 and w34397;
w34399 <= not w34123 and not w34398;
w34400 <= not w17769 and not w34399;
w34401 <= not pi0630 and w33955;
w34402 <= not w15342 and w34115;
w34403 <= w15342 and w33822;
w34404 <= not w34402 and not w34403;
w34405 <= not w18122 and not w34404;
w34406 <= pi0630 and w33951;
w34407 <= not w34401 and not w34406;
w34408 <= not w34405 and w34407;
w34409 <= pi0787 and not w34408;
w34410 <= not w34400 and not w34409;
w34411 <= pi0644 and w34410;
w34412 <= pi0715 and not w33959;
w34413 <= not w34411 and w34412;
w34414 <= w15367 and not w33822;
w34415 <= not w15367 and w34404;
w34416 <= not w34414 and not w34415;
w34417 <= pi0644 and not w34416;
w34418 <= not pi0644 and not w33822;
w34419 <= not pi0715 and not w34418;
w34420 <= not w34417 and w34419;
w34421 <= pi1160 and not w34420;
w34422 <= not w34413 and w34421;
w34423 <= pi0644 and w33958;
w34424 <= not pi0644 and w34410;
w34425 <= not pi0715 and not w34423;
w34426 <= not w34424 and w34425;
w34427 <= not pi0644 and not w34416;
w34428 <= pi0644 and not w33822;
w34429 <= pi0715 and not w34428;
w34430 <= not w34427 and w34429;
w34431 <= not pi1160 and not w34430;
w34432 <= not w34426 and w34431;
w34433 <= not w34422 and not w34432;
w34434 <= pi0790 and not w34433;
w34435 <= not pi0790 and w34410;
w34436 <= not w34434 and not w34435;
w34437 <= w4989 and not w34436;
w34438 <= not pi0222 and not w4989;
w34439 <= not w34437 and not w34438;
w34440 <= not pi0299 and not w14555;
w34441 <= pi0039 and not w34440;
w34442 <= not w14608 and w34441;
w34443 <= w12436 and not w15710;
w34444 <= not w34442 and w34443;
w34445 <= w16154 and not w34444;
w34446 <= pi0223 and not w34445;
w34447 <= not w16712 and not w34446;
w34448 <= w14638 and not w34446;
w34449 <= pi0223 and not w134;
w34450 <= pi0680 and pi0681;
w34451 <= w14481 and not w34450;
w34452 <= not pi0223 and not w14481;
w34453 <= pi0223 and w14498;
w34454 <= not pi0299 and not w34453;
w34455 <= not w34451 and w34454;
w34456 <= not w34452 and w34455;
w34457 <= pi0223 and w14507;
w34458 <= w14486 and not w34450;
w34459 <= not pi0223 and not w14486;
w34460 <= pi0299 and not w34457;
w34461 <= not w34458 and w34460;
w34462 <= not w34459 and w34461;
w34463 <= not pi0039 and not w34456;
w34464 <= not w34462 and w34463;
w34465 <= pi0681 and w14302;
w34466 <= w166 and not w34465;
w34467 <= not w14253 and w34450;
w34468 <= w3768 and w34467;
w34469 <= pi0681 and w14266;
w34470 <= not w3768 and w34469;
w34471 <= not w166 and not w34468;
w34472 <= not w34470 and w34471;
w34473 <= not w34466 and not w34472;
w34474 <= not pi0223 and not w34473;
w34475 <= pi0681 and not w33882;
w34476 <= not w14552 and not w34475;
w34477 <= w3768 and not w34476;
w34478 <= pi0681 and not w14381;
w34479 <= not w14532 and not w34478;
w34480 <= not w3768 and not w34479;
w34481 <= pi0223 and not w34477;
w34482 <= not w34480 and w34481;
w34483 <= not pi0299 and not w34482;
w34484 <= not w34474 and w34483;
w34485 <= not pi0223 and pi0681;
w34486 <= w14307 and w34485;
w34487 <= w3805 and w34476;
w34488 <= not w3805 and w34479;
w34489 <= pi0223 and not w34487;
w34490 <= not w34488 and w34489;
w34491 <= pi0215 and not w34486;
w34492 <= not w34490 and w34491;
w34493 <= pi0223 and not w14216;
w34494 <= w1011 and not w34493;
w34495 <= not w34465 and w34494;
w34496 <= pi0681 and not w33846;
w34497 <= not w3805 and not w14580;
w34498 <= not w34496 and w34497;
w34499 <= pi0681 and not w14349;
w34500 <= w3805 and not w14573;
w34501 <= not w34499 and w34500;
w34502 <= pi0223 and not w34498;
w34503 <= not w34501 and w34502;
w34504 <= not w3805 and not w34469;
w34505 <= w3805 and not w34467;
w34506 <= not pi0223 and not w34504;
w34507 <= not w34505 and w34506;
w34508 <= not w1011 and not w34507;
w34509 <= not w34503 and w34508;
w34510 <= not w34495 and not w34509;
w34511 <= not pi0215 and not w34510;
w34512 <= pi0299 and not w34492;
w34513 <= not w34511 and w34512;
w34514 <= pi0039 and not w34484;
w34515 <= not w34513 and w34514;
w34516 <= not w34464 and not w34515;
w34517 <= not pi0038 and not w34516;
w34518 <= pi0681 and w14209;
w34519 <= pi0223 and not w14204;
w34520 <= pi0038 and not w34518;
w34521 <= not w34519 and w34520;
w34522 <= w134 and not w34521;
w34523 <= not w34517 and w34522;
w34524 <= not w34449 and not w34523;
w34525 <= not pi0778 and not w34524;
w34526 <= pi0625 and w34524;
w34527 <= not pi0625 and not w34446;
w34528 <= pi1153 and not w34527;
w34529 <= not w34526 and w34528;
w34530 <= not pi0625 and w34524;
w34531 <= pi0625 and not w34446;
w34532 <= not pi1153 and not w34531;
w34533 <= not w34530 and w34532;
w34534 <= not w34529 and not w34533;
w34535 <= pi0778 and not w34534;
w34536 <= not w34525 and not w34535;
w34537 <= not w14638 and w34536;
w34538 <= not w34448 and not w34537;
w34539 <= not w14202 and w34538;
w34540 <= w14202 and w34446;
w34541 <= not w34539 and not w34540;
w34542 <= not w14198 and w34541;
w34543 <= not w14194 and w34542;
w34544 <= not w34447 and not w34543;
w34545 <= not w16705 and not w34544;
w34546 <= w15419 and not w34446;
w34547 <= not w34545 and not w34546;
w34548 <= not pi0787 and w34547;
w34549 <= not pi0647 and not w34547;
w34550 <= pi0647 and not w34446;
w34551 <= not pi1157 and not w34550;
w34552 <= not w34549 and w34551;
w34553 <= pi0647 and not w34547;
w34554 <= not pi0647 and not w34446;
w34555 <= pi1157 and not w34554;
w34556 <= not w34553 and w34555;
w34557 <= not w34552 and not w34556;
w34558 <= pi0787 and not w34557;
w34559 <= not w34548 and not w34558;
w34560 <= not pi0644 and w34559;
w34561 <= not pi0630 and w34556;
w34562 <= w15532 and not w34446;
w34563 <= w14680 and not w34446;
w34564 <= pi0039 and pi0223;
w34565 <= pi0038 and not w34564;
w34566 <= pi0642 and w14731;
w34567 <= w14230 and not w34566;
w34568 <= not pi0223 and not w14230;
w34569 <= not pi0039 and not w34568;
w34570 <= not w34567 and w34569;
w34571 <= w34565 and not w34570;
w34572 <= not pi0223 and pi0642;
w34573 <= w14789 and w34572;
w34574 <= not pi0299 and not w34573;
w34575 <= not pi0642 and w14789;
w34576 <= pi0223 and not w34575;
w34577 <= w14700 and w34576;
w34578 <= w34574 and not w34577;
w34579 <= w14794 and w34572;
w34580 <= pi0299 and not w34579;
w34581 <= w3753 and w14793;
w34582 <= pi0223 and not w14687;
w34583 <= not w34581 and w34582;
w34584 <= w34580 and not w34583;
w34585 <= not pi0039 and not w34584;
w34586 <= not w34578 and w34585;
w34587 <= w33460 and not w34566;
w34588 <= pi0642 and not w14732;
w34589 <= w33988 and not w34588;
w34590 <= not w34587 and not w34589;
w34591 <= pi0681 and w34590;
w34592 <= w3757 and w34567;
w34593 <= w14360 and w34592;
w34594 <= not w3757 and not w34590;
w34595 <= not pi0681 and not w34593;
w34596 <= not w34594 and w34595;
w34597 <= not w34591 and not w34596;
w34598 <= w3768 and w34597;
w34599 <= not pi0642 and not w14377;
w34600 <= pi0642 and not w14746;
w34601 <= not w34599 and not w34600;
w34602 <= not w3757 and w34601;
w34603 <= pi0642 and not w14745;
w34604 <= w3757 and not w34603;
w34605 <= not w14284 and w34604;
w34606 <= not pi0681 and not w34605;
w34607 <= not w34602 and w34606;
w34608 <= pi0681 and not w34601;
w34609 <= not w34607 and not w34608;
w34610 <= not w3768 and w34609;
w34611 <= pi0223 and not w34610;
w34612 <= not w34598 and w34611;
w34613 <= pi0642 and w14798;
w34614 <= w166 and not w34613;
w34615 <= not w3757 and w34613;
w34616 <= not pi0681 and not w34615;
w34617 <= pi0642 and w3757;
w34618 <= w14809 and w34617;
w34619 <= w34616 and not w34618;
w34620 <= pi0681 and not w34613;
w34621 <= not w34619 and not w34620;
w34622 <= w3768 and w34621;
w34623 <= not w14262 and w34566;
w34624 <= pi0681 and not w34623;
w34625 <= w14938 and w34617;
w34626 <= not w3757 and w34623;
w34627 <= not pi0681 and not w34625;
w34628 <= not w34626 and w34627;
w34629 <= not w34624 and not w34628;
w34630 <= not w3768 and w34629;
w34631 <= not w166 and not w34622;
w34632 <= not w34630 and w34631;
w34633 <= not pi0223 and not w34614;
w34634 <= not w34632 and w34633;
w34635 <= not pi0299 and not w34612;
w34636 <= not w34634 and w34635;
w34637 <= w14799 and w34617;
w34638 <= w34616 and not w34637;
w34639 <= w14286 and w34606;
w34640 <= not w34638 and not w34639;
w34641 <= pi0642 and w14800;
w34642 <= pi0681 and not w34641;
w34643 <= w34640 and not w34642;
w34644 <= pi0947 and not w34643;
w34645 <= w3805 and not w34638;
w34646 <= w34613 and w34645;
w34647 <= not w18486 and w34643;
w34648 <= not pi0947 and not w34646;
w34649 <= not w34647 and w34648;
w34650 <= not pi0223 and not w34644;
w34651 <= not w34649 and w34650;
w34652 <= not w3805 and w34609;
w34653 <= w3805 and w34597;
w34654 <= pi0223 and not w34652;
w34655 <= not w34653 and w34654;
w34656 <= not w34651 and not w34655;
w34657 <= pi0215 and not w34656;
w34658 <= w34494 and not w34613;
w34659 <= pi0947 and not w34629;
w34660 <= w18486 and w34621;
w34661 <= not w18486 and w34629;
w34662 <= not pi0947 and not w34660;
w34663 <= not w34661 and w34662;
w34664 <= not pi0223 and not w34659;
w34665 <= not w34663 and w34664;
w34666 <= pi0642 and not w14717;
w34667 <= not pi0642 and not w14265;
w34668 <= not w34666 and not w34667;
w34669 <= pi0681 and not w34668;
w34670 <= not w3757 and w34668;
w34671 <= w14577 and not w34566;
w34672 <= not pi0681 and not w34671;
w34673 <= not w34670 and w34672;
w34674 <= not w3805 and not w34673;
w34675 <= not w34669 and w34674;
w34676 <= w3754 and not w34588;
w34677 <= not w14333 and w34676;
w34678 <= not w34587 and not w34677;
w34679 <= pi0681 and w34678;
w34680 <= not w3757 and not w34678;
w34681 <= not w14727 and not w33457;
w34682 <= w3757 and not w34681;
w34683 <= not pi0681 and not w34682;
w34684 <= not w34680 and w34683;
w34685 <= w3805 and not w34684;
w34686 <= not w34679 and w34685;
w34687 <= pi0223 and not w34675;
w34688 <= not w34686 and w34687;
w34689 <= not w1011 and not w34665;
w34690 <= not w34688 and w34689;
w34691 <= not pi0215 and not w34658;
w34692 <= not w34690 and w34691;
w34693 <= pi0299 and not w34657;
w34694 <= not w34692 and w34693;
w34695 <= pi0039 and not w34636;
w34696 <= not w34694 and w34695;
w34697 <= not pi0038 and not w34586;
w34698 <= not w34696 and w34697;
w34699 <= w134 and not w34571;
w34700 <= not w34698 and w34699;
w34701 <= not w34449 and not w34700;
w34702 <= not w14680 and w34701;
w34703 <= not w34563 and not w34702;
w34704 <= not pi0785 and w34703;
w34705 <= pi0609 and not w34703;
w34706 <= not pi0609 and not w34446;
w34707 <= pi1155 and not w34706;
w34708 <= not w34705 and w34707;
w34709 <= not pi0609 and not w34703;
w34710 <= pi0609 and not w34446;
w34711 <= not pi1155 and not w34710;
w34712 <= not w34709 and w34711;
w34713 <= not w34708 and not w34712;
w34714 <= pi0785 and not w34713;
w34715 <= not w34704 and not w34714;
w34716 <= not pi0781 and not w34715;
w34717 <= pi0618 and w34715;
w34718 <= not pi0618 and not w34446;
w34719 <= pi1154 and not w34718;
w34720 <= not w34717 and w34719;
w34721 <= not pi0618 and w34715;
w34722 <= pi0618 and not w34446;
w34723 <= not pi1154 and not w34722;
w34724 <= not w34721 and w34723;
w34725 <= not w34720 and not w34724;
w34726 <= pi0781 and not w34725;
w34727 <= not w34716 and not w34726;
w34728 <= not pi0789 and not w34727;
w34729 <= pi0619 and w34727;
w34730 <= not pi0619 and not w34446;
w34731 <= pi1159 and not w34730;
w34732 <= not w34729 and w34731;
w34733 <= not pi0619 and w34727;
w34734 <= pi0619 and not w34446;
w34735 <= not pi1159 and not w34734;
w34736 <= not w34733 and w34735;
w34737 <= not w34732 and not w34736;
w34738 <= pi0789 and not w34737;
w34739 <= not w34728 and not w34738;
w34740 <= not w15532 and w34739;
w34741 <= not w34562 and not w34740;
w34742 <= not w15342 and w34741;
w34743 <= w15342 and w34446;
w34744 <= not w34742 and not w34743;
w34745 <= not w18122 and not w34744;
w34746 <= pi0630 and w34552;
w34747 <= not w34561 and not w34746;
w34748 <= not w34745 and w34747;
w34749 <= pi0787 and not w34748;
w34750 <= pi0628 and not w34446;
w34751 <= not pi0628 and not w34544;
w34752 <= w15340 and not w34750;
w34753 <= not w34751 and w34752;
w34754 <= not w18133 and w34741;
w34755 <= not pi0628 and not w34446;
w34756 <= pi0628 and not w34544;
w34757 <= w15339 and not w34755;
w34758 <= not w34756 and w34757;
w34759 <= not w34753 and not w34758;
w34760 <= not w34754 and w34759;
w34761 <= pi0792 and not w34760;
w34762 <= w14198 and not w34446;
w34763 <= not w34542 and not w34762;
w34764 <= w15434 and not w34763;
w34765 <= not pi0626 and w34446;
w34766 <= pi0626 and not w34739;
w34767 <= w14191 and not w34765;
w34768 <= not w34766 and w34767;
w34769 <= pi0626 and w34446;
w34770 <= not pi0626 and not w34739;
w34771 <= w14192 and not w34769;
w34772 <= not w34770 and w34771;
w34773 <= not w34764 and not w34768;
w34774 <= not w34772 and w34773;
w34775 <= pi0788 and not w34774;
w34776 <= pi0609 and w34536;
w34777 <= not w34450 and w34566;
w34778 <= not pi0642 and not w14899;
w34779 <= w34450 and not w34778;
w34780 <= not w34125 and w34779;
w34781 <= not w34777 and not w34780;
w34782 <= not w34450 and w34567;
w34783 <= pi0642 and w15056;
w34784 <= not w34778 and not w34783;
w34785 <= w14230 and not w34784;
w34786 <= w34450 and w34785;
w34787 <= pi0223 and not w34782;
w34788 <= not w34786 and w34787;
w34789 <= w34781 and not w34788;
w34790 <= w34569 and not w34789;
w34791 <= w34565 and not w34790;
w34792 <= w15181 and w34485;
w34793 <= w15180 and not w34450;
w34794 <= not w34291 and w34576;
w34795 <= not w34793 and w34794;
w34796 <= w34574 and not w34792;
w34797 <= not w34795 and w34796;
w34798 <= w15186 and w34485;
w34799 <= w15185 and not w34450;
w34800 <= pi0223 and not w34581;
w34801 <= not w34301 and w34800;
w34802 <= not w34799 and w34801;
w34803 <= w34580 and not w34798;
w34804 <= not w34802 and w34803;
w34805 <= not pi0039 and not w34797;
w34806 <= not w34804 and w34805;
w34807 <= not w34450 and not w34591;
w34808 <= not w14213 and w34785;
w34809 <= not w3754 and not w34808;
w34810 <= pi0680 and not w34809;
w34811 <= pi0642 and not w15067;
w34812 <= not pi0614 and w14906;
w34813 <= not w34811 and not w34812;
w34814 <= not pi0616 and not w34813;
w34815 <= w34810 and not w34814;
w34816 <= not w34807 and not w34815;
w34817 <= not w34596 and not w34816;
w34818 <= w3805 and not w34817;
w34819 <= not pi0680 and w34601;
w34820 <= pi0642 and not w34151;
w34821 <= not w3754 and w14888;
w34822 <= pi0680 and not w14892;
w34823 <= not w34820 and w34822;
w34824 <= not w34821 and w34823;
w34825 <= pi0681 and not w34824;
w34826 <= not w34819 and w34825;
w34827 <= not w34607 and not w34826;
w34828 <= not w3805 and not w34827;
w34829 <= pi0223 and not w34828;
w34830 <= not w34818 and w34829;
w34831 <= not pi0680 and not w34613;
w34832 <= not w14899 and not w34811;
w34833 <= w33460 and not w34832;
w34834 <= pi0680 and not w34833;
w34835 <= pi0642 and not w15111;
w34836 <= w3754 and not w34835;
w34837 <= not w15018 and w34836;
w34838 <= w34834 and not w34837;
w34839 <= not w34831 and not w34838;
w34840 <= pi0681 and not w34839;
w34841 <= w34645 and not w34840;
w34842 <= not w34450 and not w34642;
w34843 <= not pi0642 and not w3754;
w34844 <= not w15013 and w34843;
w34845 <= w15017 and w15122;
w34846 <= w14730 and not w34845;
w34847 <= pi0642 and w34170;
w34848 <= pi0680 and not w34844;
w34849 <= not w34847 and w34848;
w34850 <= not w34846 and w34849;
w34851 <= not w34842 and not w34850;
w34852 <= not w3805 and w34640;
w34853 <= not w34851 and w34852;
w34854 <= not pi0223 and not w34841;
w34855 <= not w34853 and w34854;
w34856 <= pi0215 and not w34855;
w34857 <= not w34830 and w34856;
w34858 <= not w34450 and not w34679;
w34859 <= not w14922 and not w34811;
w34860 <= w3754 and not w34859;
w34861 <= w34810 and not w34860;
w34862 <= not w34858 and not w34861;
w34863 <= w34685 and not w34862;
w34864 <= not w34450 and not w34669;
w34865 <= pi0642 and not w34201;
w34866 <= w14730 and not w34194;
w34867 <= w34196 and w34843;
w34868 <= pi0680 and not w34865;
w34869 <= not w34866 and w34868;
w34870 <= not w34867 and w34869;
w34871 <= not w34864 and not w34870;
w34872 <= w34674 and not w34871;
w34873 <= pi0223 and not w34872;
w34874 <= not w34863 and w34873;
w34875 <= not pi0642 and not w14977;
w34876 <= w34836 and not w34875;
w34877 <= w34834 and not w34876;
w34878 <= not w34831 and not w34877;
w34879 <= pi0681 and not w34878;
w34880 <= not w34619 and not w34879;
w34881 <= w3805 and not w34880;
w34882 <= not w34450 and not w34624;
w34883 <= pi0642 and w15141;
w34884 <= not w14985 and w34843;
w34885 <= pi0680 and not w34883;
w34886 <= not w14993 and w34885;
w34887 <= not w34884 and w34886;
w34888 <= not w34882 and not w34887;
w34889 <= not w34628 and not w34888;
w34890 <= not w3805 and not w34889;
w34891 <= not pi0223 and not w34881;
w34892 <= not w34890 and w34891;
w34893 <= not w1011 and not w34874;
w34894 <= not w34892 and w34893;
w34895 <= w14216 and not w34781;
w34896 <= not pi0223 and w34895;
w34897 <= w34494 and not w34788;
w34898 <= not w34896 and w34897;
w34899 <= not pi0215 and not w34898;
w34900 <= not w34894 and w34899;
w34901 <= pi0299 and not w34857;
w34902 <= not w34900 and w34901;
w34903 <= w3768 and w34817;
w34904 <= not w3768 and w34827;
w34905 <= pi0223 and not w34904;
w34906 <= not w34903 and w34905;
w34907 <= w166 and not w34895;
w34908 <= not w3768 and w34889;
w34909 <= w3768 and w34880;
w34910 <= not w166 and not w34908;
w34911 <= not w34909 and w34910;
w34912 <= not pi0223 and not w34907;
w34913 <= not w34911 and w34912;
w34914 <= not pi0299 and not w34906;
w34915 <= not w34913 and w34914;
w34916 <= pi0039 and not w34915;
w34917 <= not w34902 and w34916;
w34918 <= not pi0038 and not w34806;
w34919 <= not w34917 and w34918;
w34920 <= w134 and not w34791;
w34921 <= not w34919 and w34920;
w34922 <= not w34449 and not w34921;
w34923 <= not pi0625 and w34922;
w34924 <= pi0625 and w34701;
w34925 <= not pi1153 and not w34924;
w34926 <= not w34923 and w34925;
w34927 <= not pi0608 and not w34926;
w34928 <= not w34529 and w34927;
w34929 <= not pi0625 and w34701;
w34930 <= pi0625 and w34922;
w34931 <= pi1153 and not w34929;
w34932 <= not w34930 and w34931;
w34933 <= pi0608 and not w34932;
w34934 <= not w34533 and w34933;
w34935 <= not w34928 and not w34934;
w34936 <= pi0778 and not w34935;
w34937 <= not pi0778 and w34922;
w34938 <= not w34936 and not w34937;
w34939 <= not pi0609 and not w34938;
w34940 <= not pi1155 and not w34776;
w34941 <= not w34939 and w34940;
w34942 <= not pi0660 and not w34708;
w34943 <= not w34941 and w34942;
w34944 <= not pi0609 and w34536;
w34945 <= pi0609 and not w34938;
w34946 <= pi1155 and not w34944;
w34947 <= not w34945 and w34946;
w34948 <= pi0660 and not w34712;
w34949 <= not w34947 and w34948;
w34950 <= not w34943 and not w34949;
w34951 <= pi0785 and not w34950;
w34952 <= not pi0785 and not w34938;
w34953 <= not w34951 and not w34952;
w34954 <= not pi0618 and not w34953;
w34955 <= pi0618 and not w34538;
w34956 <= not pi1154 and not w34955;
w34957 <= not w34954 and w34956;
w34958 <= not pi0627 and not w34720;
w34959 <= not w34957 and w34958;
w34960 <= pi0618 and not w34953;
w34961 <= not pi0618 and not w34538;
w34962 <= pi1154 and not w34961;
w34963 <= not w34960 and w34962;
w34964 <= pi0627 and not w34724;
w34965 <= not w34963 and w34964;
w34966 <= not w34959 and not w34965;
w34967 <= pi0781 and not w34966;
w34968 <= not pi0781 and not w34953;
w34969 <= not w34967 and not w34968;
w34970 <= not pi0789 and w34969;
w34971 <= not pi0619 and not w34969;
w34972 <= pi0619 and w34541;
w34973 <= not pi1159 and not w34972;
w34974 <= not w34971 and w34973;
w34975 <= not pi0648 and not w34732;
w34976 <= not w34974 and w34975;
w34977 <= not pi0619 and w34541;
w34978 <= pi0619 and not w34969;
w34979 <= pi1159 and not w34977;
w34980 <= not w34978 and w34979;
w34981 <= pi0648 and not w34736;
w34982 <= not w34980 and w34981;
w34983 <= pi0789 and not w34976;
w34984 <= not w34982 and w34983;
w34985 <= w15533 and not w34970;
w34986 <= not w34984 and w34985;
w34987 <= not w34775 and not w34986;
w34988 <= not w34761 and not w34987;
w34989 <= w17927 and w34760;
w34990 <= not w17769 and not w34989;
w34991 <= not w34988 and w34990;
w34992 <= not w34749 and not w34991;
w34993 <= pi0644 and w34992;
w34994 <= pi0715 and not w34560;
w34995 <= not w34993 and w34994;
w34996 <= w15367 and not w34446;
w34997 <= not w15367 and w34744;
w34998 <= not w34996 and not w34997;
w34999 <= pi0644 and not w34998;
w35000 <= not pi0644 and not w34446;
w35001 <= not pi0715 and not w35000;
w35002 <= not w34999 and w35001;
w35003 <= pi1160 and not w35002;
w35004 <= not w34995 and w35003;
w35005 <= pi0644 and w34559;
w35006 <= not pi0644 and w34992;
w35007 <= not pi0715 and not w35005;
w35008 <= not w35006 and w35007;
w35009 <= not pi0644 and not w34998;
w35010 <= pi0644 and not w34446;
w35011 <= pi0715 and not w35010;
w35012 <= not w35009 and w35011;
w35013 <= not pi1160 and not w35012;
w35014 <= not w35008 and w35013;
w35015 <= not w35004 and not w35014;
w35016 <= pi0790 and not w35015;
w35017 <= not pi0790 and w34992;
w35018 <= not w35016 and not w35017;
w35019 <= w4989 and not w35018;
w35020 <= not pi0223 and not w4989;
w35021 <= not w35019 and not w35020;
w35022 <= pi0224 and not w33821;
w35023 <= not w16712 and not w35022;
w35024 <= pi0224 and not w134;
w35025 <= pi0224 and not w14204;
w35026 <= pi0038 and not w35025;
w35027 <= pi0662 and w14209;
w35028 <= w35026 and not w35027;
w35029 <= pi0662 and pi0680;
w35030 <= w14481 and not w35029;
w35031 <= not pi0224 and not w14481;
w35032 <= pi0224 and w14498;
w35033 <= not pi0299 and not w35032;
w35034 <= not w35030 and w35033;
w35035 <= not w35031 and w35034;
w35036 <= pi0224 and w14507;
w35037 <= w14486 and not w35029;
w35038 <= not pi0224 and not w14486;
w35039 <= pi0299 and not w35036;
w35040 <= not w35037 and w35039;
w35041 <= not w35038 and w35040;
w35042 <= not pi0039 and not w35035;
w35043 <= not w35041 and w35042;
w35044 <= pi0662 and w14218;
w35045 <= not w3756 and not w33846;
w35046 <= w14581 and not w35045;
w35047 <= not w3768 and w35046;
w35048 <= pi0662 and not w14349;
w35049 <= not pi0662 and not w14574;
w35050 <= not w35048 and not w35049;
w35051 <= w3768 and w35050;
w35052 <= pi0224 and not w35047;
w35053 <= not w35051 and w35052;
w35054 <= pi0662 and w14266;
w35055 <= not w3768 and not w35054;
w35056 <= not w14253 and w35029;
w35057 <= w3768 and not w35056;
w35058 <= w3373 and not w35055;
w35059 <= not w35057 and w35058;
w35060 <= not pi0223 and not w35044;
w35061 <= not w35059 and w35060;
w35062 <= not w35053 and w35061;
w35063 <= not pi0224 and pi0662;
w35064 <= w14292 and w35063;
w35065 <= not pi0662 and not w14553;
w35066 <= pi0662 and not w33882;
w35067 <= not w35065 and not w35066;
w35068 <= w3768 and w35067;
w35069 <= not pi0662 and not w14533;
w35070 <= pi0662 and not w14381;
w35071 <= not w35069 and not w35070;
w35072 <= not w3768 and w35071;
w35073 <= pi0224 and not w35068;
w35074 <= not w35072 and w35073;
w35075 <= pi0223 and not w35064;
w35076 <= not w35074 and w35075;
w35077 <= not pi0299 and not w35076;
w35078 <= not w35062 and w35077;
w35079 <= pi0224 and not w14216;
w35080 <= w1011 and not w35079;
w35081 <= w14221 and w35029;
w35082 <= w35080 and not w35081;
w35083 <= not w3805 and w35046;
w35084 <= w3805 and w35050;
w35085 <= pi0224 and not w35083;
w35086 <= not w35084 and w35085;
w35087 <= not w3805 and not w35054;
w35088 <= w3805 and not w35056;
w35089 <= not pi0224 and not w35087;
w35090 <= not w35088 and w35089;
w35091 <= not w1011 and not w35090;
w35092 <= not w35086 and w35091;
w35093 <= not w35082 and not w35092;
w35094 <= not pi0215 and not w35093;
w35095 <= w14307 and w35063;
w35096 <= w3805 and w35067;
w35097 <= not w3805 and w35071;
w35098 <= pi0224 and not w35096;
w35099 <= not w35097 and w35098;
w35100 <= pi0215 and not w35095;
w35101 <= not w35099 and w35100;
w35102 <= pi0299 and not w35101;
w35103 <= not w35094 and w35102;
w35104 <= pi0039 and not w35078;
w35105 <= not w35103 and w35104;
w35106 <= not w35043 and not w35105;
w35107 <= not pi0038 and not w35106;
w35108 <= w134 and not w35028;
w35109 <= not w35107 and w35108;
w35110 <= not w35024 and not w35109;
w35111 <= not pi0778 and not w35110;
w35112 <= pi0625 and w35110;
w35113 <= not pi0625 and not w35022;
w35114 <= pi1153 and not w35113;
w35115 <= not w35112 and w35114;
w35116 <= not pi0625 and w35110;
w35117 <= pi0625 and not w35022;
w35118 <= not pi1153 and not w35117;
w35119 <= not w35116 and w35118;
w35120 <= not w35115 and not w35119;
w35121 <= pi0778 and not w35120;
w35122 <= not w35111 and not w35121;
w35123 <= not w14638 and not w35122;
w35124 <= w14638 and w35022;
w35125 <= not w35123 and not w35124;
w35126 <= not w14202 and not w35125;
w35127 <= w14202 and w35022;
w35128 <= not w35126 and not w35127;
w35129 <= not w14198 and w35128;
w35130 <= not w14194 and w35129;
w35131 <= not w35023 and not w35130;
w35132 <= not w16705 and not w35131;
w35133 <= w15419 and not w35022;
w35134 <= not w35132 and not w35133;
w35135 <= not pi0787 and w35134;
w35136 <= not pi0647 and not w35134;
w35137 <= pi0647 and not w35022;
w35138 <= not pi1157 and not w35137;
w35139 <= not w35136 and w35138;
w35140 <= pi0647 and not w35134;
w35141 <= not pi0647 and not w35022;
w35142 <= pi1157 and not w35141;
w35143 <= not w35140 and w35142;
w35144 <= not w35139 and not w35143;
w35145 <= pi0787 and not w35144;
w35146 <= not w35135 and not w35145;
w35147 <= not pi0644 and w35146;
w35148 <= pi0628 and not w35022;
w35149 <= not pi0628 and not w35131;
w35150 <= w15340 and not w35148;
w35151 <= not w35149 and w35150;
w35152 <= w15532 and not w35022;
w35153 <= pi0614 and w14843;
w35154 <= w35026 and not w35153;
w35155 <= pi0614 and w14789;
w35156 <= not pi0224 and w35155;
w35157 <= not pi0614 and w14789;
w35158 <= pi0224 and not w35157;
w35159 <= w14700 and w35158;
w35160 <= not pi0299 and not w35156;
w35161 <= not w35159 and w35160;
w35162 <= pi0614 and w14794;
w35163 <= pi0224 and w14685;
w35164 <= w35162 and not w35163;
w35165 <= pi0224 and not w14504;
w35166 <= not w35164 and not w35165;
w35167 <= pi0299 and w35166;
w35168 <= not pi0039 and not w35161;
w35169 <= not w35167 and w35168;
w35170 <= pi0614 and not w33974;
w35171 <= not pi0224 and w35170;
w35172 <= not w14306 and w35171;
w35173 <= pi0614 and not w14746;
w35174 <= not w33589 and not w35173;
w35175 <= not pi0680 and not w35174;
w35176 <= pi0680 and not w14750;
w35177 <= not w33591 and w35176;
w35178 <= not w35175 and not w35177;
w35179 <= w14220 and not w35178;
w35180 <= not w14220 and not w35174;
w35181 <= not w35179 and not w35180;
w35182 <= not w3805 and w35181;
w35183 <= pi0614 and w14731;
w35184 <= w14216 and not w35183;
w35185 <= not w3755 and not w35184;
w35186 <= not w14365 and not w35185;
w35187 <= not w14220 and not w35186;
w35188 <= not pi0680 and not w35186;
w35189 <= pi0680 and w35183;
w35190 <= not w14536 and not w35189;
w35191 <= not w35188 and w35190;
w35192 <= w14220 and not w35191;
w35193 <= not w35187 and not w35192;
w35194 <= w3805 and w35193;
w35195 <= pi0224 and not w35182;
w35196 <= not w35194 and w35195;
w35197 <= not w35172 and not w35196;
w35198 <= pi0215 and not w35197;
w35199 <= w14562 and w14731;
w35200 <= w35080 and not w35199;
w35201 <= pi0614 and not w14717;
w35202 <= not pi0614 and pi0616;
w35203 <= w14262 and w35202;
w35204 <= not w3760 and w14335;
w35205 <= w3754 and not w14260;
w35206 <= not w35204 and w35205;
w35207 <= not w35201 and not w35203;
w35208 <= not w35206 and w35207;
w35209 <= not w14220 and not w35208;
w35210 <= not pi0680 and not w35208;
w35211 <= pi0614 and w14938;
w35212 <= pi0680 and not w35211;
w35213 <= w14244 and w35212;
w35214 <= not w35189 and not w35213;
w35215 <= not w35210 and w35214;
w35216 <= w14220 and not w35215;
w35217 <= not w35209 and not w35216;
w35218 <= not w3805 and w35217;
w35219 <= not w14338 and not w35185;
w35220 <= not w14220 and not w35219;
w35221 <= not pi0680 and not w35219;
w35222 <= not w14558 and not w35189;
w35223 <= not w35221 and w35222;
w35224 <= w14220 and not w35223;
w35225 <= not w35220 and not w35224;
w35226 <= w3805 and w35225;
w35227 <= pi0224 and not w35218;
w35228 <= not w35226 and w35227;
w35229 <= not w14262 and w35183;
w35230 <= not pi0680 and not w35229;
w35231 <= not w35212 and not w35230;
w35232 <= w14220 and not w35231;
w35233 <= not w14220 and not w35229;
w35234 <= not w35232 and not w35233;
w35235 <= not w3805 and not w35234;
w35236 <= pi0614 and not w34026;
w35237 <= w3805 and not w35236;
w35238 <= not pi0224 and not w35237;
w35239 <= not w35235 and w35238;
w35240 <= not w1011 and not w35239;
w35241 <= not w35228 and w35240;
w35242 <= not pi0215 and not w35200;
w35243 <= not w35241 and w35242;
w35244 <= pi0299 and not w35198;
w35245 <= not w35243 and w35244;
w35246 <= not w14287 and w35171;
w35247 <= not w3768 and w35181;
w35248 <= w3768 and w35193;
w35249 <= pi0224 and not w35247;
w35250 <= not w35248 and w35249;
w35251 <= pi0223 and not w35246;
w35252 <= not w35250 and w35251;
w35253 <= pi0614 and w14831;
w35254 <= w3768 and not w35236;
w35255 <= not w3768 and not w35234;
w35256 <= w3373 and not w35254;
w35257 <= not w35255 and w35256;
w35258 <= not w3768 and w35217;
w35259 <= w3768 and w35225;
w35260 <= pi0224 and not w35258;
w35261 <= not w35259 and w35260;
w35262 <= not pi0223 and not w35253;
w35263 <= not w35257 and w35262;
w35264 <= not w35261 and w35263;
w35265 <= not w35252 and not w35264;
w35266 <= not pi0299 and not w35265;
w35267 <= pi0039 and not w35245;
w35268 <= not w35266 and w35267;
w35269 <= not pi0038 and not w35169;
w35270 <= not w35268 and w35269;
w35271 <= w134 and not w35154;
w35272 <= not w35270 and w35271;
w35273 <= not w35024 and not w35272;
w35274 <= not w14680 and not w35273;
w35275 <= w14680 and w35022;
w35276 <= not w35274 and not w35275;
w35277 <= not pi0785 and not w35276;
w35278 <= pi0609 and w35276;
w35279 <= not pi0609 and not w35022;
w35280 <= pi1155 and not w35279;
w35281 <= not w35278 and w35280;
w35282 <= not pi0609 and w35276;
w35283 <= pi0609 and not w35022;
w35284 <= not pi1155 and not w35283;
w35285 <= not w35282 and w35284;
w35286 <= not w35281 and not w35285;
w35287 <= pi0785 and not w35286;
w35288 <= not w35277 and not w35287;
w35289 <= not pi0781 and not w35288;
w35290 <= pi0618 and w35288;
w35291 <= not pi0618 and not w35022;
w35292 <= pi1154 and not w35291;
w35293 <= not w35290 and w35292;
w35294 <= not pi0618 and w35288;
w35295 <= pi0618 and not w35022;
w35296 <= not pi1154 and not w35295;
w35297 <= not w35294 and w35296;
w35298 <= not w35293 and not w35297;
w35299 <= pi0781 and not w35298;
w35300 <= not w35289 and not w35299;
w35301 <= not pi0789 and not w35300;
w35302 <= pi0619 and w35300;
w35303 <= not pi0619 and not w35022;
w35304 <= pi1159 and not w35303;
w35305 <= not w35302 and w35304;
w35306 <= not pi0619 and w35300;
w35307 <= pi0619 and not w35022;
w35308 <= not pi1159 and not w35307;
w35309 <= not w35306 and w35308;
w35310 <= not w35305 and not w35309;
w35311 <= pi0789 and not w35310;
w35312 <= not w35301 and not w35311;
w35313 <= not w15532 and w35312;
w35314 <= not w35152 and not w35313;
w35315 <= not w18133 and w35314;
w35316 <= not pi0628 and not w35022;
w35317 <= pi0628 and not w35131;
w35318 <= w15339 and not w35316;
w35319 <= not w35317 and w35318;
w35320 <= not w35151 and not w35319;
w35321 <= not w35315 and w35320;
w35322 <= pi0792 and not w35321;
w35323 <= pi0609 and w35122;
w35324 <= pi0662 and w14918;
w35325 <= w14204 and w35324;
w35326 <= w35154 and not w35325;
w35327 <= w15180 and w35029;
w35328 <= not w35155 and not w35327;
w35329 <= not pi0224 and not w35328;
w35330 <= w15180 and not w35029;
w35331 <= not w34291 and w35158;
w35332 <= not w35330 and w35331;
w35333 <= not w35329 and not w35332;
w35334 <= not pi0299 and not w35333;
w35335 <= not w35029 and w35166;
w35336 <= not pi0614 and w14794;
w35337 <= not w34301 and not w35336;
w35338 <= pi0224 and not w35337;
w35339 <= not pi0224 and not w15185;
w35340 <= not w35162 and w35339;
w35341 <= not w35338 and not w35340;
w35342 <= w35029 and not w35341;
w35343 <= pi0299 and not w35335;
w35344 <= not w35342 and w35343;
w35345 <= not w35334 and not w35344;
w35346 <= not pi0039 and not w35345;
w35347 <= w14970 and w35029;
w35348 <= not w35199 and not w35347;
w35349 <= not pi0224 and not w35348;
w35350 <= not pi0222 and w35349;
w35351 <= not w14970 and w35202;
w35352 <= not w34183 and not w35351;
w35353 <= pi0680 and not w35352;
w35354 <= not w34238 and not w35199;
w35355 <= not w35353 and not w35354;
w35356 <= pi0662 and not w35355;
w35357 <= not pi0662 and not w35236;
w35358 <= not w35356 and not w35357;
w35359 <= w3768 and not w35358;
w35360 <= not pi0662 and not w14219;
w35361 <= not w35229 and w35360;
w35362 <= not pi0614 and w14997;
w35363 <= pi0614 and not w15141;
w35364 <= pi0680 and not w35363;
w35365 <= not w35362 and w35364;
w35366 <= not w35230 and not w35365;
w35367 <= pi0662 and not w35366;
w35368 <= not w35232 and not w35361;
w35369 <= not w35367 and w35368;
w35370 <= not w3768 and not w35369;
w35371 <= w3373 and not w35359;
w35372 <= not w35370 and w35371;
w35373 <= not w35219 and w35360;
w35374 <= not pi0614 and not w21618;
w35375 <= pi0614 and not w34125;
w35376 <= not w35374 and not w35375;
w35377 <= not w14213 and w35376;
w35378 <= pi0616 and not w35377;
w35379 <= pi0614 and not w15067;
w35380 <= not w14924 and not w35379;
w35381 <= not pi0616 and not w35380;
w35382 <= not w35378 and not w35381;
w35383 <= pi0680 and not w35382;
w35384 <= not w35221 and not w35383;
w35385 <= pi0662 and not w35384;
w35386 <= not w35224 and not w35373;
w35387 <= not w35385 and w35386;
w35388 <= w3768 and w35387;
w35389 <= not w35208 and w35360;
w35390 <= pi0614 and not w34201;
w35391 <= w34196 and w35202;
w35392 <= not w35390 and not w35391;
w35393 <= not w34199 and w35392;
w35394 <= pi0680 and not w35393;
w35395 <= not w35210 and not w35394;
w35396 <= pi0662 and not w35395;
w35397 <= not w35216 and not w35389;
w35398 <= not w35396 and w35397;
w35399 <= not w3768 and w35398;
w35400 <= pi0224 and not w35399;
w35401 <= not w35388 and w35400;
w35402 <= not pi0223 and not w35350;
w35403 <= not w35372 and w35402;
w35404 <= not w35401 and w35403;
w35405 <= pi0680 and not w15008;
w35406 <= not w35199 and not w35405;
w35407 <= not w35353 and not w35406;
w35408 <= pi0662 and not w35407;
w35409 <= not pi0662 and not w35170;
w35410 <= not w35408 and not w35409;
w35411 <= not pi0224 and not w35410;
w35412 <= not w35186 and w35360;
w35413 <= not w14908 and not w35379;
w35414 <= not pi0616 and not w35413;
w35415 <= not w35378 and not w35414;
w35416 <= pi0680 and not w35415;
w35417 <= not w35188 and not w35416;
w35418 <= pi0662 and not w35417;
w35419 <= not w35192 and not w35412;
w35420 <= not w35418 and w35419;
w35421 <= pi0224 and w35420;
w35422 <= w3768 and not w35411;
w35423 <= not w35421 and w35422;
w35424 <= not w35174 and w35360;
w35425 <= pi0614 and not w34151;
w35426 <= w14893 and not w35425;
w35427 <= pi0680 and not w35426;
w35428 <= not w35175 and not w35427;
w35429 <= pi0662 and not w35428;
w35430 <= not w35179 and not w35424;
w35431 <= not w35429 and w35430;
w35432 <= pi0224 and w35431;
w35433 <= not w14286 and w35170;
w35434 <= not pi0662 and not w35433;
w35435 <= pi0614 and not pi0680;
w35436 <= w14800 and w35435;
w35437 <= pi0614 and w34170;
w35438 <= not pi0614 and w15014;
w35439 <= pi0680 and not w35437;
w35440 <= not w35438 and w35439;
w35441 <= not w15020 and w35440;
w35442 <= pi0662 and not w35436;
w35443 <= not w35441 and w35442;
w35444 <= not w35434 and not w35443;
w35445 <= not pi0224 and not w35444;
w35446 <= not w3768 and not w35445;
w35447 <= not w35432 and w35446;
w35448 <= pi0223 and not w35447;
w35449 <= not w35423 and w35448;
w35450 <= not w35404 and not w35449;
w35451 <= not pi0299 and not w35450;
w35452 <= not w3805 and not w35431;
w35453 <= w3805 and not w35420;
w35454 <= pi0224 and not w35452;
w35455 <= not w35453 and w35454;
w35456 <= w3805 and w35410;
w35457 <= not w3805 and w35444;
w35458 <= not pi0224 and not w35457;
w35459 <= not w35456 and w35458;
w35460 <= pi0215 and not w35459;
w35461 <= not w35455 and w35460;
w35462 <= w35029 and w35376;
w35463 <= not w35029 and not w35183;
w35464 <= w14230 and w35463;
w35465 <= pi0224 and not w35464;
w35466 <= not w35462 and w35465;
w35467 <= w35080 and not w35466;
w35468 <= not w35349 and w35467;
w35469 <= not pi0224 and not w35358;
w35470 <= pi0224 and w35387;
w35471 <= w3805 and not w35469;
w35472 <= not w35470 and w35471;
w35473 <= not pi0224 and not w35369;
w35474 <= pi0224 and w35398;
w35475 <= not w3805 and not w35473;
w35476 <= not w35474 and w35475;
w35477 <= not w1011 and not w35472;
w35478 <= not w35476 and w35477;
w35479 <= not pi0215 and not w35468;
w35480 <= not w35478 and w35479;
w35481 <= pi0299 and not w35461;
w35482 <= not w35480 and w35481;
w35483 <= pi0039 and not w35451;
w35484 <= not w35482 and w35483;
w35485 <= not pi0038 and not w35346;
w35486 <= not w35484 and w35485;
w35487 <= w134 and not w35326;
w35488 <= not w35486 and w35487;
w35489 <= not w35024 and not w35488;
w35490 <= not pi0625 and w35489;
w35491 <= pi0625 and w35273;
w35492 <= not pi1153 and not w35491;
w35493 <= not w35490 and w35492;
w35494 <= not pi0608 and not w35115;
w35495 <= not w35493 and w35494;
w35496 <= not pi0625 and w35273;
w35497 <= pi0625 and w35489;
w35498 <= pi1153 and not w35496;
w35499 <= not w35497 and w35498;
w35500 <= pi0608 and not w35119;
w35501 <= not w35499 and w35500;
w35502 <= not w35495 and not w35501;
w35503 <= pi0778 and not w35502;
w35504 <= not pi0778 and w35489;
w35505 <= not w35503 and not w35504;
w35506 <= not pi0609 and not w35505;
w35507 <= not pi1155 and not w35323;
w35508 <= not w35506 and w35507;
w35509 <= not pi0660 and not w35281;
w35510 <= not w35508 and w35509;
w35511 <= not pi0609 and w35122;
w35512 <= pi0609 and not w35505;
w35513 <= pi1155 and not w35511;
w35514 <= not w35512 and w35513;
w35515 <= pi0660 and not w35285;
w35516 <= not w35514 and w35515;
w35517 <= not w35510 and not w35516;
w35518 <= pi0785 and not w35517;
w35519 <= not pi0785 and not w35505;
w35520 <= not w35518 and not w35519;
w35521 <= not pi0618 and not w35520;
w35522 <= pi0618 and w35125;
w35523 <= not pi1154 and not w35522;
w35524 <= not w35521 and w35523;
w35525 <= not pi0627 and not w35293;
w35526 <= not w35524 and w35525;
w35527 <= not pi0618 and w35125;
w35528 <= pi0618 and not w35520;
w35529 <= pi1154 and not w35527;
w35530 <= not w35528 and w35529;
w35531 <= pi0627 and not w35297;
w35532 <= not w35530 and w35531;
w35533 <= not w35526 and not w35532;
w35534 <= pi0781 and not w35533;
w35535 <= not pi0781 and not w35520;
w35536 <= not w35534 and not w35535;
w35537 <= not pi0789 and w35536;
w35538 <= not pi0619 and not w35536;
w35539 <= pi0619 and w35128;
w35540 <= not pi1159 and not w35539;
w35541 <= not w35538 and w35540;
w35542 <= not pi0648 and not w35305;
w35543 <= not w35541 and w35542;
w35544 <= pi0619 and not w35536;
w35545 <= not pi0619 and w35128;
w35546 <= pi1159 and not w35545;
w35547 <= not w35544 and w35546;
w35548 <= pi0648 and not w35309;
w35549 <= not w35547 and w35548;
w35550 <= pi0789 and not w35543;
w35551 <= not w35549 and w35550;
w35552 <= w15533 and not w35537;
w35553 <= not w35551 and w35552;
w35554 <= w14198 and not w35022;
w35555 <= not w35129 and not w35554;
w35556 <= w15434 and not w35555;
w35557 <= not pi0626 and w35022;
w35558 <= pi0626 and not w35312;
w35559 <= w14191 and not w35557;
w35560 <= not w35558 and w35559;
w35561 <= pi0626 and w35022;
w35562 <= not pi0626 and not w35312;
w35563 <= w14192 and not w35561;
w35564 <= not w35562 and w35563;
w35565 <= not w35556 and not w35560;
w35566 <= not w35564 and w35565;
w35567 <= pi0788 and not w35566;
w35568 <= not w17927 and not w35567;
w35569 <= not w35553 and w35568;
w35570 <= not w35322 and not w35569;
w35571 <= not w17769 and not w35570;
w35572 <= not pi0630 and w35143;
w35573 <= not w15342 and w35314;
w35574 <= w15342 and w35022;
w35575 <= not w35573 and not w35574;
w35576 <= not w18122 and not w35575;
w35577 <= pi0630 and w35139;
w35578 <= not w35572 and not w35577;
w35579 <= not w35576 and w35578;
w35580 <= pi0787 and not w35579;
w35581 <= not w35571 and not w35580;
w35582 <= pi0644 and w35581;
w35583 <= pi0715 and not w35147;
w35584 <= not w35582 and w35583;
w35585 <= w15367 and not w35022;
w35586 <= not w15367 and w35575;
w35587 <= not w35585 and not w35586;
w35588 <= pi0644 and not w35587;
w35589 <= not pi0644 and not w35022;
w35590 <= not pi0715 and not w35589;
w35591 <= not w35588 and w35590;
w35592 <= pi1160 and not w35591;
w35593 <= not w35584 and w35592;
w35594 <= pi0644 and w35146;
w35595 <= not pi0644 and w35581;
w35596 <= not pi0715 and not w35594;
w35597 <= not w35595 and w35596;
w35598 <= not pi0644 and not w35587;
w35599 <= pi0644 and not w35022;
w35600 <= pi0715 and not w35599;
w35601 <= not w35598 and w35600;
w35602 <= not pi1160 and not w35601;
w35603 <= not w35597 and w35602;
w35604 <= not w35593 and not w35603;
w35605 <= pi0790 and not w35604;
w35606 <= not pi0790 and w35581;
w35607 <= not w35605 and not w35606;
w35608 <= w4989 and not w35607;
w35609 <= not pi0224 and not w4989;
w35610 <= not w35608 and not w35609;
w35611 <= w110 and w188;
w35612 <= w893 and w35611;
w35613 <= not pi0062 and w35612;
w35614 <= not w891 and not w35613;
w35615 <= pi0062 and w35612;
w35616 <= w97 and w35611;
w35617 <= pi0054 and not w35616;
w35618 <= pi0092 and w96;
w35619 <= w35611 and w35618;
w35620 <= not w3732 and w3826;
w35621 <= not pi0137 and not w35620;
w35622 <= w4864 and not w35621;
w35623 <= pi0075 and not w35622;
w35624 <= pi0087 and w35611;
w35625 <= w3849 and not w35621;
w35626 <= pi0038 and not pi0137;
w35627 <= pi0039 and w110;
w35628 <= not w304 and not w542;
w35629 <= pi0137 and not w35628;
w35630 <= not w303 and not w35629;
w35631 <= not pi0332 and not w35630;
w35632 <= w80 and w8980;
w35633 <= w301 and not w35632;
w35634 <= not pi0137 and w276;
w35635 <= not w35633 and w35634;
w35636 <= w731 and not w8980;
w35637 <= not w466 and w35636;
w35638 <= w309 and not w35637;
w35639 <= w307 and not w35638;
w35640 <= not w275 and not w35639;
w35641 <= not pi0095 and not w35640;
w35642 <= w651 and not w35641;
w35643 <= pi0332 and not w35635;
w35644 <= not w35642 and w35643;
w35645 <= not w35631 and not w35644;
w35646 <= pi0210 and not w35645;
w35647 <= w485 and not w35633;
w35648 <= pi1093 and not w35647;
w35649 <= w485 and w496;
w35650 <= w80 and not w5018;
w35651 <= not w523 and w35650;
w35652 <= not pi0032 and not w35651;
w35653 <= w35649 and not w35652;
w35654 <= not pi1093 and not w35653;
w35655 <= not w496 and w35647;
w35656 <= w8979 and w35650;
w35657 <= w35649 and w35656;
w35658 <= not w35655 and not w35657;
w35659 <= w35654 and w35658;
w35660 <= not w35648 and not w35659;
w35661 <= w9112 and not w35660;
w35662 <= not w484 and not w35639;
w35663 <= not pi0095 and not w35662;
w35664 <= not w304 and not w35663;
w35665 <= pi0137 and not w35664;
w35666 <= not w496 and w586;
w35667 <= w35654 and not w35666;
w35668 <= not w560 and w35650;
w35669 <= not pi0032 and not w35668;
w35670 <= w35649 and not w35669;
w35671 <= pi1093 and not w35666;
w35672 <= not w35670 and w35671;
w35673 <= not w35667 and not w35672;
w35674 <= w9080 and not w35673;
w35675 <= w35658 and w35674;
w35676 <= not w35661 and not w35675;
w35677 <= not w35665 and w35676;
w35678 <= pi0332 and not w35677;
w35679 <= not w304 and not w549;
w35680 <= pi0137 and not w35679;
w35681 <= pi1093 and not w586;
w35682 <= not w35667 and not w35681;
w35683 <= w9112 and not w35682;
w35684 <= not w35674 and not w35683;
w35685 <= not w35680 and w35684;
w35686 <= not pi0332 and not w35685;
w35687 <= not w35678 and not w35686;
w35688 <= not w203 and w35687;
w35689 <= not pi0137 and not w35647;
w35690 <= not w35665 and not w35689;
w35691 <= pi0332 and not w35690;
w35692 <= not w587 and not w35680;
w35693 <= not pi0332 and not w35692;
w35694 <= not w35691 and not w35693;
w35695 <= w203 and w35694;
w35696 <= not pi0210 and not w35688;
w35697 <= not w35695 and w35696;
w35698 <= pi0299 and not w35646;
w35699 <= not w35697 and w35698;
w35700 <= pi0198 and not w35645;
w35701 <= w3823 and w35694;
w35702 <= not w3823 and w35687;
w35703 <= not pi0198 and not w35701;
w35704 <= not w35702 and w35703;
w35705 <= not pi0299 and not w35700;
w35706 <= not w35704 and w35705;
w35707 <= not w35699 and not w35706;
w35708 <= not pi0039 and not w35707;
w35709 <= not pi0038 and not w35627;
w35710 <= not w35708 and w35709;
w35711 <= w3700 and not w35626;
w35712 <= not w35710 and w35711;
w35713 <= not w35625 and not w35712;
w35714 <= not pi0087 and not w35713;
w35715 <= not pi0075 and not w35624;
w35716 <= not w35714 and w35715;
w35717 <= not pi0092 and not w35623;
w35718 <= not w35716 and w35717;
w35719 <= not pi0054 and not w35619;
w35720 <= not w35718 and w35719;
w35721 <= not pi0074 and not w35617;
w35722 <= not w35720 and w35721;
w35723 <= pi0074 and w3691;
w35724 <= w35611 and w35723;
w35725 <= not pi0055 and not w35724;
w35726 <= not w35722 and w35725;
w35727 <= w4911 and not w35726;
w35728 <= pi0056 and w99;
w35729 <= w35611 and w35728;
w35730 <= not w35727 and not w35729;
w35731 <= not pi0062 and not w35730;
w35732 <= w891 and not w35615;
w35733 <= not w35731 and w35732;
w35734 <= not w3683 and not w35614;
w35735 <= not w35733 and w35734;
w35736 <= pi0228 and pi0231;
w35737 <= not w4923 and not w35736;
w35738 <= pi0056 and not w35737;
w35739 <= pi0055 and not w35736;
w35740 <= not w4927 and not w35736;
w35741 <= pi0074 and not w35740;
w35742 <= pi0054 and not w35736;
w35743 <= not w11534 and not w35736;
w35744 <= pi0075 and not w35743;
w35745 <= pi0087 and not w35736;
w35746 <= not w4919 and w35745;
w35747 <= not w11538 and not w35736;
w35748 <= pi0100 and not w35747;
w35749 <= not w293 and not w686;
w35750 <= not pi0070 and not w35749;
w35751 <= not pi0051 and not w35750;
w35752 <= w311 and not w35751;
w35753 <= w731 and not w35752;
w35754 <= w309 and not w35753;
w35755 <= w307 and not w35754;
w35756 <= not w3739 and not w35755;
w35757 <= not pi0095 and not w35756;
w35758 <= w305 and not w35757;
w35759 <= not pi0039 and not w35758;
w35760 <= not pi0038 and not w965;
w35761 <= not w35759 and w35760;
w35762 <= not pi0228 and w35761;
w35763 <= not w35736 and not w35762;
w35764 <= not pi0100 and not w35763;
w35765 <= not pi0087 and not w35748;
w35766 <= not w35764 and w35765;
w35767 <= not pi0075 and not w35746;
w35768 <= not w35766 and w35767;
w35769 <= not pi0092 and not w35744;
w35770 <= not w35768 and w35769;
w35771 <= pi0092 and not w35736;
w35772 <= not w4932 and w35771;
w35773 <= not w35770 and not w35772;
w35774 <= not pi0054 and not w35773;
w35775 <= not pi0074 and not w35742;
w35776 <= not w35774 and w35775;
w35777 <= not pi0055 and not w35741;
w35778 <= not w35776 and w35777;
w35779 <= not pi0056 and not w35739;
w35780 <= not w35778 and w35779;
w35781 <= not pi0062 and not w35738;
w35782 <= not w35780 and w35781;
w35783 <= pi0062 and not w35736;
w35784 <= not w4920 and w35783;
w35785 <= not w35782 and not w35784;
w35786 <= w891 and not w35785;
w35787 <= not w891 and not w35736;
w35788 <= not w35786 and not w35787;
w35789 <= w10643 and not w10679;
w35790 <= w4043 and w35789;
w35791 <= not w3958 and not w35790;
w35792 <= pi1093 and not w35791;
w35793 <= w271 and w3983;
w35794 <= not pi0091 and not w324;
w35795 <= w35793 and not w35794;
w35796 <= not pi0072 and not w35795;
w35797 <= w8585 and w35793;
w35798 <= not w4980 and w35797;
w35799 <= not w6466 and w35796;
w35800 <= not w35798 and w35799;
w35801 <= w4043 and not w35800;
w35802 <= not w35792 and not w35801;
w35803 <= w35796 and not w35797;
w35804 <= w4043 and not w35803;
w35805 <= w7637 and not w35804;
w35806 <= not w495 and w8585;
w35807 <= w317 and w8594;
w35808 <= w8592 and w35807;
w35809 <= w35794 and not w35806;
w35810 <= not w35808 and w35809;
w35811 <= w35793 and not w35810;
w35812 <= not pi0072 and not w35811;
w35813 <= w4043 and not w35812;
w35814 <= pi0829 and not w3778;
w35815 <= not w35813 and w35814;
w35816 <= not w35802 and not w35805;
w35817 <= not w35815 and w35816;
w35818 <= not pi0039 and not w35817;
w35819 <= w9034 and not w35818;
w35820 <= not pi0039 and pi0228;
w35821 <= not w8983 and not w8988;
w35822 <= pi0039 and not w35821;
w35823 <= w3954 and w35822;
w35824 <= not w493 and not w6467;
w35825 <= not pi0032 and w7798;
w35826 <= not w35824 and w35825;
w35827 <= w530 and w35826;
w35828 <= not w9050 and w35827;
w35829 <= not w35823 and not w35828;
w35830 <= w7763 and not w35829;
w35831 <= not w35820 and not w35830;
w35832 <= not w3699 and w7760;
w35833 <= pi0120 and w3781;
w35834 <= w14215 and not w35833;
w35835 <= not w33240 and not w35834;
w35836 <= not w3768 and not w35835;
w35837 <= not w3761 and w14215;
w35838 <= not w35834 and not w35837;
w35839 <= w3768 and not w35838;
w35840 <= pi0223 and not w35836;
w35841 <= not w35839 and w35840;
w35842 <= w166 and w14215;
w35843 <= not w3776 and w5080;
w35844 <= w14224 and w35843;
w35845 <= w14212 and not w35843;
w35846 <= pi1091 and not w35844;
w35847 <= not w35845 and w35846;
w35848 <= w3946 and w14224;
w35849 <= not w3946 and w14212;
w35850 <= not pi1091 and not w35848;
w35851 <= not w35849 and w35850;
w35852 <= not w35847 and not w35851;
w35853 <= not pi0120 and not w35852;
w35854 <= not w14214 and not w35853;
w35855 <= not w3790 and w35854;
w35856 <= not w33240 and not w35855;
w35857 <= not w3768 and w35856;
w35858 <= w3761 and w35854;
w35859 <= not w35837 and not w35858;
w35860 <= w3768 and w35859;
w35861 <= not w166 and not w35857;
w35862 <= not w35860 and w35861;
w35863 <= not pi0223 and not w35842;
w35864 <= not w35862 and w35863;
w35865 <= not pi0299 and not w35841;
w35866 <= not w35864 and w35865;
w35867 <= not w3805 and not w35835;
w35868 <= w3805 and not w35838;
w35869 <= pi0215 and not w35867;
w35870 <= not w35868 and w35869;
w35871 <= not w3805 and w35856;
w35872 <= w3805 and w35859;
w35873 <= not w1011 and not w35871;
w35874 <= not w35872 and w35873;
w35875 <= not pi0215 and not w14388;
w35876 <= not w35874 and w35875;
w35877 <= pi0299 and not w35870;
w35878 <= not w35876 and w35877;
w35879 <= not w35866 and not w35878;
w35880 <= pi0039 and not w35879;
w35881 <= w3733 and w14417;
w35882 <= not w14419 and w35881;
w35883 <= not pi0040 and not w35882;
w35884 <= w7852 and not w35883;
w35885 <= pi0252 and not w35884;
w35886 <= w3840 and not w14416;
w35887 <= not w35885 and w35886;
w35888 <= not w3840 and w14429;
w35889 <= not pi1093 and not w35887;
w35890 <= not w35888 and w35889;
w35891 <= not w3732 and not w3950;
w35892 <= not w4980 and w14429;
w35893 <= not w14446 and not w35892;
w35894 <= w35891 and not w35893;
w35895 <= pi0829 and pi1091;
w35896 <= w14470 and w35895;
w35897 <= not pi0824 and not w35896;
w35898 <= pi0824 and not w14465;
w35899 <= not w3950 and not w35897;
w35900 <= not w35898 and w35899;
w35901 <= not w14429 and not w35900;
w35902 <= w35895 and w35897;
w35903 <= not w35898 and not w35902;
w35904 <= w495 and not w3950;
w35905 <= not w35903 and w35904;
w35906 <= not w35891 and not w35901;
w35907 <= not w35905 and w35906;
w35908 <= pi1093 and not w35894;
w35909 <= not w35907 and w35908;
w35910 <= not pi0039 and not w35890;
w35911 <= not w35909 and w35910;
w35912 <= not pi0038 and not w35880;
w35913 <= not w35911 and w35912;
w35914 <= w35832 and not w35913;
w35915 <= not pi0081 and not w428;
w35916 <= w4006 and not w35915;
w35917 <= w25 and not w35916;
w35918 <= w436 and not w35917;
w35919 <= w348 and not w35918;
w35920 <= w440 and not w35919;
w35921 <= w282 and not w35920;
w35922 <= not w285 and not w35921;
w35923 <= not pi0086 and not w35922;
w35924 <= w346 and not w35923;
w35925 <= w344 and not w35924;
w35926 <= not w339 and not w35925;
w35927 <= not pi0108 and not w35926;
w35928 <= w338 and not w35927;
w35929 <= w452 and not w35928;
w35930 <= not w329 and not w35929;
w35931 <= w328 and not w35930;
w35932 <= w327 and not w35931;
w35933 <= w320 and not w35932;
w35934 <= w671 and not w35933;
w35935 <= w67 and not w35934;
w35936 <= w13198 and not w35935;
w35937 <= not pi0070 and not w35936;
w35938 <= not w662 and not w35937;
w35939 <= not pi0051 and not w35938;
w35940 <= w311 and not w35939;
w35941 <= w731 and not w35940;
w35942 <= w309 and not w35941;
w35943 <= not pi1082 and w306;
w35944 <= not pi0032 and not w35943;
w35945 <= not w35942 and w35944;
w35946 <= not w975 and not w35945;
w35947 <= not pi0095 and not w35946;
w35948 <= not w304 and not w35947;
w35949 <= not pi0039 and not w35948;
w35950 <= not w4870 and not w4872;
w35951 <= w495 and w3780;
w35952 <= w3944 and w35951;
w35953 <= not w35950 and w35952;
w35954 <= w3748 and w8932;
w35955 <= not w35953 and w35954;
w35956 <= not w965 and not w35955;
w35957 <= not w35949 and w35956;
w35958 <= not pi0038 and not w35957;
w35959 <= w3700 and not w35958;
w35960 <= not pi0087 and not w3849;
w35961 <= not w35959 and w35960;
w35962 <= not w3695 and not w35961;
w35963 <= w132 and not w35962;
w35964 <= w4869 and not w35963;
w35965 <= not pi0054 and not w35964;
w35966 <= not w4904 and not w35965;
w35967 <= w6442 and not w35966;
w35968 <= w13275 and not w35967;
w35969 <= not pi0056 and not w35968;
w35970 <= not w3690 and not w35969;
w35971 <= not pi0062 and not w35970;
w35972 <= not w3862 and not w35971;
w35973 <= w891 and not w35972;
w35974 <= w3686 and not w35973;
w35975 <= not pi0230 and not pi0233;
w35976 <= not pi0212 and not pi0214;
w35977 <= not pi0211 and not w35976;
w35978 <= pi0219 and not w35977;
w35979 <= not w4989 and not w35978;
w35980 <= pi1142 and not w8049;
w35981 <= pi0211 and pi1143;
w35982 <= not pi0211 and pi1144;
w35983 <= not w35981 and not w35982;
w35984 <= not pi0212 and pi0214;
w35985 <= pi0212 and not pi0214;
w35986 <= not w35984 and not w35985;
w35987 <= not w35983 and not w35986;
w35988 <= not pi0211 and pi1143;
w35989 <= w8406 and w35988;
w35990 <= not w35987 and not w35989;
w35991 <= not pi0219 and not w35990;
w35992 <= not w35980 and not w35991;
w35993 <= w35979 and not w35992;
w35994 <= pi0299 and not w35983;
w35995 <= pi0199 and pi1142;
w35996 <= not pi0200 and not w35995;
w35997 <= not pi0199 and pi1144;
w35998 <= w35996 and not w35997;
w35999 <= not pi0199 and pi1143;
w36000 <= pi0200 and not w35999;
w36001 <= not w35998 and not w36000;
w36002 <= not pi0299 and not w36001;
w36003 <= not pi0207 and not w36002;
w36004 <= pi0207 and not pi0299;
w36005 <= w35996 and not w35999;
w36006 <= not pi0199 and pi1142;
w36007 <= pi0200 and not w36006;
w36008 <= w36004 and not w36007;
w36009 <= not w36005 and w36008;
w36010 <= not w36003 and not w36009;
w36011 <= pi0208 and not w36010;
w36012 <= pi0207 and not pi0208;
w36013 <= w36001 and w36012;
w36014 <= not w36011 and not w36013;
w36015 <= not pi0299 and not w36014;
w36016 <= not pi0214 and not w36015;
w36017 <= not w35994 and w36016;
w36018 <= pi0211 and pi1142;
w36019 <= not w35988 and not w36018;
w36020 <= pi0299 and not w36019;
w36021 <= pi0214 and not w36020;
w36022 <= not w36015 and w36021;
w36023 <= pi0212 and not w36022;
w36024 <= not w36017 and w36023;
w36025 <= not w35994 and not w36015;
w36026 <= not pi0212 and not w36016;
w36027 <= not w36025 and w36026;
w36028 <= not pi0219 and not w36024;
w36029 <= not w36027 and w36028;
w36030 <= not w35977 and w36015;
w36031 <= not pi0299 and w36014;
w36032 <= pi0299 and not pi1142;
w36033 <= w35977 and not w36032;
w36034 <= not w36031 and w36033;
w36035 <= pi0219 and not w36030;
w36036 <= not w36034 and w36035;
w36037 <= w4989 and not w36036;
w36038 <= not w36029 and w36037;
w36039 <= not w35993 and not w36038;
w36040 <= pi0213 and w36039;
w36041 <= not pi0211 and pi1157;
w36042 <= pi0211 and pi1156;
w36043 <= not w36041 and not w36042;
w36044 <= pi0214 and not w36043;
w36045 <= not pi0212 and not w36044;
w36046 <= not pi0211 and pi1156;
w36047 <= pi0211 and pi1155;
w36048 <= not w36046 and not w36047;
w36049 <= not pi0214 and not w36048;
w36050 <= not pi0211 and pi1155;
w36051 <= pi0211 and pi1154;
w36052 <= not w36050 and not w36051;
w36053 <= pi0214 and not w36052;
w36054 <= not w36049 and not w36053;
w36055 <= pi0212 and w36054;
w36056 <= not w36045 and not w36055;
w36057 <= not pi0219 and not w36056;
w36058 <= not pi0211 and pi1154;
w36059 <= not pi0214 and not w36058;
w36060 <= not pi0211 and pi1153;
w36061 <= w8406 and not w36060;
w36062 <= not pi0211 and pi0214;
w36063 <= pi1155 and w36062;
w36064 <= not pi0212 and not w36063;
w36065 <= not w36059 and not w36061;
w36066 <= not w36064 and w36065;
w36067 <= pi0219 and not w36066;
w36068 <= not w4989 and not w36067;
w36069 <= not w36057 and w36068;
w36070 <= not pi0213 and not w36069;
w36071 <= not pi0219 and pi0299;
w36072 <= w36056 and w36071;
w36073 <= pi0299 and pi1155;
w36074 <= w35984 and w36073;
w36075 <= pi0299 and pi1153;
w36076 <= pi0214 and not w36075;
w36077 <= pi0299 and pi1154;
w36078 <= not pi0214 and not w36077;
w36079 <= pi0212 and not w36076;
w36080 <= not w36078 and w36079;
w36081 <= not w36074 and not w36080;
w36082 <= not pi0211 and pi0219;
w36083 <= not w36081 and w36082;
w36084 <= not w36072 and not w36083;
w36085 <= not w36015 and w36084;
w36086 <= w4989 and not w36085;
w36087 <= w36070 and not w36086;
w36088 <= pi0209 and not w36087;
w36089 <= not w36040 and w36088;
w36090 <= not pi0211 and w8406;
w36091 <= pi0299 and not pi1143;
w36092 <= not pi0200 and pi1155;
w36093 <= pi0199 and w36092;
w36094 <= not pi0299 and w36093;
w36095 <= not pi1156 and not w36094;
w36096 <= not pi0299 and not w9007;
w36097 <= pi1156 and not w36093;
w36098 <= w36096 and w36097;
w36099 <= not w36095 and not w36098;
w36100 <= pi0207 and w36099;
w36101 <= not pi0299 and not w36100;
w36102 <= not pi0208 and not w36101;
w36103 <= not pi1157 and w36102;
w36104 <= not w36091 and w36103;
w36105 <= not pi0208 and pi1157;
w36106 <= pi0299 and pi1143;
w36107 <= not pi1155 and not w8373;
w36108 <= pi0200 and not pi0299;
w36109 <= pi1155 and not w36108;
w36110 <= not w36107 and not w36109;
w36111 <= pi0199 and not pi1155;
w36112 <= pi0199 and pi0200;
w36113 <= not pi0299 and not w36112;
w36114 <= pi1156 and not w36111;
w36115 <= w36113 and w36114;
w36116 <= w36110 and not w36115;
w36117 <= pi0207 and not w36091;
w36118 <= not w36116 and w36117;
w36119 <= not w36106 and not w36118;
w36120 <= w36105 and not w36119;
w36121 <= pi1153 and not w36113;
w36122 <= pi1154 and not w36121;
w36123 <= w8947 and w36092;
w36124 <= not w8372 and not w36112;
w36125 <= not pi1153 and not w8947;
w36126 <= pi1154 and w36124;
w36127 <= not w36125 and w36126;
w36128 <= not w36123 and not w36127;
w36129 <= w36122 and not w36128;
w36130 <= not pi0199 and not pi1155;
w36131 <= not pi0200 and not pi0299;
w36132 <= pi0199 and not pi1153;
w36133 <= w36131 and not w36132;
w36134 <= not pi1154 and not w36130;
w36135 <= w36133 and w36134;
w36136 <= not w36129 and not w36135;
w36137 <= pi0207 and w36136;
w36138 <= not w36106 and w36137;
w36139 <= not pi0199 and pi1155;
w36140 <= w36108 and w36139;
w36141 <= not pi1154 and not w36140;
w36142 <= not w36106 and w36141;
w36143 <= not pi1155 and w36106;
w36144 <= not pi0299 and not w36124;
w36145 <= pi1155 and not w36144;
w36146 <= not w36091 and w36145;
w36147 <= not pi0200 and not pi1155;
w36148 <= w8936 and w36147;
w36149 <= pi1154 and not w36148;
w36150 <= not w36143 and w36149;
w36151 <= not w36146 and w36150;
w36152 <= not pi1156 and not w36142;
w36153 <= not w36151 and w36152;
w36154 <= pi0200 and not w36139;
w36155 <= not pi0299 and not w36154;
w36156 <= pi1154 and not w36155;
w36157 <= not w36106 and w36156;
w36158 <= pi1155 and not w8936;
w36159 <= not w36107 and not w36158;
w36160 <= not w36091 and not w36159;
w36161 <= not pi1154 and not w36160;
w36162 <= pi1156 and not w36157;
w36163 <= not w36161 and w36162;
w36164 <= not w36153 and not w36163;
w36165 <= not pi0207 and w36164;
w36166 <= pi0208 and not w36138;
w36167 <= not w36165 and w36166;
w36168 <= not w36104 and not w36120;
w36169 <= not w36167 and w36168;
w36170 <= w36090 and w36169;
w36171 <= not w8406 and not w35976;
w36172 <= pi0211 and not w36169;
w36173 <= pi0299 and not pi1144;
w36174 <= w36103 and not w36173;
w36175 <= pi0299 and pi1144;
w36176 <= pi0207 and not w36173;
w36177 <= not w36116 and w36176;
w36178 <= not w36175 and not w36177;
w36179 <= w36105 and not w36178;
w36180 <= w36137 and not w36175;
w36181 <= w36141 and not w36175;
w36182 <= not pi1155 and w36175;
w36183 <= w36145 and not w36173;
w36184 <= w36149 and not w36182;
w36185 <= not w36183 and w36184;
w36186 <= not pi1156 and not w36181;
w36187 <= not w36185 and w36186;
w36188 <= w36156 and not w36175;
w36189 <= not w36159 and not w36173;
w36190 <= not pi1154 and not w36189;
w36191 <= pi1156 and not w36188;
w36192 <= not w36190 and w36191;
w36193 <= not w36187 and not w36192;
w36194 <= not pi0207 and w36193;
w36195 <= pi0208 and not w36180;
w36196 <= not w36194 and w36195;
w36197 <= not w36174 and not w36179;
w36198 <= not w36196 and w36197;
w36199 <= not pi0211 and not w36198;
w36200 <= w36171 and not w36172;
w36201 <= not w36199 and w36200;
w36202 <= not w36170 and not w36201;
w36203 <= not pi0219 and not w36202;
w36204 <= not pi0299 and w36124;
w36205 <= not w36147 and w36204;
w36206 <= not w36095 and w36205;
w36207 <= pi0207 and w36206;
w36208 <= not pi0208 and not w36207;
w36209 <= w8373 and not w36154;
w36210 <= not w36141 and w36209;
w36211 <= pi0200 and not pi1155;
w36212 <= w8947 and not w36211;
w36213 <= pi1156 and w36212;
w36214 <= not w36210 and not w36213;
w36215 <= not pi0207 and w36214;
w36216 <= not w36137 and not w36215;
w36217 <= pi0208 and not w36216;
w36218 <= not w36208 and not w36217;
w36219 <= not pi1157 and not w36218;
w36220 <= not pi1156 and not w36111;
w36221 <= w36131 and w36220;
w36222 <= not w36115 and not w36221;
w36223 <= pi0207 and not w36222;
w36224 <= not pi0208 and not w36223;
w36225 <= not w36217 and not w36224;
w36226 <= pi1157 and not w36225;
w36227 <= not w36219 and not w36226;
w36228 <= not pi0219 and not w35976;
w36229 <= not w35977 and not w36228;
w36230 <= not w36227 and w36229;
w36231 <= not pi1157 and not w36102;
w36232 <= not pi1156 and not w36110;
w36233 <= w8936 and not w36092;
w36234 <= pi1156 and not w36233;
w36235 <= not w36232 and not w36234;
w36236 <= pi0207 and w36235;
w36237 <= not pi0207 and not pi0299;
w36238 <= not pi0208 and not w36237;
w36239 <= not w36236 and w36238;
w36240 <= pi1157 and not w36239;
w36241 <= not w36032 and not w36231;
w36242 <= not w36240 and w36241;
w36243 <= pi0299 and pi1142;
w36244 <= pi1153 and w36148;
w36245 <= pi1153 and not w36108;
w36246 <= not pi1153 and not w8373;
w36247 <= not w36245 and not w36246;
w36248 <= pi1155 and not w36247;
w36249 <= not w36244 and not w36248;
w36250 <= not pi1154 and not w36249;
w36251 <= not w36132 and w36204;
w36252 <= not w36158 and not w36251;
w36253 <= pi1154 and not w36252;
w36254 <= not w36250 and not w36253;
w36255 <= not pi0299 and not w36254;
w36256 <= pi0207 and not w36243;
w36257 <= not w36255 and w36256;
w36258 <= not w36140 and not w36243;
w36259 <= not pi1154 and not pi1156;
w36260 <= not w36258 and w36259;
w36261 <= pi1156 and not w36159;
w36262 <= pi0199 and not pi0200;
w36263 <= not pi0299 and not w36262;
w36264 <= not pi1155 and not w36263;
w36265 <= not w36145 and not w36264;
w36266 <= pi1154 and not w36265;
w36267 <= not w36261 and not w36266;
w36268 <= not w36032 and not w36267;
w36269 <= not pi0207 and not w36260;
w36270 <= not w36268 and w36269;
w36271 <= pi0208 and not w36270;
w36272 <= not w36257 and w36271;
w36273 <= not w8049 and not w36229;
w36274 <= not w36242 and w36273;
w36275 <= not w36272 and w36274;
w36276 <= w4989 and not w36275;
w36277 <= not w36230 and w36276;
w36278 <= not w36203 and w36277;
w36279 <= pi0213 and not w35993;
w36280 <= not w36278 and w36279;
w36281 <= pi0211 and not w36227;
w36282 <= not pi0214 and not w36227;
w36283 <= not pi0212 and not w36282;
w36284 <= not pi0207 and not w36073;
w36285 <= not pi0208 and not w36284;
w36286 <= not w8947 and not w36109;
w36287 <= pi1156 and not w36286;
w36288 <= not pi1156 and not w36108;
w36289 <= not w36264 and w36288;
w36290 <= not w36287 and not w36289;
w36291 <= pi0207 and w36290;
w36292 <= pi1157 and w36285;
w36293 <= not w36291 and w36292;
w36294 <= not pi1155 and not w8947;
w36295 <= not pi0299 and w36095;
w36296 <= not w36144 and not w36294;
w36297 <= not w36295 and w36296;
w36298 <= w36285 and w36297;
w36299 <= pi0207 and w36254;
w36300 <= w36214 and w36284;
w36301 <= pi0208 and not w36300;
w36302 <= not w36299 and w36301;
w36303 <= not w36293 and not w36298;
w36304 <= not w36302 and w36303;
w36305 <= w36062 and w36304;
w36306 <= w36283 and not w36305;
w36307 <= not pi0211 and not pi0214;
w36308 <= pi0299 and not pi1154;
w36309 <= pi1157 and not w36308;
w36310 <= w36239 and w36309;
w36311 <= w36214 and not w36266;
w36312 <= not pi0207 and not w36311;
w36313 <= not pi0299 and w36252;
w36314 <= pi1154 and not w36313;
w36315 <= not w36135 and not w36314;
w36316 <= pi0207 and not w36315;
w36317 <= not w36312 and not w36316;
w36318 <= pi0208 and not w36317;
w36319 <= not w36077 and not w36207;
w36320 <= not pi0208 and not w36319;
w36321 <= not pi1157 and w36320;
w36322 <= not w36310 and not w36321;
w36323 <= not w36318 and w36322;
w36324 <= w36307 and w36323;
w36325 <= pi1153 and not w36263;
w36326 <= w36128 and not w36325;
w36327 <= pi0207 and not w36326;
w36328 <= pi0299 and not pi1155;
w36329 <= pi1155 and not w36096;
w36330 <= not w36328 and not w36329;
w36331 <= w36267 and w36330;
w36332 <= pi0299 and not pi1153;
w36333 <= not pi0207 and not w36332;
w36334 <= not w36331 and w36333;
w36335 <= not w36327 and not w36334;
w36336 <= pi0208 and not w36335;
w36337 <= not w36231 and not w36332;
w36338 <= not w36240 and w36337;
w36339 <= w36062 and not w36336;
w36340 <= not w36338 and w36339;
w36341 <= pi0212 and not w36324;
w36342 <= not w36340 and w36341;
w36343 <= not w36306 and not w36342;
w36344 <= not w36281 and not w36343;
w36345 <= pi0219 and not w36344;
w36346 <= not w8047 and not w36307;
w36347 <= not w36304 and w36346;
w36348 <= w8047 and not w36323;
w36349 <= not w36095 and w36102;
w36350 <= pi0299 and pi1156;
w36351 <= not w36223 and not w36350;
w36352 <= w36105 and not w36351;
w36353 <= pi0207 and not w36136;
w36354 <= not w36210 and not w36261;
w36355 <= not pi0207 and not w36354;
w36356 <= pi0207 and w36350;
w36357 <= not w36355 and not w36356;
w36358 <= not w36353 and w36357;
w36359 <= pi0208 and not w36358;
w36360 <= not w36349 and not w36352;
w36361 <= not w36359 and w36360;
w36362 <= w36307 and not w36361;
w36363 <= not w36347 and not w36362;
w36364 <= not w36348 and w36363;
w36365 <= pi0212 and not w36364;
w36366 <= pi0211 and not w36361;
w36367 <= not pi0207 and w36331;
w36368 <= w36004 and w36326;
w36369 <= pi0208 and not w36368;
w36370 <= not w36367 and w36369;
w36371 <= w36240 and not w36370;
w36372 <= not pi0211 and not w36371;
w36373 <= not w36219 and w36372;
w36374 <= pi0214 and not w36366;
w36375 <= not w36373 and w36374;
w36376 <= w36283 and not w36375;
w36377 <= not pi0219 and not w36365;
w36378 <= not w36376 and w36377;
w36379 <= w4989 and not w36378;
w36380 <= not w36345 and w36379;
w36381 <= w36070 and not w36380;
w36382 <= not pi0209 and not w36280;
w36383 <= not w36381 and w36382;
w36384 <= not w36089 and not w36383;
w36385 <= pi0230 and not w36384;
w36386 <= not w35975 and not w36385;
w36387 <= not w8050 and w36214;
w36388 <= not pi0207 and not pi0208;
w36389 <= not w8050 and not w36388;
w36390 <= not pi0199 and w36147;
w36391 <= not pi1154 and not w36123;
w36392 <= w36113 and not w36390;
w36393 <= not w36391 and w36392;
w36394 <= pi0207 and w36393;
w36395 <= not w36389 and not w36394;
w36396 <= not w36387 and not w36395;
w36397 <= not w35977 and w36396;
w36398 <= pi0219 and not w36397;
w36399 <= not pi0207 and w36077;
w36400 <= pi0207 and not w36311;
w36401 <= not w36399 and not w36400;
w36402 <= not pi0208 and not w36401;
w36403 <= not pi1155 and w8372;
w36404 <= not w36112 and not w36403;
w36405 <= not pi0299 and not w36404;
w36406 <= not w36391 and not w36405;
w36407 <= pi0207 and w36406;
w36408 <= not w36312 and not w36407;
w36409 <= pi0208 and not w36408;
w36410 <= not w36402 and not w36409;
w36411 <= not pi0211 and not w36410;
w36412 <= not w35976 and w36411;
w36413 <= w36398 and not w36412;
w36414 <= not pi0214 and not w36396;
w36415 <= not pi0212 and not w36414;
w36416 <= pi0207 and not w36354;
w36417 <= not w36350 and not w36416;
w36418 <= not pi0208 and not w36417;
w36419 <= w36357 and not w36394;
w36420 <= pi0208 and not w36419;
w36421 <= not w36418 and not w36420;
w36422 <= not pi0211 and not w36421;
w36423 <= not w36073 and w36214;
w36424 <= w36285 and not w36423;
w36425 <= pi0207 and not w36073;
w36426 <= not w36393 and w36425;
w36427 <= pi0208 and not w36426;
w36428 <= not w36300 and w36427;
w36429 <= not w36424 and not w36428;
w36430 <= pi0211 and not w36429;
w36431 <= not w36422 and not w36430;
w36432 <= pi0214 and w36431;
w36433 <= w36415 and not w36432;
w36434 <= pi0211 and not w36410;
w36435 <= not pi0211 and not w36429;
w36436 <= pi0214 and not w36435;
w36437 <= not w36434 and w36436;
w36438 <= not pi0214 and w36431;
w36439 <= pi0212 and not w36437;
w36440 <= not w36438 and w36439;
w36441 <= not pi0219 and not w36433;
w36442 <= not w36440 and w36441;
w36443 <= w33382 and not w36413;
w36444 <= not w36442 and w36443;
w36445 <= pi0211 and pi1153;
w36446 <= not w36058 and not w36445;
w36447 <= not w8406 and w36446;
w36448 <= w36228 and not w36447;
w36449 <= not w36061 and w36448;
w36450 <= not w4989 and w36449;
w36451 <= not pi1152 and not w36450;
w36452 <= pi0207 and w36330;
w36453 <= w36267 and w36452;
w36454 <= w36238 and not w36453;
w36455 <= w36004 and not w36406;
w36456 <= pi0208 and not w36455;
w36457 <= not w36367 and w36456;
w36458 <= not w36454 and not w36457;
w36459 <= not w36332 and not w36458;
w36460 <= pi0211 and w36459;
w36461 <= not w36411 and not w36460;
w36462 <= pi0214 and w36461;
w36463 <= w36415 and not w36462;
w36464 <= not pi0219 and not w36463;
w36465 <= not pi0214 and not w36461;
w36466 <= not pi0211 and not w36459;
w36467 <= pi0214 and not w36466;
w36468 <= pi0211 and not w36396;
w36469 <= w36467 and not w36468;
w36470 <= not w36465 and not w36469;
w36471 <= pi0212 and not w36470;
w36472 <= w36464 and not w36471;
w36473 <= pi0219 and not w36396;
w36474 <= w4989 and not w36473;
w36475 <= not w36472 and w36474;
w36476 <= w36451 and not w36475;
w36477 <= pi1153 and not w36307;
w36478 <= not w36059 and not w36062;
w36479 <= not w36477 and not w36478;
w36480 <= pi0212 and not w36479;
w36481 <= w35984 and not w36446;
w36482 <= not pi0219 and not w36481;
w36483 <= not w36480 and w36482;
w36484 <= w35979 and not w36483;
w36485 <= pi1152 and not w36484;
w36486 <= not w36458 and w36467;
w36487 <= not w36465 and not w36486;
w36488 <= pi0212 and not w36487;
w36489 <= w36464 and not w36488;
w36490 <= w35977 and not w36458;
w36491 <= w36398 and not w36490;
w36492 <= w4989 and not w36491;
w36493 <= not w36489 and w36492;
w36494 <= w36485 and not w36493;
w36495 <= not pi0213 and not w36476;
w36496 <= not w36494 and w36495;
w36497 <= pi0209 and not w36444;
w36498 <= not w36496 and w36497;
w36499 <= not pi0199 and pi1153;
w36500 <= pi0200 and w36499;
w36501 <= not pi0299 and w36500;
w36502 <= not pi1154 and not w36501;
w36503 <= pi1154 and w36108;
w36504 <= not w36499 and w36503;
w36505 <= not w36502 and not w36504;
w36506 <= w36263 and not w36505;
w36507 <= w36238 and not w36506;
w36508 <= not pi0200 and not pi1153;
w36509 <= not pi0199 and not w36508;
w36510 <= not pi0299 and not w36509;
w36511 <= not w36262 and w36510;
w36512 <= pi0207 and w36511;
w36513 <= not pi0207 and w36506;
w36514 <= pi0208 and not w36512;
w36515 <= not w36513 and w36514;
w36516 <= not w36507 and not w36515;
w36517 <= not pi0211 and w36516;
w36518 <= not pi0299 and w8372;
w36519 <= not pi1153 and not w36518;
w36520 <= w36122 and not w36519;
w36521 <= not pi0199 and not pi1153;
w36522 <= w36204 and not w36521;
w36523 <= not w36520 and not w36522;
w36524 <= not w8050 and w36523;
w36525 <= not pi1153 and w8372;
w36526 <= w36113 and not w36525;
w36527 <= w8050 and not w36526;
w36528 <= not w36388 and not w36527;
w36529 <= not w36524 and w36528;
w36530 <= pi0211 and not w36529;
w36531 <= not w36517 and not w36530;
w36532 <= not w35976 and w36531;
w36533 <= pi0219 and not w35976;
w36534 <= pi0219 and not w36529;
w36535 <= not w36533 and not w36534;
w36536 <= not w36532 and not w36535;
w36537 <= w4989 and not w36536;
w36538 <= not pi0207 and w36075;
w36539 <= not pi1153 and not w36131;
w36540 <= not w36144 and not w36539;
w36541 <= pi1154 and not w8936;
w36542 <= not w36539 and w36541;
w36543 <= not w36540 and not w36542;
w36544 <= pi0207 and not w36543;
w36545 <= not w36538 and not w36544;
w36546 <= not pi0208 and not w36545;
w36547 <= not pi0207 and not w36543;
w36548 <= not pi0299 and w36112;
w36549 <= pi0207 and not w36548;
w36550 <= not w36246 and w36549;
w36551 <= not w36547 and not w36550;
w36552 <= pi0208 and not w36551;
w36553 <= not w36546 and not w36552;
w36554 <= not pi0211 and not w36553;
w36555 <= pi0211 and not w36516;
w36556 <= pi0214 and not w36554;
w36557 <= not w36555 and w36556;
w36558 <= pi0207 and not w36523;
w36559 <= not w36077 and not w36558;
w36560 <= not pi0208 and not w36559;
w36561 <= pi0207 and not w36511;
w36562 <= not w36308 and w36561;
w36563 <= pi1154 and not w8373;
w36564 <= not w36520 and not w36563;
w36565 <= not w36522 and w36564;
w36566 <= not pi0207 and not w36565;
w36567 <= not w36562 and not w36566;
w36568 <= pi0208 and not w36567;
w36569 <= not w36560 and not w36568;
w36570 <= not pi0211 and not w36569;
w36571 <= pi0211 and not w36553;
w36572 <= not w36570 and not w36571;
w36573 <= not pi0214 and w36572;
w36574 <= pi0212 and not w36557;
w36575 <= not w36573 and w36574;
w36576 <= not pi0214 and not w36529;
w36577 <= not pi0212 and not w36576;
w36578 <= pi0214 and w36572;
w36579 <= w36577 and not w36578;
w36580 <= not pi0219 and not w36575;
w36581 <= not w36579 and w36580;
w36582 <= w36537 and not w36581;
w36583 <= w36485 and not w36582;
w36584 <= pi0200 and not pi1153;
w36585 <= w8947 and not w36584;
w36586 <= pi1154 and not w36585;
w36587 <= not w36502 and not w36586;
w36588 <= w36389 and w36587;
w36589 <= pi0208 and w36004;
w36590 <= pi1153 and not w8373;
w36591 <= w36589 and w36590;
w36592 <= not w36588 and not w36591;
w36593 <= pi0219 and w36592;
w36594 <= w4989 and not w36593;
w36595 <= pi1153 and not pi1154;
w36596 <= not w36096 and w36595;
w36597 <= not w36542 and not w36596;
w36598 <= pi0207 and not w36597;
w36599 <= not w36538 and not w36598;
w36600 <= not pi0208 and not w36599;
w36601 <= not pi0207 and not w36597;
w36602 <= pi0207 and not w8373;
w36603 <= pi1153 and w36602;
w36604 <= not w36601 and not w36603;
w36605 <= pi0208 and not w36604;
w36606 <= not w36600 and not w36605;
w36607 <= w36090 and w36606;
w36608 <= pi1153 and not w8936;
w36609 <= not w36246 and not w36608;
w36610 <= pi1154 and not w36609;
w36611 <= not w36501 and not w36610;
w36612 <= pi0207 and not w36611;
w36613 <= not w36399 and not w36612;
w36614 <= not pi0208 and not w36613;
w36615 <= not pi0299 and not pi1153;
w36616 <= not w8373 and not w36615;
w36617 <= not w36308 and w36616;
w36618 <= pi0207 and not w36617;
w36619 <= not pi0207 and w36611;
w36620 <= pi0208 and not w36618;
w36621 <= not w36619 and w36620;
w36622 <= not w36614 and not w36621;
w36623 <= not pi0211 and w36622;
w36624 <= pi0211 and w36606;
w36625 <= not w36623 and not w36624;
w36626 <= w36171 and not w36625;
w36627 <= not w36607 and not w36626;
w36628 <= not pi0219 and not w36627;
w36629 <= not w36062 and not w36171;
w36630 <= w36592 and w36629;
w36631 <= w36594 and not w36630;
w36632 <= not w36628 and w36631;
w36633 <= w36451 and not w36632;
w36634 <= not w36583 and not w36633;
w36635 <= not pi0213 and w36634;
w36636 <= not pi1152 and w4989;
w36637 <= w35976 and not w36592;
w36638 <= not pi0299 and not w36500;
w36639 <= not pi1154 and not w36638;
w36640 <= not w36328 and w36639;
w36641 <= not w36294 and w36610;
w36642 <= not w36640 and not w36641;
w36643 <= pi0207 and w36642;
w36644 <= w36285 and not w36643;
w36645 <= not pi0207 and w36642;
w36646 <= not w36328 and w36616;
w36647 <= pi0207 and not w36646;
w36648 <= pi0208 and not w36647;
w36649 <= not w36645 and w36648;
w36650 <= not w36644 and not w36649;
w36651 <= not pi0211 and w36650;
w36652 <= pi0211 and w36622;
w36653 <= w8406 and not w36651;
w36654 <= not w36652 and w36653;
w36655 <= not pi0211 and not w36350;
w36656 <= w36592 and w36655;
w36657 <= pi0211 and w36650;
w36658 <= not w35986 and not w36656;
w36659 <= not w36657 and w36658;
w36660 <= not w36654 and not w36659;
w36661 <= not pi0219 and not w36660;
w36662 <= pi0211 and w36592;
w36663 <= w36533 and not w36662;
w36664 <= not w36623 and w36663;
w36665 <= not w36637 and not w36664;
w36666 <= not w36661 and w36665;
w36667 <= w36636 and not w36666;
w36668 <= not w35977 and w36529;
w36669 <= not w35976 and w36570;
w36670 <= not w36668 and not w36669;
w36671 <= pi0219 and not w36670;
w36672 <= not pi0212 and w36576;
w36673 <= pi0211 and not w36569;
w36674 <= not pi0199 and not pi1154;
w36675 <= not pi0200 and w36674;
w36676 <= w36237 and w36675;
w36677 <= w36285 and not w36506;
w36678 <= not w36515 and not w36677;
w36679 <= not w36328 and not w36676;
w36680 <= not w36678 and w36679;
w36681 <= not pi0211 and w36680;
w36682 <= w8406 and not w36681;
w36683 <= not w36673 and w36682;
w36684 <= not pi0208 and not w36350;
w36685 <= not w36558 and w36684;
w36686 <= pi0299 and not pi1156;
w36687 <= w36561 and not w36686;
w36688 <= not w36350 and w36523;
w36689 <= not pi0207 and not w36688;
w36690 <= pi0208 and not w36687;
w36691 <= not w36689 and w36690;
w36692 <= not pi0211 and not w36685;
w36693 <= not w36691 and w36692;
w36694 <= pi0211 and w36680;
w36695 <= not w35986 and not w36693;
w36696 <= not w36694 and w36695;
w36697 <= not pi0219 and not w36672;
w36698 <= not w36696 and w36697;
w36699 <= not w36683 and w36698;
w36700 <= not w36671 and not w36699;
w36701 <= pi1152 and w4989;
w36702 <= not w36700 and w36701;
w36703 <= not w36667 and not w36702;
w36704 <= pi0213 and not w36703;
w36705 <= not pi0209 and not w36704;
w36706 <= not w36635 and w36705;
w36707 <= not w36498 and not w36706;
w36708 <= pi0219 and not w36058;
w36709 <= pi0212 and not w36054;
w36710 <= pi0214 and not w36048;
w36711 <= not pi0212 and w36710;
w36712 <= not pi0219 and not w36711;
w36713 <= not w36709 and w36712;
w36714 <= pi0213 and not w36708;
w36715 <= w35979 and w36714;
w36716 <= not w36713 and w36715;
w36717 <= not w36707 and not w36716;
w36718 <= pi0230 and not w36717;
w36719 <= not pi0230 and pi0234;
w36720 <= not w36718 and not w36719;
w36721 <= pi0219 and not w36050;
w36722 <= pi0219 and not w36171;
w36723 <= not pi0212 and w36044;
w36724 <= not pi0214 and not w36043;
w36725 <= not w36710 and not w36724;
w36726 <= pi0212 and not w36725;
w36727 <= not pi0219 and not w36726;
w36728 <= not w36723 and w36727;
w36729 <= not w36721 and not w36722;
w36730 <= not w4989 and w36729;
w36731 <= not w36728 and w36730;
w36732 <= pi0208 and pi1157;
w36733 <= not w36213 and not w36329;
w36734 <= pi0207 and not w36733;
w36735 <= not pi0207 and not w36290;
w36736 <= not w36734 and not w36735;
w36737 <= w36732 and not w36736;
w36738 <= not pi0207 and w36297;
w36739 <= not w36734 and not w36738;
w36740 <= pi0208 and not w36739;
w36741 <= not w36298 and not w36740;
w36742 <= not pi1157 and not w36741;
w36743 <= not w36293 and not w36737;
w36744 <= not w36742 and w36743;
w36745 <= pi0211 and not w36744;
w36746 <= not pi1156 and w36140;
w36747 <= not w36261 and not w36746;
w36748 <= pi0207 and not w36747;
w36749 <= not w36221 and not w36234;
w36750 <= not pi0207 and not w36749;
w36751 <= not w36748 and not w36750;
w36752 <= w36732 and not w36751;
w36753 <= not pi0207 and w36099;
w36754 <= not w36748 and not w36753;
w36755 <= pi0208 and not w36754;
w36756 <= not w36349 and not w36755;
w36757 <= not pi1157 and not w36756;
w36758 <= not w36352 and not w36752;
w36759 <= not w36757 and w36758;
w36760 <= not pi0211 and not w36759;
w36761 <= w8406 and not w36745;
w36762 <= not w36760 and w36761;
w36763 <= w8050 and not w36213;
w36764 <= not w36746 and w36763;
w36765 <= not pi0207 and not w36206;
w36766 <= not w36764 and not w36765;
w36767 <= not w36208 and w36766;
w36768 <= not pi1157 and not w36767;
w36769 <= not pi0207 and w36222;
w36770 <= not w36764 and not w36769;
w36771 <= not w36224 and w36770;
w36772 <= pi1157 and not w36771;
w36773 <= not w36768 and not w36772;
w36774 <= w35976 and not w36773;
w36775 <= pi0211 and not w36759;
w36776 <= not pi0207 and w36235;
w36777 <= pi0208 and not w36776;
w36778 <= not w36261 and w36452;
w36779 <= w36777 and not w36778;
w36780 <= not w36239 and not w36779;
w36781 <= pi1157 and w36780;
w36782 <= not pi0211 and not w36768;
w36783 <= not w36781 and w36782;
w36784 <= w36171 and not w36783;
w36785 <= not w36775 and w36784;
w36786 <= not w36774 and not w36785;
w36787 <= not w36762 and w36786;
w36788 <= not pi0219 and not w36787;
w36789 <= not pi0211 and w36744;
w36790 <= pi0211 and not w36773;
w36791 <= not w35986 and not w36790;
w36792 <= not w36789 and w36791;
w36793 <= w35986 and w36773;
w36794 <= pi0219 and not w36793;
w36795 <= not w36792 and w36794;
w36796 <= pi0209 and not w36795;
w36797 <= not w36788 and w36796;
w36798 <= not w36254 and w36285;
w36799 <= not pi0207 and w36254;
w36800 <= pi0208 and not w36643;
w36801 <= not w36799 and w36800;
w36802 <= not w36798 and not w36801;
w36803 <= pi0211 and not w36802;
w36804 <= w8050 and not w36587;
w36805 <= not w36136 and not w36388;
w36806 <= not w8050 and not w36805;
w36807 <= not w36804 and not w36806;
w36808 <= not w36350 and not w36807;
w36809 <= not pi0211 and not w36808;
w36810 <= w8406 and not w36803;
w36811 <= not w36809 and w36810;
w36812 <= w35976 and not w36807;
w36813 <= w36238 and not w36368;
w36814 <= w36237 and w36326;
w36815 <= not w36610 and not w36639;
w36816 <= pi0207 and w36815;
w36817 <= pi0208 and not w36814;
w36818 <= not w36816 and w36817;
w36819 <= not w36813 and not w36818;
w36820 <= pi1157 and not w36819;
w36821 <= not pi1157 and w36807;
w36822 <= not pi0211 and not w36820;
w36823 <= not w36821 and w36822;
w36824 <= pi0211 and w36808;
w36825 <= not w36823 and not w36824;
w36826 <= w36171 and not w36825;
w36827 <= not w36811 and not w36812;
w36828 <= not w36826 and w36827;
w36829 <= not pi0219 and not w36828;
w36830 <= not pi0211 and w36802;
w36831 <= pi0211 and not w36807;
w36832 <= not w35986 and not w36831;
w36833 <= not w36830 and w36832;
w36834 <= w35986 and w36807;
w36835 <= pi0219 and not w36834;
w36836 <= not w36833 and w36835;
w36837 <= not pi0209 and not w36836;
w36838 <= not w36829 and w36837;
w36839 <= not w36797 and not w36838;
w36840 <= w4989 and not w36839;
w36841 <= pi0213 and not w36731;
w36842 <= not w36840 and w36841;
w36843 <= pi0219 and not w36060;
w36844 <= not w4989 and not w36843;
w36845 <= not w36052 and w36171;
w36846 <= w8406 and not w36446;
w36847 <= not pi0219 and not w36845;
w36848 <= not w36846 and w36847;
w36849 <= not w36722 and w36844;
w36850 <= not w36848 and w36849;
w36851 <= pi1157 and not w36780;
w36852 <= pi0299 and not pi1157;
w36853 <= not w36757 and not w36852;
w36854 <= not w36851 and w36853;
w36855 <= not w36332 and not w36854;
w36856 <= not pi0211 and not w36855;
w36857 <= w36791 and not w36856;
w36858 <= w36794 and not w36857;
w36859 <= not w36141 and not w36330;
w36860 <= not w36213 and not w36859;
w36861 <= pi0207 and not w36860;
w36862 <= pi1154 and not w36098;
w36863 <= not w36205 and not w36862;
w36864 <= not pi0207 and not w36295;
w36865 <= not w36863 and w36864;
w36866 <= not w36861 and not w36865;
w36867 <= pi0208 and not w36866;
w36868 <= not w36320 and not w36867;
w36869 <= not pi1157 and not w36868;
w36870 <= w36309 and not w36780;
w36871 <= not w36869 and not w36870;
w36872 <= not pi0211 and not w36871;
w36873 <= pi0211 and w36855;
w36874 <= w8406 and not w36872;
w36875 <= not w36873 and w36874;
w36876 <= pi0211 and w36871;
w36877 <= not w36789 and not w36876;
w36878 <= w36171 and not w36877;
w36879 <= not w36774 and not w36878;
w36880 <= not w36875 and w36879;
w36881 <= not pi0219 and not w36880;
w36882 <= not w36858 and not w36881;
w36883 <= pi0209 and not w36882;
w36884 <= not w36327 and not w36538;
w36885 <= not pi0208 and not w36884;
w36886 <= not pi0207 and not w36326;
w36887 <= not w36598 and not w36886;
w36888 <= pi0208 and not w36887;
w36889 <= not w36885 and not w36888;
w36890 <= not pi0211 and w36889;
w36891 <= w36832 and not w36890;
w36892 <= w36835 and not w36891;
w36893 <= not w36316 and not w36399;
w36894 <= not pi0208 and not w36893;
w36895 <= not pi0207 and not w36315;
w36896 <= not w36612 and not w36895;
w36897 <= pi0208 and not w36896;
w36898 <= not w36894 and not w36897;
w36899 <= pi0211 and w36898;
w36900 <= not w36830 and not w36899;
w36901 <= not w35986 and not w36900;
w36902 <= not pi0211 and not w36898;
w36903 <= pi0211 and not w36889;
w36904 <= w8406 and not w36903;
w36905 <= not w36902 and w36904;
w36906 <= not w36812 and not w36905;
w36907 <= not w36901 and w36906;
w36908 <= not pi0219 and not w36907;
w36909 <= not w36892 and not w36908;
w36910 <= not pi0209 and not w36909;
w36911 <= w4989 and not w36910;
w36912 <= not w36883 and w36911;
w36913 <= not pi0213 and not w36850;
w36914 <= not w36912 and w36913;
w36915 <= not w36842 and not w36914;
w36916 <= pi0230 and not w36915;
w36917 <= not pi0230 and not pi0235;
w36918 <= not w36916 and not w36917;
w36919 <= not pi0100 and w35761;
w36920 <= w35960 and not w36919;
w36921 <= not w3695 and not w36920;
w36922 <= not pi0075 and not w36921;
w36923 <= not w4865 and not w36922;
w36924 <= not pi0092 and not w36923;
w36925 <= w11217 and not w36924;
w36926 <= not pi0074 and not w36925;
w36927 <= w3694 and not w36926;
w36928 <= not pi0056 and not w36927;
w36929 <= not w3690 and not w36928;
w36930 <= not pi0062 and not w36929;
w36931 <= w11225 and not w36930;
w36932 <= pi0211 and pi1157;
w36933 <= not pi0211 and pi1158;
w36934 <= not w36932 and not w36933;
w36935 <= w35984 and not w36934;
w36936 <= w36727 and not w36935;
w36937 <= not pi0219 and not w4989;
w36938 <= w35984 and w36046;
w36939 <= not w4989 and w36938;
w36940 <= not w36937 and not w36939;
w36941 <= pi0214 and w36058;
w36942 <= pi1155 and w36307;
w36943 <= not w36941 and not w36942;
w36944 <= pi0212 and not w36943;
w36945 <= not w4989 and w36944;
w36946 <= w36940 and not w36945;
w36947 <= not w36936 and not w36946;
w36948 <= not pi0213 and not w36947;
w36949 <= w36071 and not w36936;
w36950 <= pi0199 and pi1143;
w36951 <= not pi0200 and not w36950;
w36952 <= not w35997 and w36951;
w36953 <= not w36000 and w36589;
w36954 <= not w36952 and w36953;
w36955 <= pi0200 and not w35997;
w36956 <= not pi0199 and pi1145;
w36957 <= w36951 and not w36956;
w36958 <= w36389 and not w36955;
w36959 <= not w36957 and w36958;
w36960 <= not w36954 and not w36959;
w36961 <= not pi0299 and not w36960;
w36962 <= w35984 and w36350;
w36963 <= pi0214 and not w36077;
w36964 <= not pi0214 and not w36073;
w36965 <= pi0212 and not w36963;
w36966 <= not w36964 and w36965;
w36967 <= not w36962 and not w36966;
w36968 <= w36082 and not w36967;
w36969 <= not w36961 and not w36968;
w36970 <= not w36949 and w36969;
w36971 <= w4989 and not w36970;
w36972 <= w36948 and not w36971;
w36973 <= pi0219 and not w35988;
w36974 <= w8406 and w35983;
w36975 <= not pi0211 and pi1145;
w36976 <= pi0211 and pi1144;
w36977 <= not w36975 and not w36976;
w36978 <= not w8406 and w36977;
w36979 <= not w35976 and not w36974;
w36980 <= not w36978 and w36979;
w36981 <= not pi0219 and not w36980;
w36982 <= w35979 and not w36973;
w36983 <= not w36981 and w36982;
w36984 <= w36071 and w36980;
w36985 <= pi0299 and w36533;
w36986 <= w35988 and w36985;
w36987 <= not w36961 and not w36986;
w36988 <= not w36984 and w36987;
w36989 <= w4989 and not w36988;
w36990 <= not w36983 and not w36989;
w36991 <= pi0213 and w36990;
w36992 <= pi0209 and not w36972;
w36993 <= not w36991 and w36992;
w36994 <= w36012 and w36131;
w36995 <= pi1158 and w36518;
w36996 <= not pi0199 and not pi1158;
w36997 <= pi1156 and not w36996;
w36998 <= not w36995 and not w36997;
w36999 <= w36994 and not w36998;
w37000 <= pi0207 and w36214;
w37001 <= pi0208 and not w36765;
w37002 <= not w37000 and w37001;
w37003 <= not w36999 and not w37002;
w37004 <= not pi1157 and not w37003;
w37005 <= pi1156 and w36262;
w37006 <= not pi0200 and not pi1158;
w37007 <= not pi0199 and not w37006;
w37008 <= not w37005 and not w37007;
w37009 <= w36004 and not w37008;
w37010 <= not pi0208 and w37009;
w37011 <= pi0208 and not w36769;
w37012 <= not w37000 and w37011;
w37013 <= not w37010 and not w37012;
w37014 <= pi1157 and not w37013;
w37015 <= not w37004 and not w37014;
w37016 <= not w35977 and w37015;
w37017 <= not pi0200 and pi0207;
w37018 <= not w36998 and w37017;
w37019 <= not pi1157 and not w37018;
w37020 <= pi1156 and not w36548;
w37021 <= not pi1158 and not w36204;
w37022 <= w37020 and not w37021;
w37023 <= not w37007 and not w37022;
w37024 <= w36004 and not w37023;
w37025 <= not pi0208 and not w37019;
w37026 <= w37024 and w37025;
w37027 <= not pi0208 and not w37026;
w37028 <= not w36106 and w37027;
w37029 <= not pi0299 and not w36099;
w37030 <= not pi0200 and pi1157;
w37031 <= not pi0199 and w37030;
w37032 <= w37029 and not w37031;
w37033 <= not pi0207 and not w36091;
w37034 <= not w37032 and w37033;
w37035 <= pi0207 and not w36164;
w37036 <= pi0208 and not w37034;
w37037 <= not w37035 and w37036;
w37038 <= not w37028 and not w37037;
w37039 <= w35977 and not w37038;
w37040 <= not w37016 and not w37039;
w37041 <= pi0219 and not w37040;
w37042 <= not pi0214 and w37015;
w37043 <= not pi0212 and not w37042;
w37044 <= pi0299 and not pi1145;
w37045 <= not pi0207 and not w37044;
w37046 <= not w37032 and w37045;
w37047 <= pi0299 and pi1145;
w37048 <= w36141 and not w37047;
w37049 <= not w36265 and not w37044;
w37050 <= pi1154 and not w37049;
w37051 <= not pi1156 and not w37048;
w37052 <= not w37050 and w37051;
w37053 <= w36156 and not w37047;
w37054 <= not w36159 and not w37044;
w37055 <= not pi1154 and not w37054;
w37056 <= pi1156 and not w37053;
w37057 <= not w37055 and w37056;
w37058 <= not w37052 and not w37057;
w37059 <= pi0207 and not w37058;
w37060 <= pi0208 and not w37046;
w37061 <= not w37059 and w37060;
w37062 <= w36204 and not w36288;
w37063 <= pi1157 and not w36995;
w37064 <= not w37062 and w37063;
w37065 <= pi0207 and not w37064;
w37066 <= not pi0299 and w37005;
w37067 <= not pi1157 and not w36995;
w37068 <= not w37066 and w37067;
w37069 <= w37065 and not w37068;
w37070 <= not pi0208 and not w37047;
w37071 <= not w37069 and w37070;
w37072 <= not w37061 and not w37071;
w37073 <= not pi0211 and not w37072;
w37074 <= not w36175 and w37027;
w37075 <= not pi0207 and not w36173;
w37076 <= not w37032 and w37075;
w37077 <= pi0207 and not w36193;
w37078 <= pi0208 and not w37076;
w37079 <= not w37077 and w37078;
w37080 <= not w37074 and not w37079;
w37081 <= pi0211 and not w37080;
w37082 <= not w37073 and not w37081;
w37083 <= pi0214 and not w37082;
w37084 <= w37043 and not w37083;
w37085 <= not pi0211 and w37080;
w37086 <= pi0211 and w37038;
w37087 <= pi0214 and not w37085;
w37088 <= not w37086 and w37087;
w37089 <= not pi0214 and not w37082;
w37090 <= pi0212 and not w37088;
w37091 <= not w37089 and w37090;
w37092 <= not pi0219 and not w37084;
w37093 <= not w37091 and w37092;
w37094 <= w4989 and not w37041;
w37095 <= not w37093 and w37094;
w37096 <= pi0213 and not w36983;
w37097 <= not w37095 and w37096;
w37098 <= not w36416 and not w36750;
w37099 <= w36732 and not w37098;
w37100 <= not w36350 and not w37009;
w37101 <= w36105 and not w37100;
w37102 <= w36684 and not w37018;
w37103 <= pi0208 and not w36753;
w37104 <= not w36416 and w37103;
w37105 <= not pi1157 and not w37102;
w37106 <= not w37104 and w37105;
w37107 <= not w37099 and not w37101;
w37108 <= not w37106 and w37107;
w37109 <= w35984 and w37108;
w37110 <= pi0207 and not w36423;
w37111 <= not w36735 and not w37110;
w37112 <= w36732 and not w37111;
w37113 <= not w36073 and not w37024;
w37114 <= w36105 and not w37113;
w37115 <= not w36738 and not w37110;
w37116 <= pi0208 and not w37115;
w37117 <= not pi0208 and w36073;
w37118 <= not w36999 and not w37117;
w37119 <= not w37116 and w37118;
w37120 <= not pi1157 and not w37119;
w37121 <= not w37112 and not w37114;
w37122 <= not w37120 and w37121;
w37123 <= not pi0214 and not w37122;
w37124 <= not pi0207 and not w36235;
w37125 <= not w36308 and w37124;
w37126 <= pi1157 and not w37125;
w37127 <= not pi1157 and not w36999;
w37128 <= not w36865 and w37127;
w37129 <= not w37126 and not w37128;
w37130 <= pi0208 and not w36400;
w37131 <= not w37129 and w37130;
w37132 <= w37024 and not w37127;
w37133 <= not pi0208 and not w36077;
w37134 <= not w37132 and w37133;
w37135 <= pi0214 and not w37134;
w37136 <= not w37131 and w37135;
w37137 <= pi0212 and not w37136;
w37138 <= not w37123 and w37137;
w37139 <= not w37109 and not w37138;
w37140 <= not pi0211 and not w37139;
w37141 <= not w37016 and not w37140;
w37142 <= pi0219 and not w37141;
w37143 <= not pi0299 and w37008;
w37144 <= w36238 and not w37143;
w37145 <= not w36453 and w36777;
w37146 <= not w37144 and not w37145;
w37147 <= pi1157 and not w37146;
w37148 <= not w37004 and not w37147;
w37149 <= pi0211 and w37148;
w37150 <= w36004 and w37005;
w37151 <= not pi0299 and not w36602;
w37152 <= pi1158 and not w37151;
w37153 <= not pi0208 and not w37150;
w37154 <= not w37152 and w37153;
w37155 <= not pi1158 and w36214;
w37156 <= pi1158 and w36331;
w37157 <= pi0207 and not w37155;
w37158 <= not w37156 and w37157;
w37159 <= pi0299 and not pi1158;
w37160 <= not pi0207 and not w37159;
w37161 <= not w37029 and w37160;
w37162 <= pi0208 and not w37161;
w37163 <= not w37158 and w37162;
w37164 <= not pi1157 and not w37154;
w37165 <= not w37163 and w37164;
w37166 <= w37124 and not w37159;
w37167 <= not w37158 and not w37166;
w37168 <= w36732 and not w37167;
w37169 <= not w37065 and not w37152;
w37170 <= w36105 and not w37169;
w37171 <= not pi0211 and not w37170;
w37172 <= not w37165 and w37171;
w37173 <= not w37168 and w37172;
w37174 <= not w37149 and not w37173;
w37175 <= pi0214 and not w37174;
w37176 <= w37043 and not w37175;
w37177 <= w36346 and not w37108;
w37178 <= w8047 and not w37122;
w37179 <= w36307 and not w37148;
w37180 <= not w37177 and not w37178;
w37181 <= not w37179 and w37180;
w37182 <= pi0212 and not w37181;
w37183 <= not pi0219 and not w37182;
w37184 <= not w37176 and w37183;
w37185 <= w4989 and not w37142;
w37186 <= not w37184 and w37185;
w37187 <= w36948 and not w37186;
w37188 <= not pi0209 and not w37097;
w37189 <= not w37187 and w37188;
w37190 <= not w36993 and not w37189;
w37191 <= pi0230 and not w37190;
w37192 <= not pi0230 and not pi0237;
w37193 <= not w37191 and not w37192;
w37194 <= not pi0211 and not pi1153;
w37195 <= pi0219 and w37194;
w37196 <= w35979 and not w37195;
w37197 <= not w36848 and w37196;
w37198 <= not pi1151 and w4989;
w37199 <= w8372 and w36389;
w37200 <= not pi0299 and not w37199;
w37201 <= not w10624 and not w37200;
w37202 <= w36389 and w36518;
w37203 <= not pi0214 and not w37202;
w37204 <= not pi0212 and w37203;
w37205 <= w37201 and not w37204;
w37206 <= pi1153 and w37205;
w37207 <= not w36228 and not w37206;
w37208 <= w36445 and not w37200;
w37209 <= pi1153 and w37202;
w37210 <= not w36077 and not w37209;
w37211 <= not pi0211 and not w37210;
w37212 <= w8406 and not w37208;
w37213 <= not w37211 and w37212;
w37214 <= pi0299 and not w36052;
w37215 <= not w35986 and not w37214;
w37216 <= not w37209 and w37215;
w37217 <= not w37213 and not w37216;
w37218 <= not pi0219 and not w37217;
w37219 <= w37198 and not w37207;
w37220 <= not w37218 and w37219;
w37221 <= not w8050 and w36131;
w37222 <= not w36388 and w37221;
w37223 <= w36124 and w36589;
w37224 <= not w37222 and not w37223;
w37225 <= not w36525 and not w37224;
w37226 <= not pi0214 and not w37225;
w37227 <= not pi0212 and not w37226;
w37228 <= w36131 and not w36521;
w37229 <= not pi1153 and not w36263;
w37230 <= not w36245 and not w37229;
w37231 <= pi1155 and not w37230;
w37232 <= not w37228 and not w37231;
w37233 <= w36004 and not w36124;
w37234 <= pi0208 and not w37233;
w37235 <= not w36285 and not w37234;
w37236 <= not w37232 and not w37235;
w37237 <= not w37223 and not w37236;
w37238 <= not pi0299 and not w37237;
w37239 <= pi0214 and not w37214;
w37240 <= not w37238 and w37239;
w37241 <= w37227 and not w37240;
w37242 <= not w36077 and w36346;
w37243 <= not w37225 and w37242;
w37244 <= w36307 and w37237;
w37245 <= not pi0299 and not w37017;
w37246 <= not pi0208 and not w37245;
w37247 <= pi0200 and w36237;
w37248 <= w37234 and not w37247;
w37249 <= not w37246 and not w37248;
w37250 <= not w36246 and not w37249;
w37251 <= w8047 and not w37250;
w37252 <= pi0212 and not w37243;
w37253 <= not w37251 and w37252;
w37254 <= not w37244 and w37253;
w37255 <= not pi0219 and not w37254;
w37256 <= not w37241 and w37255;
w37257 <= pi1151 and w4989;
w37258 <= not pi0211 and not w37249;
w37259 <= pi0211 and not w37224;
w37260 <= not w37258 and not w37259;
w37261 <= not w36246 and not w37260;
w37262 <= w35976 and not w37225;
w37263 <= w37261 and not w37262;
w37264 <= pi0219 and not w37263;
w37265 <= w37257 and not w37264;
w37266 <= not w37256 and w37265;
w37267 <= not pi1152 and not w37220;
w37268 <= not w37266 and w37267;
w37269 <= not w9008 and not w36608;
w37270 <= pi0207 and not w37269;
w37271 <= not w36538 and not w37270;
w37272 <= not pi0208 and not w37271;
w37273 <= pi0200 and pi0207;
w37274 <= not pi0199 and not w37273;
w37275 <= not pi0299 and not w37274;
w37276 <= pi0208 and not w37275;
w37277 <= not pi0207 and w8372;
w37278 <= not pi0299 and not w37277;
w37279 <= not pi1153 and not w37278;
w37280 <= w37276 and not w37279;
w37281 <= not w37272 and not w37280;
w37282 <= pi0211 and not w37281;
w37283 <= not pi0207 and not w36510;
w37284 <= not w36602 and not w37283;
w37285 <= pi0208 and not w37284;
w37286 <= w36238 and not w36510;
w37287 <= not w37285 and not w37286;
w37288 <= not pi0211 and not w36308;
w37289 <= not w37287 and w37288;
w37290 <= not w37282 and not w37289;
w37291 <= w8406 and not w37290;
w37292 <= pi0299 and w36052;
w37293 <= not w35986 and not w37287;
w37294 <= not w37292 and w37293;
w37295 <= not w37291 and not w37294;
w37296 <= not pi0219 and not w37295;
w37297 <= not w8050 and w36508;
w37298 <= not w36389 and not w37017;
w37299 <= w8947 and not w37298;
w37300 <= not w37297 and w37299;
w37301 <= not pi0211 and w36075;
w37302 <= not w35976 and w37301;
w37303 <= not w37300 and not w37302;
w37304 <= not w36228 and not w37303;
w37305 <= not w37296 and not w37304;
w37306 <= w37198 and not w37305;
w37307 <= w36004 and w36124;
w37308 <= pi0208 and w36113;
w37309 <= not w37277 and w37308;
w37310 <= not w37307 and not w37309;
w37311 <= not pi0214 and w37310;
w37312 <= not w37209 and w37311;
w37313 <= not pi0212 and not w37312;
w37314 <= not pi0214 and w37313;
w37315 <= w36511 and not w36549;
w37316 <= pi0208 and not w37315;
w37317 <= w36238 and not w36512;
w37318 <= not w37316 and not w37317;
w37319 <= not pi0211 and not w37318;
w37320 <= not w36328 and w37319;
w37321 <= pi0211 and not w37318;
w37322 <= not w36308 and w37321;
w37323 <= not w37320 and not w37322;
w37324 <= not w35986 and not w37323;
w37325 <= not w37208 and w37310;
w37326 <= not w37289 and w37325;
w37327 <= w8406 and not w37326;
w37328 <= not pi0219 and not w37314;
w37329 <= not w37327 and w37328;
w37330 <= not w37324 and w37329;
w37331 <= pi0219 and w37310;
w37332 <= not w37206 and w37331;
w37333 <= w37257 and not w37332;
w37334 <= not w37330 and w37333;
w37335 <= pi1152 and not w37334;
w37336 <= not w37306 and w37335;
w37337 <= not w37268 and not w37336;
w37338 <= not pi0209 and not w37337;
w37339 <= w36204 and w36595;
w37340 <= w8050 and not w37339;
w37341 <= not w36520 and w37340;
w37342 <= not w36806 and not w37341;
w37343 <= not pi0214 and not w37342;
w37344 <= not pi0212 and w37343;
w37345 <= pi0211 and w37342;
w37346 <= pi1153 and not w36144;
w37347 <= not w36520 and not w37346;
w37348 <= pi0207 and not w37347;
w37349 <= not w36886 and not w37348;
w37350 <= pi0208 and not w37349;
w37351 <= not w36885 and not w37350;
w37352 <= not pi0211 and not w37351;
w37353 <= not w37345 and not w37352;
w37354 <= w36533 and w37353;
w37355 <= not w36113 and w36647;
w37356 <= not pi1154 and not w36615;
w37357 <= not w36144 and w37356;
w37358 <= pi0207 and not w37357;
w37359 <= w36564 and w37358;
w37360 <= pi0208 and not w37359;
w37361 <= not w37355 and w37360;
w37362 <= not w36799 and w37361;
w37363 <= not w36798 and not w37362;
w37364 <= not pi0211 and not w37363;
w37365 <= w36564 and not w37339;
w37366 <= pi0207 and not w37365;
w37367 <= not w36895 and not w37366;
w37368 <= pi0208 and not w37367;
w37369 <= not w36894 and not w37368;
w37370 <= pi0211 and not w37369;
w37371 <= w35984 and not w37364;
w37372 <= not w37370 and w37371;
w37373 <= w8047 and not w37351;
w37374 <= w36307 and not w37363;
w37375 <= w36346 and not w37369;
w37376 <= pi0212 and not w37373;
w37377 <= not w37374 and w37376;
w37378 <= not w37375 and w37377;
w37379 <= not w37372 and not w37378;
w37380 <= not pi0219 and not w37379;
w37381 <= w4989 and not w37344;
w37382 <= not w37354 and w37381;
w37383 <= not w37380 and w37382;
w37384 <= pi0209 and not w37383;
w37385 <= not w37338 and not w37384;
w37386 <= not w37197 and not w37385;
w37387 <= pi0213 and not w37386;
w37388 <= not pi0211 and w36171;
w37389 <= pi1153 and w37388;
w37390 <= w36937 and w37389;
w37391 <= not pi1151 and not w37390;
w37392 <= pi0219 and not w37202;
w37393 <= w4989 and not w37392;
w37394 <= not w10624 and not w37209;
w37395 <= pi0212 and not w37203;
w37396 <= not w37394 and w37395;
w37397 <= not pi0219 and not w37396;
w37398 <= w37203 and w37206;
w37399 <= w35984 and w37301;
w37400 <= not w37202 and not w37399;
w37401 <= w37397 and w37400;
w37402 <= not w37398 and w37401;
w37403 <= w37206 and w37393;
w37404 <= not w37402 and w37403;
w37405 <= w37391 and not w37404;
w37406 <= w8049 and not w37389;
w37407 <= w35979 and not w37406;
w37408 <= pi1151 and not w37407;
w37409 <= not pi0214 and w37261;
w37410 <= not w37225 and w37394;
w37411 <= pi0214 and not w37410;
w37412 <= pi0212 and not w37411;
w37413 <= not w37409 and w37412;
w37414 <= not pi0212 and not w37263;
w37415 <= not w37413 and not w37414;
w37416 <= not pi0219 and not w37415;
w37417 <= not pi0211 and pi0299;
w37418 <= not w37209 and not w37417;
w37419 <= not w37225 and w37418;
w37420 <= not w37262 and not w37419;
w37421 <= pi0219 and not w37420;
w37422 <= w4989 and not w37421;
w37423 <= not w37416 and w37422;
w37424 <= w37408 and not w37423;
w37425 <= not pi1152 and not w37405;
w37426 <= not w37424 and w37425;
w37427 <= not w8048 and w36228;
w37428 <= not w4989 and w37427;
w37429 <= not w8406 and not w37194;
w37430 <= not w36090 and not w37429;
w37431 <= w37428 and not w37430;
w37432 <= not w8049 and w35979;
w37433 <= pi1151 and not w37432;
w37434 <= not w37431 and w37433;
w37435 <= not w37209 and w37310;
w37436 <= not w37319 and w37435;
w37437 <= pi0214 and w37436;
w37438 <= not w37312 and not w37437;
w37439 <= not pi0212 and not w37438;
w37440 <= not w37436 and not w37439;
w37441 <= pi0219 and not w37440;
w37442 <= w4989 and not w37441;
w37443 <= pi1153 and not w37200;
w37444 <= not w37321 and not w37443;
w37445 <= pi0214 and w37310;
w37446 <= w37444 and w37445;
w37447 <= w37313 and not w37446;
w37448 <= pi0214 and w37318;
w37449 <= w37311 and w37444;
w37450 <= pi0212 and not w37448;
w37451 <= not w37449 and w37450;
w37452 <= not pi0219 and not w37447;
w37453 <= not w37451 and w37452;
w37454 <= w37442 and not w37453;
w37455 <= w37434 and not w37454;
w37456 <= not pi1151 and not w37431;
w37457 <= pi0219 and not w37300;
w37458 <= w4989 and not w37457;
w37459 <= not pi0211 and w37281;
w37460 <= w37293 and not w37459;
w37461 <= not w36171 and w37300;
w37462 <= pi0299 and w36090;
w37463 <= not pi0219 and not w37462;
w37464 <= not w37461 and w37463;
w37465 <= not w37460 and w37464;
w37466 <= w37458 and not w37465;
w37467 <= w37456 and not w37466;
w37468 <= pi1152 and not w37467;
w37469 <= not w37455 and w37468;
w37470 <= not w37426 and not w37469;
w37471 <= not pi0209 and w37470;
w37472 <= not pi0219 and w36171;
w37473 <= not w37342 and not w37472;
w37474 <= w37353 and w37472;
w37475 <= w4989 and not w37473;
w37476 <= not w37474 and w37475;
w37477 <= w37391 and not w37476;
w37478 <= not w36814 and w37360;
w37479 <= not w36813 and not w37478;
w37480 <= not pi0211 and not w37479;
w37481 <= not w37345 and not w37480;
w37482 <= not w35976 and w37481;
w37483 <= not w37344 and not w37482;
w37484 <= pi0219 and not w37483;
w37485 <= w4989 and not w37484;
w37486 <= pi0214 and w37353;
w37487 <= not w37343 and not w37486;
w37488 <= not pi0212 and not w37487;
w37489 <= not pi0214 and not w37353;
w37490 <= pi0211 and not w37479;
w37491 <= not pi0211 and w37342;
w37492 <= not w37490 and not w37491;
w37493 <= pi0214 and not w37492;
w37494 <= pi0212 and not w37489;
w37495 <= not w37493 and w37494;
w37496 <= not w37488 and not w37495;
w37497 <= not pi0219 and not w37496;
w37498 <= w37485 and not w37497;
w37499 <= w37408 and not w37498;
w37500 <= not pi1152 and not w37477;
w37501 <= not w37499 and w37500;
w37502 <= not w37352 and not w37490;
w37503 <= not pi0214 and not w37502;
w37504 <= pi0214 and not w37481;
w37505 <= not w37503 and not w37504;
w37506 <= pi0212 and not w37505;
w37507 <= pi0214 and w37502;
w37508 <= not pi0212 and not w37343;
w37509 <= not w37507 and w37508;
w37510 <= not pi0219 and not w37509;
w37511 <= not w37506 and w37510;
w37512 <= pi0219 and not w37342;
w37513 <= w4989 and not w37512;
w37514 <= not w37511 and w37513;
w37515 <= w37456 and not w37514;
w37516 <= pi0214 and not w37479;
w37517 <= not w37503 and not w37516;
w37518 <= pi0212 and not w37517;
w37519 <= w37510 and not w37518;
w37520 <= w37485 and not w37519;
w37521 <= w37434 and not w37520;
w37522 <= pi1152 and not w37515;
w37523 <= not w37521 and w37522;
w37524 <= pi0209 and not w37501;
w37525 <= not w37523 and w37524;
w37526 <= not pi0213 and not w37471;
w37527 <= not w37525 and w37526;
w37528 <= not w37387 and not w37527;
w37529 <= pi0230 and not w37528;
w37530 <= not pi0230 and pi0238;
w37531 <= not w37529 and not w37530;
w37532 <= w36012 and not w36214;
w37533 <= pi0212 and not w37532;
w37534 <= w4989 and not w37533;
w37535 <= not pi0214 and w37532;
w37536 <= not pi0212 and not w37535;
w37537 <= not pi0219 and w37536;
w37538 <= pi0299 and pi1158;
w37539 <= not w36012 and w37538;
w37540 <= not pi0208 and w37158;
w37541 <= not w37539 and not w37540;
w37542 <= not pi0211 and not w37541;
w37543 <= not pi1157 and not w37532;
w37544 <= pi0208 and pi0299;
w37545 <= pi1157 and not w37544;
w37546 <= not w36454 and w37545;
w37547 <= pi0211 and not w37543;
w37548 <= not w37546 and w37547;
w37549 <= not w37542 and not w37548;
w37550 <= pi0214 and not w37549;
w37551 <= w37537 and not w37550;
w37552 <= pi0219 and w37536;
w37553 <= pi0211 and not w37532;
w37554 <= pi0214 and not w37553;
w37555 <= not w36418 and w36655;
w37556 <= w37554 and not w37555;
w37557 <= w37552 and not w37556;
w37558 <= not pi0209 and w37534;
w37559 <= not w37557 and w37558;
w37560 <= not w37551 and w37559;
w37561 <= not pi0219 and not w36935;
w37562 <= not w36940 and not w37561;
w37563 <= w37010 and not w37127;
w37564 <= not pi0214 and w37563;
w37565 <= not pi0212 and not w37564;
w37566 <= not pi0219 and w37565;
w37567 <= not w37144 and w37545;
w37568 <= not w37127 and not w37567;
w37569 <= pi0211 and not w37568;
w37570 <= pi0208 and not w37538;
w37571 <= not w36105 and not w37570;
w37572 <= not w37154 and w37571;
w37573 <= w37171 and not w37572;
w37574 <= pi0214 and not w37569;
w37575 <= not w37573 and w37574;
w37576 <= w37566 and not w37575;
w37577 <= pi0212 and not w37563;
w37578 <= w4989 and not w37577;
w37579 <= pi0219 and w37565;
w37580 <= pi0211 and not w37563;
w37581 <= w36655 and not w37563;
w37582 <= pi0214 and not w37581;
w37583 <= not w37580 and w37582;
w37584 <= w37579 and not w37583;
w37585 <= pi0209 and w37578;
w37586 <= not w37584 and w37585;
w37587 <= not w37576 and w37586;
w37588 <= pi0213 and not w37562;
w37589 <= not w37587 and w37588;
w37590 <= not w37560 and w37589;
w37591 <= not w4989 and not w36708;
w37592 <= w35984 and not w36712;
w37593 <= w37591 and w37592;
w37594 <= pi0211 and not w36073;
w37595 <= not w37026 and w37594;
w37596 <= w37582 and not w37595;
w37597 <= w37566 and not w37596;
w37598 <= not pi0211 and not w36077;
w37599 <= not w37026 and w37598;
w37600 <= pi0214 and not w37580;
w37601 <= not w37599 and w37600;
w37602 <= w37579 and not w37601;
w37603 <= w37578 and not w37597;
w37604 <= not w37602 and w37603;
w37605 <= pi0209 and not w37604;
w37606 <= not w36077 and not w36402;
w37607 <= w37554 and not w37606;
w37608 <= w37552 and not w37607;
w37609 <= not w36424 and w37594;
w37610 <= pi0214 and not w37609;
w37611 <= not w37555 and w37610;
w37612 <= w37537 and not w37611;
w37613 <= w37534 and not w37612;
w37614 <= not w37608 and w37613;
w37615 <= not pi0209 and not w37614;
w37616 <= not w37605 and not w37615;
w37617 <= not pi0213 and not w37593;
w37618 <= not w37616 and w37617;
w37619 <= not w37590 and not w37618;
w37620 <= pi0230 and not w37619;
w37621 <= not pi0230 and not pi0239;
w37622 <= not w37620 and not w37621;
w37623 <= w4989 and w37299;
w37624 <= not w37393 and not w37623;
w37625 <= not pi0214 and not w37299;
w37626 <= not pi0212 and not w37625;
w37627 <= w8947 and w36012;
w37628 <= not pi0299 and not w37627;
w37629 <= not w37276 and w37628;
w37630 <= pi0214 and w37629;
w37631 <= w37626 and not w37630;
w37632 <= not pi0219 and not w37631;
w37633 <= pi0211 and w37299;
w37634 <= not pi0211 and not w37629;
w37635 <= pi0214 and not w37633;
w37636 <= not w37634 and w37635;
w37637 <= pi0212 and not w37636;
w37638 <= not w37629 and w37637;
w37639 <= w37632 and not w37638;
w37640 <= not w37624 and not w37639;
w37641 <= not w37428 and not w37640;
w37642 <= not pi1147 and w37641;
w37643 <= not pi0211 and not w4989;
w37644 <= not w36937 and not w37643;
w37645 <= not w35976 and not w37644;
w37646 <= pi0299 and not w35976;
w37647 <= w4989 and not w35978;
w37648 <= w37646 and w37647;
w37649 <= w36113 and not w36388;
w37650 <= w4989 and w37649;
w37651 <= not w37648 and not w37650;
w37652 <= not w37645 and w37651;
w37653 <= pi1147 and w37652;
w37654 <= pi1149 and not w37653;
w37655 <= not w37642 and w37654;
w37656 <= pi0211 and w35984;
w37657 <= pi0212 and w36346;
w37658 <= not w37656 and not w37657;
w37659 <= w36937 and not w37658;
w37660 <= not w36389 and not w36602;
w37661 <= not w8050 and w36096;
w37662 <= not w37660 and not w37661;
w37663 <= w37278 and w37662;
w37664 <= pi0299 and w8047;
w37665 <= not w37663 and not w37664;
w37666 <= not pi0212 and not w37665;
w37667 <= not pi0219 and not w37666;
w37668 <= not pi0299 and not w37662;
w37669 <= pi0214 and not w37668;
w37670 <= not pi0214 and w37663;
w37671 <= not pi0212 and not w37670;
w37672 <= not w37669 and w37671;
w37673 <= not pi0211 and not w37668;
w37674 <= not w37663 and not w37673;
w37675 <= pi0214 and not w37674;
w37676 <= pi0212 and not w37675;
w37677 <= not pi0214 and not w37668;
w37678 <= w37676 and not w37677;
w37679 <= not w37672 and not w37678;
w37680 <= not w10624 and not w37663;
w37681 <= not w37669 and w37680;
w37682 <= pi0212 and not w37681;
w37683 <= w37679 and w37682;
w37684 <= w37667 and not w37683;
w37685 <= pi0219 and not w37663;
w37686 <= w4989 and not w37685;
w37687 <= not w37684 and w37686;
w37688 <= not w37659 and not w37687;
w37689 <= not pi1147 and w37688;
w37690 <= w4989 and not w37310;
w37691 <= pi0212 and not w36307;
w37692 <= not pi0219 and not w37656;
w37693 <= not w37691 and w37692;
w37694 <= w35979 and not w37693;
w37695 <= w37648 and not w37693;
w37696 <= not w37690 and not w37694;
w37697 <= not w37695 and w37696;
w37698 <= pi1147 and w37697;
w37699 <= not pi1149 and not w37698;
w37700 <= not w37689 and w37699;
w37701 <= not w37655 and not w37700;
w37702 <= pi1148 and not w37701;
w37703 <= w14042 and w37199;
w37704 <= not pi0219 and not w14042;
w37705 <= w37388 and w37704;
w37706 <= not w37703 and not w37705;
w37707 <= not pi1147 and w37706;
w37708 <= w8049 and not w37388;
w37709 <= w35979 and not w37708;
w37710 <= not pi0211 and not w37224;
w37711 <= pi0211 and not w37249;
w37712 <= pi0214 and not w37711;
w37713 <= not w37710 and w37712;
w37714 <= w8406 and not w37713;
w37715 <= not pi0214 and w37224;
w37716 <= not pi0212 and not w37715;
w37717 <= pi0214 and w37260;
w37718 <= w37716 and not w37717;
w37719 <= not pi0219 and not w37718;
w37720 <= pi0212 and not w37713;
w37721 <= not w37260 and w37720;
w37722 <= w37719 and not w37721;
w37723 <= not w37714 and w37722;
w37724 <= pi0212 and not w37260;
w37725 <= pi0219 and not w37724;
w37726 <= not w37718 and w37725;
w37727 <= w4989 and not w37726;
w37728 <= not w37723 and w37727;
w37729 <= not w37709 and not w37728;
w37730 <= pi1147 and w37729;
w37731 <= pi1149 and not w37707;
w37732 <= not w37730 and w37731;
w37733 <= not pi0212 and not w37664;
w37734 <= w37310 and w37733;
w37735 <= w37310 and not w37417;
w37736 <= not w37311 and not w37735;
w37737 <= not pi0214 and w10624;
w37738 <= pi0212 and not w37737;
w37739 <= not w37736 and w37738;
w37740 <= not w37734 and not w37739;
w37741 <= not pi0219 and not w37740;
w37742 <= w36263 and not w37273;
w37743 <= pi0208 and not w37742;
w37744 <= not pi0199 and not w37743;
w37745 <= not w37310 and not w37744;
w37746 <= not pi0299 and not w37745;
w37747 <= not pi0219 and w37746;
w37748 <= not w37741 and not w37747;
w37749 <= not pi0211 and not w37748;
w37750 <= not w10624 and w37445;
w37751 <= not pi0214 and w37735;
w37752 <= pi0212 and not w37751;
w37753 <= not w37750 and w37752;
w37754 <= not pi0212 and w37736;
w37755 <= not pi0219 and not w37754;
w37756 <= not w37753 and w37755;
w37757 <= pi0219 and not w37417;
w37758 <= w37647 and not w37757;
w37759 <= not w37690 and not w37758;
w37760 <= not w37756 and not w37759;
w37761 <= not w37746 and w37760;
w37762 <= not w37749 and w37761;
w37763 <= not w37432 and not w37762;
w37764 <= pi1147 and not pi1149;
w37765 <= not w37763 and w37764;
w37766 <= not w37732 and not w37765;
w37767 <= not pi1148 and not w37766;
w37768 <= not w37702 and not w37767;
w37769 <= pi0213 and not w37768;
w37770 <= w8409 and w36228;
w37771 <= not w4989 and w37770;
w37772 <= not pi0211 and pi1146;
w37773 <= pi0211 and pi1145;
w37774 <= not w37772 and not w37773;
w37775 <= pi0214 and not w37774;
w37776 <= pi0211 and pi1146;
w37777 <= not pi0214 and w37776;
w37778 <= not w37775 and not w37777;
w37779 <= pi0212 and not w37778;
w37780 <= w35984 and w37776;
w37781 <= not w37779 and not w37780;
w37782 <= not w36533 and w37781;
w37783 <= not w4989 and w36975;
w37784 <= not w36937 and not w37783;
w37785 <= not w37782 and not w37784;
w37786 <= pi1147 and not w37771;
w37787 <= not w37785 and w37786;
w37788 <= not pi0211 and w37047;
w37789 <= pi0219 and not w37788;
w37790 <= w37647 and not w37789;
w37791 <= not w37690 and not w37790;
w37792 <= w35976 and not w37310;
w37793 <= not pi0219 and not w37792;
w37794 <= pi0299 and not w37774;
w37795 <= w37310 and not w37794;
w37796 <= w8406 and not w37795;
w37797 <= pi0299 and pi1146;
w37798 <= pi0211 and w37797;
w37799 <= not w37417 and not w37798;
w37800 <= w37310 and w37799;
w37801 <= w36171 and not w37800;
w37802 <= w37793 and not w37796;
w37803 <= not w37801 and w37802;
w37804 <= not w37791 and not w37803;
w37805 <= w37787 and not w37804;
w37806 <= w4989 and w37663;
w37807 <= not pi1147 and not w37785;
w37808 <= pi0219 and w37790;
w37809 <= pi0299 and not w37781;
w37810 <= w33677 and w37809;
w37811 <= not w37808 and not w37810;
w37812 <= w37807 and w37811;
w37813 <= not w37806 and w37812;
w37814 <= pi1148 and not w37805;
w37815 <= not w37813 and w37814;
w37816 <= w36975 and w36985;
w37817 <= not w36228 and w37745;
w37818 <= not pi1146 and w10624;
w37819 <= w36171 and not w37818;
w37820 <= not w37796 and not w37819;
w37821 <= not pi0219 and not w37746;
w37822 <= not w37820 and w37821;
w37823 <= not w37816 and not w37817;
w37824 <= not w37822 and w37823;
w37825 <= w4989 and not w37824;
w37826 <= w37787 and not w37825;
w37827 <= not pi1148 and not w37812;
w37828 <= not w37826 and w37827;
w37829 <= not w37815 and not w37828;
w37830 <= not pi1149 and not w37829;
w37831 <= pi0219 and w37224;
w37832 <= w4989 and not w37831;
w37833 <= not w37790 and not w37832;
w37834 <= not pi0299 and w37248;
w37835 <= not w36994 and not w37834;
w37836 <= not w37797 and w37835;
w37837 <= pi0211 and not w37836;
w37838 <= not w37258 and not w37837;
w37839 <= pi0214 and w37838;
w37840 <= w37716 and not w37839;
w37841 <= pi0214 and not w37794;
w37842 <= w37835 and w37841;
w37843 <= not pi0214 and w37838;
w37844 <= pi0212 and not w37842;
w37845 <= not w37843 and w37844;
w37846 <= not pi0219 and not w37840;
w37847 <= not w37845 and w37846;
w37848 <= not w37833 and not w37847;
w37849 <= w37787 and not w37848;
w37850 <= not w37703 and w37812;
w37851 <= not pi1148 and not w37850;
w37852 <= not w37849 and w37851;
w37853 <= pi0219 and not w37649;
w37854 <= w4989 and not w37853;
w37855 <= pi0211 and not w37649;
w37856 <= pi0214 and pi0299;
w37857 <= not w37649 and not w37856;
w37858 <= not pi0212 and not w37857;
w37859 <= not w37855 and w37858;
w37860 <= not pi0299 and not w37649;
w37861 <= pi0212 and not w37860;
w37862 <= pi0299 and w37691;
w37863 <= w37861 and not w37862;
w37864 <= not pi0219 and not w37859;
w37865 <= not w37863 and w37864;
w37866 <= w37854 and not w37865;
w37867 <= w37787 and w37811;
w37868 <= not w37866 and w37867;
w37869 <= not w35977 and w37299;
w37870 <= not w35976 and w37634;
w37871 <= pi0219 and not w37869;
w37872 <= not w37870 and w37871;
w37873 <= w4989 and not w37872;
w37874 <= w8947 and w37873;
w37875 <= not w37790 and not w37874;
w37876 <= not w37299 and not w37798;
w37877 <= w37626 and not w37876;
w37878 <= pi0212 and not w37629;
w37879 <= not w37299 and w37778;
w37880 <= w37878 and not w37879;
w37881 <= not pi0219 and not w37877;
w37882 <= not w37880 and w37881;
w37883 <= not w37875 and not w37882;
w37884 <= w37807 and not w37883;
w37885 <= pi1148 and not w37868;
w37886 <= not w37884 and w37885;
w37887 <= not w37852 and not w37886;
w37888 <= pi1149 and not w37887;
w37889 <= not w37830 and not w37888;
w37890 <= not pi0213 and not w37889;
w37891 <= pi0209 and not w37890;
w37892 <= not w37769 and w37891;
w37893 <= pi0200 and not w36956;
w37894 <= pi0199 and pi1145;
w37895 <= not pi0200 and not w37894;
w37896 <= not pi0199 and pi1146;
w37897 <= w37895 and not w37896;
w37898 <= w36004 and not w37893;
w37899 <= not w37897 and w37898;
w37900 <= not w36389 and not w37899;
w37901 <= pi0200 and not w37896;
w37902 <= not pi0299 and not w37901;
w37903 <= not w37895 and w37902;
w37904 <= not w8050 and not w37903;
w37905 <= not w37900 and not w37904;
w37906 <= w35976 and w37905;
w37907 <= pi0219 and not w37906;
w37908 <= not w35976 and w37905;
w37909 <= not w35977 and not w37908;
w37910 <= w36262 and not w37894;
w37911 <= w37902 and not w37910;
w37912 <= not pi0207 and w37911;
w37913 <= w37895 and w37912;
w37914 <= not w37797 and not w37899;
w37915 <= not w37912 and w37914;
w37916 <= pi0208 and not w37915;
w37917 <= not w37913 and w37916;
w37918 <= w36012 and w37903;
w37919 <= not w37917 and not w37918;
w37920 <= not pi0299 and not w37919;
w37921 <= not pi0211 and not w37047;
w37922 <= not w37920 and w37921;
w37923 <= not w37909 and not w37922;
w37924 <= w37907 and not w37923;
w37925 <= not w37798 and not w37905;
w37926 <= not pi0214 and not w37905;
w37927 <= not pi0212 and not w37926;
w37928 <= not w37925 and w37927;
w37929 <= not pi0219 and not w37928;
w37930 <= w37841 and not w37920;
w37931 <= not pi0214 and w37925;
w37932 <= pi0212 and not w37931;
w37933 <= not w37930 and w37932;
w37934 <= w37929 and not w37933;
w37935 <= w4989 and not w37924;
w37936 <= not w37934 and w37935;
w37937 <= w37807 and not w37936;
w37938 <= not w8050 and not w37911;
w37939 <= not w37900 and not w37938;
w37940 <= not w35977 and w37939;
w37941 <= pi0219 and not w37940;
w37942 <= w36012 and w37911;
w37943 <= not w37916 and not w37942;
w37944 <= not pi0299 and w37943;
w37945 <= not pi0211 and not w37944;
w37946 <= not w37044 and w37945;
w37947 <= not w35976 and w37946;
w37948 <= w37941 and not w37947;
w37949 <= not w37939 and not w37945;
w37950 <= not pi0214 and not w37939;
w37951 <= not pi0212 and not w37950;
w37952 <= not w37949 and w37951;
w37953 <= pi0211 and not w37944;
w37954 <= not w37044 and w37953;
w37955 <= w37841 and w37943;
w37956 <= w8047 and not w37944;
w37957 <= not w37955 and not w37956;
w37958 <= not w37954 and not w37957;
w37959 <= not pi0214 and w37799;
w37960 <= w37943 and w37959;
w37961 <= pi0212 and not w37960;
w37962 <= not w37958 and w37961;
w37963 <= w37929 and not w37952;
w37964 <= not w37962 and w37963;
w37965 <= w4989 and not w37948;
w37966 <= not w37964 and w37965;
w37967 <= w37787 and not w37966;
w37968 <= not w37937 and not w37967;
w37969 <= not pi0213 and w37968;
w37970 <= pi1147 and not w37694;
w37971 <= not w35976 and w37945;
w37972 <= w37941 and not w37971;
w37973 <= w4989 and not w37972;
w37974 <= not pi0299 and w37919;
w37975 <= pi0214 and not w37974;
w37976 <= not w37953 and not w37975;
w37977 <= pi0212 and not w37976;
w37978 <= not pi0219 and not w37939;
w37979 <= not w37956 and w37978;
w37980 <= not w37977 and w37979;
w37981 <= w37973 and not w37980;
w37982 <= w37970 and not w37981;
w37983 <= not w37906 and w37980;
w37984 <= pi0219 and not w37905;
w37985 <= pi0214 and w37949;
w37986 <= not w37974 and not w37985;
w37987 <= pi0212 and not w37986;
w37988 <= not pi0214 and w37905;
w37989 <= not pi0212 and not w37988;
w37990 <= not w37975 and w37989;
w37991 <= not w37987 and not w37990;
w37992 <= not pi0219 and not w37991;
w37993 <= w4989 and not w37984;
w37994 <= not w37992 and w37993;
w37995 <= not w37983 and w37994;
w37996 <= not pi1147 and not w37659;
w37997 <= not w37995 and w37996;
w37998 <= not pi1149 and not w37982;
w37999 <= not w37997 and w37998;
w38000 <= not w37646 and w37978;
w38001 <= w37973 and not w38000;
w38002 <= pi1147 and not w37645;
w38003 <= not w38001 and w38002;
w38004 <= not pi1147 and not w37428;
w38005 <= not w37994 and w38004;
w38006 <= pi1149 and not w38003;
w38007 <= not w38005 and w38006;
w38008 <= pi1148 and not w38007;
w38009 <= not w37999 and w38008;
w38010 <= not pi1147 and w4989;
w38011 <= w37905 and w38010;
w38012 <= pi0214 and not w37939;
w38013 <= not w37953 and w38012;
w38014 <= not w37945 and w37950;
w38015 <= pi0212 and not w38013;
w38016 <= not w38014 and w38015;
w38017 <= not pi0219 and not w37952;
w38018 <= not w38016 and w38017;
w38019 <= w37981 and not w38018;
w38020 <= not w37432 and not w38019;
w38021 <= pi1147 and not w38020;
w38022 <= not w38011 and not w38021;
w38023 <= not pi1149 and not w38022;
w38024 <= w37973 and not w38018;
w38025 <= not w37709 and not w38024;
w38026 <= pi1147 and not w38025;
w38027 <= not pi1147 and w37770;
w38028 <= not w38011 and not w38027;
w38029 <= w14042 and w37770;
w38030 <= w37919 and w38029;
w38031 <= not w38028 and not w38030;
w38032 <= not w38026 and not w38031;
w38033 <= pi1149 and not w38032;
w38034 <= not pi1148 and not w38033;
w38035 <= not w38023 and w38034;
w38036 <= pi0213 and not w38009;
w38037 <= not w38035 and w38036;
w38038 <= not pi0209 and not w37969;
w38039 <= not w38037 and w38038;
w38040 <= not w37892 and not w38039;
w38041 <= pi0230 and not w38040;
w38042 <= not pi0230 and not pi0240;
w38043 <= not w38041 and not w38042;
w38044 <= pi0213 and not w37470;
w38045 <= w37198 and w37209;
w38046 <= w36071 and w37388;
w38047 <= not w37225 and not w38046;
w38048 <= not w4989 and not w37770;
w38049 <= pi1151 and not w38048;
w38050 <= not w38047 and w38049;
w38051 <= not w38045 and not w38050;
w38052 <= not pi1152 and not w38051;
w38053 <= not w37318 and w37770;
w38054 <= w37435 and not w38053;
w38055 <= pi1152 and not w38054;
w38056 <= w4989 and not w38055;
w38057 <= w38049 and not w38056;
w38058 <= pi1152 and w37198;
w38059 <= w37300 and w38058;
w38060 <= not w38052 and not w38059;
w38061 <= not w38057 and w38060;
w38062 <= not pi1150 and not w38061;
w38063 <= pi1151 and not w37428;
w38064 <= pi0219 and not w37209;
w38065 <= w4989 and not w38064;
w38066 <= not w37690 and not w38065;
w38067 <= w37313 and not w37448;
w38068 <= not pi0219 and not w38067;
w38069 <= not pi0214 and w37318;
w38070 <= pi0212 and not w38069;
w38071 <= not w37437 and w38070;
w38072 <= w38068 and not w38071;
w38073 <= pi1152 and not w38072;
w38074 <= not pi0299 and not w37250;
w38075 <= not pi0214 and w37249;
w38076 <= pi0212 and not w38075;
w38077 <= not w37717 and w38076;
w38078 <= not w37227 and not w38077;
w38079 <= not w38074 and not w38078;
w38080 <= not pi0219 and not w38079;
w38081 <= not pi1152 and not w37831;
w38082 <= not w38080 and w38081;
w38083 <= not w38073 and not w38082;
w38084 <= not w38066 and not w38083;
w38085 <= w38063 and not w38084;
w38086 <= not pi1151 and not w37659;
w38087 <= not pi0212 and not w37200;
w38088 <= not w37203 and w38087;
w38089 <= not w37417 and w38088;
w38090 <= not pi0219 and not w38089;
w38091 <= pi0214 and not w37201;
w38092 <= not pi0211 and w37203;
w38093 <= pi0212 and not w37200;
w38094 <= not w38092 and w38093;
w38095 <= not w38091 and w38094;
w38096 <= w38090 and not w38095;
w38097 <= not w37209 and w37397;
w38098 <= not pi0299 and w38097;
w38099 <= not w38096 and not w38098;
w38100 <= w38065 and w38099;
w38101 <= not pi1152 and not w38100;
w38102 <= not w37300 and not w38099;
w38103 <= w37458 and not w38102;
w38104 <= pi1152 and not w38103;
w38105 <= not w38101 and not w38104;
w38106 <= w38086 and not w38105;
w38107 <= pi1150 and not w38106;
w38108 <= not w38085 and w38107;
w38109 <= not w38062 and not w38108;
w38110 <= not pi1149 and not w38109;
w38111 <= pi1151 and not w37709;
w38112 <= not pi0214 and not w37419;
w38113 <= w37412 and not w38112;
w38114 <= not pi0212 and not w37420;
w38115 <= not w38113 and not w38114;
w38116 <= not pi0219 and not w38115;
w38117 <= not pi1152 and w37422;
w38118 <= not w38116 and w38117;
w38119 <= not w36346 and not w37318;
w38120 <= pi0212 and w37435;
w38121 <= not w38119 and w38120;
w38122 <= not w37439 and not w38121;
w38123 <= not pi0219 and not w38122;
w38124 <= pi1152 and not w38123;
w38125 <= w37442 and w38124;
w38126 <= w38111 and not w38118;
w38127 <= not w38125 and w38126;
w38128 <= not pi1151 and not w37432;
w38129 <= not w37758 and not w38065;
w38130 <= not w38097 and not w38129;
w38131 <= not pi1152 and w38130;
w38132 <= not w37458 and w38129;
w38133 <= not w37300 and w37397;
w38134 <= pi1152 and not w38132;
w38135 <= not w38133 and w38134;
w38136 <= w38128 and not w38131;
w38137 <= not w38135 and w38136;
w38138 <= not pi1150 and not w38137;
w38139 <= not w38127 and w38138;
w38140 <= not pi1151 and not w37694;
w38141 <= w8406 and w37287;
w38142 <= not w37204 and not w37394;
w38143 <= not w8406 and not w37300;
w38144 <= not w38142 and w38143;
w38145 <= not w38141 and not w38144;
w38146 <= not pi0219 and not w38145;
w38147 <= not w38132 and not w38146;
w38148 <= pi1152 and not w38147;
w38149 <= w38101 and not w38130;
w38150 <= not w38148 and not w38149;
w38151 <= w38140 and not w38150;
w38152 <= pi0212 and not w37318;
w38153 <= w38068 and not w38152;
w38154 <= pi1152 and not w38153;
w38155 <= w37442 and w38154;
w38156 <= pi1151 and not w37645;
w38157 <= not w37262 and not w38074;
w38158 <= not pi0219 and not w38157;
w38159 <= w38117 and not w38158;
w38160 <= w38156 and not w38159;
w38161 <= not w38155 and w38160;
w38162 <= pi1150 and not w38151;
w38163 <= not w38161 and w38162;
w38164 <= not w38139 and not w38163;
w38165 <= pi1149 and not w38164;
w38166 <= not w38110 and not w38165;
w38167 <= not pi0213 and not w38166;
w38168 <= pi0209 and not w38044;
w38169 <= not w38167 and w38168;
w38170 <= not pi1150 and pi1151;
w38171 <= not w37706 and w38170;
w38172 <= not w37687 and w38086;
w38173 <= not w37640 and w38063;
w38174 <= pi1150 and not w38173;
w38175 <= not w38172 and w38174;
w38176 <= not pi1149 and not w38171;
w38177 <= not w38175 and w38176;
w38178 <= w37651 and w38156;
w38179 <= not pi1151 and w37697;
w38180 <= pi1150 and not w38178;
w38181 <= not w38179 and w38180;
w38182 <= not w37762 and w38128;
w38183 <= not w37728 and w38111;
w38184 <= not pi1150 and not w38182;
w38185 <= not w38183 and w38184;
w38186 <= pi1149 and not w38181;
w38187 <= not w38185 and w38186;
w38188 <= not w38177 and not w38187;
w38189 <= not pi0213 and w38188;
w38190 <= not w37716 and not w37720;
w38191 <= not w36332 and w37258;
w38192 <= not w37259 and not w38191;
w38193 <= not w37714 and w38192;
w38194 <= not w38190 and not w38193;
w38195 <= not pi0219 and not w38194;
w38196 <= w37727 and not w38195;
w38197 <= w37408 and not w38196;
w38198 <= pi0299 and w37194;
w38199 <= not w37745 and not w38046;
w38200 <= w4989 and not w38199;
w38201 <= not w38198 and w38200;
w38202 <= w37391 and not w38201;
w38203 <= not pi1152 and not w38202;
w38204 <= not w38197 and w38203;
w38205 <= not w37713 and not w37715;
w38206 <= not pi0219 and not w37862;
w38207 <= not w37263 and w38206;
w38208 <= not w38205 and w38207;
w38209 <= w37727 and not w38208;
w38210 <= w37434 and not w38209;
w38211 <= not w37646 and not w37745;
w38212 <= not w36204 and w37430;
w38213 <= not w38211 and not w38212;
w38214 <= not pi0219 and not w38213;
w38215 <= pi0219 and not w37745;
w38216 <= w4989 and not w38215;
w38217 <= not w38214 and w38216;
w38218 <= w37456 and not w38217;
w38219 <= pi1152 and not w38218;
w38220 <= not w38210 and w38219;
w38221 <= not pi1150 and not w38220;
w38222 <= not w38204 and w38221;
w38223 <= not pi0219 and not w37649;
w38224 <= not w37862 and w38223;
w38225 <= not pi1153 and w38224;
w38226 <= pi0299 and w8048;
w38227 <= not pi0219 and not w38226;
w38228 <= w37758 and not w38227;
w38229 <= not w37866 and not w38228;
w38230 <= not w38225 and not w38229;
w38231 <= w37408 and not w38230;
w38232 <= pi1153 and w38046;
w38233 <= w37391 and not w38232;
w38234 <= not pi1152 and not w38233;
w38235 <= not pi1151 and not w37690;
w38236 <= not pi1152 and not w38235;
w38237 <= not w38234 and not w38236;
w38238 <= not w38231 and not w38237;
w38239 <= not pi0211 and w38224;
w38240 <= not w37651 and not w38239;
w38241 <= w37434 and not w38240;
w38242 <= not w38230 and w38241;
w38243 <= w4989 and not w37331;
w38244 <= w8406 and not w37735;
w38245 <= not pi0299 and w37310;
w38246 <= not w35986 and not w38198;
w38247 <= not w38245 and w38246;
w38248 <= w37793 and not w38244;
w38249 <= not w38247 and w38248;
w38250 <= w38243 and not w38249;
w38251 <= w37456 and not w38250;
w38252 <= pi1152 and not w38251;
w38253 <= not w38242 and w38252;
w38254 <= pi1150 and not w38238;
w38255 <= not w38253 and w38254;
w38256 <= pi1149 and not w38255;
w38257 <= not w38222 and w38256;
w38258 <= pi0219 and not w37205;
w38259 <= w4989 and not w38258;
w38260 <= not w37402 and w38259;
w38261 <= w37408 and not w38260;
w38262 <= w38234 and not w38261;
w38263 <= pi0299 and w37427;
w38264 <= not w37430 and w38263;
w38265 <= w37456 and not w38264;
w38266 <= w38090 and not w38094;
w38267 <= w38259 and not w38266;
w38268 <= w37434 and not w38260;
w38269 <= not w38267 and w38268;
w38270 <= pi1152 and not w38265;
w38271 <= not w38269 and w38270;
w38272 <= not pi1150 and not w38262;
w38273 <= not w38271 and w38272;
w38274 <= not w37472 and w37663;
w38275 <= not w36332 and not w37668;
w38276 <= not pi0211 and not w38275;
w38277 <= w37472 and not w37674;
w38278 <= not w38276 and w38277;
w38279 <= not w38274 and not w38278;
w38280 <= w4989 and not w38279;
w38281 <= w37391 and not w38280;
w38282 <= pi0211 and not w37629;
w38283 <= not w8936 and w36238;
w38284 <= not w37276 and not w38283;
w38285 <= not pi0211 and not w36332;
w38286 <= not w38284 and w38285;
w38287 <= not w38282 and not w38286;
w38288 <= not w37299 and not w38282;
w38289 <= pi0214 and w38288;
w38290 <= w37625 and not w37634;
w38291 <= pi0212 and not w38290;
w38292 <= not w38289 and w38291;
w38293 <= not w38287 and w38292;
w38294 <= not w37633 and not w38286;
w38295 <= w37626 and not w38294;
w38296 <= not pi0219 and not w38295;
w38297 <= not w38293 and w38296;
w38298 <= w37873 and not w38297;
w38299 <= w37408 and not w38298;
w38300 <= not pi1152 and not w38281;
w38301 <= not w38299 and w38300;
w38302 <= pi0214 and w38287;
w38303 <= w37626 and not w38302;
w38304 <= not pi0214 and w38287;
w38305 <= w37878 and not w38304;
w38306 <= not pi0219 and not w38303;
w38307 <= not w38305 and w38306;
w38308 <= w37873 and not w38307;
w38309 <= w37434 and not w38308;
w38310 <= not w37668 and not w38198;
w38311 <= pi0214 and w38310;
w38312 <= w37671 and not w38311;
w38313 <= not pi0214 and w38310;
w38314 <= w37676 and not w38313;
w38315 <= not w38312 and not w38314;
w38316 <= not pi0219 and not w38315;
w38317 <= w37686 and not w38316;
w38318 <= w37456 and not w38317;
w38319 <= pi1152 and not w38309;
w38320 <= not w38318 and w38319;
w38321 <= pi1150 and not w38301;
w38322 <= not w38320 and w38321;
w38323 <= not pi1149 and not w38273;
w38324 <= not w38322 and w38323;
w38325 <= not w38257 and not w38324;
w38326 <= pi0213 and not w38325;
w38327 <= not pi0209 and not w38189;
w38328 <= not w38326 and w38327;
w38329 <= not w38169 and not w38328;
w38330 <= pi0230 and not w38329;
w38331 <= not pi0230 and not pi0241;
w38332 <= not w38330 and not w38331;
w38333 <= not pi0230 and not pi0242;
w38334 <= pi0219 and not w35982;
w38335 <= pi0214 and not w36977;
w38336 <= not pi0214 and not w37774;
w38337 <= not w38335 and not w38336;
w38338 <= pi0212 and not w38337;
w38339 <= not pi0212 and w37775;
w38340 <= not pi0219 and not w38339;
w38341 <= not w38338 and w38340;
w38342 <= w35979 and not w38334;
w38343 <= not w38341 and w38342;
w38344 <= pi0199 and pi1144;
w38345 <= not pi0200 and not w38344;
w38346 <= not w37896 and w38345;
w38347 <= not pi0299 and not w37893;
w38348 <= not w38346 and w38347;
w38349 <= w36389 and w38348;
w38350 <= not pi0207 and not w38348;
w38351 <= not pi0299 and not w36955;
w38352 <= not w36956 and w38345;
w38353 <= w38351 and not w38352;
w38354 <= pi0207 and not w38353;
w38355 <= pi0208 and not w38350;
w38356 <= not w38354 and w38355;
w38357 <= not w38349 and not w38356;
w38358 <= not pi0214 and w38357;
w38359 <= not pi0212 and not w38358;
w38360 <= w36012 and w38348;
w38361 <= not w37797 and not w38360;
w38362 <= not w38356 and w38361;
w38363 <= not pi0211 and not w38362;
w38364 <= not w37047 and not w38360;
w38365 <= not w38356 and w38364;
w38366 <= pi0211 and not w38365;
w38367 <= not w38363 and not w38366;
w38368 <= pi0214 and w38367;
w38369 <= w38359 and not w38368;
w38370 <= not pi0211 and not w38365;
w38371 <= not w36175 and not w38360;
w38372 <= not w38356 and w38371;
w38373 <= pi0211 and not w38372;
w38374 <= pi0214 and not w38370;
w38375 <= not w38373 and w38374;
w38376 <= not pi0214 and w38367;
w38377 <= pi0212 and not w38375;
w38378 <= not w38376 and w38377;
w38379 <= not pi0219 and not w38369;
w38380 <= not w38378 and w38379;
w38381 <= not w35977 and not w38357;
w38382 <= pi0219 and not w38381;
w38383 <= w35977 and not w38372;
w38384 <= w38382 and not w38383;
w38385 <= w4989 and not w38384;
w38386 <= not w38380 and w38385;
w38387 <= not w38343 and not w38386;
w38388 <= pi0213 and w38387;
w38389 <= w35976 and not w38349;
w38390 <= pi0211 and not w38349;
w38391 <= w35977 and not w36243;
w38392 <= not w38360 and w38391;
w38393 <= not w38390 and not w38392;
w38394 <= pi0219 and not w38393;
w38395 <= w8406 and not w36020;
w38396 <= not w35994 and w36171;
w38397 <= not w38395 and not w38396;
w38398 <= not pi0219 and not w38360;
w38399 <= not w38397 and w38398;
w38400 <= not w38389 and not w38399;
w38401 <= not w38394 and w38400;
w38402 <= not w38356 and not w38401;
w38403 <= w4989 and not w38402;
w38404 <= not pi0213 and not w35993;
w38405 <= not w38403 and w38404;
w38406 <= not w38388 and not w38405;
w38407 <= pi0209 and not w38406;
w38408 <= not pi0213 and not w36039;
w38409 <= pi0219 and w35976;
w38410 <= not w38334 and not w38409;
w38411 <= not w38341 and w38410;
w38412 <= pi0299 and not w38411;
w38413 <= w4989 and not w38412;
w38414 <= not w36031 and w38413;
w38415 <= not w38343 and not w38414;
w38416 <= pi0213 and not w38415;
w38417 <= not pi0209 and not w38416;
w38418 <= not w38408 and w38417;
w38419 <= not w38407 and not w38418;
w38420 <= pi0230 and not w38419;
w38421 <= not w38333 and not w38420;
w38422 <= pi0253 and pi0254;
w38423 <= pi0267 and w38422;
w38424 <= not pi0263 and w38423;
w38425 <= not pi0083 and not pi0085;
w38426 <= pi0314 and not w38425;
w38427 <= pi0802 and w38426;
w38428 <= pi0276 and w38427;
w38429 <= not pi1091 and w38428;
w38430 <= pi0271 and w38429;
w38431 <= pi0273 and w38430;
w38432 <= pi0243 and w38431;
w38433 <= not pi1091 and not w38428;
w38434 <= pi0271 and not w38433;
w38435 <= not pi1091 and not w38434;
w38436 <= pi0273 and not w38435;
w38437 <= not pi1091 and not w38436;
w38438 <= not pi0243 and w38437;
w38439 <= pi0243 and not pi1091;
w38440 <= w36041 and not w38439;
w38441 <= not w38429 and w38440;
w38442 <= not w38432 and not w38441;
w38443 <= not w38438 and w38442;
w38444 <= pi0219 and not w38443;
w38445 <= not w36042 and not w36050;
w38446 <= pi1091 and w38445;
w38447 <= not pi0081 and w38425;
w38448 <= pi0314 and not w38447;
w38449 <= pi0802 and w38448;
w38450 <= pi0276 and w38449;
w38451 <= not pi1091 and w38450;
w38452 <= pi0271 and w38451;
w38453 <= pi0273 and w38452;
w38454 <= not w38436 and not w38453;
w38455 <= w38439 and w38454;
w38456 <= not pi0243 and w38453;
w38457 <= not pi0219 and not w38446;
w38458 <= not w38456 and w38457;
w38459 <= not w38455 and w38458;
w38460 <= not w38444 and not w38459;
w38461 <= w38424 and not w38460;
w38462 <= not pi0243 and not pi1091;
w38463 <= not pi0219 and not w38445;
w38464 <= pi1157 and w36082;
w38465 <= not w38463 and not w38464;
w38466 <= pi1091 and not w38465;
w38467 <= not w38462 and not w38466;
w38468 <= not w38424 and not w38467;
w38469 <= not w4989 and not w38468;
w38470 <= not w38461 and w38469;
w38471 <= pi0272 and pi0283;
w38472 <= pi0275 and w38471;
w38473 <= pi0268 and w38472;
w38474 <= not pi0299 and pi1091;
w38475 <= w36404 and w38474;
w38476 <= not w38462 and not w38475;
w38477 <= pi1156 and not w38476;
w38478 <= pi1091 and not w36518;
w38479 <= w37020 and w38478;
w38480 <= not w38477 and not w38479;
w38481 <= not pi0299 and w36262;
w38482 <= pi1091 and not w38481;
w38483 <= not w38439 and not w38482;
w38484 <= not pi1155 and not w38462;
w38485 <= not w38439 and not w38484;
w38486 <= w36131 and w38485;
w38487 <= not w38483 and not w38486;
w38488 <= not pi1156 and not w38487;
w38489 <= w38480 and not w38488;
w38490 <= pi1157 and not w38489;
w38491 <= not w38478 and w38485;
w38492 <= not pi1156 and not w38491;
w38493 <= pi1155 and not w38439;
w38494 <= pi0199 and pi1091;
w38495 <= not pi0299 and w38494;
w38496 <= w38493 and not w38495;
w38497 <= pi1156 and not w38496;
w38498 <= not pi1155 and not w38439;
w38499 <= not w9007 and w38474;
w38500 <= w38498 and not w38499;
w38501 <= w38497 and not w38500;
w38502 <= not pi1157 and not w38492;
w38503 <= not w38501 and w38502;
w38504 <= not w38490 and not w38503;
w38505 <= pi0211 and not w38504;
w38506 <= pi1091 and not w9008;
w38507 <= w38498 and not w38506;
w38508 <= not w38496 and not w38507;
w38509 <= pi0200 and not pi1156;
w38510 <= w38474 and w38509;
w38511 <= not w38508 and not w38510;
w38512 <= not pi1157 and not w38511;
w38513 <= w38476 and w38497;
w38514 <= pi0200 and pi1091;
w38515 <= not pi0299 and w38514;
w38516 <= w38493 and not w38515;
w38517 <= not pi1155 and w38483;
w38518 <= not pi1156 and not w38516;
w38519 <= not w38517 and w38518;
w38520 <= not w38513 and not w38519;
w38521 <= pi1157 and not w38520;
w38522 <= not pi0211 and not w38512;
w38523 <= not w38521 and w38522;
w38524 <= not w38505 and not w38523;
w38525 <= not pi0219 and not w38524;
w38526 <= w36932 and not w38477;
w38527 <= not w38488 and w38526;
w38528 <= pi0299 and pi1091;
w38529 <= w38511 and not w38528;
w38530 <= not pi1157 and not w38529;
w38531 <= pi1091 and w36263;
w38532 <= w38498 and not w38531;
w38533 <= not w38516 and not w38532;
w38534 <= not pi1156 and not w38533;
w38535 <= w36041 and not w38534;
w38536 <= w38480 and w38535;
w38537 <= pi0219 and not w38527;
w38538 <= not w38530 and not w38536;
w38539 <= w38537 and w38538;
w38540 <= not w38525 and not w38539;
w38541 <= not w38424 and not w38540;
w38542 <= pi0199 and not w38437;
w38543 <= not pi1091 and w38454;
w38544 <= not pi0199 and not w38543;
w38545 <= not w38542 and not w38544;
w38546 <= not pi0200 and not w38451;
w38547 <= not w38545 and not w38546;
w38548 <= not pi0299 and not w38547;
w38549 <= pi0299 and w38437;
w38550 <= not w38453 and w38549;
w38551 <= not w38548 and not w38550;
w38552 <= not pi0243 and not w38551;
w38553 <= not pi0200 and not w38437;
w38554 <= w38451 and not w38545;
w38555 <= not pi0299 and not w38554;
w38556 <= not w38553 and w38555;
w38557 <= pi0299 and not w38431;
w38558 <= not w38556 and not w38557;
w38559 <= pi0243 and w38558;
w38560 <= not w38552 and not w38559;
w38561 <= pi1155 and not w38560;
w38562 <= not w38544 and w38548;
w38563 <= not w38549 and not w38562;
w38564 <= not pi0243 and not w38563;
w38565 <= not w38542 and w38555;
w38566 <= w38558 and not w38565;
w38567 <= pi0243 and w38566;
w38568 <= not w38564 and not w38567;
w38569 <= not w38561 and w38568;
w38570 <= not pi1156 and not w38569;
w38571 <= not w38553 and w38565;
w38572 <= not w38549 and not w38571;
w38573 <= not pi0243 and w38572;
w38574 <= not w38542 and w38548;
w38575 <= not w38544 and w38556;
w38576 <= not w38557 and not w38575;
w38577 <= not w38574 and w38576;
w38578 <= pi0243 and not w38577;
w38579 <= not w38573 and not w38578;
w38580 <= not pi1155 and not w38564;
w38581 <= pi1155 and not w38552;
w38582 <= pi0243 and w38576;
w38583 <= w38581 and not w38582;
w38584 <= not w38580 and not w38583;
w38585 <= not w38579 and not w38584;
w38586 <= pi1156 and not w38585;
w38587 <= w36932 and not w38570;
w38588 <= not w38586 and w38587;
w38589 <= not w38544 and w38555;
w38590 <= w38559 and not w38589;
w38591 <= not w38549 and not w38574;
w38592 <= not pi0243 and not w38591;
w38593 <= pi1155 and not w38592;
w38594 <= not w38590 and w38593;
w38595 <= not w38555 and not w38557;
w38596 <= w38462 and not w38595;
w38597 <= not pi1155 and not w38596;
w38598 <= pi0243 and w38595;
w38599 <= w38597 and not w38598;
w38600 <= not pi1156 and not w38599;
w38601 <= not w38594 and w38600;
w38602 <= not w38557 and not w38589;
w38603 <= pi1155 and w38602;
w38604 <= not w38548 and w38602;
w38605 <= not w38603 and not w38604;
w38606 <= pi0243 and not w38605;
w38607 <= pi0299 and not w38453;
w38608 <= not w38556 and not w38607;
w38609 <= not pi1155 and w38608;
w38610 <= not w38451 and w38609;
w38611 <= not w38549 and not w38565;
w38612 <= not pi0243 and not w38611;
w38613 <= not w38610 and w38612;
w38614 <= not w38606 and not w38613;
w38615 <= pi1156 and not w38614;
w38616 <= not pi1157 and not w38601;
w38617 <= not w38615 and w38616;
w38618 <= not w38549 and not w38556;
w38619 <= pi0243 and not w38618;
w38620 <= not w38557 and not w38562;
w38621 <= not pi0243 and not w38620;
w38622 <= pi0243 and not w38565;
w38623 <= not pi1155 and not w38622;
w38624 <= not w38621 and w38623;
w38625 <= not w38548 and not w38557;
w38626 <= not pi0243 and pi1155;
w38627 <= w38625 and w38626;
w38628 <= not pi1156 and not w38627;
w38629 <= not w38619 and w38628;
w38630 <= not w38624 and w38629;
w38631 <= not w38577 and w38619;
w38632 <= pi1155 and not w38631;
w38633 <= w38573 and w38625;
w38634 <= w38632 and not w38633;
w38635 <= not w38571 and not w38607;
w38636 <= not w38439 and not w38635;
w38637 <= not w38564 and not w38636;
w38638 <= not w38579 and w38637;
w38639 <= not pi1155 and not w38638;
w38640 <= not w38634 and not w38639;
w38641 <= pi1156 and not w38640;
w38642 <= w36041 and not w38630;
w38643 <= not w38641 and w38642;
w38644 <= not w38588 and not w38617;
w38645 <= not w38643 and w38644;
w38646 <= pi0219 and not w38645;
w38647 <= not w38555 and not w38607;
w38648 <= not pi1155 and w38647;
w38649 <= not w38580 and not w38648;
w38650 <= pi0243 and w38608;
w38651 <= not w38565 and w38650;
w38652 <= not w38649 and not w38651;
w38653 <= not pi1156 and not w38652;
w38654 <= not w38548 and not w38607;
w38655 <= not pi0243 and w38654;
w38656 <= not w38550 and not w38556;
w38657 <= pi0243 and not w38656;
w38658 <= not w38655 and not w38657;
w38659 <= w38653 and w38658;
w38660 <= not w38550 and not w38575;
w38661 <= pi1155 and w38660;
w38662 <= not w38632 and not w38661;
w38663 <= not w38571 and w38655;
w38664 <= not w38662 and not w38663;
w38665 <= not w38562 and not w38571;
w38666 <= not w38550 and w38665;
w38667 <= not pi0243 and not w38666;
w38668 <= not w38574 and not w38607;
w38669 <= pi0243 and not w38575;
w38670 <= w38668 and w38669;
w38671 <= not w38667 and not w38670;
w38672 <= not pi1155 and not w38671;
w38673 <= not w38664 and not w38672;
w38674 <= pi1156 and not w38673;
w38675 <= pi1157 and not w38659;
w38676 <= not w38674 and w38675;
w38677 <= not pi1155 and w38656;
w38678 <= not w38654 and w38677;
w38679 <= not w38550 and not w38589;
w38680 <= pi0243 and not w38679;
w38681 <= not w38565 and not w38607;
w38682 <= not pi0243 and w38681;
w38683 <= not w38680 and not w38682;
w38684 <= pi1156 and not w38610;
w38685 <= w38683 and w38684;
w38686 <= not w38678 and w38685;
w38687 <= pi0243 and w38647;
w38688 <= not w38597 and not w38648;
w38689 <= not w38687 and not w38688;
w38690 <= not pi1156 and not w38689;
w38691 <= w38658 and w38683;
w38692 <= pi1155 and not w38691;
w38693 <= w38690 and not w38692;
w38694 <= not pi1157 and not w38686;
w38695 <= not w38693 and w38694;
w38696 <= not pi0211 and not w38695;
w38697 <= not w38676 and w38696;
w38698 <= w38581 and not w38650;
w38699 <= w38493 and w38542;
w38700 <= not w38698 and not w38699;
w38701 <= w38690 and w38700;
w38702 <= not pi1157 and not w38685;
w38703 <= not w38701 and w38702;
w38704 <= w38653 and not w38698;
w38705 <= not w38636 and w38673;
w38706 <= pi1156 and not w38705;
w38707 <= pi1157 and not w38704;
w38708 <= not w38706 and w38707;
w38709 <= pi0211 and not w38703;
w38710 <= not w38708 and w38709;
w38711 <= not pi0219 and not w38697;
w38712 <= not w38710 and w38711;
w38713 <= w38424 and not w38646;
w38714 <= not w38712 and w38713;
w38715 <= w4989 and not w38541;
w38716 <= not w38714 and w38715;
w38717 <= not w38470 and w38473;
w38718 <= not w38716 and w38717;
w38719 <= w4989 and w38540;
w38720 <= not w4989 and w38467;
w38721 <= not w38473 and not w38720;
w38722 <= not w38719 and w38721;
w38723 <= not pi0230 and not w38722;
w38724 <= not w38718 and w38723;
w38725 <= not w14042 and not w38465;
w38726 <= pi0199 and not w37030;
w38727 <= not w36403 and not w38509;
w38728 <= not w38726 and w38727;
w38729 <= w14042 and w38728;
w38730 <= pi0230 and not w38725;
w38731 <= not w38729 and w38730;
w38732 <= not w38724 and not w38731;
w38733 <= not pi0230 and not pi0244;
w38734 <= pi0213 and not w37968;
w38735 <= not pi0211 and not w36106;
w38736 <= not w37920 and w38735;
w38737 <= not w37909 and not w38736;
w38738 <= w37907 and not w38737;
w38739 <= not w36173 and w37953;
w38740 <= not w37946 and not w38739;
w38741 <= not w37974 and not w38740;
w38742 <= pi0214 and not w38741;
w38743 <= w37927 and not w38742;
w38744 <= w35983 and w37856;
w38745 <= not pi0214 and w38740;
w38746 <= pi0212 and not w38744;
w38747 <= not w38745 and w38746;
w38748 <= not w37974 and w38747;
w38749 <= not pi0219 and not w38743;
w38750 <= not w38748 and w38749;
w38751 <= w38010 and not w38738;
w38752 <= not w38750 and w38751;
w38753 <= pi0299 and w36973;
w38754 <= pi0214 and w38740;
w38755 <= w37951 and not w38754;
w38756 <= not w37944 and w38747;
w38757 <= not pi0219 and not w38755;
w38758 <= not w38756 and w38757;
w38759 <= pi1147 and not w38753;
w38760 <= w37973 and w38759;
w38761 <= not w38758 and w38760;
w38762 <= not pi0213 and not w36983;
w38763 <= not w38761 and w38762;
w38764 <= not w38752 and w38763;
w38765 <= not w38734 and not w38764;
w38766 <= pi0209 and not w38765;
w38767 <= not pi0213 and not w36990;
w38768 <= w37807 and not w37810;
w38769 <= not w37787 and not w38768;
w38770 <= not w8406 and w37799;
w38771 <= w8406 and not w37794;
w38772 <= w37807 and not w37809;
w38773 <= w36228 and not w38770;
w38774 <= not w38771 and w38773;
w38775 <= not w38772 and w38774;
w38776 <= not w36961 and not w37816;
w38777 <= not w38775 and w38776;
w38778 <= w4989 and not w38777;
w38779 <= not w38769 and not w38778;
w38780 <= pi0213 and not w38779;
w38781 <= not pi0209 and not w38767;
w38782 <= not w38780 and w38781;
w38783 <= not w38766 and not w38782;
w38784 <= pi0230 and not w38783;
w38785 <= not w38733 and not w38784;
w38786 <= not pi0213 and not w38387;
w38787 <= pi1146 and w37432;
w38788 <= not pi1147 and not w38787;
w38789 <= w37428 and not w37708;
w38790 <= w38788 and not w38789;
w38791 <= not w35976 and w38363;
w38792 <= w38382 and not w38791;
w38793 <= w4989 and not w38792;
w38794 <= pi0214 and not w37798;
w38795 <= not pi0299 and not w38367;
w38796 <= w38794 and not w38795;
w38797 <= pi0212 and not w38796;
w38798 <= not pi0299 and w38365;
w38799 <= not pi0211 and not w38798;
w38800 <= w38357 and not w38799;
w38801 <= not pi0214 and w38800;
w38802 <= w38797 and not w38801;
w38803 <= w38359 and not w38800;
w38804 <= not pi0219 and not w38803;
w38805 <= not w38802 and w38804;
w38806 <= w38793 and not w38805;
w38807 <= w38790 and not w38806;
w38808 <= pi1147 and not w37428;
w38809 <= not w38787 and w38808;
w38810 <= pi0211 and not w38362;
w38811 <= not w38799 and not w38810;
w38812 <= pi0214 and not w38811;
w38813 <= not pi0214 and not w38798;
w38814 <= not w38812 and not w38813;
w38815 <= pi0212 and not w38814;
w38816 <= w38359 and not w38798;
w38817 <= not pi0219 and not w38816;
w38818 <= not w38815 and w38817;
w38819 <= w38793 and not w38818;
w38820 <= w38809 and not w38819;
w38821 <= pi1148 and not w38807;
w38822 <= not w38820 and w38821;
w38823 <= not w37970 and not w38809;
w38824 <= not w10624 and w38357;
w38825 <= not pi0214 and not w38824;
w38826 <= not w38812 and not w38825;
w38827 <= pi0212 and not w38826;
w38828 <= w38359 and not w38824;
w38829 <= not pi0219 and not w38828;
w38830 <= not w38827 and w38829;
w38831 <= w38793 and not w38830;
w38832 <= not w38823 and not w38831;
w38833 <= not w38358 and w38797;
w38834 <= not pi0212 and not w38357;
w38835 <= not pi0219 and not w38834;
w38836 <= not w38833 and w38835;
w38837 <= w38793 and not w38836;
w38838 <= w38788 and not w38837;
w38839 <= not pi1148 and not w38832;
w38840 <= not w38838 and w38839;
w38841 <= not w38822 and not w38840;
w38842 <= pi0213 and not w38841;
w38843 <= not pi0209 and not w38786;
w38844 <= not w38842 and w38843;
w38845 <= pi0199 and pi1146;
w38846 <= w36262 and not w38845;
w38847 <= w36113 and not w38846;
w38848 <= not w8050 and not w38847;
w38849 <= w37902 and not w38846;
w38850 <= pi0207 and w38849;
w38851 <= not w36389 and not w38850;
w38852 <= not w38848 and not w38851;
w38853 <= not w35977 and w38852;
w38854 <= pi0219 and not w38853;
w38855 <= w36012 and w38847;
w38856 <= pi0208 and w38849;
w38857 <= not pi0200 and not w38845;
w38858 <= w36113 and not w38857;
w38859 <= not pi0207 and w38858;
w38860 <= not w37797 and not w38859;
w38861 <= not w38850 and w38860;
w38862 <= pi0208 and not w38861;
w38863 <= not pi0299 and w38862;
w38864 <= not w38855 and not w38856;
w38865 <= not w38863 and w38864;
w38866 <= not w37797 and w38865;
w38867 <= w35977 and not w38866;
w38868 <= w38854 and not w38867;
w38869 <= not pi0214 and not w38852;
w38870 <= not pi0212 and not w38869;
w38871 <= not pi0299 and w38865;
w38872 <= w38870 and not w38871;
w38873 <= not pi0219 and not w38872;
w38874 <= pi0212 and not w38871;
w38875 <= w8047 and w38866;
w38876 <= w38874 and not w38875;
w38877 <= w38873 and not w38876;
w38878 <= w4989 and not w38868;
w38879 <= not w38877 and w38878;
w38880 <= w38809 and not w38879;
w38881 <= not pi0208 and w37797;
w38882 <= w37902 and not w38857;
w38883 <= pi0207 and w38882;
w38884 <= pi1146 and not w36263;
w38885 <= not w38883 and not w38884;
w38886 <= pi0208 and not w38885;
w38887 <= not pi0207 and not w38856;
w38888 <= w37221 and not w38846;
w38889 <= not w38887 and w38888;
w38890 <= not w38881 and not w38886;
w38891 <= not w38889 and w38890;
w38892 <= not pi0299 and not w38891;
w38893 <= not pi0214 and not w38892;
w38894 <= not pi0212 and not w38893;
w38895 <= not w8050 and not w37222;
w38896 <= w38882 and not w38895;
w38897 <= pi0211 and not w38896;
w38898 <= not pi0299 and not w38882;
w38899 <= not w38891 and not w38898;
w38900 <= not pi0299 and not w38899;
w38901 <= not pi0211 and w38900;
w38902 <= not w38897 and not w38901;
w38903 <= not w38892 and not w38902;
w38904 <= w38894 and not w38903;
w38905 <= not pi0219 and not w38904;
w38906 <= w38794 and not w38892;
w38907 <= not pi0214 and w38903;
w38908 <= pi0212 and not w38907;
w38909 <= not w38906 and w38908;
w38910 <= w38905 and not w38909;
w38911 <= not w35977 and w38892;
w38912 <= pi0219 and not w38911;
w38913 <= w35977 and not w38891;
w38914 <= w38912 and not w38913;
w38915 <= w4989 and not w38914;
w38916 <= not w38910 and w38915;
w38917 <= w38790 and not w38916;
w38918 <= pi1148 and not w38880;
w38919 <= not w38917 and w38918;
w38920 <= not w38226 and not w38892;
w38921 <= not w38885 and not w38920;
w38922 <= not pi0219 and not w38921;
w38923 <= pi0219 and not w38896;
w38924 <= not w36533 and not w38923;
w38925 <= not w35976 and not w38897;
w38926 <= w38899 and w38925;
w38927 <= not w38924 and not w38926;
w38928 <= w4989 and not w38927;
w38929 <= not w38922 and w38928;
w38930 <= w38788 and not w38929;
w38931 <= not w8050 and not w38858;
w38932 <= not w38851 and not w38931;
w38933 <= not w10624 and not w38932;
w38934 <= pi0214 and not w38933;
w38935 <= not pi0214 and w38932;
w38936 <= not pi0212 and not w38935;
w38937 <= not w38934 and w38936;
w38938 <= not pi0214 and not w38933;
w38939 <= w36012 and w38858;
w38940 <= not w38881 and not w38939;
w38941 <= not w38862 and w38940;
w38942 <= not pi0299 and w38941;
w38943 <= pi0214 and not w38942;
w38944 <= not pi0211 and not w38871;
w38945 <= not w38852 and not w38944;
w38946 <= w38943 and not w38945;
w38947 <= pi0212 and not w38946;
w38948 <= not w38938 and w38947;
w38949 <= not w38937 and not w38948;
w38950 <= not pi0219 and not w38949;
w38951 <= not pi1146 and not w36346;
w38952 <= w37862 and not w38951;
w38953 <= w38950 and not w38952;
w38954 <= not w35976 and w38932;
w38955 <= not w35977 and not w38954;
w38956 <= not w38941 and not w38955;
w38957 <= not pi0212 and w38935;
w38958 <= pi0219 and not w38957;
w38959 <= not w38956 and w38958;
w38960 <= w4989 and not w38959;
w38961 <= not w38953 and w38960;
w38962 <= not w38823 and not w38961;
w38963 <= not pi1148 and not w38930;
w38964 <= not w38962 and w38963;
w38965 <= not w38919 and not w38964;
w38966 <= pi0213 and not w38965;
w38967 <= pi1147 and w4989;
w38968 <= not w36175 and w38865;
w38969 <= w35977 and not w38968;
w38970 <= w38854 and not w38969;
w38971 <= not w37794 and w38865;
w38972 <= pi0214 and w38971;
w38973 <= w38870 and not w38972;
w38974 <= pi0299 and not w38337;
w38975 <= w38865 and not w38974;
w38976 <= pi0212 and not w38975;
w38977 <= not pi0219 and not w38976;
w38978 <= not w38973 and w38977;
w38979 <= w38967 and not w38970;
w38980 <= not w38978 and w38979;
w38981 <= not pi0299 and w38891;
w38982 <= w35977 and not w38981;
w38983 <= not w36173 and w38982;
w38984 <= w38912 and not w38983;
w38985 <= not w37794 and not w38892;
w38986 <= w38894 and not w38985;
w38987 <= not w38892 and not w38974;
w38988 <= pi0212 and not w38987;
w38989 <= not pi0219 and not w38988;
w38990 <= not w38986 and w38989;
w38991 <= w38010 and not w38984;
w38992 <= not w38990 and w38991;
w38993 <= pi1148 and not w38343;
w38994 <= not w38980 and w38993;
w38995 <= not w38992 and w38994;
w38996 <= not w38942 and w38976;
w38997 <= w38943 and not w38971;
w38998 <= not w38935 and not w38997;
w38999 <= not pi0212 and not w38998;
w39000 <= not pi0219 and not w38996;
w39001 <= not w38999 and w39000;
w39002 <= not w38942 and not w38968;
w39003 <= not pi0211 and not w39002;
w39004 <= not w38955 and not w39003;
w39005 <= w38958 and not w39004;
w39006 <= w38967 and not w39001;
w39007 <= not w39005 and w39006;
w39008 <= not w38898 and w38988;
w39009 <= not pi0214 and w38896;
w39010 <= pi0214 and not w38900;
w39011 <= not w38985 and w39010;
w39012 <= not w39009 and not w39011;
w39013 <= not pi0212 and not w39012;
w39014 <= not pi0219 and not w39008;
w39015 <= not w39013 and w39014;
w39016 <= not w36173 and not w38900;
w39017 <= not pi0211 and not w39016;
w39018 <= w38925 and not w39017;
w39019 <= not w38924 and not w39018;
w39020 <= w38010 and not w39019;
w39021 <= not w39015 and w39020;
w39022 <= not pi1148 and not w38343;
w39023 <= not w39007 and w39022;
w39024 <= not w39021 and w39023;
w39025 <= not pi0213 and not w38995;
w39026 <= not w39024 and w39025;
w39027 <= pi0209 and not w39026;
w39028 <= not w38966 and w39027;
w39029 <= not w38844 and not w39028;
w39030 <= pi0230 and not w39029;
w39031 <= not pi0230 and not pi0245;
w39032 <= not w39030 and not w39031;
w39033 <= not pi1150 and w37697;
w39034 <= pi1150 and w37652;
w39035 <= pi1149 and not w39033;
w39036 <= not w39034 and w39035;
w39037 <= not pi1150 and w37763;
w39038 <= pi1150 and w37729;
w39039 <= not pi1149 and not w39037;
w39040 <= not w39038 and w39039;
w39041 <= not w39036 and not w39040;
w39042 <= pi1148 and not w39041;
w39043 <= not pi1150 and w37688;
w39044 <= pi1150 and w37641;
w39045 <= pi1149 and not w39044;
w39046 <= not w39043 and w39045;
w39047 <= not pi1149 and pi1150;
w39048 <= not w37706 and w39047;
w39049 <= not w39046 and not w39048;
w39050 <= not pi1148 and not w39049;
w39051 <= not w39042 and not w39050;
w39052 <= pi0213 and not w39051;
w39053 <= not w37747 and not w37756;
w39054 <= w38790 and not w39053;
w39055 <= not w38790 and not w38809;
w39056 <= pi0219 and not w37797;
w39057 <= w37647 and not w39056;
w39058 <= w37690 and not w37744;
w39059 <= not w39057 and not w39058;
w39060 <= not w37746 and not w37818;
w39061 <= w35986 and not w39060;
w39062 <= not w38211 and not w39061;
w39063 <= not pi0219 and not w39062;
w39064 <= not w39059 and not w39063;
w39065 <= not w39055 and not w39064;
w39066 <= not pi1150 and not w39054;
w39067 <= not w39065 and w39066;
w39068 <= not w37832 and not w39057;
w39069 <= not pi0214 and w37260;
w39070 <= pi0214 and not w37710;
w39071 <= not w37837 and w39070;
w39072 <= pi0212 and not w39069;
w39073 <= not w39071 and w39072;
w39074 <= w37719 and not w39073;
w39075 <= not w39068 and not w39074;
w39076 <= w38790 and not w39075;
w39077 <= not w37839 and w38076;
w39078 <= not pi0212 and not w37224;
w39079 <= not pi0219 and not w39078;
w39080 <= not w38088 and w39079;
w39081 <= not w39077 and w39080;
w39082 <= not w39068 and not w39081;
w39083 <= w38809 and not w39082;
w39084 <= pi1150 and not w39076;
w39085 <= not w39083 and w39084;
w39086 <= not w39067 and not w39085;
w39087 <= pi1148 and not w39086;
w39088 <= pi1150 and w37202;
w39089 <= pi0299 and w37656;
w39090 <= not pi0219 and not w39089;
w39091 <= not w38952 and w39090;
w39092 <= not w39088 and w39091;
w39093 <= not w38823 and w39092;
w39094 <= not pi0219 and not w37776;
w39095 <= not w38227 and not w39094;
w39096 <= w39057 and w39095;
w39097 <= w38788 and not w39096;
w39098 <= not w38823 and not w39057;
w39099 <= not w39097 and not w39098;
w39100 <= pi1150 and w37703;
w39101 <= not w39099 and not w39100;
w39102 <= not pi1148 and not w39093;
w39103 <= not w39101 and w39102;
w39104 <= not w39087 and not w39103;
w39105 <= not pi1149 and not w39104;
w39106 <= not pi1146 and w37685;
w39107 <= w37647 and not w37668;
w39108 <= not w37686 and not w39107;
w39109 <= w37776 and w37856;
w39110 <= not w37663 and not w39109;
w39111 <= w37684 and w39110;
w39112 <= not w39106 and not w39108;
w39113 <= not w39111 and w39112;
w39114 <= not w38823 and not w39113;
w39115 <= not w37665 and not w38087;
w39116 <= not pi0219 and not w39115;
w39117 <= not w39108 and not w39116;
w39118 <= not pi1146 and not w37663;
w39119 <= w39117 and not w39118;
w39120 <= w38788 and not w39119;
w39121 <= not pi1150 and not w39120;
w39122 <= not w39114 and w39121;
w39123 <= not w37874 and not w39057;
w39124 <= not w37625 and not w38288;
w39125 <= not pi0214 and w38288;
w39126 <= w37637 and not w39125;
w39127 <= not pi0219 and not w39126;
w39128 <= not w39124 and w39127;
w39129 <= not pi0212 and w39124;
w39130 <= w39127 and not w39129;
w39131 <= not pi0299 and w37276;
w39132 <= not w37627 and not w37797;
w39133 <= not w39131 and w39132;
w39134 <= w39130 and w39133;
w39135 <= not w39123 and not w39128;
w39136 <= not w39134 and w39135;
w39137 <= not w37623 and not w39136;
w39138 <= w37626 and not w37636;
w39139 <= not pi0219 and not w39138;
w39140 <= not w38292 and w39139;
w39141 <= w37873 and not w39140;
w39142 <= not w39137 and w39141;
w39143 <= w38788 and not w39142;
w39144 <= not w38823 and not w39136;
w39145 <= pi1150 and not w39144;
w39146 <= not w39143 and w39145;
w39147 <= not pi1148 and not w39146;
w39148 <= not w39122 and w39147;
w39149 <= not w37690 and not w39057;
w39150 <= w37310 and w38794;
w39151 <= w37752 and not w39150;
w39152 <= not w37735 and w37753;
w39153 <= not w37740 and not w39152;
w39154 <= not w38790 and not w39153;
w39155 <= w37755 and not w39151;
w39156 <= not w39154 and w39155;
w39157 <= not w39149 and not w39156;
w39158 <= not w39055 and not w39157;
w39159 <= not pi1150 and not w39158;
w39160 <= not w37866 and not w39096;
w39161 <= w38790 and w39160;
w39162 <= pi0214 and w37855;
w39163 <= w37861 and not w39162;
w39164 <= not pi0219 and not w37858;
w39165 <= not w39163 and w39164;
w39166 <= w37854 and not w39165;
w39167 <= pi1146 and w37648;
w39168 <= w38809 and not w39167;
w39169 <= not w39166 and w39168;
w39170 <= pi1150 and not w39169;
w39171 <= not w39161 and w39170;
w39172 <= pi1148 and not w39171;
w39173 <= not w39159 and w39172;
w39174 <= pi1149 and not w39173;
w39175 <= not w39148 and w39174;
w39176 <= not w39105 and not w39175;
w39177 <= not pi0213 and not w39176;
w39178 <= pi0209 and not w39052;
w39179 <= not w39177 and w39178;
w39180 <= not pi0213 and not w38965;
w39181 <= pi0219 and not w38932;
w39182 <= w38967 and not w39181;
w39183 <= not w38950 and w39182;
w39184 <= not pi0212 and not w39009;
w39185 <= not w10624 and not w38896;
w39186 <= pi0214 and not w39185;
w39187 <= w39184 and not w39186;
w39188 <= not pi0214 and not w39185;
w39189 <= pi0214 and w38902;
w39190 <= pi0212 and not w39189;
w39191 <= not w39188 and w39190;
w39192 <= not w39187 and not w39191;
w39193 <= not pi0219 and not w39192;
w39194 <= w38010 and not w38923;
w39195 <= not w39193 and w39194;
w39196 <= not pi1150 and not w37659;
w39197 <= not w39183 and w39196;
w39198 <= not w39195 and w39197;
w39199 <= w38936 and not w38943;
w39200 <= not pi0214 and not w38942;
w39201 <= w38947 and not w39200;
w39202 <= not w39199 and not w39201;
w39203 <= not pi0219 and not w39202;
w39204 <= not w39181 and not w39203;
w39205 <= pi1147 and not w39204;
w39206 <= not w39010 and w39184;
w39207 <= not pi0214 and not w38900;
w39208 <= w39190 and not w39207;
w39209 <= not w39206 and not w39208;
w39210 <= not pi0219 and not w39209;
w39211 <= not w38923 and not w39210;
w39212 <= not pi1147 and not w39211;
w39213 <= w4989 and not w39205;
w39214 <= not w39212 and w39213;
w39215 <= pi1150 and not w37428;
w39216 <= not w39214 and w39215;
w39217 <= not w39198 and not w39216;
w39218 <= pi1149 and not w39217;
w39219 <= pi1150 and w37770;
w39220 <= w38896 and not w39219;
w39221 <= not pi1147 and not w39220;
w39222 <= pi1147 and not w38932;
w39223 <= w4989 and not w39221;
w39224 <= not w39222 and w39223;
w39225 <= not pi1147 and w38899;
w39226 <= w14042 and not w39225;
w39227 <= w39219 and not w39226;
w39228 <= not pi1149 and not w39224;
w39229 <= not w39227 and w39228;
w39230 <= not w39218 and not w39229;
w39231 <= not pi1148 and not w39230;
w39232 <= not w35976 and w38944;
w39233 <= w38854 and not w39232;
w39234 <= w38967 and not w39233;
w39235 <= pi0214 and not w10624;
w39236 <= w38865 and w39235;
w39237 <= pi0212 and not w39236;
w39238 <= not w38869 and w39237;
w39239 <= not pi0212 and w38852;
w39240 <= not pi0219 and not w39239;
w39241 <= not w39238 and w39240;
w39242 <= w39234 and not w39241;
w39243 <= w38912 and not w38982;
w39244 <= w38010 and not w39243;
w39245 <= not pi0219 and w38920;
w39246 <= w39244 and not w39245;
w39247 <= not pi1150 and not w37432;
w39248 <= not w39242 and w39247;
w39249 <= not w39246 and w39248;
w39250 <= not w38892 and w39185;
w39251 <= pi0214 and w39250;
w39252 <= w38908 and not w39251;
w39253 <= w38905 and not w39252;
w39254 <= w39244 and not w39253;
w39255 <= not pi0214 and w38945;
w39256 <= w39237 and not w39255;
w39257 <= w38870 and not w38945;
w39258 <= not pi0219 and not w39257;
w39259 <= not w39256 and w39258;
w39260 <= w39234 and not w39259;
w39261 <= pi1150 and not w37709;
w39262 <= not w39260 and w39261;
w39263 <= not w39254 and w39262;
w39264 <= not pi1149 and not w39249;
w39265 <= not w39263 and w39264;
w39266 <= pi0057 and w36229;
w39267 <= not w3868 and not w36229;
w39268 <= w38873 and not w38874;
w39269 <= not w39233 and not w39268;
w39270 <= w3868 and w39269;
w39271 <= not pi0057 and pi1147;
w39272 <= not w39267 and w39271;
w39273 <= not w39270 and w39272;
w39274 <= w3868 and not w36228;
w39275 <= w38911 and w39274;
w39276 <= not w36229 and not w38981;
w39277 <= not pi0057 and not pi1147;
w39278 <= not w39267 and w39277;
w39279 <= not w39276 and w39278;
w39280 <= not w39275 and w39279;
w39281 <= not w39266 and not w39280;
w39282 <= not w39273 and w39281;
w39283 <= pi1150 and not w39282;
w39284 <= w38894 and not w39251;
w39285 <= not w39010 and w39250;
w39286 <= pi0212 and not w39285;
w39287 <= not pi0219 and not w39284;
w39288 <= not w39286 and w39287;
w39289 <= w39244 and not w39288;
w39290 <= not w38239 and w38967;
w39291 <= w39269 and w39290;
w39292 <= not pi1150 and not w37694;
w39293 <= not w39291 and w39292;
w39294 <= not w39289 and w39293;
w39295 <= pi1149 and not w39294;
w39296 <= not w39283 and w39295;
w39297 <= pi1148 and not w39296;
w39298 <= not w39265 and w39297;
w39299 <= pi0213 and not w39298;
w39300 <= not w39231 and w39299;
w39301 <= not pi0209 and not w39180;
w39302 <= not w39300 and w39301;
w39303 <= not w39179 and not w39302;
w39304 <= pi0230 and not w39303;
w39305 <= not pi0230 and not pi0246;
w39306 <= not w39304 and not w39305;
w39307 <= pi0213 and w38188;
w39308 <= pi1151 and not w37694;
w39309 <= w37873 and not w39128;
w39310 <= w39308 and not w39309;
w39311 <= w37667 and not w37682;
w39312 <= not w39108 and not w39311;
w39313 <= not w37694 and not w39312;
w39314 <= not pi1151 and w39313;
w39315 <= pi1147 and not w39310;
w39316 <= not w39314 and w39315;
w39317 <= not pi1147 and not w38172;
w39318 <= pi1151 and not w37659;
w39319 <= not w37624 and not w39130;
w39320 <= w39318 and not w39319;
w39321 <= w39317 and not w39320;
w39322 <= not pi1149 and not w39316;
w39323 <= not w39321 and w39322;
w39324 <= pi1147 and not w38178;
w39325 <= not w37645 and not w37648;
w39326 <= w38235 and w39325;
w39327 <= w39324 and not w39326;
w39328 <= not pi1151 and not w37428;
w39329 <= w37755 and not w39152;
w39330 <= w38243 and not w39329;
w39331 <= not w37741 and w38243;
w39332 <= not w39330 and not w39331;
w39333 <= w39328 and w39332;
w39334 <= w38063 and not w39166;
w39335 <= not pi1147 and not w39334;
w39336 <= not w39333 and w39335;
w39337 <= pi1149 and not w39327;
w39338 <= not w39336 and w39337;
w39339 <= pi1150 and not w39338;
w39340 <= not w39323 and w39339;
w39341 <= not w37658 and w37704;
w39342 <= not pi1151 and not w39341;
w39343 <= not pi1147 and not w39342;
w39344 <= w37393 and not w38096;
w39345 <= w39318 and not w39344;
w39346 <= w39343 and not w39345;
w39347 <= not w38267 and w39308;
w39348 <= not w37695 and w38140;
w39349 <= pi1147 and not w39348;
w39350 <= not w39347 and w39349;
w39351 <= not pi1149 and not w39346;
w39352 <= not w39350 and w39351;
w39353 <= pi0212 and not w37249;
w39354 <= w39080 and not w39353;
w39355 <= w37727 and not w39354;
w39356 <= w38156 and not w39355;
w39357 <= pi1147 and not w39356;
w39358 <= w35986 and not w37736;
w39359 <= not w37746 and w38216;
w39360 <= not w39358 and w39359;
w39361 <= not pi1151 and not w37645;
w39362 <= not w39360 and w39361;
w39363 <= not w37761 and w39362;
w39364 <= w39357 and not w39363;
w39365 <= w39328 and not w39360;
w39366 <= not w38077 and w39080;
w39367 <= w37832 and not w39366;
w39368 <= not w37428 and not w39367;
w39369 <= pi1151 and w39368;
w39370 <= not pi1147 and not w39365;
w39371 <= not w39369 and w39370;
w39372 <= pi1149 and not w39371;
w39373 <= not w39364 and w39372;
w39374 <= not pi1150 and not w39352;
w39375 <= not w39373 and w39374;
w39376 <= not w39340 and not w39375;
w39377 <= pi1148 and not w39376;
w39378 <= not pi1151 and not w37806;
w39379 <= not pi1147 and not w39378;
w39380 <= pi1151 and not w37623;
w39381 <= w39379 and not w39380;
w39382 <= not w39140 and w39309;
w39383 <= w37433 and not w39382;
w39384 <= not w37432 and not w39117;
w39385 <= not pi1151 and w39384;
w39386 <= pi1147 and not w39385;
w39387 <= not w39383 and w39386;
w39388 <= pi1150 and not w39381;
w39389 <= not w39387 and w39388;
w39390 <= not pi1147 and pi1151;
w39391 <= w37703 and w39390;
w39392 <= not w37202 and w38227;
w39393 <= w38259 and not w39392;
w39394 <= w37433 and not w39393;
w39395 <= w38128 and not w38228;
w39396 <= pi1147 and not w39395;
w39397 <= not w39394 and w39396;
w39398 <= not pi1150 and not w39391;
w39399 <= not w39397 and w39398;
w39400 <= not w39389 and not w39399;
w39401 <= not pi1149 and not w39400;
w39402 <= not pi1151 and not w37771;
w39403 <= not w38200 and w39402;
w39404 <= not w37722 and w37832;
w39405 <= not w37771 and not w39404;
w39406 <= pi1151 and w39405;
w39407 <= not pi1147 and not w39403;
w39408 <= not w39406 and w39407;
w39409 <= pi1147 and not w38183;
w39410 <= not pi1151 and not w37709;
w39411 <= not w37761 and w39410;
w39412 <= w39409 and not w39411;
w39413 <= not pi1150 and not w39408;
w39414 <= not w39412 and w39413;
w39415 <= w38111 and w38229;
w39416 <= pi1147 and not w39415;
w39417 <= not w37709 and not w37760;
w39418 <= not pi1151 and w39417;
w39419 <= w39416 and not w39418;
w39420 <= not w39330 and w39402;
w39421 <= pi1151 and not w37771;
w39422 <= not w37866 and w39421;
w39423 <= not pi1147 and not w39422;
w39424 <= not w39420 and w39423;
w39425 <= pi1150 and not w39419;
w39426 <= not w39424 and w39425;
w39427 <= not w39414 and not w39426;
w39428 <= pi1149 and not w39427;
w39429 <= not pi1148 and not w39401;
w39430 <= not w39428 and w39429;
w39431 <= not w39377 and not w39430;
w39432 <= not pi0213 and not w39431;
w39433 <= pi0209 and not w39307;
w39434 <= not w39432 and w39433;
w39435 <= not pi0213 and not w37768;
w39436 <= not w39330 and w39421;
w39437 <= pi1147 and not w38235;
w39438 <= not w39436 and w39437;
w39439 <= w4989 and not w38274;
w39440 <= not w38277 and w39439;
w39441 <= not w38048 and not w39440;
w39442 <= w39379 and w39441;
w39443 <= not pi1150 and not w39442;
w39444 <= not w39438 and w39443;
w39445 <= w38063 and w39332;
w39446 <= w38086 and not w39331;
w39447 <= pi1147 and not w39446;
w39448 <= not w39445 and w39447;
w39449 <= w37679 and w37686;
w39450 <= w38063 and not w39449;
w39451 <= w39317 and not w39450;
w39452 <= pi1150 and not w39448;
w39453 <= not w39451 and w39452;
w39454 <= not w39444 and not w39453;
w39455 <= not pi1149 and not w39454;
w39456 <= w38128 and not w39382;
w39457 <= not w37709 and not w39141;
w39458 <= pi1151 and w39457;
w39459 <= not pi1147 and not w39458;
w39460 <= not w39456 and w39459;
w39461 <= not w37650 and w39395;
w39462 <= w39416 and not w39461;
w39463 <= not pi1150 and not w39462;
w39464 <= not w39460 and w39463;
w39465 <= not w37694 and not w38240;
w39466 <= not pi1151 and w39465;
w39467 <= w39324 and not w39466;
w39468 <= w38140 and not w39309;
w39469 <= w37632 and not w37878;
w39470 <= w37873 and not w39469;
w39471 <= w38156 and not w39470;
w39472 <= not pi1147 and not w39471;
w39473 <= not w39468 and w39472;
w39474 <= pi1150 and not w39467;
w39475 <= not w39473 and w39474;
w39476 <= not w39464 and not w39475;
w39477 <= pi1149 and not w39476;
w39478 <= pi1148 and not w39477;
w39479 <= not w39455 and w39478;
w39480 <= not w14042 and w37427;
w39481 <= pi1151 and not w39480;
w39482 <= w39343 and not w39481;
w39483 <= w38063 and not w39360;
w39484 <= w37748 and w38216;
w39485 <= not w37659 and not w39484;
w39486 <= not pi1151 and w39485;
w39487 <= pi1147 and not w39483;
w39488 <= not w39486 and w39487;
w39489 <= pi1150 and not w39482;
w39490 <= not w39488 and w39489;
w39491 <= w37705 and w39390;
w39492 <= not w37771 and not w38200;
w39493 <= not pi1151 and not w39058;
w39494 <= pi1147 and not w39493;
w39495 <= not w39492 and w39494;
w39496 <= not pi1150 and not w39491;
w39497 <= not w39495 and w39496;
w39498 <= not w39490 and not w39497;
w39499 <= not pi1149 and not w39498;
w39500 <= w37205 and w37393;
w39501 <= not w8406 and w39500;
w39502 <= not w39393 and not w39501;
w39503 <= w38111 and w39502;
w39504 <= w38128 and not w39393;
w39505 <= not pi1147 and not w39504;
w39506 <= not w39503 and w39505;
w39507 <= not pi0219 and not w38094;
w39508 <= not w38205 and w39507;
w39509 <= w37727 and not w39508;
w39510 <= not w37723 and w39509;
w39511 <= w38128 and not w39510;
w39512 <= w39409 and not w39511;
w39513 <= not pi1150 and not w39506;
w39514 <= not w39512 and w39513;
w39515 <= w38156 and not w39500;
w39516 <= not w38267 and w39515;
w39517 <= w38140 and not w38267;
w39518 <= not pi1147 and not w39516;
w39519 <= not w39517 and w39518;
w39520 <= not w37694 and not w39509;
w39521 <= not pi1151 and w39520;
w39522 <= w39357 and not w39521;
w39523 <= pi1150 and not w39519;
w39524 <= not w39522 and w39523;
w39525 <= not w39514 and not w39524;
w39526 <= pi1149 and not w39525;
w39527 <= not pi1148 and not w39499;
w39528 <= not w39526 and w39527;
w39529 <= not w39479 and not w39528;
w39530 <= pi0213 and not w39529;
w39531 <= not pi0209 and not w39435;
w39532 <= not w39530 and w39531;
w39533 <= not w39434 and not w39532;
w39534 <= pi0230 and not w39533;
w39535 <= not pi0230 and not pi0247;
w39536 <= not w39534 and not w39535;
w39537 <= not pi1151 and not w37705;
w39538 <= not w37703 and w39537;
w39539 <= pi1152 and not w39538;
w39540 <= not w38173 and w39539;
w39541 <= pi1151 and not pi1152;
w39542 <= not w37688 and w39541;
w39543 <= not pi1150 and not w39540;
w39544 <= not w39542 and w39543;
w39545 <= pi1151 and w37697;
w39546 <= not pi1152 and not w39545;
w39547 <= not w38182 and w39546;
w39548 <= pi1152 and not w38178;
w39549 <= not w37728 and w39410;
w39550 <= w39548 and not w39549;
w39551 <= pi1150 and not w39547;
w39552 <= not w39550 and w39551;
w39553 <= not w39544 and not w39552;
w39554 <= pi0213 and w39553;
w39555 <= pi1152 and not w39517;
w39556 <= not w39310 and w39555;
w39557 <= pi1151 and w39313;
w39558 <= not pi1152 and not w39348;
w39559 <= not w39557 and w39558;
w39560 <= not pi1150 and not w39556;
w39561 <= not w39559 and w39560;
w39562 <= not w39355 and w39361;
w39563 <= w39548 and not w39562;
w39564 <= pi1151 and not w37690;
w39565 <= w39325 and w39564;
w39566 <= not pi1152 and not w39565;
w39567 <= not w39363 and w39566;
w39568 <= pi1150 and not w39567;
w39569 <= not w39563 and w39568;
w39570 <= pi1148 and not w39561;
w39571 <= not w39569 and w39570;
w39572 <= not w37687 and w39318;
w39573 <= not pi1152 and not w39572;
w39574 <= not w39342 and w39573;
w39575 <= w38086 and not w39344;
w39576 <= pi1152 and not w39575;
w39577 <= not w39320 and w39576;
w39578 <= not pi1150 and not w39577;
w39579 <= not w39574 and w39578;
w39580 <= not pi1151 and w39368;
w39581 <= pi1152 and not w39334;
w39582 <= not w39580 and w39581;
w39583 <= not pi1152 and not w39365;
w39584 <= not w39445 and w39583;
w39585 <= pi1150 and not w39582;
w39586 <= not w39584 and w39585;
w39587 <= not pi1148 and not w39586;
w39588 <= not w39579 and w39587;
w39589 <= not w39571 and not w39588;
w39590 <= pi1149 and not w39589;
w39591 <= not pi1152 and not w39403;
w39592 <= not w39436 and w39591;
w39593 <= not pi1151 and w39405;
w39594 <= pi1152 and not w39422;
w39595 <= not w39593 and w39594;
w39596 <= pi1150 and not w39592;
w39597 <= not w39595 and w39596;
w39598 <= w37806 and w39541;
w39599 <= not pi1151 and not w37703;
w39600 <= pi1152 and not w39380;
w39601 <= not w39599 and w39600;
w39602 <= not pi1150 and not w39598;
w39603 <= not w39601 and w39602;
w39604 <= not w39597 and not w39603;
w39605 <= not pi1148 and not w39604;
w39606 <= pi1152 and not w39549;
w39607 <= not w39415 and w39606;
w39608 <= pi1151 and w39417;
w39609 <= not pi1152 and not w39411;
w39610 <= not w39608 and w39609;
w39611 <= not w39607 and not w39610;
w39612 <= pi1150 and not w39611;
w39613 <= pi1151 and w39384;
w39614 <= not w39395 and not w39613;
w39615 <= not pi1152 and not w39614;
w39616 <= not w39383 and not w39504;
w39617 <= pi1152 and not w39616;
w39618 <= not pi1150 and not w39615;
w39619 <= not w39617 and w39618;
w39620 <= pi1148 and not w39619;
w39621 <= not w39612 and w39620;
w39622 <= not pi1149 and not w39605;
w39623 <= not w39621 and w39622;
w39624 <= not w39590 and not w39623;
w39625 <= not pi0213 and not w39624;
w39626 <= pi0209 and not w39554;
w39627 <= not w39625 and w39626;
w39628 <= not pi0213 and not w39051;
w39629 <= w39341 and w39541;
w39630 <= pi1152 and not w39481;
w39631 <= not w39537 and w39630;
w39632 <= not pi1150 and not w39629;
w39633 <= not w39631 and w39632;
w39634 <= not pi1152 and not w39504;
w39635 <= not w39347 and w39634;
w39636 <= w39410 and w39502;
w39637 <= pi1152 and not w39516;
w39638 <= not w39636 and w39637;
w39639 <= pi1150 and not w39635;
w39640 <= not w39638 and w39639;
w39641 <= not pi1149 and not w39633;
w39642 <= not w39640 and w39641;
w39643 <= not pi1151 and w39457;
w39644 <= pi1152 and not w39471;
w39645 <= not w39643 and w39644;
w39646 <= not pi1152 and not w39310;
w39647 <= not w39456 and w39646;
w39648 <= pi1150 and not w39645;
w39649 <= not w39647 and w39648;
w39650 <= not w39378 and w39573;
w39651 <= not pi1151 and not w39441;
w39652 <= pi1152 and not w39651;
w39653 <= not w39450 and w39652;
w39654 <= not pi1150 and not w39653;
w39655 <= not w39650 and w39654;
w39656 <= pi1149 and not w39649;
w39657 <= not w39655 and w39656;
w39658 <= not pi1148 and not w39642;
w39659 <= not w39657 and w39658;
w39660 <= w39318 and not w39331;
w39661 <= w38236 and not w39660;
w39662 <= pi1152 and not w39420;
w39663 <= not w39445 and w39662;
w39664 <= not pi1150 and not w39661;
w39665 <= not w39663 and w39664;
w39666 <= pi1151 and w39465;
w39667 <= not pi1152 and not w39461;
w39668 <= not w39666 and w39667;
w39669 <= w38229 and w39410;
w39670 <= w39548 and not w39669;
w39671 <= pi1150 and not w39668;
w39672 <= not w39670 and w39671;
w39673 <= pi1149 and not w39672;
w39674 <= not w39665 and w39673;
w39675 <= pi1151 and w39485;
w39676 <= not pi1152 and not w39493;
w39677 <= not w39675 and w39676;
w39678 <= pi1152 and not w39403;
w39679 <= not w39483 and w39678;
w39680 <= not pi1150 and not w39679;
w39681 <= not w39677 and w39680;
w39682 <= not w39356 and w39606;
w39683 <= pi1151 and w39520;
w39684 <= not pi1152 and not w39511;
w39685 <= not w39683 and w39684;
w39686 <= pi1150 and not w39682;
w39687 <= not w39685 and w39686;
w39688 <= not pi1149 and not w39681;
w39689 <= not w39687 and w39688;
w39690 <= pi1148 and not w39674;
w39691 <= not w39689 and w39690;
w39692 <= pi0213 and not w39659;
w39693 <= not w39691 and w39692;
w39694 <= not pi0209 and not w39628;
w39695 <= not w39693 and w39694;
w39696 <= not w39627 and not w39695;
w39697 <= pi0230 and not w39696;
w39698 <= not pi0230 and not pi0248;
w39699 <= not w39697 and not w39698;
w39700 <= not pi0213 and w39553;
w39701 <= pi0057 and not w36449;
w39702 <= not w3868 and w36449;
w39703 <= not w37301 and w37445;
w39704 <= pi0299 and w36446;
w39705 <= not w38245 and not w39704;
w39706 <= not pi0214 and not w39705;
w39707 <= pi0212 and not w39703;
w39708 <= not w39706 and w39707;
w39709 <= pi0214 and not w39705;
w39710 <= not pi0212 and not w37311;
w39711 <= not w39709 and w39710;
w39712 <= not pi0219 and not w39708;
w39713 <= not w39711 and w39712;
w39714 <= w3868 and not w37331;
w39715 <= not w39713 and w39714;
w39716 <= not pi0057 and pi1151;
w39717 <= not w39702 and w39716;
w39718 <= not w39715 and w39717;
w39719 <= not w37746 and not w39704;
w39720 <= not w37311 and w39719;
w39721 <= not pi0212 and not w39720;
w39722 <= not pi0214 and w39719;
w39723 <= not w37417 and not w37745;
w39724 <= pi0214 and not w38198;
w39725 <= not w39723 and w39724;
w39726 <= pi0212 and not w39725;
w39727 <= not w39722 and w39726;
w39728 <= not w39721 and not w39727;
w39729 <= not pi0219 and not w39728;
w39730 <= w3868 and not w38215;
w39731 <= not w39729 and w39730;
w39732 <= not pi0057 and not pi1151;
w39733 <= not w39702 and w39732;
w39734 <= not w39731 and w39733;
w39735 <= not w39701 and not w39718;
w39736 <= not w39734 and w39735;
w39737 <= not pi1152 and not w39736;
w39738 <= pi0299 and not w36446;
w39739 <= not w8406 and w39738;
w39740 <= not w36480 and not w39739;
w39741 <= w37646 and not w39740;
w39742 <= w38223 and not w39741;
w39743 <= not w37758 and not w37854;
w39744 <= pi1151 and not w39743;
w39745 <= not w39742 and w39744;
w39746 <= w38088 and not w39704;
w39747 <= not w37249 and not w39704;
w39748 <= not pi0214 and not w39747;
w39749 <= w37712 and not w38191;
w39750 <= pi0212 and not w39748;
w39751 <= not w39749 and w39750;
w39752 <= w39079 and not w39746;
w39753 <= not w39751 and w39752;
w39754 <= not pi1151 and not w39753;
w39755 <= w37727 and w39754;
w39756 <= w36485 and not w39745;
w39757 <= not w39755 and w39756;
w39758 <= pi1150 and not w39757;
w39759 <= not w39737 and w39758;
w39760 <= not pi0212 and w37299;
w39761 <= w37625 and not w39738;
w39762 <= pi0212 and not w39761;
w39763 <= not w38302 and w39762;
w39764 <= not pi0219 and not w39760;
w39765 <= not w39746 and w39764;
w39766 <= not w39763 and w39765;
w39767 <= w37257 and not w37872;
w39768 <= not w39766 and w39767;
w39769 <= not pi1151 and w39393;
w39770 <= not w37301 and not w39739;
w39771 <= w36448 and w37198;
w39772 <= not w39770 and w39771;
w39773 <= w36485 and not w39772;
w39774 <= not w39769 and w39773;
w39775 <= not w39768 and w39774;
w39776 <= w8406 and w38276;
w39777 <= w36629 and not w37663;
w39778 <= not w36308 and w37673;
w39779 <= pi0211 and w38275;
w39780 <= w36171 and not w39778;
w39781 <= not w39779 and w39780;
w39782 <= not w39776 and not w39777;
w39783 <= not w39781 and w39782;
w39784 <= not pi0219 and not w39783;
w39785 <= pi1151 and w37686;
w39786 <= not w39784 and w39785;
w39787 <= w36451 and not w39772;
w39788 <= not w39786 and w39787;
w39789 <= not pi1150 and not w39775;
w39790 <= not w39788 and w39789;
w39791 <= not w39759 and not w39790;
w39792 <= pi0213 and not w39791;
w39793 <= not pi0209 and not w39792;
w39794 <= not w39700 and w39793;
w39795 <= pi0213 and w36634;
w39796 <= not w8047 and not w36592;
w39797 <= w36238 and not w36816;
w39798 <= pi0207 and not w36332;
w39799 <= not w36590 and w39798;
w39800 <= not pi0207 and w36815;
w39801 <= pi0208 and not w39799;
w39802 <= not w39800 and w39801;
w39803 <= not w39797 and not w39802;
w39804 <= pi0211 and not w39803;
w39805 <= pi0214 and w39804;
w39806 <= not w39796 and not w39805;
w39807 <= not pi0212 and not w39806;
w39808 <= not pi0219 and not w39807;
w39809 <= not pi0211 and w39803;
w39810 <= not w36662 and not w39809;
w39811 <= pi0214 and not w39810;
w39812 <= not pi0211 and not w36592;
w39813 <= not pi0214 and not w39812;
w39814 <= not w39804 and w39813;
w39815 <= pi0212 and not w39814;
w39816 <= not w39811 and w39815;
w39817 <= w39808 and not w39816;
w39818 <= w36594 and not w39817;
w39819 <= w39318 and not w39818;
w39820 <= not w36592 and w36636;
w39821 <= not w39541 and not w39820;
w39822 <= not w39819 and not w39821;
w39823 <= not w36529 and not w37472;
w39824 <= not w36531 and w37472;
w39825 <= w4989 and not w39823;
w39826 <= not w39824 and w39825;
w39827 <= w39402 and not w39826;
w39828 <= pi0214 and w36516;
w39829 <= w36577 and not w39828;
w39830 <= not pi0219 and not w39829;
w39831 <= pi0214 and not w36531;
w39832 <= not pi0214 and w36516;
w39833 <= pi0212 and not w39832;
w39834 <= not w39831 and w39833;
w39835 <= w39830 and not w39834;
w39836 <= w4989 and not w36534;
w39837 <= not w39835 and w39836;
w39838 <= w38063 and not w39837;
w39839 <= pi1152 and not w39827;
w39840 <= not w39838 and w39839;
w39841 <= not w39822 and not w39840;
w39842 <= not pi1150 and not w39841;
w39843 <= not w35976 and w39810;
w39844 <= pi0219 and not w36637;
w39845 <= not w39843 and w39844;
w39846 <= w4989 and not w39845;
w39847 <= pi0212 and not w39806;
w39848 <= not pi0212 and not w36592;
w39849 <= not pi0219 and not w39848;
w39850 <= not w39847 and w39849;
w39851 <= w39846 and not w39850;
w39852 <= w38128 and not w39851;
w39853 <= pi0214 and w39803;
w39854 <= w39815 and not w39853;
w39855 <= w39808 and not w39854;
w39856 <= w39846 and not w39855;
w39857 <= w39308 and not w39856;
w39858 <= not pi1152 and not w39852;
w39859 <= not w39857 and w39858;
w39860 <= pi0212 and not w36516;
w39861 <= w39830 and not w39860;
w39862 <= w36537 and not w39861;
w39863 <= w38156 and not w39862;
w39864 <= not w36576 and not w39831;
w39865 <= not pi0212 and not w39864;
w39866 <= not pi0211 and w36529;
w39867 <= not w36555 and not w39866;
w39868 <= pi0214 and not w39867;
w39869 <= not pi0214 and w36531;
w39870 <= pi0212 and not w39868;
w39871 <= not w39869 and w39870;
w39872 <= not w39865 and not w39871;
w39873 <= not pi0219 and not w39872;
w39874 <= w36537 and not w39873;
w39875 <= w39410 and not w39874;
w39876 <= pi1152 and not w39863;
w39877 <= not w39875 and w39876;
w39878 <= not w39859 and not w39877;
w39879 <= pi1150 and not w39878;
w39880 <= not w39842 and not w39879;
w39881 <= not pi0213 and not w39880;
w39882 <= pi0209 and not w39795;
w39883 <= not w39881 and w39882;
w39884 <= not w39794 and not w39883;
w39885 <= pi0230 and not w39884;
w39886 <= not pi0230 and not pi0249;
w39887 <= not w39885 and not w39886;
w39888 <= w94 and w9076;
w39889 <= not w3849 and not w39888;
w39890 <= not pi0075 and not w39889;
w39891 <= w4896 and w6529;
w39892 <= not w39890 and not w39891;
w39893 <= not pi0087 and not pi0250;
w39894 <= w6444 and w39893;
w39895 <= not w39892 and w39894;
w39896 <= pi0897 and w8372;
w39897 <= not pi0476 and w9007;
w39898 <= not w39896 and not w39897;
w39899 <= not pi0200 and pi1053;
w39900 <= pi0200 and pi1039;
w39901 <= not pi0199 and not w39899;
w39902 <= not w39900 and w39901;
w39903 <= not w39898 and not w39902;
w39904 <= pi0251 and w39898;
w39905 <= not w39903 and not w39904;
w39906 <= not w8546 and w9115;
w39907 <= not w3761 and w9115;
w39908 <= not pi0979 and not pi0984;
w39909 <= pi1001 and w39908;
w39910 <= w3749 and w39909;
w39911 <= not w3776 and w39910;
w39912 <= w3943 and w39911;
w39913 <= not pi0252 and not w39912;
w39914 <= pi1092 and not pi1093;
w39915 <= not w39913 and w39914;
w39916 <= w3955 and not w39915;
w39917 <= w3954 and w39915;
w39918 <= not w39916 and not w39917;
w39919 <= w3761 and w39918;
w39920 <= not w39907 and not w39919;
w39921 <= w3805 and not w39920;
w39922 <= not w3790 and w39918;
w39923 <= w3790 and w9115;
w39924 <= not w39922 and not w39923;
w39925 <= not w3805 and not w39924;
w39926 <= pi0299 and not w39921;
w39927 <= not w39925 and w39926;
w39928 <= w3768 and not w39920;
w39929 <= not w3768 and not w39924;
w39930 <= not pi0299 and not w39928;
w39931 <= not w39929 and w39930;
w39932 <= w8546 and not w39927;
w39933 <= not w39931 and w39932;
w39934 <= not w5206 and not w39906;
w39935 <= not w39933 and w39934;
w39936 <= pi0057 and w9114;
w39937 <= w8545 and w39910;
w39938 <= w18693 and w39937;
w39939 <= w3780 and w39938;
w39940 <= not w35950 and w39939;
w39941 <= w3943 and w39940;
w39942 <= not pi0252 and not w39941;
w39943 <= not pi0057 and pi1092;
w39944 <= not w39942 and w39943;
w39945 <= w5206 and not w39936;
w39946 <= not w39944 and w39945;
w39947 <= not w39935 and not w39946;
w39948 <= not w10624 and not w36071;
w39949 <= not w36263 and w39948;
w39950 <= w4989 and w39949;
w39951 <= pi0219 and w37643;
w39952 <= not w39950 and not w39951;
w39953 <= pi1153 and not w39952;
w39954 <= not pi1151 and not w39953;
w39955 <= w8407 and w36247;
w39956 <= pi0211 and not w36133;
w39957 <= not w39955 and not w39956;
w39958 <= not w36108 and not w36125;
w39959 <= w36082 and not w39958;
w39960 <= w4989 and not w39959;
w39961 <= w39957 and w39960;
w39962 <= not w9009 and w36844;
w39963 <= pi1151 and not w39962;
w39964 <= not w39961 and w39963;
w39965 <= not w39954 and not w39964;
w39966 <= not pi1152 and not w39965;
w39967 <= w36082 and w37346;
w39968 <= not pi1151 and not w9010;
w39969 <= not w36251 and w39968;
w39970 <= not w39967 and w39969;
w39971 <= not w8947 and not w36071;
w39972 <= not w36131 and not w37417;
w39973 <= pi1153 and not w39972;
w39974 <= pi1151 and w39971;
w39975 <= not w39973 and w39974;
w39976 <= w4989 and not w39975;
w39977 <= not w39970 and w39976;
w39978 <= not pi1151 and w8407;
w39979 <= not w36843 and not w39978;
w39980 <= not w4989 and w39979;
w39981 <= pi1152 and not w39980;
w39982 <= not w39977 and w39981;
w39983 <= not w39966 and not w39982;
w39984 <= pi0230 and not w39983;
w39985 <= not pi0253 and not pi1091;
w39986 <= not w4989 and not w39985;
w39987 <= pi0211 and pi1091;
w39988 <= pi1091 and not pi1153;
w39989 <= pi0219 and w39988;
w39990 <= not w39987 and not w39989;
w39991 <= w39986 and w39990;
w39992 <= pi1091 and not w39957;
w39993 <= not pi1153 and not w38478;
w39994 <= pi1153 and not w38515;
w39995 <= w36082 and not w39994;
w39996 <= not w39993 and w39995;
w39997 <= not w39992 and not w39996;
w39998 <= pi0253 and not w39997;
w39999 <= not w10627 and not w39973;
w40000 <= pi1091 and not w39999;
w40001 <= not pi0253 and not w40000;
w40002 <= w4989 and not w40001;
w40003 <= not w39998 and w40002;
w40004 <= pi1151 and not w39991;
w40005 <= not w40003 and w40004;
w40006 <= pi0253 and not pi1091;
w40007 <= pi0219 and pi1091;
w40008 <= not w36060 and w40007;
w40009 <= w39986 and not w40008;
w40010 <= pi0219 and w40009;
w40011 <= pi1091 and pi1153;
w40012 <= w39950 and w40011;
w40013 <= not pi1151 and not w40006;
w40014 <= not w40012 and w40013;
w40015 <= not w40010 and w40014;
w40016 <= not w40005 and not w40015;
w40017 <= not pi1152 and not w40016;
w40018 <= not pi0211 and pi1091;
w40019 <= not pi0219 and w40018;
w40020 <= w40009 and not w40019;
w40021 <= w9009 and w38474;
w40022 <= not w36251 and w40021;
w40023 <= not pi1153 and not w38506;
w40024 <= not w36124 and w38474;
w40025 <= pi1153 and not w40024;
w40026 <= w36082 and not w40025;
w40027 <= not w40023 and w40026;
w40028 <= pi0253 and not w40022;
w40029 <= not w40027 and w40028;
w40030 <= pi1091 and w37346;
w40031 <= pi1091 and w36108;
w40032 <= w36521 and w40031;
w40033 <= w36082 and not w40032;
w40034 <= not w40030 and w40033;
w40035 <= pi1091 and w36251;
w40036 <= pi0211 and not w38528;
w40037 <= not w40035 and w40036;
w40038 <= not pi0253 and not w40034;
w40039 <= not w40037 and w40038;
w40040 <= not w40029 and not w40039;
w40041 <= not w9009 and not w36082;
w40042 <= not w40006 and w40041;
w40043 <= not w40035 and w40042;
w40044 <= w37198 and not w40043;
w40045 <= not w40040 and w40044;
w40046 <= w39972 and not w40006;
w40047 <= not w39988 and not w40046;
w40048 <= w39971 and not w40047;
w40049 <= w4989 and not w39985;
w40050 <= not w40048 and w40049;
w40051 <= not w40009 and not w40050;
w40052 <= pi1151 and not w40051;
w40053 <= pi1152 and not w40020;
w40054 <= not w40052 and w40053;
w40055 <= not w40045 and w40054;
w40056 <= not w38473 and not w40055;
w40057 <= not w40017 and w40056;
w40058 <= w38551 and w38635;
w40059 <= pi1153 and not w40058;
w40060 <= not pi1153 and not w38681;
w40061 <= not pi0219 and not w40060;
w40062 <= not w40059 and w40061;
w40063 <= not pi1153 and not w38611;
w40064 <= not w38550 and not w38574;
w40065 <= not pi0211 and w38607;
w40066 <= w40064 and not w40065;
w40067 <= w38563 and not w38571;
w40068 <= w40066 and w40067;
w40069 <= pi1153 and not w40068;
w40070 <= pi0219 and not w40063;
w40071 <= not w40069 and w40070;
w40072 <= pi0253 and not w40062;
w40073 <= not w40071 and w40072;
w40074 <= not w38556 and w38611;
w40075 <= not pi0211 and w40074;
w40076 <= not w38576 and not w40075;
w40077 <= pi1153 and not w40076;
w40078 <= not w38602 and not w40077;
w40079 <= pi0219 and w40078;
w40080 <= not pi1153 and w38679;
w40081 <= pi1153 and w38660;
w40082 <= not pi0219 and not w40080;
w40083 <= not w40081 and w40082;
w40084 <= not pi0253 and not w40083;
w40085 <= not w40079 and w40084;
w40086 <= not w40073 and not w40085;
w40087 <= w4989 and not w40086;
w40088 <= not pi0219 and not w38543;
w40089 <= not pi0211 and not w38453;
w40090 <= w40088 and not w40089;
w40091 <= not pi0219 and not w40090;
w40092 <= not w4989 and w40091;
w40093 <= not w38437 and w40092;
w40094 <= not w38431 and not w40008;
w40095 <= not w40088 and w40094;
w40096 <= pi0253 and not w40095;
w40097 <= not pi0219 and not w38453;
w40098 <= pi0211 and w38431;
w40099 <= not pi0211 and not w38437;
w40100 <= pi0219 and not w40098;
w40101 <= not w40099 and w40100;
w40102 <= not w40008 and not w40097;
w40103 <= not w40101 and w40102;
w40104 <= not pi0253 and not w40103;
w40105 <= not w4989 and not w40096;
w40106 <= not w40104 and w40105;
w40107 <= pi1151 and not w40093;
w40108 <= not w40106 and w40107;
w40109 <= not w40087 and w40108;
w40110 <= not w38635 and not w40075;
w40111 <= w40088 and not w40110;
w40112 <= not w38550 and not w38562;
w40113 <= not pi1153 and not w40112;
w40114 <= not w38665 and not w40113;
w40115 <= w40111 and not w40114;
w40116 <= pi0219 and w38572;
w40117 <= not w38620 and w40069;
w40118 <= w40116 and not w40117;
w40119 <= not w40115 and not w40118;
w40120 <= pi0253 and not w40119;
w40121 <= not w38575 and w40066;
w40122 <= not w40113 and w40121;
w40123 <= not pi0219 and not w40122;
w40124 <= pi0219 and w38574;
w40125 <= not w40123 and not w40124;
w40126 <= not w40079 and w40125;
w40127 <= not pi0253 and not w40126;
w40128 <= w4989 and not w40120;
w40129 <= not w40127 and w40128;
w40130 <= not pi1151 and not w40129;
w40131 <= not w40109 and not w40130;
w40132 <= w40097 and not w40099;
w40133 <= w40088 and not w40132;
w40134 <= pi0219 and not w38437;
w40135 <= not w4989 and not w40134;
w40136 <= not w40133 and w40135;
w40137 <= not w38437 and w40136;
w40138 <= not w40106 and not w40137;
w40139 <= not w40131 and w40138;
w40140 <= pi1152 and not w40139;
w40141 <= pi0219 and not w40078;
w40142 <= not w40083 and w40111;
w40143 <= not w40141 and not w40142;
w40144 <= not w38556 and not w40143;
w40145 <= not pi0253 and not w40144;
w40146 <= pi1153 and not w38551;
w40147 <= w40066 and w40088;
w40148 <= not w40146 and w40147;
w40149 <= not pi1153 and not w38591;
w40150 <= not w38625 and not w40068;
w40151 <= pi1153 and w40150;
w40152 <= pi0219 and not w40149;
w40153 <= not w40151 and w40152;
w40154 <= not w40148 and not w40153;
w40155 <= pi0253 and not w40154;
w40156 <= w4989 and not w40155;
w40157 <= not w40145 and w40156;
w40158 <= w40108 and not w40157;
w40159 <= not pi1091 and not w38602;
w40160 <= not pi1153 and not w40159;
w40161 <= not w38620 and not w40068;
w40162 <= not pi0219 and w40112;
w40163 <= not w40160 and not w40162;
w40164 <= w40161 and w40163;
w40165 <= pi0253 and not w40164;
w40166 <= not w38565 and w40141;
w40167 <= not pi1153 and not w38647;
w40168 <= not w38556 and not w40167;
w40169 <= not pi0219 and w38681;
w40170 <= w40168 and w40169;
w40171 <= not pi0253 and not w40170;
w40172 <= not w40166 and w40171;
w40173 <= w4989 and not w40165;
w40174 <= not w40172 and w40173;
w40175 <= not pi1151 and not w40106;
w40176 <= not w40174 and w40175;
w40177 <= not pi1152 and not w40176;
w40178 <= not w40158 and w40177;
w40179 <= not w40140 and not w40178;
w40180 <= w38473 and not w40179;
w40181 <= not pi0230 and not w40057;
w40182 <= not w40180 and w40181;
w40183 <= not w39984 and not w40182;
w40184 <= not pi0219 and not w36445;
w40185 <= not w36708 and not w40184;
w40186 <= not w4989 and w40185;
w40187 <= pi1154 and w36540;
w40188 <= not w36596 and not w40187;
w40189 <= w9009 and not w40188;
w40190 <= pi0299 and w36082;
w40191 <= not w9009 and w36522;
w40192 <= not w40190 and not w40191;
w40193 <= not w36502 and not w40192;
w40194 <= not w40189 and not w40193;
w40195 <= w4989 and not w40194;
w40196 <= not pi1152 and not w40186;
w40197 <= not w40195 and w40196;
w40198 <= w9009 and not w36445;
w40199 <= w37591 and not w40198;
w40200 <= not pi0200 and pi1154;
w40201 <= w8936 and not w40200;
w40202 <= w36539 and not w37417;
w40203 <= not w40201 and not w40202;
w40204 <= not pi0219 and not w40203;
w40205 <= not w36121 and not w36539;
w40206 <= w36051 and not w40205;
w40207 <= not pi1154 and not w36585;
w40208 <= not w36504 and not w40207;
w40209 <= not w40206 and w40208;
w40210 <= pi0219 and not w40209;
w40211 <= w4989 and not w40204;
w40212 <= not w40210 and w40211;
w40213 <= pi1152 and not w40199;
w40214 <= not w40212 and w40213;
w40215 <= not w40197 and not w40214;
w40216 <= pi0230 and not w40215;
w40217 <= not pi0254 and not pi1091;
w40218 <= pi1091 and not w40185;
w40219 <= not w4989 and not w40217;
w40220 <= not w40218 and w40219;
w40221 <= not w4989 and w40019;
w40222 <= not w40220 and not w40221;
w40223 <= pi1153 and not w38495;
w40224 <= not pi1154 and not w40223;
w40225 <= not pi0211 and w36246;
w40226 <= not w39993 and w40224;
w40227 <= not w40225 and w40226;
w40228 <= pi1091 and w36051;
w40229 <= not w36131 and w40228;
w40230 <= not w36608 and w40229;
w40231 <= not w40227 and not w40230;
w40232 <= not pi0219 and not w40231;
w40233 <= pi1154 and w40018;
w40234 <= not w40007 and not w40233;
w40235 <= not w40209 and not w40234;
w40236 <= not w40232 and not w40235;
w40237 <= pi0254 and not w40236;
w40238 <= pi1154 and not w39972;
w40239 <= pi0219 and not w36585;
w40240 <= not w40238 and w40239;
w40241 <= not w40204 and not w40240;
w40242 <= not pi0254 and not w40241;
w40243 <= not w40217 and not w40242;
w40244 <= not w40237 and w40243;
w40245 <= w4989 and w40244;
w40246 <= pi1152 and w40222;
w40247 <= not w40245 and w40246;
w40248 <= w38481 and w39988;
w40249 <= not w40030 and not w40248;
w40250 <= pi0211 and not w40224;
w40251 <= not w40249 and w40250;
w40252 <= w9008 and w40011;
w40253 <= not pi1154 and not w40252;
w40254 <= pi1091 and w36522;
w40255 <= pi1154 and not w40254;
w40256 <= not pi0211 and not w40253;
w40257 <= not w40255 and w40256;
w40258 <= not w40251 and not w40257;
w40259 <= not pi0219 and not w40258;
w40260 <= pi0211 and w40255;
w40261 <= pi1091 and w37229;
w40262 <= w36058 and not w40261;
w40263 <= not w40030 and w40262;
w40264 <= pi0219 and not w40253;
w40265 <= not w40263 and w40264;
w40266 <= not w40260 and w40265;
w40267 <= not w40259 and not w40266;
w40268 <= not pi0254 and not w40267;
w40269 <= not pi1153 and not w38482;
w40270 <= not w40025 and not w40269;
w40271 <= pi1091 and not pi1154;
w40272 <= w36096 and w40271;
w40273 <= not w40270 and not w40272;
w40274 <= w9009 and not w40273;
w40275 <= pi1091 and not w9009;
w40276 <= not w36501 and w40275;
w40277 <= not pi1154 and not w40276;
w40278 <= w38531 and w40026;
w40279 <= pi1091 and not w36204;
w40280 <= not w40270 and not w40279;
w40281 <= w40041 and not w40280;
w40282 <= pi1154 and not w40278;
w40283 <= not w40281 and w40282;
w40284 <= not w40277 and not w40283;
w40285 <= pi0254 and not w40274;
w40286 <= not w40284 and w40285;
w40287 <= not w40268 and not w40286;
w40288 <= w4989 and not w40287;
w40289 <= not pi1152 and not w40220;
w40290 <= not w40288 and w40289;
w40291 <= not w38473 and not w40247;
w40292 <= not w40290 and w40291;
w40293 <= pi1091 and w36708;
w40294 <= not pi0211 and not w38429;
w40295 <= w40134 and not w40294;
w40296 <= not pi0219 and w38453;
w40297 <= not w40295 and not w40296;
w40298 <= w9009 and w39988;
w40299 <= pi0254 and not w40298;
w40300 <= not w40293 and w40299;
w40301 <= w40297 and w40300;
w40302 <= not w40011 and w40132;
w40303 <= not pi0254 and not w40293;
w40304 <= not w40101 and w40303;
w40305 <= not w40302 and w40304;
w40306 <= pi0253 and not w40301;
w40307 <= not w40305 and w40306;
w40308 <= pi0253 and not w4989;
w40309 <= w40222 and not w40308;
w40310 <= not w40307 and not w40309;
w40311 <= not pi0253 and not w40244;
w40312 <= pi1154 and not w38548;
w40313 <= w40066 and w40312;
w40314 <= not w40059 and w40313;
w40315 <= not pi1153 and w40122;
w40316 <= not w38681 and not w40315;
w40317 <= not pi1154 and not w40316;
w40318 <= pi0254 and not w40314;
w40319 <= not w40317 and w40318;
w40320 <= pi0211 and w38607;
w40321 <= not w38556 and not w40320;
w40322 <= not pi1153 and not w40321;
w40323 <= not w38575 and w38591;
w40324 <= pi1154 and w40323;
w40325 <= not w38679 and not w40324;
w40326 <= not pi0254 and not w40322;
w40327 <= not w40325 and w40326;
w40328 <= not w40319 and not w40327;
w40329 <= not pi0219 and not w40328;
w40330 <= pi1154 and not w40069;
w40331 <= not w40150 and w40330;
w40332 <= pi1153 and not w38611;
w40333 <= not pi1154 and not w40149;
w40334 <= not w40332 and w40333;
w40335 <= pi0254 and not w40334;
w40336 <= not w40331 and w40335;
w40337 <= not w40063 and w40323;
w40338 <= w36058 and not w40337;
w40339 <= not w38553 and w40338;
w40340 <= not pi1153 and not w38595;
w40341 <= w38604 and not w40340;
w40342 <= not pi1154 and not w40341;
w40343 <= not w38556 and w38602;
w40344 <= w40342 and not w40343;
w40345 <= pi1153 and w38576;
w40346 <= w36051 and not w38558;
w40347 <= not w40345 and w40346;
w40348 <= not pi0254 and not w40347;
w40349 <= not w40339 and w40348;
w40350 <= not w40344 and w40349;
w40351 <= not w40336 and not w40350;
w40352 <= pi0219 and not w40351;
w40353 <= pi0253 and not w40352;
w40354 <= not w40329 and w40353;
w40355 <= w4989 and not w40311;
w40356 <= not w40354 and w40355;
w40357 <= pi1152 and not w40310;
w40358 <= not w40356 and w40357;
w40359 <= not w40220 and not w40308;
w40360 <= not w40133 and w40301;
w40361 <= not w40091 and w40305;
w40362 <= pi0253 and not w40360;
w40363 <= not w40361 and w40362;
w40364 <= not w40359 and not w40363;
w40365 <= not pi0253 and w40287;
w40366 <= w36058 and not w38620;
w40367 <= not pi1153 and w38563;
w40368 <= not pi1154 and not w38566;
w40369 <= not pi1154 and not w40368;
w40370 <= not w40067 and not w40367;
w40371 <= not w40369 and w40370;
w40372 <= pi0219 and not w40366;
w40373 <= not w40371 and w40372;
w40374 <= pi1154 and w38562;
w40375 <= w40110 and not w40367;
w40376 <= not pi0219 and not w40374;
w40377 <= not w40375 and w40376;
w40378 <= not w40373 and not w40377;
w40379 <= pi0254 and not w40378;
w40380 <= w38577 and not w40063;
w40381 <= w36051 and not w40380;
w40382 <= pi0219 and not w40338;
w40383 <= not w40342 and w40382;
w40384 <= not w40381 and w40383;
w40385 <= pi1154 and w38574;
w40386 <= not w38607 and not w40385;
w40387 <= not pi0211 and not w40386;
w40388 <= not w38548 and w38679;
w40389 <= not w40167 and w40388;
w40390 <= not pi1154 and not w40389;
w40391 <= not w38556 and w38681;
w40392 <= pi1154 and not w40391;
w40393 <= not w40389 and w40392;
w40394 <= not pi0219 and not w40387;
w40395 <= not w40390 and w40394;
w40396 <= not w40393 and w40395;
w40397 <= not pi0254 and not w40396;
w40398 <= not w40384 and w40397;
w40399 <= not w40379 and not w40398;
w40400 <= pi0253 and not w40399;
w40401 <= w4989 and not w40365;
w40402 <= not w40400 and w40401;
w40403 <= not pi1152 and not w40364;
w40404 <= not w40402 and w40403;
w40405 <= w38473 and not w40404;
w40406 <= not w40358 and w40405;
w40407 <= not pi0230 and not w40292;
w40408 <= not w40406 and w40407;
w40409 <= not w40216 and not w40408;
w40410 <= not pi0200 and pi1049;
w40411 <= pi0200 and pi1036;
w40412 <= not w40410 and not w40411;
w40413 <= not w39898 and w40412;
w40414 <= not pi0255 and w39898;
w40415 <= not w40413 and not w40414;
w40416 <= not pi0200 and pi1048;
w40417 <= pi0200 and pi1070;
w40418 <= not w40416 and not w40417;
w40419 <= not w39898 and w40418;
w40420 <= not pi0256 and w39898;
w40421 <= not w40419 and not w40420;
w40422 <= not pi0200 and pi1084;
w40423 <= pi0200 and pi1065;
w40424 <= not w40422 and not w40423;
w40425 <= not w39898 and w40424;
w40426 <= not pi0257 and w39898;
w40427 <= not w40425 and not w40426;
w40428 <= not pi0200 and pi1072;
w40429 <= pi0200 and pi1062;
w40430 <= not w40428 and not w40429;
w40431 <= not w39898 and w40430;
w40432 <= not pi0258 and w39898;
w40433 <= not w40431 and not w40432;
w40434 <= not pi0200 and pi1059;
w40435 <= pi0200 and pi1069;
w40436 <= not w40434 and not w40435;
w40437 <= not w39898 and w40436;
w40438 <= not pi0259 and w39898;
w40439 <= not w40437 and not w40438;
w40440 <= not pi0200 and pi1044;
w40441 <= pi0200 and pi1067;
w40442 <= not pi0199 and not w40440;
w40443 <= not w40441 and w40442;
w40444 <= not w39898 and not w40443;
w40445 <= pi0260 and w39898;
w40446 <= not w40444 and not w40445;
w40447 <= not pi0200 and pi1037;
w40448 <= pi0200 and pi1040;
w40449 <= not pi0199 and not w40447;
w40450 <= not w40448 and w40449;
w40451 <= not w39898 and not w40450;
w40452 <= pi0261 and w39898;
w40453 <= not w40451 and not w40452;
w40454 <= pi1093 and pi1142;
w40455 <= not pi0262 and not pi1093;
w40456 <= not w40454 and not w40455;
w40457 <= not pi0228 and not w40456;
w40458 <= not pi0123 and not pi1142;
w40459 <= pi0123 and pi0262;
w40460 <= pi0228 and not w40458;
w40461 <= not w40459 and w40460;
w40462 <= not w40457 and not w40461;
w40463 <= not pi0228 and not pi1093;
w40464 <= pi0123 and pi0228;
w40465 <= not w40463 and not w40464;
w40466 <= not pi0262 and not w40465;
w40467 <= not w38263 and not w40466;
w40468 <= pi0199 and w40465;
w40469 <= w36004 and not w40468;
w40470 <= w40467 and not w40469;
w40471 <= not w40462 and not w40470;
w40472 <= not pi0207 and w40466;
w40473 <= not pi0208 and not w40472;
w40474 <= not w38263 and not w40473;
w40475 <= not w40471 and not w40474;
w40476 <= not w37274 and w40465;
w40477 <= not pi0299 and not w40476;
w40478 <= not w40462 and w40477;
w40479 <= pi0299 and not w40467;
w40480 <= pi0208 and not w40478;
w40481 <= not w40479 and w40480;
w40482 <= w4989 and not w40481;
w40483 <= not w40475 and w40482;
w40484 <= not w37427 and w40465;
w40485 <= not w4989 and not w40462;
w40486 <= not w40484 and w40485;
w40487 <= not w40483 and not w40486;
w40488 <= not w38478 and not w40271;
w40489 <= not pi1156 and not w36140;
w40490 <= not w40488 and w40489;
w40491 <= pi1155 and not w36548;
w40492 <= w38515 and not w40491;
w40493 <= not pi1154 and w40279;
w40494 <= not w40492 and not w40493;
w40495 <= not w38528 and w40494;
w40496 <= w36042 and not w40495;
w40497 <= not pi1154 and not w36265;
w40498 <= w36108 and not w36139;
w40499 <= pi1154 and not w40498;
w40500 <= pi1091 and w36046;
w40501 <= not w40499 and w40500;
w40502 <= not w40497 and w40501;
w40503 <= pi0219 and not w40490;
w40504 <= not w40502 and w40503;
w40505 <= not w40496 and w40504;
w40506 <= not pi0211 and not w40494;
w40507 <= w36131 and not w36674;
w40508 <= w39987 and not w40507;
w40509 <= not w36329 and w40508;
w40510 <= not w40506 and not w40509;
w40511 <= pi1156 and not w40510;
w40512 <= not w36329 and not w40488;
w40513 <= pi0211 and w40512;
w40514 <= not w36140 and not w36563;
w40515 <= w40018 and w40514;
w40516 <= not w40513 and not w40515;
w40517 <= not pi1156 and not w40516;
w40518 <= not pi0219 and not w40517;
w40519 <= not w40511 and w40518;
w40520 <= not w40505 and not w40519;
w40521 <= not pi0263 and not w40520;
w40522 <= not pi1154 and w36209;
w40523 <= pi1154 and not w36154;
w40524 <= pi1156 and not w40523;
w40525 <= not pi0299 and not w40524;
w40526 <= not w37417 and not w40522;
w40527 <= not w40525 and w40526;
w40528 <= pi1156 and not w40527;
w40529 <= not w40514 and w40525;
w40530 <= pi0219 and not w40529;
w40531 <= not w40528 and w40530;
w40532 <= not w36211 and w37062;
w40533 <= not w36563 and not w40532;
w40534 <= not pi0211 and not w40533;
w40535 <= not pi1156 and w40512;
w40536 <= not w36131 and not w36158;
w40537 <= pi1154 and not w40536;
w40538 <= not w36107 and w40497;
w40539 <= pi1156 and not w40537;
w40540 <= not w40538 and w40539;
w40541 <= pi0211 and not w40535;
w40542 <= not w40540 and w40541;
w40543 <= not pi0219 and not w40534;
w40544 <= not w40542 and w40543;
w40545 <= pi0263 and pi1091;
w40546 <= not w40531 and w40545;
w40547 <= not w40544 and w40546;
w40548 <= not w40521 and not w40547;
w40549 <= w4989 and w40548;
w40550 <= pi0219 and not w36046;
w40551 <= not pi0219 and not w36047;
w40552 <= not w36058 and w40551;
w40553 <= not w40550 and not w40552;
w40554 <= pi1091 and not w40553;
w40555 <= pi0263 and not pi1091;
w40556 <= not w40554 and not w40555;
w40557 <= not w4989 and not w40556;
w40558 <= not w38473 and not w40557;
w40559 <= not w40549 and w40558;
w40560 <= pi1091 and w40550;
w40561 <= pi0211 and w38437;
w40562 <= not pi0211 and not w40271;
w40563 <= not w36047 and not w40562;
w40564 <= not w40561 and w40563;
w40565 <= not w38453 and not w40564;
w40566 <= not pi0219 and not w40565;
w40567 <= not pi0263 and not w40295;
w40568 <= not w40566 and w40567;
w40569 <= not w36047 and not w40233;
w40570 <= not w40561 and not w40569;
w40571 <= w40097 and not w40570;
w40572 <= pi0263 and not w40101;
w40573 <= not w40571 and w40572;
w40574 <= not w40568 and not w40573;
w40575 <= w38423 and not w40560;
w40576 <= not w40574 and w40575;
w40577 <= not w38423 and w40556;
w40578 <= not w4989 and not w40577;
w40579 <= not w40576 and w40578;
w40580 <= not w38423 and not w40548;
w40581 <= pi1155 and not w38681;
w40582 <= pi1154 and not w40581;
w40583 <= w38668 and w40582;
w40584 <= not pi1155 and w40159;
w40585 <= pi1155 and not w38572;
w40586 <= not pi1154 and not w40585;
w40587 <= not w40584 and w40586;
w40588 <= not w38679 and w40584;
w40589 <= pi1155 and not w38635;
w40590 <= not pi1154 and not w40589;
w40591 <= not w40588 and w40590;
w40592 <= not pi1156 and not w40591;
w40593 <= not w40583 and not w40587;
w40594 <= w40592 and w40593;
w40595 <= not pi1155 and w38563;
w40596 <= not w38607 and w38665;
w40597 <= not w40595 and not w40596;
w40598 <= not pi1154 and not w40597;
w40599 <= pi1156 and not w40598;
w40600 <= w38563 and w40586;
w40601 <= not w38546 and w40583;
w40602 <= not w40600 and not w40601;
w40603 <= w40599 and w40602;
w40604 <= not pi0211 and not w40594;
w40605 <= not w40603 and w40604;
w40606 <= w38551 and w40582;
w40607 <= w40599 and not w40606;
w40608 <= w40064 and w40582;
w40609 <= w40592 and not w40608;
w40610 <= pi0211 and not w40607;
w40611 <= not w40609 and w40610;
w40612 <= not pi0219 and not w40605;
w40613 <= not w40611 and w40612;
w40614 <= pi1155 and w38571;
w40615 <= pi1154 and w38591;
w40616 <= not w40614 and w40615;
w40617 <= not w38548 and w40616;
w40618 <= not w40600 and not w40617;
w40619 <= w36042 and not w40618;
w40620 <= not w40587 and not w40616;
w40621 <= not pi1156 and not w40620;
w40622 <= not pi1154 and w38602;
w40623 <= not w38625 and not w40622;
w40624 <= w36046 and not w40614;
w40625 <= not w40623 and w40624;
w40626 <= pi0219 and not w40625;
w40627 <= not w40619 and w40626;
w40628 <= not w40621 and w40627;
w40629 <= not pi0263 and not w40628;
w40630 <= not w40613 and w40629;
w40631 <= not w38603 and not w38618;
w40632 <= pi1154 and not w40631;
w40633 <= pi1155 and not w40323;
w40634 <= not pi1155 and not w40074;
w40635 <= not pi1154 and not w40633;
w40636 <= not w40634 and w40635;
w40637 <= w36046 and not w40632;
w40638 <= not w40636 and w40637;
w40639 <= not w38577 and not w40385;
w40640 <= not w40631 and not w40639;
w40641 <= w36042 and not w40640;
w40642 <= not w38589 and w40640;
w40643 <= not pi1156 and not w40642;
w40644 <= pi0219 and not w40638;
w40645 <= not w40641 and w40644;
w40646 <= not w40643 and w40645;
w40647 <= pi1154 and not w38661;
w40648 <= not w38609 and w40647;
w40649 <= not pi1154 and not w38648;
w40650 <= pi1155 and w40388;
w40651 <= w40649 and not w40650;
w40652 <= not w38677 and w40647;
w40653 <= not pi1156 and not w40374;
w40654 <= not w40652 and w40653;
w40655 <= not pi1156 and not w40654;
w40656 <= not w40651 and not w40655;
w40657 <= pi1156 and w40391;
w40658 <= not w40656 and not w40657;
w40659 <= not w40648 and not w40658;
w40660 <= pi0211 and not w40659;
w40661 <= not w38589 and w38654;
w40662 <= pi1155 and w40661;
w40663 <= w40649 and not w40662;
w40664 <= not w40391 and w40663;
w40665 <= pi1156 and not w40664;
w40666 <= not w40652 and w40665;
w40667 <= w40654 and not w40663;
w40668 <= not pi0211 and not w40666;
w40669 <= not w40667 and w40668;
w40670 <= not pi0219 and not w40669;
w40671 <= not w40660 and w40670;
w40672 <= pi0263 and not w40646;
w40673 <= not w40671 and w40672;
w40674 <= w38423 and not w40630;
w40675 <= not w40673 and w40674;
w40676 <= w4989 and not w40580;
w40677 <= not w40675 and w40676;
w40678 <= w38473 and not w40579;
w40679 <= not w40677 and w40678;
w40680 <= not pi0230 and not w40559;
w40681 <= not w40679 and w40680;
w40682 <= not w4989 and w40553;
w40683 <= not w36141 and w36212;
w40684 <= not pi1156 and not w40683;
w40685 <= w36155 and not w36675;
w40686 <= not w40684 and w40685;
w40687 <= pi1156 and w37417;
w40688 <= pi0219 and not w40687;
w40689 <= not w40686 and w40688;
w40690 <= not w36073 and not w40686;
w40691 <= pi0211 and not w40690;
w40692 <= w40543 and not w40691;
w40693 <= w4989 and not w40689;
w40694 <= not w40692 and w40693;
w40695 <= pi0230 and not w40682;
w40696 <= not w40694 and w40695;
w40697 <= not w40681 and not w40696;
w40698 <= pi1091 and pi1143;
w40699 <= not pi0200 and w40698;
w40700 <= not pi0796 and w38426;
w40701 <= pi0264 and not w38426;
w40702 <= not pi1091 and not w40700;
w40703 <= not w40701 and w40702;
w40704 <= pi0199 and not w40699;
w40705 <= not w40703 and w40704;
w40706 <= pi1091 and pi1141;
w40707 <= not pi0796 and w38448;
w40708 <= pi0264 and not w38448;
w40709 <= not pi1091 and not w40707;
w40710 <= not w40708 and w40709;
w40711 <= not w40706 and not w40710;
w40712 <= not pi0200 and not w40711;
w40713 <= pi1091 and pi1142;
w40714 <= not w40710 and not w40713;
w40715 <= pi0200 and not w40714;
w40716 <= not pi0199 and not w40712;
w40717 <= not w40715 and w40716;
w40718 <= w14042 and not w40705;
w40719 <= not w40717 and w40718;
w40720 <= pi0219 and not w40018;
w40721 <= not w36973 and not w40720;
w40722 <= not w40703 and not w40721;
w40723 <= not pi0211 and not w40711;
w40724 <= pi0211 and not w40714;
w40725 <= not pi0219 and not w40723;
w40726 <= not w40724 and w40725;
w40727 <= not w14042 and not w40722;
w40728 <= not w40726 and w40727;
w40729 <= not w40719 and not w40728;
w40730 <= not pi0230 and not w40729;
w40731 <= not pi0211 and pi1141;
w40732 <= not pi0219 and not w36018;
w40733 <= not w40731 and w40732;
w40734 <= not w36973 and not w40733;
w40735 <= not w14042 and not w40734;
w40736 <= not pi0199 and pi1141;
w40737 <= w36951 and not w40736;
w40738 <= not w36007 and not w40737;
w40739 <= w14042 and not w40738;
w40740 <= pi0230 and not w40735;
w40741 <= not w40739 and w40740;
w40742 <= not w40730 and not w40741;
w40743 <= pi1091 and pi1144;
w40744 <= not pi0200 and w40743;
w40745 <= not pi0819 and w38426;
w40746 <= pi0265 and not w38426;
w40747 <= not pi1091 and not w40745;
w40748 <= not w40746 and w40747;
w40749 <= pi0199 and not w40744;
w40750 <= not w40748 and w40749;
w40751 <= not pi0819 and w38448;
w40752 <= pi0265 and not w38448;
w40753 <= not pi1091 and not w40751;
w40754 <= not w40752 and w40753;
w40755 <= not w40713 and not w40754;
w40756 <= not pi0200 and not w40755;
w40757 <= not w40698 and not w40754;
w40758 <= pi0200 and not w40757;
w40759 <= not pi0199 and not w40756;
w40760 <= not w40758 and w40759;
w40761 <= w14042 and not w40750;
w40762 <= not w40760 and w40761;
w40763 <= not w38334 and not w40720;
w40764 <= not w40748 and not w40763;
w40765 <= not pi0211 and not w40755;
w40766 <= pi0211 and not w40757;
w40767 <= not pi0219 and not w40765;
w40768 <= not w40766 and w40767;
w40769 <= not w14042 and not w40764;
w40770 <= not w40768 and w40769;
w40771 <= not w40762 and not w40770;
w40772 <= not pi0230 and not w40771;
w40773 <= not pi0211 and pi1142;
w40774 <= not pi0219 and not w35981;
w40775 <= not w40773 and w40774;
w40776 <= not w38334 and not w40775;
w40777 <= not w14042 and not w40776;
w40778 <= not w36006 and w38345;
w40779 <= not w36000 and not w40778;
w40780 <= w14042 and not w40779;
w40781 <= pi0230 and not w40777;
w40782 <= not w40780 and w40781;
w40783 <= not w40772 and not w40782;
w40784 <= not pi0211 and pi1136;
w40785 <= pi0219 and not w40784;
w40786 <= pi0211 and not pi1135;
w40787 <= not w40785 and not w40786;
w40788 <= not w8407 and w40787;
w40789 <= not w4989 and w40788;
w40790 <= pi0299 and w40788;
w40791 <= not pi0199 and pi1135;
w40792 <= pi0200 and not w40791;
w40793 <= pi0199 and pi1136;
w40794 <= not pi0200 and not w40793;
w40795 <= not pi0299 and not w40792;
w40796 <= not w40794 and w40795;
w40797 <= not w40790 and not w40796;
w40798 <= w4989 and not w40797;
w40799 <= pi0230 and not w40789;
w40800 <= not w40798 and w40799;
w40801 <= not w40720 and not w40785;
w40802 <= not pi0266 and not w38426;
w40803 <= not pi0948 and w38426;
w40804 <= not pi1091 and not w40802;
w40805 <= not w40803 and w40804;
w40806 <= not w40801 and not w40805;
w40807 <= not w14042 and not w40806;
w40808 <= not pi0266 and not w38448;
w40809 <= not pi0948 and w38448;
w40810 <= not pi1091 and not w40808;
w40811 <= not w40809 and w40810;
w40812 <= not pi0219 and not w40811;
w40813 <= pi1135 and w39987;
w40814 <= w40812 and not w40813;
w40815 <= w40807 and not w40814;
w40816 <= not pi0199 and not w40811;
w40817 <= pi1091 and pi1136;
w40818 <= pi0199 and not w40805;
w40819 <= not w40817 and w40818;
w40820 <= not w40816 and not w40819;
w40821 <= not pi0200 and w40820;
w40822 <= pi1091 and pi1135;
w40823 <= w40816 and not w40822;
w40824 <= pi0200 and not w40818;
w40825 <= not w40823 and w40824;
w40826 <= not w40821 and not w40825;
w40827 <= w14042 and not w40826;
w40828 <= not pi0230 and not w40815;
w40829 <= not w40827 and w40828;
w40830 <= not w40800 and not w40829;
w40831 <= not pi1134 and not w40830;
w40832 <= w36262 and not w40793;
w40833 <= not w40792 and not w40832;
w40834 <= w14042 and w40833;
w40835 <= not w14042 and w40787;
w40836 <= pi0230 and not w40834;
w40837 <= not w40835 and w40836;
w40838 <= pi1091 and not w40786;
w40839 <= w40812 and not w40838;
w40840 <= w40807 and not w40839;
w40841 <= not pi0199 and pi1091;
w40842 <= not w40820 and not w40841;
w40843 <= not pi0200 and not w40842;
w40844 <= not w40825 and not w40843;
w40845 <= w14042 and not w40844;
w40846 <= not pi0230 and not w40840;
w40847 <= not w40845 and w40846;
w40848 <= not w40837 and not w40847;
w40849 <= pi1134 and not w40848;
w40850 <= not w40831 and not w40849;
w40851 <= pi1155 and not w39994;
w40852 <= not w40269 and w40851;
w40853 <= not pi1155 and not w36590;
w40854 <= pi1091 and w40853;
w40855 <= not w40852 and not w40854;
w40856 <= not pi1154 and not w40855;
w40857 <= w40279 and w40851;
w40858 <= not pi1155 and not w40223;
w40859 <= not w40023 and w40858;
w40860 <= not w40857 and not w40859;
w40861 <= pi1154 and not w40860;
w40862 <= not pi0219 and not w40856;
w40863 <= not w40861 and w40862;
w40864 <= pi1153 and w36518;
w40865 <= w40271 and not w40864;
w40866 <= not w37231 and w40865;
w40867 <= pi1091 and w40491;
w40868 <= not w39993 and w40867;
w40869 <= pi1154 and not w40868;
w40870 <= not pi0299 and w36509;
w40871 <= pi1091 and not w40870;
w40872 <= w40869 and w40871;
w40873 <= pi0219 and not w40866;
w40874 <= not w40872 and w40873;
w40875 <= not w40863 and not w40874;
w40876 <= not pi0211 and not w40875;
w40877 <= pi1155 and w36526;
w40878 <= pi1154 and not w40877;
w40879 <= not pi1155 and not w36510;
w40880 <= not w36145 and not w40879;
w40881 <= not w10625 and not w40880;
w40882 <= pi1091 and w40878;
w40883 <= not w40881 and w40882;
w40884 <= not w36264 and not w38482;
w40885 <= w40865 and not w40884;
w40886 <= pi0211 and not w40885;
w40887 <= not w40883 and w40886;
w40888 <= not w40876 and not w40887;
w40889 <= pi0267 and not w40888;
w40890 <= w36131 and w40011;
w40891 <= not w40248 and not w40890;
w40892 <= not w40853 and not w40891;
w40893 <= pi0211 and not pi1154;
w40894 <= not w40892 and w40893;
w40895 <= pi1091 and not pi1155;
w40896 <= not w36510 and w40895;
w40897 <= w36051 and not w40896;
w40898 <= not w40868 and w40897;
w40899 <= not pi1154 and w36108;
w40900 <= not w36233 and not w40899;
w40901 <= not w36246 and w40900;
w40902 <= pi1091 and w40901;
w40903 <= not pi0211 and not w40902;
w40904 <= not pi0219 and not w40898;
w40905 <= not w40903 and w40904;
w40906 <= w40870 and w40895;
w40907 <= w40869 and not w40906;
w40908 <= w40491 and w40878;
w40909 <= not w40907 and not w40908;
w40910 <= pi0211 and not w40909;
w40911 <= pi1154 and not w40907;
w40912 <= not w36264 and w40271;
w40913 <= not w37230 and w40912;
w40914 <= not pi0211 and not w40913;
w40915 <= not w40911 and w40914;
w40916 <= pi0219 and not w40910;
w40917 <= not w40915 and w40916;
w40918 <= not w40905 and not w40917;
w40919 <= not pi0267 and not w40894;
w40920 <= not w40918 and w40919;
w40921 <= not w40889 and not w40920;
w40922 <= w4989 and w40921;
w40923 <= not pi0219 and not w36051;
w40924 <= not w36060 and w40923;
w40925 <= not w36721 and not w40924;
w40926 <= pi1091 and not w40925;
w40927 <= not pi0267 and not pi1091;
w40928 <= not w40926 and not w40927;
w40929 <= not w4989 and not w40928;
w40930 <= not w38473 and not w40929;
w40931 <= not w40922 and w40930;
w40932 <= not pi0267 and not w38543;
w40933 <= not w40101 and w40932;
w40934 <= pi0267 and w40297;
w40935 <= w38422 and not w40933;
w40936 <= not w40934 and w40935;
w40937 <= not w38422 and w40927;
w40938 <= not w40926 and not w40937;
w40939 <= not w40936 and w40938;
w40940 <= not w4989 and not w40939;
w40941 <= not w38422 and not w40921;
w40942 <= not w40340 and w40343;
w40943 <= w40368 and not w40942;
w40944 <= pi1154 and pi1155;
w40945 <= not w38577 and w40944;
w40946 <= not w40345 and w40945;
w40947 <= not w40943 and not w40946;
w40948 <= pi0211 and not w40947;
w40949 <= pi1153 and w38618;
w40950 <= w36050 and not w40074;
w40951 <= not w40949 and w40950;
w40952 <= not w40324 and w40951;
w40953 <= w38602 and w40312;
w40954 <= not pi1155 and not w40953;
w40955 <= not w40942 and w40954;
w40956 <= not pi0267 and not w40955;
w40957 <= not w40952 and w40956;
w40958 <= not w40948 and w40957;
w40959 <= pi1155 and not w40146;
w40960 <= w38571 and not w40622;
w40961 <= w40959 and not w40960;
w40962 <= not w40161 and w40961;
w40963 <= not w40064 and not w40080;
w40964 <= w38572 and not w40963;
w40965 <= pi1154 and not w40964;
w40966 <= not pi1154 and not w38591;
w40967 <= not w40160 and w40966;
w40968 <= not pi1155 and not w40967;
w40969 <= not w40965 and w40968;
w40970 <= pi0267 and not w40962;
w40971 <= not w40969 and w40970;
w40972 <= not w40958 and not w40971;
w40973 <= pi0219 and not w40972;
w40974 <= not pi1155 and not w40388;
w40975 <= not w40942 and w40974;
w40976 <= w38635 and not w40964;
w40977 <= w40633 and not w40976;
w40978 <= pi1154 and not w40977;
w40979 <= not pi1154 and not w40060;
w40980 <= pi1155 and not w40979;
w40981 <= w38608 and not w40980;
w40982 <= not w40978 and not w40981;
w40983 <= pi0211 and not w40975;
w40984 <= not w40982 and w40983;
w40985 <= not w40391 and not w40949;
w40986 <= pi1155 and not w40985;
w40987 <= pi1153 and not w38679;
w40988 <= not pi1155 and not w40987;
w40989 <= w40168 and w40988;
w40990 <= not pi1154 and not w40986;
w40991 <= not w40989 and w40990;
w40992 <= not pi1153 and not w40661;
w40993 <= w40988 and not w40992;
w40994 <= pi1154 and not w40662;
w40995 <= not w40986 and w40994;
w40996 <= not w40993 and w40995;
w40997 <= not pi0211 and not w40991;
w40998 <= not w40996 and w40997;
w40999 <= not pi0267 and not w40998;
w41000 <= not w40984 and w40999;
w41001 <= not pi1153 and w38656;
w41002 <= not w38681 and not w41001;
w41003 <= not pi1155 and w38635;
w41004 <= not w41002 and w41003;
w41005 <= w40596 and w40959;
w41006 <= pi1154 and not w41004;
w41007 <= not w41005 and w41006;
w41008 <= not pi1154 and not w40080;
w41009 <= not w38668 and w41008;
w41010 <= not pi1155 and not w41009;
w41011 <= not w38551 and w41008;
w41012 <= not w41010 and w41011;
w41013 <= not w41007 and not w41012;
w41014 <= pi0211 and not w41013;
w41015 <= pi1154 and w41002;
w41016 <= w41010 and not w41015;
w41017 <= pi1154 and w38571;
w41018 <= not w38654 and not w40367;
w41019 <= pi1155 and not w41017;
w41020 <= not w41018 and w41019;
w41021 <= not pi0211 and not w41020;
w41022 <= not w41016 and w41021;
w41023 <= pi0267 and not w41022;
w41024 <= not w41014 and w41023;
w41025 <= not pi0219 and not w41024;
w41026 <= not w41000 and w41025;
w41027 <= not w40973 and not w41026;
w41028 <= w38422 and not w41027;
w41029 <= w4989 and not w40941;
w41030 <= not w41028 and w41029;
w41031 <= w38473 and not w40940;
w41032 <= not w41030 and w41031;
w41033 <= not pi0230 and not w40931;
w41034 <= not w41032 and w41033;
w41035 <= pi0219 and not w36526;
w41036 <= not pi1155 and w40864;
w41037 <= not pi1154 and not w41036;
w41038 <= not w36510 and not w41037;
w41039 <= pi1155 and w37228;
w41040 <= not w41038 and not w41039;
w41041 <= not w41035 and not w41040;
w41042 <= pi0211 and not w41041;
w41043 <= not pi0199 and pi1154;
w41044 <= pi0200 and not w41043;
w41045 <= not w36294 and not w36525;
w41046 <= not w41044 and w41045;
w41047 <= not w36073 and not w41046;
w41048 <= pi0219 and not w41047;
w41049 <= not pi0219 and w40901;
w41050 <= not pi0211 and not w41049;
w41051 <= not w41048 and w41050;
w41052 <= w4989 and not w41051;
w41053 <= not w41042 and w41052;
w41054 <= not w4989 and w40925;
w41055 <= pi0230 and not w41054;
w41056 <= not w41053 and w41055;
w41057 <= not w41034 and not w41056;
w41058 <= pi0268 and pi1152;
w41059 <= not pi0211 and not w14042;
w41060 <= w4989 and w36131;
w41061 <= not w41059 and not w41060;
w41062 <= not pi1151 and w41061;
w41063 <= not pi0199 and w14042;
w41064 <= not w37704 and not w41063;
w41065 <= pi1152 and not w41061;
w41066 <= w41064 and not w41065;
w41067 <= pi1150 and not w41062;
w41068 <= not w41066 and w41067;
w41069 <= not w41058 and w41068;
w41070 <= not pi1151 and w39952;
w41071 <= w4989 and not w9011;
w41072 <= not w4989 and w9009;
w41073 <= not w41071 and not w41072;
w41074 <= pi1151 and not w41073;
w41075 <= not pi1152 and not w41074;
w41076 <= not w14042 and w40041;
w41077 <= w4989 and w36144;
w41078 <= not w41076 and not w41077;
w41079 <= pi1151 and not w41078;
w41080 <= pi1152 and w41079;
w41081 <= not pi1150 and not w41070;
w41082 <= not w41075 and w41081;
w41083 <= not w41080 and w41082;
w41084 <= not w41069 and not w41083;
w41085 <= pi1091 and not w41084;
w41086 <= pi1152 and w41068;
w41087 <= pi1091 and not w41086;
w41088 <= pi0268 and not w41087;
w41089 <= not w41085 and not w41088;
w41090 <= not w38472 and not w41089;
w41091 <= not w40090 and w40135;
w41092 <= not w38575 and w40147;
w41093 <= pi0219 and not w40076;
w41094 <= not w38574 and w41093;
w41095 <= not w41092 and not w41094;
w41096 <= w4989 and not w40068;
w41097 <= w41095 and w41096;
w41098 <= not w41091 and not w41097;
w41099 <= not pi1151 and not w41098;
w41100 <= w4989 and not w40169;
w41101 <= pi0219 and w38611;
w41102 <= w41100 and not w41101;
w41103 <= w40135 and not w40296;
w41104 <= not w41102 and not w41103;
w41105 <= pi1151 and not w41104;
w41106 <= not w41099 and not w41105;
w41107 <= pi0268 and not w41106;
w41108 <= not w4989 and not w40101;
w41109 <= not w40132 and w41108;
w41110 <= not w4989 and not w40295;
w41111 <= not w40088 and w41110;
w41112 <= w41109 and not w41111;
w41113 <= pi0219 and not w38557;
w41114 <= not w40111 and not w41113;
w41115 <= not w38556 and not w41114;
w41116 <= w4989 and not w38589;
w41117 <= w41115 and w41116;
w41118 <= not w41112 and not w41117;
w41119 <= not pi1151 and w41118;
w41120 <= not w38437 and not w41104;
w41121 <= pi0219 and not w4989;
w41122 <= not w38431 and w41121;
w41123 <= not w38595 and w41100;
w41124 <= not w40097 and not w41122;
w41125 <= not w41123 and w41124;
w41126 <= not w41120 and not w41125;
w41127 <= pi1151 and w41126;
w41128 <= not pi0268 and not w41127;
w41129 <= not w41119 and w41128;
w41130 <= not w41107 and not w41129;
w41131 <= not pi1152 and not w41130;
w41132 <= not w40090 and w41110;
w41133 <= not w38625 and not w40162;
w41134 <= not w41095 and not w41133;
w41135 <= w4989 and not w41134;
w41136 <= not w38431 and not w40150;
w41137 <= w41135 and not w41136;
w41138 <= not w41132 and not w41137;
w41139 <= not pi1151 and not w41138;
w41140 <= not w38433 and w41096;
w41141 <= not w40296 and w41110;
w41142 <= not w41102 and not w41141;
w41143 <= not w41140 and w41142;
w41144 <= pi1151 and not w41143;
w41145 <= pi0268 and not w41144;
w41146 <= not w41139 and w41145;
w41147 <= not w40075 and not w41115;
w41148 <= w4989 and not w41147;
w41149 <= not w41109 and not w41148;
w41150 <= not pi1151 and not w41149;
w41151 <= not w40091 and w41108;
w41152 <= not pi0219 and w38660;
w41153 <= not w41093 and not w41152;
w41154 <= w4989 and not w41153;
w41155 <= not w41112 and not w41151;
w41156 <= not w41154 and w41155;
w41157 <= pi1151 and not w41156;
w41158 <= not pi0268 and not w41157;
w41159 <= not w41150 and w41158;
w41160 <= pi1152 and not w41159;
w41161 <= not w41146 and w41160;
w41162 <= not w41131 and not w41161;
w41163 <= pi1150 and not w41162;
w41164 <= not w40097 and w41108;
w41165 <= not pi0219 and not w38608;
w41166 <= not w38565 and not w41165;
w41167 <= w41154 and w41166;
w41168 <= not w41164 and not w41167;
w41169 <= not pi1151 and not w41168;
w41170 <= w4989 and not w41095;
w41171 <= not w41151 and not w41170;
w41172 <= pi1151 and not w41171;
w41173 <= pi1152 and not w41169;
w41174 <= not w41172 and w41173;
w41175 <= not pi1151 and w41125;
w41176 <= not w40092 and not w41122;
w41177 <= not w41135 and w41176;
w41178 <= pi1151 and w41177;
w41179 <= not pi1152 and not w41175;
w41180 <= not w41178 and w41179;
w41181 <= not w41174 and not w41180;
w41182 <= not pi0268 and not w41181;
w41183 <= pi0219 and not w40161;
w41184 <= w4989 and not w40162;
w41185 <= not w41183 and w41184;
w41186 <= not w41111 and not w41185;
w41187 <= not pi1151 and w41186;
w41188 <= not w40133 and w41110;
w41189 <= not w40111 and not w41183;
w41190 <= w38665 and not w41189;
w41191 <= w4989 and not w41190;
w41192 <= not w41188 and not w41191;
w41193 <= pi1151 and w41192;
w41194 <= pi1152 and not w41187;
w41195 <= not w41193 and w41194;
w41196 <= w38437 and not w41104;
w41197 <= not pi1151 and not w41196;
w41198 <= w4989 and not w40116;
w41199 <= not w40111 and w41198;
w41200 <= not w40136 and not w41199;
w41201 <= pi1151 and w41200;
w41202 <= not pi1152 and not w41197;
w41203 <= not w41201 and w41202;
w41204 <= pi0268 and not w41203;
w41205 <= not w41195 and w41204;
w41206 <= not pi1150 and not w41205;
w41207 <= not w41182 and w41206;
w41208 <= not w41163 and not w41207;
w41209 <= w38472 and not w41208;
w41210 <= not pi0230 and not w41090;
w41211 <= not w41209 and w41210;
w41212 <= pi0230 and not w41068;
w41213 <= not w41083 and w41212;
w41214 <= not w41211 and not w41213;
w41215 <= not pi0199 and pi1137;
w41216 <= pi0200 and not w41215;
w41217 <= pi0199 and pi1138;
w41218 <= not pi0199 and pi1136;
w41219 <= not pi0200 and not w41217;
w41220 <= not w41218 and w41219;
w41221 <= not w41216 and not w41220;
w41222 <= w14042 and not w41221;
w41223 <= not pi0211 and pi1138;
w41224 <= pi0219 and w41223;
w41225 <= pi0211 and pi1137;
w41226 <= not w40784 and not w41225;
w41227 <= not pi0219 and not w41226;
w41228 <= not w41224 and not w41227;
w41229 <= not w14042 and w41228;
w41230 <= not w41222 and not w41229;
w41231 <= pi0230 and not w41230;
w41232 <= not pi0200 and w40817;
w41233 <= pi1137 and w38514;
w41234 <= not w41232 and not w41233;
w41235 <= w41063 and w41234;
w41236 <= pi1091 and not w41226;
w41237 <= w37704 and not w41236;
w41238 <= not w41235 and not w41237;
w41239 <= not pi0817 and w38448;
w41240 <= pi0269 and not w38448;
w41241 <= not pi1091 and not w41239;
w41242 <= not w41240 and w41241;
w41243 <= not w41238 and not w41242;
w41244 <= not pi0817 and w38426;
w41245 <= pi0269 and not w38426;
w41246 <= not pi1091 and not w41244;
w41247 <= not w41245 and w41246;
w41248 <= pi1138 and w40018;
w41249 <= pi0219 and not w14042;
w41250 <= not w41248 and w41249;
w41251 <= not pi0200 and pi1091;
w41252 <= pi1138 and w41251;
w41253 <= pi0199 and not w41252;
w41254 <= w14042 and w41253;
w41255 <= not w41250 and not w41254;
w41256 <= not w41247 and not w41255;
w41257 <= not w41243 and not w41256;
w41258 <= not pi0230 and not w41257;
w41259 <= not w41231 and not w41258;
w41260 <= not pi0805 and w38426;
w41261 <= pi0270 and not w38426;
w41262 <= not pi1091 and not w41260;
w41263 <= not w41261 and w41262;
w41264 <= w40018 and w40731;
w41265 <= w41249 and not w41264;
w41266 <= not pi0200 and w40706;
w41267 <= pi0199 and not w41266;
w41268 <= w14042 and w41267;
w41269 <= not w41265 and not w41268;
w41270 <= not w41263 and not w41269;
w41271 <= not pi0805 and w38448;
w41272 <= pi0270 and not w38448;
w41273 <= not pi1091 and not w41271;
w41274 <= not w41272 and w41273;
w41275 <= not pi0211 and pi1139;
w41276 <= pi0211 and pi1140;
w41277 <= not w41275 and not w41276;
w41278 <= pi1091 and not w41277;
w41279 <= w37704 and not w41278;
w41280 <= pi1091 and pi1140;
w41281 <= pi0200 and w41280;
w41282 <= pi1139 and w41251;
w41283 <= not w41281 and not w41282;
w41284 <= w41063 and w41283;
w41285 <= not w41279 and not w41284;
w41286 <= not w41274 and not w41285;
w41287 <= not pi0230 and not w41270;
w41288 <= not w41286 and w41287;
w41289 <= pi0219 and not w40731;
w41290 <= not pi0219 and w41277;
w41291 <= not w41289 and not w41290;
w41292 <= not w14042 and not w41291;
w41293 <= not pi0199 and pi1140;
w41294 <= pi0200 and not w41293;
w41295 <= pi0199 and pi1141;
w41296 <= not pi0199 and pi1139;
w41297 <= not pi0200 and not w41295;
w41298 <= not w41296 and w41297;
w41299 <= not w41294 and not w41298;
w41300 <= w14042 and not w41299;
w41301 <= pi0230 and not w41292;
w41302 <= not w41300 and w41301;
w41303 <= not w41288 and not w41302;
w41304 <= not pi0211 and pi1147;
w41305 <= w40007 and w41304;
w41306 <= not pi0271 and not w38429;
w41307 <= not w38434 and not w41306;
w41308 <= pi0219 and not w41307;
w41309 <= not pi1091 and not w38450;
w41310 <= pi0271 and not w41309;
w41311 <= not pi0271 and not w38451;
w41312 <= not w41310 and not w41311;
w41313 <= pi1091 and pi1146;
w41314 <= not w41312 and not w41313;
w41315 <= not pi0211 and w41313;
w41316 <= not w41314 and not w41315;
w41317 <= pi1091 and w36975;
w41318 <= not pi0219 and not w41317;
w41319 <= not w41316 and w41318;
w41320 <= not w41308 and not w41319;
w41321 <= not w14042 and not w41305;
w41322 <= not w41320 and w41321;
w41323 <= pi0199 and not w41307;
w41324 <= not pi0199 and w41314;
w41325 <= not w41323 and not w41324;
w41326 <= pi0200 and not w41325;
w41327 <= pi1147 and w38494;
w41328 <= pi1091 and pi1145;
w41329 <= not pi0199 and not w41328;
w41330 <= not w41312 and w41329;
w41331 <= not w41323 and not w41330;
w41332 <= not pi0200 and not w41327;
w41333 <= not w41331 and w41332;
w41334 <= not w41326 and not w41333;
w41335 <= w14042 and not w41334;
w41336 <= not w41322 and not w41335;
w41337 <= not pi0230 and not w41336;
w41338 <= pi1147 and w39949;
w41339 <= not w37788 and not w37798;
w41340 <= not pi0219 and not w41339;
w41341 <= not pi0200 and not w36956;
w41342 <= w37902 and not w41341;
w41343 <= not w41338 and not w41340;
w41344 <= not w41342 and w41343;
w41345 <= w4989 and not w41344;
w41346 <= pi0219 and not w41304;
w41347 <= not w36975 and w39094;
w41348 <= not w41346 and not w41347;
w41349 <= not w4989 and w41348;
w41350 <= pi0230 and not w41349;
w41351 <= not w41345 and w41350;
w41352 <= not w41337 and not w41351;
w41353 <= not w4989 and w8407;
w41354 <= not w10628 and not w41353;
w41355 <= not pi1150 and w41354;
w41356 <= not w41061 and not w41355;
w41357 <= not pi1149 and not w41356;
w41358 <= pi1149 and not pi1150;
w41359 <= not w41061 and not w41358;
w41360 <= w41064 and not w41359;
w41361 <= not w41357 and not w41360;
w41362 <= pi1091 and not w41361;
w41363 <= pi1148 and not w41362;
w41364 <= pi1150 and not w39952;
w41365 <= not pi1149 and not w41364;
w41366 <= pi1091 and w41365;
w41367 <= not w14042 and w40275;
w41368 <= w4989 and w38499;
w41369 <= not w41367 and not w41368;
w41370 <= not pi1150 and w41369;
w41371 <= pi1091 and not w41078;
w41372 <= pi1150 and not w41371;
w41373 <= pi1149 and not w41370;
w41374 <= not w41372 and w41373;
w41375 <= not pi1148 and not w41366;
w41376 <= not w41374 and w41375;
w41377 <= not pi0283 and not w41363;
w41378 <= not w41376 and w41377;
w41379 <= not pi1150 and not w41196;
w41380 <= pi1150 and w41186;
w41381 <= not pi1149 and not w41379;
w41382 <= not w41380 and w41381;
w41383 <= pi1150 and w41192;
w41384 <= not pi1150 and w41200;
w41385 <= pi1149 and not w41384;
w41386 <= not w41383 and w41385;
w41387 <= not w41382 and not w41386;
w41388 <= not pi1148 and not w41387;
w41389 <= not pi1150 and w41104;
w41390 <= pi1150 and w41143;
w41391 <= pi1149 and not w41389;
w41392 <= not w41390 and w41391;
w41393 <= not pi1150 and w41098;
w41394 <= pi1150 and w41138;
w41395 <= not pi1149 and not w41393;
w41396 <= not w41394 and w41395;
w41397 <= not w41392 and not w41396;
w41398 <= pi1148 and not w41397;
w41399 <= pi0283 and not w41388;
w41400 <= not w41398 and w41399;
w41401 <= pi0272 and not w41378;
w41402 <= not w41400 and w41401;
w41403 <= not pi1150 and not w41126;
w41404 <= pi1150 and not w41156;
w41405 <= pi1149 and not w41403;
w41406 <= not w41404 and w41405;
w41407 <= pi1150 and not w41149;
w41408 <= not pi1150 and not w41118;
w41409 <= not pi1149 and not w41408;
w41410 <= not w41407 and w41409;
w41411 <= not w41406 and not w41410;
w41412 <= pi1148 and not w41411;
w41413 <= pi1150 and w41168;
w41414 <= not pi1150 and not w41125;
w41415 <= not pi1149 and not w41414;
w41416 <= not w41413 and w41415;
w41417 <= not pi1150 and not w41177;
w41418 <= pi1150 and w41171;
w41419 <= pi1149 and not w41418;
w41420 <= not w41417 and w41419;
w41421 <= not pi1148 and not w41416;
w41422 <= not w41420 and w41421;
w41423 <= not w41412 and not w41422;
w41424 <= pi0283 and not w41423;
w41425 <= w4989 and w36113;
w41426 <= not w37704 and not w41425;
w41427 <= not w41059 and w41426;
w41428 <= pi1150 and not w41427;
w41429 <= pi1149 and not w41428;
w41430 <= w41064 and w41429;
w41431 <= pi1148 and not w41357;
w41432 <= not w41430 and w41431;
w41433 <= pi1091 and w41432;
w41434 <= not pi1148 and not w41365;
w41435 <= not pi1150 and not w41073;
w41436 <= pi1150 and w41078;
w41437 <= pi1149 and not w41435;
w41438 <= not w41436 and w41437;
w41439 <= pi1091 and not w41438;
w41440 <= w41434 and w41439;
w41441 <= not pi0283 and not w41440;
w41442 <= not w41433 and w41441;
w41443 <= not pi0272 and not w41442;
w41444 <= not w41424 and w41443;
w41445 <= not pi0230 and not w41402;
w41446 <= not w41444 and w41445;
w41447 <= pi1149 and not w41078;
w41448 <= not w41429 and not w41447;
w41449 <= not w41435 and not w41448;
w41450 <= w41434 and not w41449;
w41451 <= pi0230 and not w41432;
w41452 <= not w41450 and w41451;
w41453 <= not w41446 and not w41452;
w41454 <= not pi0273 and not w38430;
w41455 <= not w38436 and not w41454;
w41456 <= pi0219 and not w41455;
w41457 <= not pi0273 and not w38452;
w41458 <= w38454 and not w41457;
w41459 <= not pi0219 and not w41315;
w41460 <= not w41458 and w41459;
w41461 <= not w41456 and not w41460;
w41462 <= not w4989 and w41461;
w41463 <= pi0299 and w41461;
w41464 <= pi0199 and not w41455;
w41465 <= not pi0200 and w41313;
w41466 <= not pi0199 and not w41465;
w41467 <= not w41458 and w41466;
w41468 <= not pi0299 and not w41464;
w41469 <= not w41467 and w41468;
w41470 <= not w41463 and not w41469;
w41471 <= not w9010 and not w38604;
w41472 <= pi1091 and not w41471;
w41473 <= w41470 and not w41472;
w41474 <= w4989 and not w41473;
w41475 <= pi1091 and w40136;
w41476 <= not w41474 and not w41475;
w41477 <= pi1147 and not w41476;
w41478 <= w38010 and not w41470;
w41479 <= not pi1148 and not w41478;
w41480 <= pi1091 and w36082;
w41481 <= not w41461 and not w41480;
w41482 <= pi0299 and not w41481;
w41483 <= w38495 and not w41326;
w41484 <= not w41469 and not w41483;
w41485 <= not w41482 and w41484;
w41486 <= w4989 and not w41485;
w41487 <= w37643 and w40007;
w41488 <= pi1148 and not w41487;
w41489 <= not w41486 and w41488;
w41490 <= not w41479 and not w41489;
w41491 <= not w41462 and not w41490;
w41492 <= not w41477 and w41491;
w41493 <= not pi0230 and not w41492;
w41494 <= pi1146 and not w38967;
w41495 <= not w41354 and w41494;
w41496 <= not pi0211 and not w37797;
w41497 <= w37704 and not w41496;
w41498 <= not pi1146 and w8372;
w41499 <= w41063 and not w41498;
w41500 <= not w41497 and not w41499;
w41501 <= pi1147 and not w41500;
w41502 <= not pi1148 and not w41495;
w41503 <= not w41501 and w41502;
w41504 <= not pi0199 and pi1147;
w41505 <= pi0200 and not w41504;
w41506 <= not w41498 and not w41505;
w41507 <= w14042 and w41506;
w41508 <= not pi1146 and w8407;
w41509 <= pi1147 and w37704;
w41510 <= not w41059 and not w41509;
w41511 <= not w41508 and not w41510;
w41512 <= pi1148 and not w41507;
w41513 <= not w41511 and w41512;
w41514 <= pi0230 and not w41503;
w41515 <= not w41513 and w41514;
w41516 <= not w41493 and not w41515;
w41517 <= not pi0200 and w41328;
w41518 <= not pi0659 and w38426;
w41519 <= pi0274 and not w38426;
w41520 <= not pi1091 and not w41518;
w41521 <= not w41519 and w41520;
w41522 <= pi0199 and not w41517;
w41523 <= not w41521 and w41522;
w41524 <= not pi0659 and w38448;
w41525 <= pi0274 and not w38448;
w41526 <= not pi1091 and not w41524;
w41527 <= not w41525 and w41526;
w41528 <= not w40743 and not w41527;
w41529 <= pi0200 and not w41528;
w41530 <= not w40698 and not w41527;
w41531 <= not pi0200 and not w41530;
w41532 <= not pi0199 and not w41529;
w41533 <= not w41531 and w41532;
w41534 <= w14042 and not w41523;
w41535 <= not w41533 and w41534;
w41536 <= pi0211 and not w41528;
w41537 <= not pi0211 and not w41530;
w41538 <= not pi0219 and not w41536;
w41539 <= not w41537 and w41538;
w41540 <= pi0219 and not w41317;
w41541 <= not w41521 and w41540;
w41542 <= not w14042 and not w41541;
w41543 <= not w41539 and w41542;
w41544 <= not pi0230 and not w41535;
w41545 <= not w41543 and w41544;
w41546 <= not w36071 and not w37788;
w41547 <= not pi0219 and not w35988;
w41548 <= not w36976 and w41547;
w41549 <= not w41546 and not w41548;
w41550 <= not w35999 and w37895;
w41551 <= w38351 and not w41550;
w41552 <= not w41549 and not w41551;
w41553 <= w4989 and not w41552;
w41554 <= not w37784 and not w41548;
w41555 <= pi0230 and not w41553;
w41556 <= not w41554 and w41555;
w41557 <= not w41545 and not w41556;
w41558 <= pi1151 and not w41061;
w41559 <= pi1149 and w41064;
w41560 <= not w41558 and w41559;
w41561 <= not pi1149 and w41079;
w41562 <= not w41560 and not w41561;
w41563 <= pi1150 and not w41562;
w41564 <= not pi1151 and w41354;
w41565 <= pi1149 and not w41061;
w41566 <= not w41564 and w41565;
w41567 <= not pi1149 and pi1151;
w41568 <= not w39952 and w41567;
w41569 <= not pi1150 and not w41568;
w41570 <= not w41566 and w41569;
w41571 <= not w41563 and not w41570;
w41572 <= pi1091 and not w41571;
w41573 <= not pi1151 and w39047;
w41574 <= not w41369 and w41573;
w41575 <= not w41572 and not w41574;
w41576 <= pi0275 and not w41575;
w41577 <= w41061 and w41358;
w41578 <= w38170 and not w39952;
w41579 <= not pi1151 and w41073;
w41580 <= pi1150 and not w41579;
w41581 <= not w41079 and w41580;
w41582 <= not pi1149 and not w41578;
w41583 <= not w41581 and w41582;
w41584 <= not w41560 and not w41577;
w41585 <= not w41583 and w41584;
w41586 <= pi1091 and w41585;
w41587 <= not pi0275 and not w41586;
w41588 <= not w38471 and not w41587;
w41589 <= not w41576 and w41588;
w41590 <= not pi1150 and w41168;
w41591 <= pi1151 and not w41418;
w41592 <= not w41590 and w41591;
w41593 <= pi1150 and not w41177;
w41594 <= not pi1151 and not w41414;
w41595 <= not w41593 and w41594;
w41596 <= not w41592 and not w41595;
w41597 <= not pi0275 and not w41596;
w41598 <= pi1150 and w41200;
w41599 <= not w41379 and not w41598;
w41600 <= not pi1151 and not w41599;
w41601 <= not pi1150 and w41186;
w41602 <= not w41383 and not w41601;
w41603 <= pi1151 and not w41602;
w41604 <= pi0275 and not w41600;
w41605 <= not w41603 and w41604;
w41606 <= not pi1149 and not w41605;
w41607 <= not w41597 and w41606;
w41608 <= pi1150 and not w41126;
w41609 <= not pi1151 and not w41608;
w41610 <= not w41408 and w41609;
w41611 <= not pi1150 and not w41149;
w41612 <= pi1151 and not w41404;
w41613 <= not w41611 and w41612;
w41614 <= not pi0275 and not w41610;
w41615 <= not w41613 and w41614;
w41616 <= pi1151 and not w41138;
w41617 <= not pi1150 and not w41099;
w41618 <= not w41616 and w41617;
w41619 <= not pi1151 and not w41104;
w41620 <= pi1150 and not w41619;
w41621 <= not w41144 and w41620;
w41622 <= pi0275 and not w41621;
w41623 <= not w41618 and w41622;
w41624 <= pi1149 and not w41615;
w41625 <= not w41623 and w41624;
w41626 <= w38471 and not w41607;
w41627 <= not w41625 and w41626;
w41628 <= not w41589 and not w41627;
w41629 <= not pi0230 and not w41628;
w41630 <= pi0230 and w41585;
w41631 <= not w41629 and not w41630;
w41632 <= not pi0276 and not w38449;
w41633 <= w41309 and not w41632;
w41634 <= not w35982 and not w37773;
w41635 <= pi1091 and not w41634;
w41636 <= w37704 and not w41635;
w41637 <= pi1145 and w38514;
w41638 <= not w40744 and not w41637;
w41639 <= w41063 and w41638;
w41640 <= not w41636 and not w41639;
w41641 <= not w41633 and not w41640;
w41642 <= not pi0276 and not w38427;
w41643 <= w38433 and not w41642;
w41644 <= w41249 and not w41315;
w41645 <= pi0199 and not w41465;
w41646 <= w14042 and w41645;
w41647 <= not w41644 and not w41646;
w41648 <= not w41643 and not w41647;
w41649 <= not pi0230 and not w41641;
w41650 <= not w41648 and w41649;
w41651 <= not w35997 and w38857;
w41652 <= not w37893 and not w41651;
w41653 <= w14042 and not w41652;
w41654 <= not pi0219 and not w41634;
w41655 <= pi1146 and w36082;
w41656 <= not w41654 and not w41655;
w41657 <= not w14042 and w41656;
w41658 <= pi0230 and not w41653;
w41659 <= not w41657 and w41658;
w41660 <= not w41650 and not w41659;
w41661 <= not pi0200 and w40713;
w41662 <= not pi0820 and w38426;
w41663 <= pi0277 and not w38426;
w41664 <= not pi1091 and not w41662;
w41665 <= not w41663 and w41664;
w41666 <= pi0199 and not w41661;
w41667 <= not w41665 and w41666;
w41668 <= not pi0820 and w38448;
w41669 <= pi0277 and not w38448;
w41670 <= not pi1091 and not w41668;
w41671 <= not w41669 and w41670;
w41672 <= not w41280 and not w41671;
w41673 <= not pi0200 and not w41672;
w41674 <= not w40706 and not w41671;
w41675 <= pi0200 and not w41674;
w41676 <= not pi0199 and not w41673;
w41677 <= not w41675 and w41676;
w41678 <= w14042 and not w41667;
w41679 <= not w41677 and w41678;
w41680 <= pi0219 and not w40773;
w41681 <= not w40720 and not w41680;
w41682 <= not w41665 and not w41681;
w41683 <= not pi0211 and not w41672;
w41684 <= pi0211 and not w41674;
w41685 <= not pi0219 and not w41683;
w41686 <= not w41684 and w41685;
w41687 <= not w14042 and not w41682;
w41688 <= not w41686 and w41687;
w41689 <= not w41679 and not w41688;
w41690 <= not pi0230 and not w41689;
w41691 <= pi0211 and pi1141;
w41692 <= not pi0211 and pi1140;
w41693 <= not pi0219 and not w41691;
w41694 <= not w41692 and w41693;
w41695 <= not w41680 and not w41694;
w41696 <= not w14042 and not w41695;
w41697 <= w35996 and not w41293;
w41698 <= pi0200 and not w40736;
w41699 <= not w41697 and not w41698;
w41700 <= w14042 and not w41699;
w41701 <= pi0230 and not w41696;
w41702 <= not w41700 and w41701;
w41703 <= not w41690 and not w41702;
w41704 <= not pi0278 and not w38426;
w41705 <= not pi0976 and w38426;
w41706 <= not pi1091 and not w41704;
w41707 <= not w41705 and w41706;
w41708 <= pi0199 and not w41707;
w41709 <= pi1091 and not pi1132;
w41710 <= pi0976 and w38448;
w41711 <= pi0278 and not w38448;
w41712 <= not pi1091 and not w41710;
w41713 <= not w41711 and w41712;
w41714 <= not w41709 and not w41713;
w41715 <= not pi0199 and not w41714;
w41716 <= not w41708 and not w41715;
w41717 <= not pi0200 and not w41716;
w41718 <= pi1091 and not pi1133;
w41719 <= not w41713 and not w41718;
w41720 <= not pi0199 and not w41719;
w41721 <= not w41708 and not w41720;
w41722 <= pi0200 and not w41721;
w41723 <= not pi0299 and not w41722;
w41724 <= not w41717 and w41723;
w41725 <= pi0219 and not w41707;
w41726 <= pi0211 and not pi1133;
w41727 <= not pi0211 and not pi1132;
w41728 <= not w41726 and not w41727;
w41729 <= pi1091 and not w41728;
w41730 <= not w41713 and not w41729;
w41731 <= not pi0219 and not w41730;
w41732 <= not w41725 and not w41731;
w41733 <= pi0299 and w41732;
w41734 <= not w41724 and not w41733;
w41735 <= w4989 and not w41734;
w41736 <= not w4989 and w41732;
w41737 <= not pi0230 and not w41736;
w41738 <= not w41735 and w41737;
w41739 <= w36937 and w41728;
w41740 <= not pi0199 and pi1132;
w41741 <= not pi0200 and not w41740;
w41742 <= not pi0199 and pi1133;
w41743 <= pi0200 and not w41742;
w41744 <= not pi0299 and not w41743;
w41745 <= not w41741 and w41744;
w41746 <= w36071 and w41728;
w41747 <= not w41745 and not w41746;
w41748 <= w4989 and not w41747;
w41749 <= pi0230 and not w41739;
w41750 <= not w41748 and w41749;
w41751 <= not w41738 and not w41750;
w41752 <= not pi1134 and not w41751;
w41753 <= w8372 and not w41740;
w41754 <= w41744 and not w41753;
w41755 <= not w40190 and not w41746;
w41756 <= not w41754 and w41755;
w41757 <= w4989 and not w41756;
w41758 <= not pi0219 and not w41728;
w41759 <= not w37644 and not w41758;
w41760 <= pi0230 and not w41757;
w41761 <= not w41759 and w41760;
w41762 <= not w38494 and w41717;
w41763 <= w41723 and not w41762;
w41764 <= w10625 and w40018;
w41765 <= not w41733 and not w41764;
w41766 <= not w41763 and w41765;
w41767 <= w4989 and not w41766;
w41768 <= not w41487 and w41737;
w41769 <= not w41767 and w41768;
w41770 <= not w41761 and not w41769;
w41771 <= pi1134 and not w41770;
w41772 <= not w41752 and not w41771;
w41773 <= not pi0279 and not w38426;
w41774 <= not pi0958 and w38426;
w41775 <= not pi1091 and not w41773;
w41776 <= not w41774 and w41775;
w41777 <= pi1135 and w41251;
w41778 <= not w41776 and not w41777;
w41779 <= pi0199 and not w41778;
w41780 <= pi0958 and w38448;
w41781 <= pi0279 and not w38448;
w41782 <= not pi1091 and not w41780;
w41783 <= not w41781 and w41782;
w41784 <= not pi1133 and w41251;
w41785 <= not pi0199 and not w41784;
w41786 <= not w41783 and w41785;
w41787 <= not w41779 and not w41786;
w41788 <= w14042 and not w41787;
w41789 <= not w38514 and w41788;
w41790 <= not w39987 and not w41718;
w41791 <= not w41783 and w41790;
w41792 <= not pi0219 and not w41791;
w41793 <= pi1135 and w40018;
w41794 <= pi0219 and not w41793;
w41795 <= not w41776 and w41794;
w41796 <= not w14042 and not w41795;
w41797 <= not w41792 and w41796;
w41798 <= not pi0230 and not w41797;
w41799 <= not w41789 and w41798;
w41800 <= pi1135 and w36082;
w41801 <= not pi0211 and not pi1133;
w41802 <= not pi0219 and not w41801;
w41803 <= not pi0211 and w41802;
w41804 <= not w41800 and not w41803;
w41805 <= not w4989 and not w41804;
w41806 <= pi0199 and pi1135;
w41807 <= not w41742 and not w41806;
w41808 <= w36131 and not w41807;
w41809 <= pi0299 and not w41804;
w41810 <= not w41808 and not w41809;
w41811 <= w4989 and not w41810;
w41812 <= pi0230 and not w41805;
w41813 <= not w41811 and w41812;
w41814 <= not w41799 and not w41813;
w41815 <= not pi1134 and not w41814;
w41816 <= not pi1133 and w8372;
w41817 <= not pi0200 and pi1135;
w41818 <= pi0199 and not w41817;
w41819 <= not w41816 and not w41818;
w41820 <= w14042 and not w41819;
w41821 <= not w41800 and not w41802;
w41822 <= not w14042 and w41821;
w41823 <= not w41820 and not w41822;
w41824 <= pi0230 and not w41823;
w41825 <= pi1091 and not w41801;
w41826 <= w37704 and w41825;
w41827 <= not w41788 and not w41826;
w41828 <= w41798 and w41827;
w41829 <= not w41824 and not w41828;
w41830 <= pi1134 and not w41829;
w41831 <= not w41815 and not w41830;
w41832 <= not pi0211 and pi1135;
w41833 <= pi0211 and pi1136;
w41834 <= not w41832 and not w41833;
w41835 <= pi1091 and w41834;
w41836 <= not pi0280 and not w38448;
w41837 <= pi0914 and w38448;
w41838 <= not pi1091 and not w41836;
w41839 <= not w41837 and w41838;
w41840 <= not w41835 and not w41839;
w41841 <= not pi0219 and not w41840;
w41842 <= not pi0211 and pi1137;
w41843 <= pi0219 and not w41842;
w41844 <= not w40720 and not w41843;
w41845 <= not pi0914 and w38426;
w41846 <= pi0280 and not w38426;
w41847 <= not pi1091 and not w41845;
w41848 <= not w41846 and w41847;
w41849 <= not w41844 and not w41848;
w41850 <= not w41841 and not w41849;
w41851 <= not w14042 and not w41850;
w41852 <= pi1137 and w41251;
w41853 <= not w41848 and not w41852;
w41854 <= pi0199 and not w41853;
w41855 <= pi0200 and pi1136;
w41856 <= pi1091 and not w41817;
w41857 <= not w41855 and w41856;
w41858 <= not pi0199 and not w41857;
w41859 <= not w41839 and w41858;
w41860 <= w14042 and not w41854;
w41861 <= not w41859 and w41860;
w41862 <= not w41851 and not w41861;
w41863 <= not pi0230 and not w41862;
w41864 <= pi0200 and not w41218;
w41865 <= pi0199 and pi1137;
w41866 <= not pi0200 and not w40791;
w41867 <= not w41865 and w41866;
w41868 <= not w41864 and not w41867;
w41869 <= w14042 and w41868;
w41870 <= not pi0219 and w41834;
w41871 <= not w41843 and not w41870;
w41872 <= not w14042 and w41871;
w41873 <= pi0230 and not w41869;
w41874 <= not w41872 and w41873;
w41875 <= not w41863 and not w41874;
w41876 <= not pi0199 and pi1138;
w41877 <= pi0200 and not w41876;
w41878 <= pi0199 and pi1139;
w41879 <= not pi0200 and not w41215;
w41880 <= not w41878 and w41879;
w41881 <= not w41877 and not w41880;
w41882 <= w14042 and not w41881;
w41883 <= pi0219 and w41275;
w41884 <= pi0211 and pi1138;
w41885 <= not w41842 and not w41884;
w41886 <= not pi0219 and not w41885;
w41887 <= not w41883 and not w41886;
w41888 <= not w14042 and w41887;
w41889 <= not w41882 and not w41888;
w41890 <= pi0230 and not w41889;
w41891 <= not pi0830 and w38448;
w41892 <= pi0281 and not w38448;
w41893 <= not pi1091 and not w41891;
w41894 <= not w41892 and w41893;
w41895 <= pi1091 and not w41885;
w41896 <= w37704 and not w41895;
w41897 <= pi1138 and w38514;
w41898 <= not w41852 and not w41897;
w41899 <= w41063 and w41898;
w41900 <= not w41896 and not w41899;
w41901 <= not w41894 and not w41900;
w41902 <= not pi0830 and w38426;
w41903 <= pi0281 and not w38426;
w41904 <= not pi1091 and not w41902;
w41905 <= not w41903 and w41904;
w41906 <= pi1139 and w40018;
w41907 <= w41249 and not w41906;
w41908 <= pi0199 and not w41282;
w41909 <= w14042 and w41908;
w41910 <= not w41907 and not w41909;
w41911 <= not w41905 and not w41910;
w41912 <= not w41901 and not w41911;
w41913 <= not pi0230 and not w41912;
w41914 <= not w41890 and not w41913;
w41915 <= pi0200 and not w41296;
w41916 <= pi0199 and pi1140;
w41917 <= not pi0200 and not w41876;
w41918 <= not w41916 and w41917;
w41919 <= not w41915 and not w41918;
w41920 <= w14042 and not w41919;
w41921 <= pi0219 and w41692;
w41922 <= pi0211 and pi1139;
w41923 <= not w41223 and not w41922;
w41924 <= not pi0219 and not w41923;
w41925 <= not w41921 and not w41924;
w41926 <= not w14042 and w41925;
w41927 <= not w41920 and not w41926;
w41928 <= pi0230 and not w41927;
w41929 <= not pi0836 and w38448;
w41930 <= pi0282 and not w38448;
w41931 <= not pi1091 and not w41929;
w41932 <= not w41930 and w41931;
w41933 <= pi1091 and not w41923;
w41934 <= w37704 and not w41933;
w41935 <= pi1139 and w38514;
w41936 <= not w41252 and not w41935;
w41937 <= w41063 and w41936;
w41938 <= not w41934 and not w41937;
w41939 <= not w41932 and not w41938;
w41940 <= not pi0836 and w38426;
w41941 <= pi0282 and not w38426;
w41942 <= not pi1091 and not w41940;
w41943 <= not w41941 and w41942;
w41944 <= pi1140 and w40018;
w41945 <= w41249 and not w41944;
w41946 <= not pi0200 and w41280;
w41947 <= pi0199 and not w41946;
w41948 <= w14042 and w41947;
w41949 <= not w41945 and not w41948;
w41950 <= not w41943 and not w41949;
w41951 <= not w41939 and not w41950;
w41952 <= not pi0230 and not w41951;
w41953 <= not w41928 and not w41952;
w41954 <= pi1147 and not w41354;
w41955 <= pi1149 and not w39952;
w41956 <= not w41954 and not w41955;
w41957 <= not pi1148 and not w41956;
w41958 <= w41447 and not w41954;
w41959 <= pi1147 and not w41064;
w41960 <= not pi1149 and w41073;
w41961 <= not w41959 and w41960;
w41962 <= pi1148 and not w41958;
w41963 <= not w41961 and w41962;
w41964 <= pi0230 and not w41957;
w41965 <= not w41963 and w41964;
w41966 <= not pi1147 and w41200;
w41967 <= pi1147 and w41104;
w41968 <= pi1148 and not w41967;
w41969 <= not w41966 and w41968;
w41970 <= pi1147 and w41098;
w41971 <= not pi1147 and not w41196;
w41972 <= not pi1148 and not w41971;
w41973 <= not w41970 and w41972;
w41974 <= not pi1149 and not w41969;
w41975 <= not w41973 and w41974;
w41976 <= not pi1147 and w41192;
w41977 <= pi1147 and w41143;
w41978 <= pi1148 and not w41977;
w41979 <= not w41976 and w41978;
w41980 <= not pi1147 and w41186;
w41981 <= pi1147 and w41138;
w41982 <= not pi1148 and not w41980;
w41983 <= not w41981 and w41982;
w41984 <= pi1149 and not w41979;
w41985 <= not w41983 and w41984;
w41986 <= pi0283 and not w41975;
w41987 <= not w41985 and w41986;
w41988 <= not pi1147 and w41168;
w41989 <= pi1147 and w41149;
w41990 <= pi1149 and not w41988;
w41991 <= not w41989 and w41990;
w41992 <= not pi1147 and not w41125;
w41993 <= pi1147 and w41118;
w41994 <= not pi1149 and not w41992;
w41995 <= not w41993 and w41994;
w41996 <= not pi1148 and not w41995;
w41997 <= not w41991 and w41996;
w41998 <= not pi1147 and w41171;
w41999 <= pi1147 and w41156;
w42000 <= pi1149 and not w41999;
w42001 <= not w41998 and w42000;
w42002 <= pi1147 and w41126;
w42003 <= not pi1147 and not w41177;
w42004 <= not pi1149 and not w42002;
w42005 <= not w42003 and w42004;
w42006 <= pi1148 and not w42001;
w42007 <= not w42005 and w42006;
w42008 <= not pi0283 and not w41997;
w42009 <= not w42007 and w42008;
w42010 <= not pi0230 and not w41987;
w42011 <= not w42009 and w42010;
w42012 <= not w41965 and not w42011;
w42013 <= not pi0284 and not w40465;
w42014 <= pi1143 and w40465;
w42015 <= not w37706 and w42014;
w42016 <= not w42013 and not w42015;
w42017 <= w135 and not w7962;
w42018 <= not w4983 and w42017;
w42019 <= pi0286 and w42018;
w42020 <= pi0288 and pi0289;
w42021 <= w42019 and w42020;
w42022 <= pi0285 and w42021;
w42023 <= pi0285 and w42017;
w42024 <= not w42021 and not w42023;
w42025 <= w4989 and not w42022;
w42026 <= not w42024 and w42025;
w42027 <= w4989 and w42021;
w42028 <= not pi0286 and w4983;
w42029 <= not pi0288 and w42028;
w42030 <= not pi0289 and w42029;
w42031 <= pi0285 and not w42030;
w42032 <= not w42027 and w42031;
w42033 <= not w42026 and not w42032;
w42034 <= not pi0793 and not w42033;
w42035 <= not pi0288 and not w4987;
w42036 <= w4983 and w42035;
w42037 <= pi0286 and not w42036;
w42038 <= not pi0286 and w42036;
w42039 <= not w4989 and not w42037;
w42040 <= not w42038 and w42039;
w42041 <= w4983 and not w42017;
w42042 <= pi0286 and not w42041;
w42043 <= not w42017 and w42028;
w42044 <= not w42042 and not w42043;
w42045 <= w42035 and not w42044;
w42046 <= not pi0286 and not w42018;
w42047 <= pi0288 and not w42019;
w42048 <= not w42046 and w42047;
w42049 <= w4989 and not w42045;
w42050 <= not w42048 and w42049;
w42051 <= not pi0793 and not w42040;
w42052 <= not w42050 and w42051;
w42053 <= not pi0287 and pi0457;
w42054 <= not pi0332 and not w42053;
w42055 <= pi0288 and not w4983;
w42056 <= not w42036 and not w42055;
w42057 <= w4989 and w42017;
w42058 <= not w42056 and w42057;
w42059 <= w42056 and not w42057;
w42060 <= not pi0793 and not w42058;
w42061 <= not w42059 and w42060;
w42062 <= pi0289 and not w42029;
w42063 <= pi0285 and not pi0289;
w42064 <= w42029 and w42063;
w42065 <= not w4989 and not w42062;
w42066 <= not w42064 and w42065;
w42067 <= not pi0289 and w42047;
w42068 <= w42043 and w42063;
w42069 <= pi0289 and not w42043;
w42070 <= not pi0288 and not w42068;
w42071 <= not w42069 and w42070;
w42072 <= not w42021 and not w42067;
w42073 <= not w42071 and w42072;
w42074 <= w4989 and not w42073;
w42075 <= not pi0793 and not w42066;
w42076 <= not w42074 and w42075;
w42077 <= not pi0290 and pi0476;
w42078 <= not pi0476 and not pi1048;
w42079 <= not w42077 and not w42078;
w42080 <= not pi0291 and pi0476;
w42081 <= not pi0476 and not pi1049;
w42082 <= not w42080 and not w42081;
w42083 <= not pi0292 and pi0476;
w42084 <= not pi0476 and not pi1084;
w42085 <= not w42083 and not w42084;
w42086 <= not pi0293 and pi0476;
w42087 <= not pi0476 and not pi1059;
w42088 <= not w42086 and not w42087;
w42089 <= not pi0294 and pi0476;
w42090 <= not pi0476 and not pi1072;
w42091 <= not w42089 and not w42090;
w42092 <= not pi0295 and pi0476;
w42093 <= not pi0476 and not pi1053;
w42094 <= not w42092 and not w42093;
w42095 <= not pi0296 and pi0476;
w42096 <= not pi0476 and not pi1037;
w42097 <= not w42095 and not w42096;
w42098 <= not pi0297 and pi0476;
w42099 <= not pi0476 and not pi1044;
w42100 <= not w42098 and not w42099;
w42101 <= not pi0478 and pi1044;
w42102 <= pi0298 and pi0478;
w42103 <= not w42101 and not w42102;
w42104 <= pi0054 and w84;
w42105 <= not pi0054 and w10716;
w42106 <= w10974 and w42105;
w42107 <= not w42104 and not w42106;
w42108 <= w184 and w6443;
w42109 <= not w42107 and w42108;
w42110 <= not pi0039 and not w42109;
w42111 <= not w8826 and not w42110;
w42112 <= pi0057 and not pi0059;
w42113 <= w7631 and w42112;
w42114 <= not pi0312 and w42113;
w42115 <= pi0300 and not w42114;
w42116 <= not pi0300 and w42114;
w42117 <= not pi0055 and not w42116;
w42118 <= not w42115 and w42117;
w42119 <= not pi0301 and w42117;
w42120 <= not pi0055 and pi0301;
w42121 <= w42116 and w42120;
w42122 <= not w42119 and not w42121;
w42123 <= w3399 and w4989;
w42124 <= not pi0222 and not pi0223;
w42125 <= pi0937 and not w42124;
w42126 <= pi0273 and w914;
w42127 <= not w42125 and not w42126;
w42128 <= w42123 and w42127;
w42129 <= not w166 and w42128;
w42130 <= w1012 and not w14042;
w42131 <= not w42128 and not w42130;
w42132 <= pi0237 and not w42131;
w42133 <= w3343 and not w14042;
w42134 <= not w42123 and not w42133;
w42135 <= not pi1148 and w42134;
w42136 <= not pi0215 and w873;
w42137 <= not pi0273 and w42136;
w42138 <= pi0833 and w5133;
w42139 <= not pi0937 and w42138;
w42140 <= not w42137 and not w42139;
w42141 <= not w14042 and not w42140;
w42142 <= not w42129 and not w42141;
w42143 <= not w42132 and w42142;
w42144 <= not w42135 and w42143;
w42145 <= not pi0478 and pi1049;
w42146 <= pi0303 and pi0478;
w42147 <= not w42145 and not w42146;
w42148 <= not pi0478 and pi1048;
w42149 <= pi0304 and pi0478;
w42150 <= not w42148 and not w42149;
w42151 <= not pi0478 and pi1084;
w42152 <= pi0305 and pi0478;
w42153 <= not w42151 and not w42152;
w42154 <= not pi0478 and pi1059;
w42155 <= pi0306 and pi0478;
w42156 <= not w42154 and not w42155;
w42157 <= not pi0478 and pi1053;
w42158 <= pi0307 and pi0478;
w42159 <= not w42157 and not w42158;
w42160 <= not pi0478 and pi1037;
w42161 <= pi0308 and pi0478;
w42162 <= not w42160 and not w42161;
w42163 <= not pi0478 and pi1072;
w42164 <= pi0309 and pi0478;
w42165 <= not w42163 and not w42164;
w42166 <= pi1147 and w42134;
w42167 <= pi0222 and not pi0934;
w42168 <= not pi0271 and w914;
w42169 <= not w42167 and not w42168;
w42170 <= w42123 and w42169;
w42171 <= not w1011 and w42133;
w42172 <= pi0934 and not w89;
w42173 <= pi0271 and w873;
w42174 <= not w42172 and not w42173;
w42175 <= w42171 and not w42174;
w42176 <= not w42130 and not w42170;
w42177 <= not w42175 and w42176;
w42178 <= not w42166 and w42177;
w42179 <= not pi0233 and not w42178;
w42180 <= w167 and w14042;
w42181 <= w42123 and not w42169;
w42182 <= w42133 and w42174;
w42183 <= pi1147 and not w42180;
w42184 <= not w42181 and w42183;
w42185 <= not w42182 and w42184;
w42186 <= not w166 and w42123;
w42187 <= not w42171 and not w42186;
w42188 <= not pi1147 and not w42187;
w42189 <= not w42177 and w42188;
w42190 <= not w42185 and not w42189;
w42191 <= pi0233 and not w42190;
w42192 <= not w42179 and not w42191;
w42193 <= not pi0055 and not pi0311;
w42194 <= not w42121 and not w42193;
w42195 <= not pi0311 and w42121;
w42196 <= not w42194 and not w42195;
w42197 <= pi0312 and not w42113;
w42198 <= not w42114 and not w42197;
w42199 <= not pi0055 and not w42198;
w42200 <= not w7951 and not w11009;
w42201 <= w3841 and not w11016;
w42202 <= w7729 and not w42201;
w42203 <= not w42200 and w42202;
w42204 <= not pi0954 and not w42203;
w42205 <= pi0313 and pi0954;
w42206 <= not w42204 and not w42205;
w42207 <= w3886 and w6443;
w42208 <= w12003 and not w42207;
w42209 <= pi0039 and not w12860;
w42210 <= not pi0039 and not w12077;
w42211 <= w171 and not w42209;
w42212 <= not w42210 and w42211;
w42213 <= not w12896 and not w42212;
w42214 <= w97 and w7726;
w42215 <= not w42213 and w42214;
w42216 <= not w42208 and not w42215;
w42217 <= w11995 and w11996;
w42218 <= not w42216 and w42217;
w42219 <= not pi0340 and w42017;
w42220 <= w4989 and w42219;
w42221 <= pi0315 and not w42220;
w42222 <= pi1080 and w42220;
w42223 <= not w42221 and not w42222;
w42224 <= pi0316 and not w42220;
w42225 <= pi1047 and w42220;
w42226 <= not w42224 and not w42225;
w42227 <= not pi0330 and w42057;
w42228 <= pi0317 and not w42227;
w42229 <= pi1078 and w42227;
w42230 <= not w42228 and not w42229;
w42231 <= not pi0341 and w42017;
w42232 <= w4989 and w42231;
w42233 <= pi0318 and not w42232;
w42234 <= pi1074 and w42232;
w42235 <= not w42233 and not w42234;
w42236 <= pi0319 and not w42232;
w42237 <= pi1072 and w42232;
w42238 <= not w42236 and not w42237;
w42239 <= pi0320 and not w42220;
w42240 <= pi1048 and w42220;
w42241 <= not w42239 and not w42240;
w42242 <= pi0321 and not w42220;
w42243 <= pi1058 and w42220;
w42244 <= not w42242 and not w42243;
w42245 <= pi0322 and not w42220;
w42246 <= pi1051 and w42220;
w42247 <= not w42245 and not w42246;
w42248 <= pi0323 and not w42220;
w42249 <= pi1065 and w42220;
w42250 <= not w42248 and not w42249;
w42251 <= pi0324 and not w42232;
w42252 <= pi1086 and w42232;
w42253 <= not w42251 and not w42252;
w42254 <= pi0325 and not w42232;
w42255 <= pi1063 and w42232;
w42256 <= not w42254 and not w42255;
w42257 <= pi0326 and not w42232;
w42258 <= pi1057 and w42232;
w42259 <= not w42257 and not w42258;
w42260 <= pi0327 and not w42220;
w42261 <= pi1040 and w42220;
w42262 <= not w42260 and not w42261;
w42263 <= pi0328 and not w42232;
w42264 <= pi1058 and w42232;
w42265 <= not w42263 and not w42264;
w42266 <= pi0329 and not w42232;
w42267 <= pi1043 and w42232;
w42268 <= not w42266 and not w42267;
w42269 <= pi1092 and not w493;
w42270 <= not w4989 and w42269;
w42271 <= not pi0330 and w42270;
w42272 <= w4989 and w42269;
w42273 <= not pi0330 and not w42017;
w42274 <= not w42219 and not w42273;
w42275 <= w42272 and not w42274;
w42276 <= not w42271 and not w42275;
w42277 <= not pi0331 and w42270;
w42278 <= not pi0331 and not w42017;
w42279 <= not w42231 and not w42278;
w42280 <= w42272 and not w42279;
w42281 <= not w42277 and not w42280;
w42282 <= w8565 and w10729;
w42283 <= not w8565 and not w10665;
w42284 <= w5008 and not w42283;
w42285 <= not pi0070 and not w42284;
w42286 <= pi0332 and w6680;
w42287 <= not w42285 and w42286;
w42288 <= not w42282 and not w42287;
w42289 <= not pi0039 and not w42288;
w42290 <= pi0039 and w7931;
w42291 <= not pi0038 and not w42290;
w42292 <= not w42289 and w42291;
w42293 <= w35832 and not w42292;
w42294 <= pi0333 and not w42232;
w42295 <= pi1040 and w42232;
w42296 <= not w42294 and not w42295;
w42297 <= pi0334 and not w42232;
w42298 <= pi1065 and w42232;
w42299 <= not w42297 and not w42298;
w42300 <= pi0335 and not w42232;
w42301 <= pi1069 and w42232;
w42302 <= not w42300 and not w42301;
w42303 <= pi0336 and not w42227;
w42304 <= pi1070 and w42227;
w42305 <= not w42303 and not w42304;
w42306 <= pi0337 and not w42227;
w42307 <= pi1044 and w42227;
w42308 <= not w42306 and not w42307;
w42309 <= pi0338 and not w42227;
w42310 <= pi1072 and w42227;
w42311 <= not w42309 and not w42310;
w42312 <= pi0339 and not w42227;
w42313 <= pi1086 and w42227;
w42314 <= not w42312 and not w42313;
w42315 <= pi0340 and w42270;
w42316 <= not pi0340 and not w42017;
w42317 <= not pi0331 and w42017;
w42318 <= w42272 and not w42316;
w42319 <= not w42317 and w42318;
w42320 <= not w42315 and not w42319;
w42321 <= not pi0341 and not w42057;
w42322 <= not w42227 and not w42321;
w42323 <= w42269 and not w42322;
w42324 <= pi0342 and not w42220;
w42325 <= pi1049 and w42220;
w42326 <= not w42324 and not w42325;
w42327 <= pi0343 and not w42220;
w42328 <= pi1062 and w42220;
w42329 <= not w42327 and not w42328;
w42330 <= pi0344 and not w42220;
w42331 <= pi1069 and w42220;
w42332 <= not w42330 and not w42331;
w42333 <= pi0345 and not w42220;
w42334 <= pi1039 and w42220;
w42335 <= not w42333 and not w42334;
w42336 <= pi0346 and not w42220;
w42337 <= pi1067 and w42220;
w42338 <= not w42336 and not w42337;
w42339 <= pi0347 and not w42220;
w42340 <= pi1055 and w42220;
w42341 <= not w42339 and not w42340;
w42342 <= pi0348 and not w42220;
w42343 <= pi1087 and w42220;
w42344 <= not w42342 and not w42343;
w42345 <= pi0349 and not w42220;
w42346 <= pi1043 and w42220;
w42347 <= not w42345 and not w42346;
w42348 <= pi0350 and not w42220;
w42349 <= pi1035 and w42220;
w42350 <= not w42348 and not w42349;
w42351 <= pi0351 and not w42220;
w42352 <= pi1079 and w42220;
w42353 <= not w42351 and not w42352;
w42354 <= pi0352 and not w42220;
w42355 <= pi1078 and w42220;
w42356 <= not w42354 and not w42355;
w42357 <= pi0353 and not w42220;
w42358 <= pi1063 and w42220;
w42359 <= not w42357 and not w42358;
w42360 <= pi0354 and not w42220;
w42361 <= pi1045 and w42220;
w42362 <= not w42360 and not w42361;
w42363 <= pi0355 and not w42220;
w42364 <= pi1084 and w42220;
w42365 <= not w42363 and not w42364;
w42366 <= pi0356 and not w42220;
w42367 <= pi1081 and w42220;
w42368 <= not w42366 and not w42367;
w42369 <= pi0357 and not w42220;
w42370 <= pi1076 and w42220;
w42371 <= not w42369 and not w42370;
w42372 <= pi0358 and not w42220;
w42373 <= pi1071 and w42220;
w42374 <= not w42372 and not w42373;
w42375 <= pi0359 and not w42220;
w42376 <= pi1068 and w42220;
w42377 <= not w42375 and not w42376;
w42378 <= pi0360 and not w42220;
w42379 <= pi1042 and w42220;
w42380 <= not w42378 and not w42379;
w42381 <= pi0361 and not w42220;
w42382 <= pi1059 and w42220;
w42383 <= not w42381 and not w42382;
w42384 <= pi0362 and not w42220;
w42385 <= pi1070 and w42220;
w42386 <= not w42384 and not w42385;
w42387 <= pi0363 and not w42227;
w42388 <= pi1049 and w42227;
w42389 <= not w42387 and not w42388;
w42390 <= pi0364 and not w42227;
w42391 <= pi1062 and w42227;
w42392 <= not w42390 and not w42391;
w42393 <= pi0365 and not w42227;
w42394 <= pi1065 and w42227;
w42395 <= not w42393 and not w42394;
w42396 <= pi0366 and not w42227;
w42397 <= pi1069 and w42227;
w42398 <= not w42396 and not w42397;
w42399 <= pi0367 and not w42227;
w42400 <= pi1039 and w42227;
w42401 <= not w42399 and not w42400;
w42402 <= pi0368 and not w42227;
w42403 <= pi1067 and w42227;
w42404 <= not w42402 and not w42403;
w42405 <= pi0369 and not w42227;
w42406 <= pi1080 and w42227;
w42407 <= not w42405 and not w42406;
w42408 <= pi0370 and not w42227;
w42409 <= pi1055 and w42227;
w42410 <= not w42408 and not w42409;
w42411 <= pi0371 and not w42227;
w42412 <= pi1051 and w42227;
w42413 <= not w42411 and not w42412;
w42414 <= pi0372 and not w42227;
w42415 <= pi1048 and w42227;
w42416 <= not w42414 and not w42415;
w42417 <= pi0373 and not w42227;
w42418 <= pi1087 and w42227;
w42419 <= not w42417 and not w42418;
w42420 <= pi0374 and not w42227;
w42421 <= pi1035 and w42227;
w42422 <= not w42420 and not w42421;
w42423 <= pi0375 and not w42227;
w42424 <= pi1047 and w42227;
w42425 <= not w42423 and not w42424;
w42426 <= pi0376 and not w42227;
w42427 <= pi1079 and w42227;
w42428 <= not w42426 and not w42427;
w42429 <= pi0377 and not w42227;
w42430 <= pi1074 and w42227;
w42431 <= not w42429 and not w42430;
w42432 <= pi0378 and not w42227;
w42433 <= pi1063 and w42227;
w42434 <= not w42432 and not w42433;
w42435 <= pi0379 and not w42227;
w42436 <= pi1045 and w42227;
w42437 <= not w42435 and not w42436;
w42438 <= pi0380 and not w42227;
w42439 <= pi1084 and w42227;
w42440 <= not w42438 and not w42439;
w42441 <= pi0381 and not w42227;
w42442 <= pi1081 and w42227;
w42443 <= not w42441 and not w42442;
w42444 <= pi0382 and not w42227;
w42445 <= pi1076 and w42227;
w42446 <= not w42444 and not w42445;
w42447 <= pi0383 and not w42227;
w42448 <= pi1071 and w42227;
w42449 <= not w42447 and not w42448;
w42450 <= pi0384 and not w42227;
w42451 <= pi1068 and w42227;
w42452 <= not w42450 and not w42451;
w42453 <= pi0385 and not w42227;
w42454 <= pi1042 and w42227;
w42455 <= not w42453 and not w42454;
w42456 <= pi0386 and not w42227;
w42457 <= pi1059 and w42227;
w42458 <= not w42456 and not w42457;
w42459 <= pi0387 and not w42227;
w42460 <= pi1053 and w42227;
w42461 <= not w42459 and not w42460;
w42462 <= pi0388 and not w42227;
w42463 <= pi1037 and w42227;
w42464 <= not w42462 and not w42463;
w42465 <= pi0389 and not w42227;
w42466 <= pi1036 and w42227;
w42467 <= not w42465 and not w42466;
w42468 <= pi0390 and not w42232;
w42469 <= pi1049 and w42232;
w42470 <= not w42468 and not w42469;
w42471 <= pi0391 and not w42232;
w42472 <= pi1062 and w42232;
w42473 <= not w42471 and not w42472;
w42474 <= pi0392 and not w42232;
w42475 <= pi1039 and w42232;
w42476 <= not w42474 and not w42475;
w42477 <= pi0393 and not w42232;
w42478 <= pi1067 and w42232;
w42479 <= not w42477 and not w42478;
w42480 <= pi0394 and not w42232;
w42481 <= pi1080 and w42232;
w42482 <= not w42480 and not w42481;
w42483 <= pi0395 and not w42232;
w42484 <= pi1055 and w42232;
w42485 <= not w42483 and not w42484;
w42486 <= pi0396 and not w42232;
w42487 <= pi1051 and w42232;
w42488 <= not w42486 and not w42487;
w42489 <= pi0397 and not w42232;
w42490 <= pi1048 and w42232;
w42491 <= not w42489 and not w42490;
w42492 <= pi0398 and not w42232;
w42493 <= pi1087 and w42232;
w42494 <= not w42492 and not w42493;
w42495 <= pi0399 and not w42232;
w42496 <= pi1047 and w42232;
w42497 <= not w42495 and not w42496;
w42498 <= pi0400 and not w42232;
w42499 <= pi1035 and w42232;
w42500 <= not w42498 and not w42499;
w42501 <= pi0401 and not w42232;
w42502 <= pi1079 and w42232;
w42503 <= not w42501 and not w42502;
w42504 <= pi0402 and not w42232;
w42505 <= pi1078 and w42232;
w42506 <= not w42504 and not w42505;
w42507 <= pi0403 and not w42232;
w42508 <= pi1045 and w42232;
w42509 <= not w42507 and not w42508;
w42510 <= pi0404 and not w42232;
w42511 <= pi1084 and w42232;
w42512 <= not w42510 and not w42511;
w42513 <= pi0405 and not w42232;
w42514 <= pi1081 and w42232;
w42515 <= not w42513 and not w42514;
w42516 <= pi0406 and not w42232;
w42517 <= pi1076 and w42232;
w42518 <= not w42516 and not w42517;
w42519 <= pi0407 and not w42232;
w42520 <= pi1071 and w42232;
w42521 <= not w42519 and not w42520;
w42522 <= pi0408 and not w42232;
w42523 <= pi1068 and w42232;
w42524 <= not w42522 and not w42523;
w42525 <= pi0409 and not w42232;
w42526 <= pi1042 and w42232;
w42527 <= not w42525 and not w42526;
w42528 <= pi0410 and not w42232;
w42529 <= pi1059 and w42232;
w42530 <= not w42528 and not w42529;
w42531 <= pi0411 and not w42232;
w42532 <= pi1053 and w42232;
w42533 <= not w42531 and not w42532;
w42534 <= pi0412 and not w42232;
w42535 <= pi1037 and w42232;
w42536 <= not w42534 and not w42535;
w42537 <= pi0413 and not w42232;
w42538 <= pi1036 and w42232;
w42539 <= not w42537 and not w42538;
w42540 <= w4989 and w42317;
w42541 <= pi0414 and not w42540;
w42542 <= pi1049 and w42540;
w42543 <= not w42541 and not w42542;
w42544 <= pi0415 and not w42540;
w42545 <= pi1062 and w42540;
w42546 <= not w42544 and not w42545;
w42547 <= pi0416 and not w42540;
w42548 <= pi1069 and w42540;
w42549 <= not w42547 and not w42548;
w42550 <= pi0417 and not w42540;
w42551 <= pi1039 and w42540;
w42552 <= not w42550 and not w42551;
w42553 <= pi0418 and not w42540;
w42554 <= pi1067 and w42540;
w42555 <= not w42553 and not w42554;
w42556 <= pi0419 and not w42540;
w42557 <= pi1080 and w42540;
w42558 <= not w42556 and not w42557;
w42559 <= pi0420 and not w42540;
w42560 <= pi1055 and w42540;
w42561 <= not w42559 and not w42560;
w42562 <= pi0421 and not w42540;
w42563 <= pi1051 and w42540;
w42564 <= not w42562 and not w42563;
w42565 <= pi0422 and not w42540;
w42566 <= pi1048 and w42540;
w42567 <= not w42565 and not w42566;
w42568 <= pi0423 and not w42540;
w42569 <= pi1087 and w42540;
w42570 <= not w42568 and not w42569;
w42571 <= pi0424 and not w42540;
w42572 <= pi1047 and w42540;
w42573 <= not w42571 and not w42572;
w42574 <= pi0425 and not w42540;
w42575 <= pi1035 and w42540;
w42576 <= not w42574 and not w42575;
w42577 <= pi0426 and not w42540;
w42578 <= pi1079 and w42540;
w42579 <= not w42577 and not w42578;
w42580 <= pi0427 and not w42540;
w42581 <= pi1078 and w42540;
w42582 <= not w42580 and not w42581;
w42583 <= pi0428 and not w42540;
w42584 <= pi1045 and w42540;
w42585 <= not w42583 and not w42584;
w42586 <= pi0429 and not w42540;
w42587 <= pi1084 and w42540;
w42588 <= not w42586 and not w42587;
w42589 <= pi0430 and not w42540;
w42590 <= pi1076 and w42540;
w42591 <= not w42589 and not w42590;
w42592 <= pi0431 and not w42540;
w42593 <= pi1071 and w42540;
w42594 <= not w42592 and not w42593;
w42595 <= pi0432 and not w42540;
w42596 <= pi1068 and w42540;
w42597 <= not w42595 and not w42596;
w42598 <= pi0433 and not w42540;
w42599 <= pi1042 and w42540;
w42600 <= not w42598 and not w42599;
w42601 <= pi0434 and not w42540;
w42602 <= pi1059 and w42540;
w42603 <= not w42601 and not w42602;
w42604 <= pi0435 and not w42540;
w42605 <= pi1053 and w42540;
w42606 <= not w42604 and not w42605;
w42607 <= pi0436 and not w42540;
w42608 <= pi1037 and w42540;
w42609 <= not w42607 and not w42608;
w42610 <= pi0437 and not w42540;
w42611 <= pi1070 and w42540;
w42612 <= not w42610 and not w42611;
w42613 <= pi0438 and not w42540;
w42614 <= pi1036 and w42540;
w42615 <= not w42613 and not w42614;
w42616 <= pi0439 and not w42227;
w42617 <= pi1057 and w42227;
w42618 <= not w42616 and not w42617;
w42619 <= pi0440 and not w42227;
w42620 <= pi1043 and w42227;
w42621 <= not w42619 and not w42620;
w42622 <= pi0441 and not w42220;
w42623 <= pi1044 and w42220;
w42624 <= not w42622 and not w42623;
w42625 <= pi0442 and not w42227;
w42626 <= pi1058 and w42227;
w42627 <= not w42625 and not w42626;
w42628 <= pi0443 and not w42540;
w42629 <= pi1044 and w42540;
w42630 <= not w42628 and not w42629;
w42631 <= pi0444 and not w42540;
w42632 <= pi1072 and w42540;
w42633 <= not w42631 and not w42632;
w42634 <= pi0445 and not w42540;
w42635 <= pi1081 and w42540;
w42636 <= not w42634 and not w42635;
w42637 <= pi0446 and not w42540;
w42638 <= pi1086 and w42540;
w42639 <= not w42637 and not w42638;
w42640 <= pi0447 and not w42227;
w42641 <= pi1040 and w42227;
w42642 <= not w42640 and not w42641;
w42643 <= pi0448 and not w42540;
w42644 <= pi1074 and w42540;
w42645 <= not w42643 and not w42644;
w42646 <= pi0449 and not w42540;
w42647 <= pi1057 and w42540;
w42648 <= not w42646 and not w42647;
w42649 <= pi0450 and not w42220;
w42650 <= pi1036 and w42220;
w42651 <= not w42649 and not w42650;
w42652 <= pi0451 and not w42540;
w42653 <= pi1063 and w42540;
w42654 <= not w42652 and not w42653;
w42655 <= pi0452 and not w42220;
w42656 <= pi1053 and w42220;
w42657 <= not w42655 and not w42656;
w42658 <= pi0453 and not w42540;
w42659 <= pi1040 and w42540;
w42660 <= not w42658 and not w42659;
w42661 <= pi0454 and not w42540;
w42662 <= pi1043 and w42540;
w42663 <= not w42661 and not w42662;
w42664 <= pi0455 and not w42220;
w42665 <= pi1037 and w42220;
w42666 <= not w42664 and not w42665;
w42667 <= pi0456 and not w42232;
w42668 <= pi1044 and w42232;
w42669 <= not w42667 and not w42668;
w42670 <= pi0594 and pi0600;
w42671 <= pi0597 and w42670;
w42672 <= pi0601 and w42671;
w42673 <= not pi0804 and not pi0810;
w42674 <= not pi0595 and w42673;
w42675 <= not pi0599 and pi0810;
w42676 <= pi0596 and not w42675;
w42677 <= pi0804 and not w42676;
w42678 <= pi0595 and pi0815;
w42679 <= not w42677 and w42678;
w42680 <= not w42674 and not w42679;
w42681 <= w42672 and not w42680;
w42682 <= pi0600 and not pi0810;
w42683 <= pi0804 and not w42682;
w42684 <= not pi0601 and not w42673;
w42685 <= not pi0815 and not w42683;
w42686 <= not w42684 and w42685;
w42687 <= not w42681 and not w42686;
w42688 <= pi0605 and not w42687;
w42689 <= pi0990 and w42670;
w42690 <= not pi0815 and w42683;
w42691 <= w42689 and w42690;
w42692 <= not w42688 and not w42691;
w42693 <= pi0821 and not w42692;
w42694 <= pi0458 and not w42220;
w42695 <= pi1072 and w42220;
w42696 <= not w42694 and not w42695;
w42697 <= pi0459 and not w42540;
w42698 <= pi1058 and w42540;
w42699 <= not w42697 and not w42698;
w42700 <= pi0460 and not w42220;
w42701 <= pi1086 and w42220;
w42702 <= not w42700 and not w42701;
w42703 <= pi0461 and not w42220;
w42704 <= pi1057 and w42220;
w42705 <= not w42703 and not w42704;
w42706 <= pi0462 and not w42220;
w42707 <= pi1074 and w42220;
w42708 <= not w42706 and not w42707;
w42709 <= pi0463 and not w42232;
w42710 <= pi1070 and w42232;
w42711 <= not w42709 and not w42710;
w42712 <= pi0464 and not w42540;
w42713 <= pi1065 and w42540;
w42714 <= not w42712 and not w42713;
w42715 <= not pi0299 and w42124;
w42716 <= not w8986 and not w42715;
w42717 <= not w8959 and not w8962;
w42718 <= not pi0243 and not w42717;
w42719 <= not pi0243 and pi1157;
w42720 <= not w42716 and not w42719;
w42721 <= not w42718 and w42720;
w42722 <= not w1034 and not w8987;
w42723 <= pi0926 and w42719;
w42724 <= not w42722 and w42723;
w42725 <= not w3399 and not w3417;
w42726 <= pi0926 and not w42725;
w42727 <= pi1157 and w42725;
w42728 <= not w42718 and not w42726;
w42729 <= not w42727 and w42728;
w42730 <= not w42721 and not w42724;
w42731 <= not w42729 and w42730;
w42732 <= w4989 and not w42731;
w42733 <= not pi0243 and w42136;
w42734 <= pi0926 and w42138;
w42735 <= pi1157 and not w3343;
w42736 <= not w4989 and not w42733;
w42737 <= not w42734 and not w42735;
w42738 <= w42736 and w42737;
w42739 <= not w42732 and not w42738;
w42740 <= not w4989 and not w42136;
w42741 <= w4989 and w42717;
w42742 <= not w42740 and not w42741;
w42743 <= not pi0943 and not w42742;
w42744 <= not w42134 and w42743;
w42745 <= pi0943 and w42187;
w42746 <= not w42743 and not w42745;
w42747 <= not pi1151 and not w42746;
w42748 <= w4989 and not w42716;
w42749 <= w89 and not w4989;
w42750 <= not w42748 and not w42749;
w42751 <= not pi0275 and not w42750;
w42752 <= not w42130 and not w42180;
w42753 <= pi0943 and pi1151;
w42754 <= not w42752 and w42753;
w42755 <= not w42744 and not w42751;
w42756 <= not w42754 and w42755;
w42757 <= not w42747 and w42756;
w42758 <= pi0040 and not pi0287;
w42759 <= w39909 and w42758;
w42760 <= not w35951 and w42759;
w42761 <= not w7728 and not w42760;
w42762 <= not pi0102 and not w10944;
w42763 <= w6460 and w7725;
w42764 <= w14410 and w42763;
w42765 <= not w42762 and w42764;
w42766 <= w14408 and w42765;
w42767 <= w42759 and not w42766;
w42768 <= not w42759 and w42766;
w42769 <= not w42767 and not w42768;
w42770 <= w5053 and not w42769;
w42771 <= not w3840 and not w42769;
w42772 <= w3840 and w42766;
w42773 <= not w42771 and not w42772;
w42774 <= not w5053 and not w42773;
w42775 <= pi1091 and not w42770;
w42776 <= not w42774 and w42775;
w42777 <= not pi1093 and not w42773;
w42778 <= not w4980 and not w42769;
w42779 <= w4980 and w42766;
w42780 <= not w42778 and not w42779;
w42781 <= pi1093 and not w42780;
w42782 <= not pi1091 and not w42777;
w42783 <= not w42781 and w42782;
w42784 <= not w42776 and not w42783;
w42785 <= w173 and w42207;
w42786 <= not w42784 and w42785;
w42787 <= not w42761 and not w42786;
w42788 <= w7763 and w8900;
w42789 <= pi0038 and not pi0039;
w42790 <= w7760 and w42789;
w42791 <= w6525 and w42790;
w42792 <= pi0468 and not w42791;
w42793 <= not w42788 and not w42792;
w42794 <= not pi0263 and not w42717;
w42795 <= not pi0263 and pi1156;
w42796 <= not w42716 and not w42795;
w42797 <= not w42794 and w42796;
w42798 <= pi0942 and w42795;
w42799 <= not w42722 and w42798;
w42800 <= pi0942 and not w42725;
w42801 <= pi1156 and w42725;
w42802 <= not w42794 and not w42800;
w42803 <= not w42801 and w42802;
w42804 <= not w42797 and not w42799;
w42805 <= not w42803 and w42804;
w42806 <= w4989 and not w42805;
w42807 <= pi1156 and not w3343;
w42808 <= pi0942 and w42138;
w42809 <= not pi0263 and w42136;
w42810 <= not w4989 and not w42809;
w42811 <= not w42807 and not w42808;
w42812 <= w42810 and w42811;
w42813 <= not w42806 and not w42812;
w42814 <= pi0267 and not w42717;
w42815 <= pi0267 and pi1155;
w42816 <= not w42716 and not w42815;
w42817 <= not w42814 and w42816;
w42818 <= pi0925 and w42815;
w42819 <= not w42722 and w42818;
w42820 <= pi0925 and not w42725;
w42821 <= pi1155 and w42725;
w42822 <= not w42814 and not w42820;
w42823 <= not w42821 and w42822;
w42824 <= not w42817 and not w42819;
w42825 <= not w42823 and w42824;
w42826 <= w4989 and not w42825;
w42827 <= pi1155 and not w3343;
w42828 <= pi0925 and w42138;
w42829 <= pi0267 and w42136;
w42830 <= not w4989 and not w42829;
w42831 <= not w42827 and not w42828;
w42832 <= w42830 and w42831;
w42833 <= not w42826 and not w42832;
w42834 <= pi0253 and not w42717;
w42835 <= pi0253 and pi1153;
w42836 <= not w42716 and not w42835;
w42837 <= not w42834 and w42836;
w42838 <= pi0941 and w42835;
w42839 <= not w42722 and w42838;
w42840 <= pi0941 and not w42725;
w42841 <= pi1153 and w42725;
w42842 <= not w42834 and not w42840;
w42843 <= not w42841 and w42842;
w42844 <= not w42837 and not w42839;
w42845 <= not w42843 and w42844;
w42846 <= w4989 and not w42845;
w42847 <= pi1153 and not w3343;
w42848 <= pi0941 and w42138;
w42849 <= pi0253 and w42136;
w42850 <= not w4989 and not w42849;
w42851 <= not w42847 and not w42848;
w42852 <= w42850 and w42851;
w42853 <= not w42846 and not w42852;
w42854 <= pi0254 and not w42717;
w42855 <= pi0254 and pi1154;
w42856 <= not w42716 and not w42855;
w42857 <= not w42854 and w42856;
w42858 <= pi0923 and w42855;
w42859 <= not w42722 and w42858;
w42860 <= pi0923 and not w42725;
w42861 <= pi1154 and w42725;
w42862 <= not w42854 and not w42860;
w42863 <= not w42861 and w42862;
w42864 <= not w42857 and not w42859;
w42865 <= not w42863 and w42864;
w42866 <= w4989 and not w42865;
w42867 <= pi1154 and not w3343;
w42868 <= pi0923 and w42138;
w42869 <= pi0254 and w42136;
w42870 <= not w4989 and not w42869;
w42871 <= not w42867 and not w42868;
w42872 <= w42870 and w42871;
w42873 <= not w42866 and not w42872;
w42874 <= not pi0922 and not w42742;
w42875 <= not w42134 and w42874;
w42876 <= pi0922 and w42187;
w42877 <= not w42874 and not w42876;
w42878 <= not pi1152 and not w42877;
w42879 <= not pi0268 and not w42750;
w42880 <= pi0922 and pi1152;
w42881 <= not w42752 and w42880;
w42882 <= not w42875 and not w42879;
w42883 <= not w42881 and w42882;
w42884 <= not w42878 and w42883;
w42885 <= not pi0931 and not w42742;
w42886 <= not w42134 and w42885;
w42887 <= pi0931 and w42187;
w42888 <= not w42885 and not w42887;
w42889 <= not pi1150 and not w42888;
w42890 <= not pi0272 and not w42750;
w42891 <= pi0931 and pi1150;
w42892 <= not w42752 and w42891;
w42893 <= not w42886 and not w42890;
w42894 <= not w42892 and w42893;
w42895 <= not w42889 and w42894;
w42896 <= not pi0936 and not w42742;
w42897 <= not w42134 and w42896;
w42898 <= pi0936 and w42187;
w42899 <= not w42896 and not w42898;
w42900 <= not pi1149 and not w42899;
w42901 <= not pi0283 and not w42750;
w42902 <= pi0936 and pi1149;
w42903 <= not w42752 and w42902;
w42904 <= not w42897 and not w42901;
w42905 <= not w42903 and w42904;
w42906 <= not w42900 and w42905;
w42907 <= pi0071 and w41072;
w42908 <= pi0071 and not w9011;
w42909 <= w9011 and w10615;
w42910 <= w7713 and not w9011;
w42911 <= w7710 and w42910;
w42912 <= not w42909 and not w42911;
w42913 <= w135 and w7725;
w42914 <= not w42912 and w42913;
w42915 <= w10613 and w42914;
w42916 <= not w42908 and not w42915;
w42917 <= w4989 and not w42916;
w42918 <= not w42907 and not w42917;
w42919 <= pi0071 and not w41354;
w42920 <= pi0481 and not w32338;
w42921 <= pi0248 and w32338;
w42922 <= not w42920 and not w42921;
w42923 <= pi0482 and not w32354;
w42924 <= pi0249 and w32354;
w42925 <= not w42923 and not w42924;
w42926 <= pi0483 and not w32478;
w42927 <= pi0242 and w32478;
w42928 <= not w42926 and not w42927;
w42929 <= pi0484 and not w32478;
w42930 <= pi0249 and w32478;
w42931 <= not w42929 and not w42930;
w42932 <= pi0485 and not w33674;
w42933 <= pi0234 and w33674;
w42934 <= not w42932 and not w42933;
w42935 <= pi0486 and not w33674;
w42936 <= pi0244 and w33674;
w42937 <= not w42935 and not w42936;
w42938 <= pi0487 and not w32338;
w42939 <= pi0246 and w32338;
w42940 <= not w42938 and not w42939;
w42941 <= pi0488 and not w32338;
w42942 <= not pi0239 and w32338;
w42943 <= not w42941 and not w42942;
w42944 <= pi0489 and not w33674;
w42945 <= pi0242 and w33674;
w42946 <= not w42944 and not w42945;
w42947 <= pi0490 and not w32478;
w42948 <= pi0241 and w32478;
w42949 <= not w42947 and not w42948;
w42950 <= pi0491 and not w32478;
w42951 <= pi0238 and w32478;
w42952 <= not w42950 and not w42951;
w42953 <= pi0492 and not w32478;
w42954 <= pi0240 and w32478;
w42955 <= not w42953 and not w42954;
w42956 <= pi0493 and not w32478;
w42957 <= pi0244 and w32478;
w42958 <= not w42956 and not w42957;
w42959 <= pi0494 and not w32478;
w42960 <= not pi0239 and w32478;
w42961 <= not w42959 and not w42960;
w42962 <= pi0495 and not w32478;
w42963 <= pi0235 and w32478;
w42964 <= not w42962 and not w42963;
w42965 <= pi0496 and not w32470;
w42966 <= pi0249 and w32470;
w42967 <= not w42965 and not w42966;
w42968 <= pi0497 and not w32470;
w42969 <= not pi0239 and w32470;
w42970 <= not w42968 and not w42969;
w42971 <= pi0498 and not w32354;
w42972 <= pi0238 and w32354;
w42973 <= not w42971 and not w42972;
w42974 <= pi0499 and not w32470;
w42975 <= pi0246 and w32470;
w42976 <= not w42974 and not w42975;
w42977 <= pi0500 and not w32470;
w42978 <= pi0241 and w32470;
w42979 <= not w42977 and not w42978;
w42980 <= pi0501 and not w32470;
w42981 <= pi0248 and w32470;
w42982 <= not w42980 and not w42981;
w42983 <= pi0502 and not w32470;
w42984 <= pi0247 and w32470;
w42985 <= not w42983 and not w42984;
w42986 <= pi0503 and not w32470;
w42987 <= pi0245 and w32470;
w42988 <= not w42986 and not w42987;
w42989 <= pi0504 and not w32463;
w42990 <= pi0242 and w32463;
w42991 <= not w42989 and not w42990;
w42992 <= not w3889 and w14042;
w42993 <= not w32458 and not w42992;
w42994 <= not pi0234 and w42993;
w42995 <= w32470 and w42994;
w42996 <= pi0505 and not w42995;
w42997 <= pi0234 and w32462;
w42998 <= not pi0505 and w32341;
w42999 <= w42997 and w42998;
w43000 <= not w42996 and not w42999;
w43001 <= pi0506 and not w32463;
w43002 <= pi0241 and w32463;
w43003 <= not w43001 and not w43002;
w43004 <= pi0507 and not w32463;
w43005 <= pi0238 and w32463;
w43006 <= not w43004 and not w43005;
w43007 <= pi0508 and not w32463;
w43008 <= pi0247 and w32463;
w43009 <= not w43007 and not w43008;
w43010 <= pi0509 and not w32463;
w43011 <= pi0245 and w32463;
w43012 <= not w43010 and not w43011;
w43013 <= pi0510 and not w32338;
w43014 <= pi0242 and w32338;
w43015 <= not w43013 and not w43014;
w43016 <= w4147 and w4989;
w43017 <= not w32332 and not w43016;
w43018 <= not pi0234 and w43017;
w43019 <= w32338 and not w43018;
w43020 <= pi0511 and not w32338;
w43021 <= not w43019 and not w43020;
w43022 <= pi0512 and not w32338;
w43023 <= pi0235 and w32338;
w43024 <= not w43022 and not w43023;
w43025 <= pi0513 and not w32338;
w43026 <= pi0244 and w32338;
w43027 <= not w43025 and not w43026;
w43028 <= pi0514 and not w32338;
w43029 <= pi0245 and w32338;
w43030 <= not w43028 and not w43029;
w43031 <= pi0515 and not w32338;
w43032 <= pi0240 and w32338;
w43033 <= not w43031 and not w43032;
w43034 <= pi0516 and not w32338;
w43035 <= pi0247 and w32338;
w43036 <= not w43034 and not w43035;
w43037 <= pi0517 and not w32338;
w43038 <= pi0238 and w32338;
w43039 <= not w43037 and not w43038;
w43040 <= w32346 and w43018;
w43041 <= pi0518 and not w43040;
w43042 <= pi0234 and w32337;
w43043 <= not pi0518 and w32341;
w43044 <= w43042 and w43043;
w43045 <= not w43041 and not w43044;
w43046 <= pi0519 and not w32346;
w43047 <= not pi0239 and w32346;
w43048 <= not w43046 and not w43047;
w43049 <= pi0520 and not w32346;
w43050 <= pi0246 and w32346;
w43051 <= not w43049 and not w43050;
w43052 <= pi0521 and not w32346;
w43053 <= pi0248 and w32346;
w43054 <= not w43052 and not w43053;
w43055 <= pi0522 and not w32346;
w43056 <= pi0238 and w32346;
w43057 <= not w43055 and not w43056;
w43058 <= w33702 and w43018;
w43059 <= pi0523 and not w43058;
w43060 <= not pi0523 and w32473;
w43061 <= w43042 and w43060;
w43062 <= not w43059 and not w43061;
w43063 <= pi0524 and not w33702;
w43064 <= not pi0239 and w33702;
w43065 <= not w43063 and not w43064;
w43066 <= pi0525 and not w33702;
w43067 <= pi0245 and w33702;
w43068 <= not w43066 and not w43067;
w43069 <= pi0526 and not w33702;
w43070 <= pi0246 and w33702;
w43071 <= not w43069 and not w43070;
w43072 <= pi0527 and not w33702;
w43073 <= pi0247 and w33702;
w43074 <= not w43072 and not w43073;
w43075 <= pi0528 and not w33702;
w43076 <= pi0249 and w33702;
w43077 <= not w43075 and not w43076;
w43078 <= pi0529 and not w33702;
w43079 <= pi0238 and w33702;
w43080 <= not w43078 and not w43079;
w43081 <= pi0530 and not w33702;
w43082 <= pi0240 and w33702;
w43083 <= not w43081 and not w43082;
w43084 <= pi0531 and not w32354;
w43085 <= pi0235 and w32354;
w43086 <= not w43084 and not w43085;
w43087 <= pi0532 and not w32354;
w43088 <= pi0247 and w32354;
w43089 <= not w43087 and not w43088;
w43090 <= pi0533 and not w32463;
w43091 <= pi0235 and w32463;
w43092 <= not w43090 and not w43091;
w43093 <= pi0534 and not w32463;
w43094 <= not pi0239 and w32463;
w43095 <= not w43093 and not w43094;
w43096 <= pi0535 and not w32463;
w43097 <= pi0240 and w32463;
w43098 <= not w43096 and not w43097;
w43099 <= pi0536 and not w32463;
w43100 <= pi0246 and w32463;
w43101 <= not w43099 and not w43100;
w43102 <= pi0537 and not w32463;
w43103 <= pi0248 and w32463;
w43104 <= not w43102 and not w43103;
w43105 <= pi0538 and not w32463;
w43106 <= pi0249 and w32463;
w43107 <= not w43105 and not w43106;
w43108 <= pi0539 and not w32470;
w43109 <= pi0242 and w32470;
w43110 <= not w43108 and not w43109;
w43111 <= pi0540 and not w32470;
w43112 <= pi0235 and w32470;
w43113 <= not w43111 and not w43112;
w43114 <= pi0541 and not w32470;
w43115 <= pi0244 and w32470;
w43116 <= not w43114 and not w43115;
w43117 <= pi0542 and not w32470;
w43118 <= pi0240 and w32470;
w43119 <= not w43117 and not w43118;
w43120 <= pi0543 and not w32470;
w43121 <= pi0238 and w32470;
w43122 <= not w43120 and not w43121;
w43123 <= w32478 and w42994;
w43124 <= pi0544 and not w43123;
w43125 <= not pi0544 and w32473;
w43126 <= w42997 and w43125;
w43127 <= not w43124 and not w43126;
w43128 <= pi0545 and not w32478;
w43129 <= pi0245 and w32478;
w43130 <= not w43128 and not w43129;
w43131 <= pi0546 and not w32478;
w43132 <= pi0246 and w32478;
w43133 <= not w43131 and not w43132;
w43134 <= pi0547 and not w32478;
w43135 <= pi0247 and w32478;
w43136 <= not w43134 and not w43135;
w43137 <= pi0548 and not w32478;
w43138 <= pi0248 and w32478;
w43139 <= not w43137 and not w43138;
w43140 <= pi0549 and not w33674;
w43141 <= pi0235 and w33674;
w43142 <= not w43140 and not w43141;
w43143 <= pi0550 and not w33674;
w43144 <= not pi0239 and w33674;
w43145 <= not w43143 and not w43144;
w43146 <= pi0551 and not w33674;
w43147 <= pi0240 and w33674;
w43148 <= not w43146 and not w43147;
w43149 <= pi0552 and not w33674;
w43150 <= pi0247 and w33674;
w43151 <= not w43149 and not w43150;
w43152 <= pi0553 and not w33674;
w43153 <= pi0241 and w33674;
w43154 <= not w43152 and not w43153;
w43155 <= pi0554 and not w33674;
w43156 <= pi0248 and w33674;
w43157 <= not w43155 and not w43156;
w43158 <= pi0555 and not w33674;
w43159 <= pi0249 and w33674;
w43160 <= not w43158 and not w43159;
w43161 <= pi0556 and not w32354;
w43162 <= pi0242 and w32354;
w43163 <= not w43161 and not w43162;
w43164 <= w32463 and w42994;
w43165 <= pi0557 and not w43164;
w43166 <= not pi0557 and w32146;
w43167 <= w42997 and w43166;
w43168 <= not w43165 and not w43167;
w43169 <= pi0558 and not w32463;
w43170 <= pi0244 and w32463;
w43171 <= not w43169 and not w43170;
w43172 <= pi0559 and not w32338;
w43173 <= pi0241 and w32338;
w43174 <= not w43172 and not w43173;
w43175 <= pi0560 and not w32354;
w43176 <= pi0240 and w32354;
w43177 <= not w43175 and not w43176;
w43178 <= pi0561 and not w32346;
w43179 <= pi0247 and w32346;
w43180 <= not w43178 and not w43179;
w43181 <= pi0562 and not w32354;
w43182 <= pi0241 and w32354;
w43183 <= not w43181 and not w43182;
w43184 <= pi0563 and not w33674;
w43185 <= pi0246 and w33674;
w43186 <= not w43184 and not w43185;
w43187 <= pi0564 and not w32354;
w43188 <= pi0246 and w32354;
w43189 <= not w43187 and not w43188;
w43190 <= pi0565 and not w32354;
w43191 <= pi0248 and w32354;
w43192 <= not w43190 and not w43191;
w43193 <= pi0566 and not w32354;
w43194 <= pi0244 and w32354;
w43195 <= not w43193 and not w43194;
w43196 <= not pi0567 and pi1092;
w43197 <= not pi1093 and w43196;
w43198 <= pi0603 and not w14680;
w43199 <= w14745 and not w17788;
w43200 <= not w17798 and w43199;
w43201 <= w43198 and w43200;
w43202 <= not pi0789 and not w43197;
w43203 <= not w43201 and w43202;
w43204 <= not pi0619 and w43201;
w43205 <= not w43197 and not w43204;
w43206 <= not pi1159 and not w43205;
w43207 <= pi0619 and w43201;
w43208 <= not w43197 and not w43207;
w43209 <= pi1159 and not w43208;
w43210 <= pi0789 and not w43206;
w43211 <= not w43209 and w43210;
w43212 <= not w43203 and not w43211;
w43213 <= pi0680 and w14389;
w43214 <= not w16709 and w43213;
w43215 <= not w43197 and not w43214;
w43216 <= w16713 and not w43215;
w43217 <= not w14197 and w43211;
w43218 <= w43216 and not w43217;
w43219 <= not w43212 and not w43218;
w43220 <= w15533 and not w43219;
w43221 <= w32920 and w43212;
w43222 <= not w14198 and w43216;
w43223 <= pi0641 and w43222;
w43224 <= not w43197 and not w43223;
w43225 <= w15428 and not w43224;
w43226 <= not pi0641 and w43222;
w43227 <= not w43197 and not w43226;
w43228 <= w15429 and not w43227;
w43229 <= not w43225 and not w43228;
w43230 <= not w43221 and w43229;
w43231 <= pi0788 and not w43230;
w43232 <= not w43220 and not w43231;
w43233 <= not w17927 and not w43232;
w43234 <= w16714 and not w43215;
w43235 <= pi0628 and w43234;
w43236 <= not w43197 and not w43235;
w43237 <= pi1156 and not w43236;
w43238 <= not w15532 and w43212;
w43239 <= w15532 and w43197;
w43240 <= not w43238 and not w43239;
w43241 <= w15417 and not w43240;
w43242 <= not pi0629 and not w43237;
w43243 <= not w43241 and w43242;
w43244 <= not pi0628 and w43234;
w43245 <= not w43197 and not w43244;
w43246 <= not pi1156 and not w43245;
w43247 <= w15416 and not w43240;
w43248 <= pi0629 and not w43246;
w43249 <= not w43247 and w43248;
w43250 <= pi0792 and not w43243;
w43251 <= not w43249 and w43250;
w43252 <= not w43233 and not w43251;
w43253 <= not pi0647 and not w43252;
w43254 <= not w15342 and not w43240;
w43255 <= w15342 and w43197;
w43256 <= not w43254 and not w43255;
w43257 <= pi0647 and not w43256;
w43258 <= not pi1157 and not w43257;
w43259 <= not w43253 and w43258;
w43260 <= not w16705 and w43234;
w43261 <= pi0647 and w43260;
w43262 <= pi1157 and not w43197;
w43263 <= not w43261 and w43262;
w43264 <= not pi0630 and not w43263;
w43265 <= not w43259 and w43264;
w43266 <= pi0647 and not w43252;
w43267 <= not pi0647 and not w43256;
w43268 <= pi1157 and not w43267;
w43269 <= not w43266 and w43268;
w43270 <= not pi0647 and w43260;
w43271 <= not pi1157 and not w43197;
w43272 <= not w43270 and w43271;
w43273 <= pi0630 and not w43272;
w43274 <= not w43269 and w43273;
w43275 <= not w43265 and not w43274;
w43276 <= pi0787 and not w43275;
w43277 <= not pi0787 and not w43252;
w43278 <= not w43276 and not w43277;
w43279 <= not pi0790 and not w43278;
w43280 <= not w16905 and w43260;
w43281 <= not w43197 and not w43280;
w43282 <= pi0644 and not w43281;
w43283 <= not pi0644 and not w43278;
w43284 <= not pi0715 and not w43282;
w43285 <= not w43283 and w43284;
w43286 <= not w15367 and w43254;
w43287 <= not pi0644 and w43286;
w43288 <= pi0715 and not w43197;
w43289 <= not w43287 and w43288;
w43290 <= not w43285 and not w43289;
w43291 <= not pi1160 and not w43290;
w43292 <= pi0644 and w43286;
w43293 <= not w43197 and not w43292;
w43294 <= not pi0715 and not w43293;
w43295 <= not pi0644 and w43281;
w43296 <= pi0644 and w43278;
w43297 <= pi0715 and not w43295;
w43298 <= not w43296 and w43297;
w43299 <= pi1160 and not w43294;
w43300 <= not w43298 and w43299;
w43301 <= pi0790 and not w43300;
w43302 <= not w43291 and w43301;
w43303 <= not w43279 and not w43302;
w43304 <= pi0230 and not w43303;
w43305 <= not pi0230 and w43196;
w43306 <= not w43304 and not w43305;
w43307 <= pi0568 and not w32354;
w43308 <= pi0245 and w32354;
w43309 <= not w43307 and not w43308;
w43310 <= pi0569 and not w32354;
w43311 <= not pi0239 and w32354;
w43312 <= not w43310 and not w43311;
w43313 <= w32354 and w43018;
w43314 <= pi0570 and not w43313;
w43315 <= not pi0570 and w32349;
w43316 <= w43042 and w43315;
w43317 <= not w43314 and not w43316;
w43318 <= pi0571 and not w33702;
w43319 <= pi0241 and w33702;
w43320 <= not w43318 and not w43319;
w43321 <= pi0572 and not w33702;
w43322 <= pi0244 and w33702;
w43323 <= not w43321 and not w43322;
w43324 <= pi0573 and not w33702;
w43325 <= pi0242 and w33702;
w43326 <= not w43324 and not w43325;
w43327 <= pi0574 and not w32346;
w43328 <= pi0241 and w32346;
w43329 <= not w43327 and not w43328;
w43330 <= pi0575 and not w33702;
w43331 <= pi0235 and w33702;
w43332 <= not w43330 and not w43331;
w43333 <= pi0576 and not w33702;
w43334 <= pi0248 and w33702;
w43335 <= not w43333 and not w43334;
w43336 <= pi0577 and not w33674;
w43337 <= pi0238 and w33674;
w43338 <= not w43336 and not w43337;
w43339 <= pi0578 and not w32346;
w43340 <= pi0249 and w32346;
w43341 <= not w43339 and not w43340;
w43342 <= pi0579 and not w32338;
w43343 <= pi0249 and w32338;
w43344 <= not w43342 and not w43343;
w43345 <= pi0580 and not w33674;
w43346 <= pi0245 and w33674;
w43347 <= not w43345 and not w43346;
w43348 <= pi0581 and not w32346;
w43349 <= pi0235 and w32346;
w43350 <= not w43348 and not w43349;
w43351 <= pi0582 and not w32346;
w43352 <= pi0240 and w32346;
w43353 <= not w43351 and not w43352;
w43354 <= pi0584 and not w32346;
w43355 <= pi0245 and w32346;
w43356 <= not w43354 and not w43355;
w43357 <= pi0585 and not w32346;
w43358 <= pi0244 and w32346;
w43359 <= not w43357 and not w43358;
w43360 <= pi0586 and not w32346;
w43361 <= pi0242 and w32346;
w43362 <= not w43360 and not w43361;
w43363 <= not pi0230 and pi0587;
w43364 <= pi0230 and w14731;
w43365 <= not w17788 and w43364;
w43366 <= not w33138 and w43365;
w43367 <= w17800 and w43366;
w43368 <= w28360 and w43367;
w43369 <= not w43363 and not w43368;
w43370 <= not pi0123 and w9936;
w43371 <= not pi0588 and not w43370;
w43372 <= not pi0591 and w43370;
w43373 <= w42269 and not w43371;
w43374 <= not w43372 and w43373;
w43375 <= not pi0204 and w42993;
w43376 <= not pi0201 and w43017;
w43377 <= pi0233 and not w43375;
w43378 <= not w43376 and w43377;
w43379 <= not pi0205 and w42993;
w43380 <= not pi0202 and w43017;
w43381 <= not pi0233 and not w43379;
w43382 <= not w43380 and w43381;
w43383 <= not w43378 and not w43382;
w43384 <= pi0237 and not w43383;
w43385 <= not pi0206 and w42993;
w43386 <= not pi0220 and w43017;
w43387 <= pi0233 and not w43385;
w43388 <= not w43386 and w43387;
w43389 <= not pi0218 and w42993;
w43390 <= not pi0203 and w43017;
w43391 <= not pi0233 and not w43389;
w43392 <= not w43390 and w43391;
w43393 <= not w43388 and not w43392;
w43394 <= not pi0237 and not w43393;
w43395 <= not w43384 and not w43394;
w43396 <= pi0588 and w43370;
w43397 <= pi0590 and not w43370;
w43398 <= w42269 and not w43396;
w43399 <= not w43397 and w43398;
w43400 <= not pi0591 and not w43370;
w43401 <= not pi0592 and w43370;
w43402 <= w42269 and not w43400;
w43403 <= not w43401 and w43402;
w43404 <= not pi0592 and not w43370;
w43405 <= not pi0590 and w43370;
w43406 <= w42269 and not w43404;
w43407 <= not w43405 and w43406;
w43408 <= pi0234 and w43017;
w43409 <= pi0518 and not w43408;
w43410 <= pi0246 and not pi0520;
w43411 <= not pi0246 and pi0520;
w43412 <= pi0249 and not pi0578;
w43413 <= not pi0249 and pi0578;
w43414 <= pi0248 and not pi0521;
w43415 <= not pi0248 and pi0521;
w43416 <= pi0241 and pi0574;
w43417 <= not pi0241 and not pi0574;
w43418 <= not w43416 and not w43417;
w43419 <= not pi0518 and not w43018;
w43420 <= not w43410 and not w43411;
w43421 <= not w43412 and not w43413;
w43422 <= not w43414 and not w43415;
w43423 <= w43421 and w43422;
w43424 <= not w43418 and w43420;
w43425 <= w43423 and w43424;
w43426 <= not w43409 and w43425;
w43427 <= not w43419 and w43426;
w43428 <= pi0582 and w43427;
w43429 <= pi0240 and not w43428;
w43430 <= not pi0582 and w43427;
w43431 <= not pi0240 and not w43430;
w43432 <= not w43429 and not w43431;
w43433 <= not pi0239 and pi0519;
w43434 <= pi0239 and not pi0519;
w43435 <= not w43433 and not w43434;
w43436 <= w43432 and not w43435;
w43437 <= pi0242 and pi0586;
w43438 <= not pi0242 and not pi0586;
w43439 <= not w43437 and not w43438;
w43440 <= w43436 and not w43439;
w43441 <= pi0235 and pi0581;
w43442 <= not pi0235 and not pi0581;
w43443 <= not w43441 and not w43442;
w43444 <= w43440 and not w43443;
w43445 <= pi0585 and w43444;
w43446 <= pi0244 and not w43445;
w43447 <= not pi0585 and w43444;
w43448 <= not pi0244 and not w43447;
w43449 <= not w43446 and not w43448;
w43450 <= pi0584 and w43449;
w43451 <= pi0245 and not w43450;
w43452 <= not pi0584 and w43449;
w43453 <= not pi0245 and not w43452;
w43454 <= not w43451 and not w43453;
w43455 <= not pi0247 and not pi0561;
w43456 <= pi0247 and pi0561;
w43457 <= not w43455 and not w43456;
w43458 <= w43454 and not w43457;
w43459 <= pi0238 and w43458;
w43460 <= pi0240 and pi0542;
w43461 <= not pi0240 and not pi0542;
w43462 <= not w43460 and not w43461;
w43463 <= not pi0248 and not pi0501;
w43464 <= pi0248 and pi0501;
w43465 <= not w43463 and not w43464;
w43466 <= pi0234 and w42993;
w43467 <= pi0505 and not w43466;
w43468 <= not pi0505 and not w42994;
w43469 <= pi0249 and not pi0496;
w43470 <= not pi0249 and pi0496;
w43471 <= not pi0246 and not pi0499;
w43472 <= pi0246 and pi0499;
w43473 <= not w43471 and not w43472;
w43474 <= not w43469 and not w43470;
w43475 <= not w43465 and w43474;
w43476 <= not w43473 and w43475;
w43477 <= not w43467 and w43476;
w43478 <= not w43468 and w43477;
w43479 <= not pi0241 and not pi0500;
w43480 <= pi0241 and pi0500;
w43481 <= not w43479 and not w43480;
w43482 <= w43478 and not w43481;
w43483 <= not w43462 and w43482;
w43484 <= pi0497 and w43483;
w43485 <= not pi0239 and not w43484;
w43486 <= not pi0497 and w43483;
w43487 <= pi0239 and not w43486;
w43488 <= not w43485 and not w43487;
w43489 <= pi0539 and w43488;
w43490 <= pi0242 and not w43489;
w43491 <= not pi0539 and w43488;
w43492 <= not pi0242 and not w43491;
w43493 <= not w43490 and not w43492;
w43494 <= pi0540 and w43493;
w43495 <= pi0235 and not w43494;
w43496 <= not pi0540 and w43493;
w43497 <= not pi0235 and not w43496;
w43498 <= not w43495 and not w43497;
w43499 <= pi0244 and pi0541;
w43500 <= not pi0244 and not pi0541;
w43501 <= not w43499 and not w43500;
w43502 <= w43498 and not w43501;
w43503 <= pi0245 and pi0503;
w43504 <= not pi0245 and not pi0503;
w43505 <= not w43503 and not w43504;
w43506 <= w43502 and not w43505;
w43507 <= not pi0502 and w43506;
w43508 <= not pi0247 and not w43507;
w43509 <= pi0502 and w43506;
w43510 <= pi0247 and not w43509;
w43511 <= not w43508 and not w43510;
w43512 <= not pi0238 and w43511;
w43513 <= pi0522 and not w43459;
w43514 <= not w43512 and w43513;
w43515 <= not w43455 and not w43508;
w43516 <= pi0502 and not w43454;
w43517 <= not pi0500 and w43482;
w43518 <= w43478 and w43480;
w43519 <= not w43427 and not w43518;
w43520 <= not w43517 and w43519;
w43521 <= not pi0582 and not w43520;
w43522 <= pi0582 and w43482;
w43523 <= not pi0240 and not w43522;
w43524 <= not w43521 and w43523;
w43525 <= not w43429 and not w43524;
w43526 <= not pi0542 and not w43525;
w43527 <= pi0582 and not w43520;
w43528 <= not pi0582 and w43482;
w43529 <= pi0240 and not w43528;
w43530 <= not w43527 and w43529;
w43531 <= not w43431 and not w43530;
w43532 <= pi0542 and not w43531;
w43533 <= not w43526 and not w43532;
w43534 <= not pi0497 and w43533;
w43535 <= pi0497 and w43432;
w43536 <= pi0239 and not w43535;
w43537 <= not w43534 and w43536;
w43538 <= not w43485 and not w43537;
w43539 <= not pi0519 and not w43538;
w43540 <= pi0497 and w43533;
w43541 <= not pi0497 and w43432;
w43542 <= not pi0239 and not w43541;
w43543 <= not w43540 and w43542;
w43544 <= not w43487 and not w43543;
w43545 <= pi0519 and not w43544;
w43546 <= not w43539 and not w43545;
w43547 <= not pi0539 and w43546;
w43548 <= pi0539 and w43436;
w43549 <= not pi0242 and not w43548;
w43550 <= not w43547 and w43549;
w43551 <= not w43490 and not w43550;
w43552 <= not pi0586 and not w43551;
w43553 <= pi0539 and w43546;
w43554 <= not pi0539 and w43436;
w43555 <= pi0242 and not w43554;
w43556 <= not w43553 and w43555;
w43557 <= not w43492 and not w43556;
w43558 <= pi0586 and not w43557;
w43559 <= not w43552 and not w43558;
w43560 <= not pi0540 and w43559;
w43561 <= pi0540 and w43440;
w43562 <= not pi0235 and not w43561;
w43563 <= not w43560 and w43562;
w43564 <= not w43495 and not w43563;
w43565 <= not pi0581 and not w43564;
w43566 <= pi0540 and w43559;
w43567 <= not pi0540 and w43440;
w43568 <= pi0235 and not w43567;
w43569 <= not w43566 and w43568;
w43570 <= not w43497 and not w43569;
w43571 <= pi0581 and not w43570;
w43572 <= not w43565 and not w43571;
w43573 <= not pi0585 and w43572;
w43574 <= pi0585 and w43498;
w43575 <= not pi0244 and not w43574;
w43576 <= not w43573 and w43575;
w43577 <= not w43446 and not w43576;
w43578 <= not pi0541 and not w43577;
w43579 <= pi0585 and w43572;
w43580 <= not pi0585 and w43498;
w43581 <= pi0244 and not w43580;
w43582 <= not w43579 and w43581;
w43583 <= not w43448 and not w43582;
w43584 <= pi0541 and not w43583;
w43585 <= not w43578 and not w43584;
w43586 <= not pi0584 and w43585;
w43587 <= pi0584 and w43502;
w43588 <= not pi0245 and not w43587;
w43589 <= not w43586 and w43588;
w43590 <= not w43451 and not w43589;
w43591 <= not pi0503 and not w43590;
w43592 <= pi0584 and w43585;
w43593 <= not pi0584 and w43502;
w43594 <= pi0245 and not w43593;
w43595 <= not w43592 and w43594;
w43596 <= not w43453 and not w43595;
w43597 <= pi0503 and not w43596;
w43598 <= not w43591 and not w43597;
w43599 <= not pi0502 and not w43598;
w43600 <= not pi0561 and not w43516;
w43601 <= not w43599 and w43600;
w43602 <= not w43515 and not w43601;
w43603 <= not w43456 and not w43510;
w43604 <= not pi0502 and not w43454;
w43605 <= pi0502 and not w43598;
w43606 <= pi0561 and not w43604;
w43607 <= not w43605 and w43606;
w43608 <= not w43603 and not w43607;
w43609 <= not w43602 and not w43608;
w43610 <= not pi0238 and w43609;
w43611 <= not pi0522 and not w43610;
w43612 <= not pi0543 and not w43514;
w43613 <= not w43611 and w43612;
w43614 <= not pi0238 and w43458;
w43615 <= pi0238 and w43511;
w43616 <= not pi0522 and not w43614;
w43617 <= not w43615 and w43616;
w43618 <= pi0238 and w43609;
w43619 <= pi0522 and not w43618;
w43620 <= pi0543 and not w43617;
w43621 <= not w43619 and w43620;
w43622 <= not w43613 and not w43621;
w43623 <= not pi0233 and not w43622;
w43624 <= pi0246 and pi0536;
w43625 <= not pi0246 and not pi0536;
w43626 <= not w43624 and not w43625;
w43627 <= not pi0557 and not w42994;
w43628 <= pi0557 and not w43466;
w43629 <= not w43626 and not w43627;
w43630 <= not w43628 and w43629;
w43631 <= not pi0538 and w43630;
w43632 <= not pi0249 and not w43631;
w43633 <= pi0538 and w43630;
w43634 <= pi0249 and not w43633;
w43635 <= not w43632 and not w43634;
w43636 <= not pi0537 and w43635;
w43637 <= not pi0248 and not w43636;
w43638 <= pi0537 and w43635;
w43639 <= pi0248 and not w43638;
w43640 <= not w43637 and not w43639;
w43641 <= pi0241 and pi0506;
w43642 <= not pi0241 and not pi0506;
w43643 <= not w43641 and not w43642;
w43644 <= w43640 and not w43643;
w43645 <= pi0240 and pi0535;
w43646 <= not pi0240 and not pi0535;
w43647 <= not w43645 and not w43646;
w43648 <= w43644 and not w43647;
w43649 <= pi0534 and w43648;
w43650 <= not pi0239 and not w43649;
w43651 <= not pi0534 and w43648;
w43652 <= pi0239 and not w43651;
w43653 <= not w43650 and not w43652;
w43654 <= pi0504 and w43653;
w43655 <= pi0242 and not w43654;
w43656 <= not pi0504 and w43653;
w43657 <= not pi0242 and not w43656;
w43658 <= not w43655 and not w43657;
w43659 <= pi0533 and w43658;
w43660 <= pi0235 and not w43659;
w43661 <= not pi0533 and w43658;
w43662 <= not pi0235 and not w43661;
w43663 <= not w43660 and not w43662;
w43664 <= pi0558 and w43663;
w43665 <= pi0244 and not w43664;
w43666 <= not pi0558 and w43663;
w43667 <= not pi0244 and not w43666;
w43668 <= not w43665 and not w43667;
w43669 <= pi0509 and w43668;
w43670 <= pi0245 and not w43669;
w43671 <= not pi0509 and w43668;
w43672 <= not pi0245 and not w43671;
w43673 <= not w43670 and not w43672;
w43674 <= pi0508 and w43673;
w43675 <= pi0247 and not w43674;
w43676 <= not pi0508 and w43673;
w43677 <= not pi0247 and not w43676;
w43678 <= not w43675 and not w43677;
w43679 <= not pi0238 and w43678;
w43680 <= pi0248 and pi0481;
w43681 <= not pi0248 and not pi0481;
w43682 <= not w43680 and not w43681;
w43683 <= pi0246 and pi0487;
w43684 <= not pi0246 and not pi0487;
w43685 <= not w43683 and not w43684;
w43686 <= not pi0511 and not w43018;
w43687 <= pi0511 and not w43408;
w43688 <= not w43685 and not w43686;
w43689 <= not w43687 and w43688;
w43690 <= not pi0249 and not pi0579;
w43691 <= pi0249 and pi0579;
w43692 <= not w43690 and not w43691;
w43693 <= w43689 and not w43692;
w43694 <= not w43682 and w43693;
w43695 <= pi0559 and w43694;
w43696 <= pi0241 and not w43695;
w43697 <= not pi0559 and w43694;
w43698 <= not pi0241 and not w43697;
w43699 <= not w43696 and not w43698;
w43700 <= pi0515 and w43699;
w43701 <= pi0240 and not w43700;
w43702 <= not pi0515 and w43699;
w43703 <= not pi0240 and not w43702;
w43704 <= not w43701 and not w43703;
w43705 <= not pi0239 and pi0488;
w43706 <= pi0239 and not pi0488;
w43707 <= not w43705 and not w43706;
w43708 <= w43704 and not w43707;
w43709 <= pi0242 and pi0510;
w43710 <= not pi0242 and not pi0510;
w43711 <= not w43709 and not w43710;
w43712 <= w43708 and not w43711;
w43713 <= pi0235 and pi0512;
w43714 <= not pi0235 and not pi0512;
w43715 <= not w43713 and not w43714;
w43716 <= w43712 and not w43715;
w43717 <= pi0244 and pi0513;
w43718 <= not pi0244 and not pi0513;
w43719 <= not w43717 and not w43718;
w43720 <= w43716 and not w43719;
w43721 <= pi0245 and pi0514;
w43722 <= not pi0245 and not pi0514;
w43723 <= not w43721 and not w43722;
w43724 <= w43720 and not w43723;
w43725 <= pi0247 and pi0516;
w43726 <= not pi0247 and not pi0516;
w43727 <= not w43725 and not w43726;
w43728 <= w43724 and not w43727;
w43729 <= pi0238 and w43728;
w43730 <= pi0517 and not w43729;
w43731 <= not w43679 and w43730;
w43732 <= not pi0579 and not w43693;
w43733 <= not w43632 and w43689;
w43734 <= pi0579 and not w43733;
w43735 <= not w43732 and not w43734;
w43736 <= not w43635 and not w43735;
w43737 <= not pi0537 and not w43736;
w43738 <= pi0537 and w43693;
w43739 <= not pi0248 and not w43738;
w43740 <= not w43737 and w43739;
w43741 <= not w43639 and not w43740;
w43742 <= not pi0481 and not w43741;
w43743 <= pi0537 and not w43736;
w43744 <= not pi0537 and w43693;
w43745 <= pi0248 and not w43744;
w43746 <= not w43743 and w43745;
w43747 <= not w43637 and not w43746;
w43748 <= pi0481 and not w43747;
w43749 <= not w43742 and not w43748;
w43750 <= not pi0559 and w43749;
w43751 <= pi0559 and w43640;
w43752 <= not pi0241 and not w43751;
w43753 <= not w43750 and w43752;
w43754 <= not w43696 and not w43753;
w43755 <= not pi0506 and not w43754;
w43756 <= pi0559 and w43749;
w43757 <= not pi0559 and w43640;
w43758 <= pi0241 and not w43757;
w43759 <= not w43756 and w43758;
w43760 <= not w43698 and not w43759;
w43761 <= pi0506 and not w43760;
w43762 <= not w43755 and not w43761;
w43763 <= not pi0515 and w43762;
w43764 <= pi0515 and w43644;
w43765 <= not pi0240 and not w43764;
w43766 <= not w43763 and w43765;
w43767 <= not w43701 and not w43766;
w43768 <= not pi0535 and not w43767;
w43769 <= pi0515 and w43762;
w43770 <= not pi0515 and w43644;
w43771 <= pi0240 and not w43770;
w43772 <= not w43769 and w43771;
w43773 <= not w43703 and not w43772;
w43774 <= pi0535 and not w43773;
w43775 <= not w43768 and not w43774;
w43776 <= not pi0534 and w43775;
w43777 <= pi0534 and w43704;
w43778 <= pi0239 and not w43777;
w43779 <= not w43776 and w43778;
w43780 <= not w43650 and not w43779;
w43781 <= not pi0488 and not w43780;
w43782 <= pi0534 and w43775;
w43783 <= not pi0534 and w43704;
w43784 <= not pi0239 and not w43783;
w43785 <= not w43782 and w43784;
w43786 <= not w43652 and not w43785;
w43787 <= pi0488 and not w43786;
w43788 <= not w43781 and not w43787;
w43789 <= not pi0504 and w43788;
w43790 <= pi0504 and w43708;
w43791 <= not pi0242 and not w43790;
w43792 <= not w43789 and w43791;
w43793 <= not w43655 and not w43792;
w43794 <= not pi0510 and not w43793;
w43795 <= pi0504 and w43788;
w43796 <= not pi0504 and w43708;
w43797 <= pi0242 and not w43796;
w43798 <= not w43795 and w43797;
w43799 <= not w43657 and not w43798;
w43800 <= pi0510 and not w43799;
w43801 <= not w43794 and not w43800;
w43802 <= not pi0533 and w43801;
w43803 <= pi0533 and w43712;
w43804 <= not pi0235 and not w43803;
w43805 <= not w43802 and w43804;
w43806 <= not w43660 and not w43805;
w43807 <= not pi0512 and not w43806;
w43808 <= pi0533 and w43801;
w43809 <= not pi0533 and w43712;
w43810 <= pi0235 and not w43809;
w43811 <= not w43808 and w43810;
w43812 <= not w43662 and not w43811;
w43813 <= pi0512 and not w43812;
w43814 <= not w43807 and not w43813;
w43815 <= not pi0558 and w43814;
w43816 <= pi0558 and w43716;
w43817 <= not pi0244 and not w43816;
w43818 <= not w43815 and w43817;
w43819 <= not w43665 and not w43818;
w43820 <= not pi0513 and not w43819;
w43821 <= pi0558 and w43814;
w43822 <= not pi0558 and w43716;
w43823 <= pi0244 and not w43822;
w43824 <= not w43821 and w43823;
w43825 <= not w43667 and not w43824;
w43826 <= pi0513 and not w43825;
w43827 <= not w43820 and not w43826;
w43828 <= not pi0509 and w43827;
w43829 <= pi0509 and w43720;
w43830 <= not pi0245 and not w43829;
w43831 <= not w43828 and w43830;
w43832 <= not w43670 and not w43831;
w43833 <= not pi0514 and not w43832;
w43834 <= pi0509 and w43827;
w43835 <= not pi0509 and w43720;
w43836 <= pi0245 and not w43835;
w43837 <= not w43834 and w43836;
w43838 <= not w43672 and not w43837;
w43839 <= pi0514 and not w43838;
w43840 <= not w43833 and not w43839;
w43841 <= not pi0508 and w43840;
w43842 <= pi0508 and w43724;
w43843 <= not pi0247 and not w43842;
w43844 <= not w43841 and w43843;
w43845 <= not w43675 and not w43844;
w43846 <= not pi0516 and not w43845;
w43847 <= pi0508 and w43840;
w43848 <= not pi0508 and w43724;
w43849 <= pi0247 and not w43848;
w43850 <= not w43847 and w43849;
w43851 <= not w43677 and not w43850;
w43852 <= pi0516 and not w43851;
w43853 <= not w43846 and not w43852;
w43854 <= not pi0238 and w43853;
w43855 <= not pi0517 and not w43854;
w43856 <= not pi0507 and not w43731;
w43857 <= not w43855 and w43856;
w43858 <= pi0238 and w43678;
w43859 <= not pi0238 and w43728;
w43860 <= not pi0517 and not w43859;
w43861 <= not w43858 and w43860;
w43862 <= pi0238 and w43853;
w43863 <= pi0517 and not w43862;
w43864 <= pi0507 and not w43861;
w43865 <= not w43863 and w43864;
w43866 <= not w43857 and not w43865;
w43867 <= pi0233 and not w43866;
w43868 <= pi0237 and not w43623;
w43869 <= not w43867 and w43868;
w43870 <= not pi0240 and not pi0492;
w43871 <= pi0240 and pi0492;
w43872 <= not w43870 and not w43871;
w43873 <= pi0241 and pi0490;
w43874 <= not pi0241 and not pi0490;
w43875 <= not w43873 and not w43874;
w43876 <= pi0248 and pi0548;
w43877 <= not pi0248 and not pi0548;
w43878 <= not w43876 and not w43877;
w43879 <= pi0249 and pi0484;
w43880 <= not pi0249 and not pi0484;
w43881 <= not w43879 and not w43880;
w43882 <= pi0246 and pi0546;
w43883 <= not pi0246 and not pi0546;
w43884 <= not w43882 and not w43883;
w43885 <= not pi0544 and not w42994;
w43886 <= pi0544 and not w43466;
w43887 <= not w43878 and not w43881;
w43888 <= not w43884 and w43887;
w43889 <= not w43885 and w43888;
w43890 <= not w43886 and w43889;
w43891 <= not w43875 and w43890;
w43892 <= not w43872 and w43891;
w43893 <= pi0494 and w43892;
w43894 <= not pi0239 and not w43893;
w43895 <= not pi0494 and w43892;
w43896 <= pi0239 and not w43895;
w43897 <= not w43894 and not w43896;
w43898 <= pi0483 and w43897;
w43899 <= pi0242 and not w43898;
w43900 <= not pi0483 and w43897;
w43901 <= not pi0242 and not w43900;
w43902 <= not w43899 and not w43901;
w43903 <= pi0495 and w43902;
w43904 <= pi0235 and not w43903;
w43905 <= not pi0495 and w43902;
w43906 <= not pi0235 and not w43905;
w43907 <= not w43904 and not w43906;
w43908 <= pi0244 and pi0493;
w43909 <= not pi0244 and not pi0493;
w43910 <= not w43908 and not w43909;
w43911 <= w43907 and not w43910;
w43912 <= pi0545 and w43911;
w43913 <= pi0245 and not w43912;
w43914 <= not pi0545 and w43911;
w43915 <= not pi0245 and not w43914;
w43916 <= not w43913 and not w43915;
w43917 <= pi0547 and w43916;
w43918 <= pi0247 and not w43917;
w43919 <= not pi0547 and w43916;
w43920 <= not pi0247 and not w43919;
w43921 <= not w43918 and not w43920;
w43922 <= not pi0238 and w43921;
w43923 <= pi0523 and not w43408;
w43924 <= pi0248 and pi0576;
w43925 <= not pi0248 and not pi0576;
w43926 <= not w43924 and not w43925;
w43927 <= pi0249 and pi0528;
w43928 <= not pi0249 and not pi0528;
w43929 <= not w43927 and not w43928;
w43930 <= pi0246 and pi0526;
w43931 <= not pi0246 and not pi0526;
w43932 <= not w43930 and not w43931;
w43933 <= not pi0523 and not w43018;
w43934 <= not w43926 and not w43929;
w43935 <= not w43932 and w43934;
w43936 <= not w43923 and w43935;
w43937 <= not w43933 and w43936;
w43938 <= pi0571 and w43937;
w43939 <= pi0241 and not w43938;
w43940 <= not pi0571 and w43937;
w43941 <= not pi0241 and not w43940;
w43942 <= not w43939 and not w43941;
w43943 <= not pi0530 and w43942;
w43944 <= not pi0240 and not w43943;
w43945 <= pi0530 and w43942;
w43946 <= pi0240 and not w43945;
w43947 <= not w43944 and not w43946;
w43948 <= not pi0239 and pi0524;
w43949 <= pi0239 and not pi0524;
w43950 <= not w43948 and not w43949;
w43951 <= w43947 and not w43950;
w43952 <= pi0242 and pi0573;
w43953 <= not pi0242 and not pi0573;
w43954 <= not w43952 and not w43953;
w43955 <= w43951 and not w43954;
w43956 <= pi0235 and pi0575;
w43957 <= not pi0235 and not pi0575;
w43958 <= not w43956 and not w43957;
w43959 <= w43955 and not w43958;
w43960 <= pi0572 and w43959;
w43961 <= pi0244 and not w43960;
w43962 <= not pi0572 and w43959;
w43963 <= not pi0244 and not w43962;
w43964 <= not w43961 and not w43963;
w43965 <= pi0245 and pi0525;
w43966 <= not pi0245 and not pi0525;
w43967 <= not w43965 and not w43966;
w43968 <= w43964 and not w43967;
w43969 <= pi0247 and pi0527;
w43970 <= not pi0247 and not pi0527;
w43971 <= not w43969 and not w43970;
w43972 <= w43968 and not w43971;
w43973 <= pi0238 and w43972;
w43974 <= pi0529 and not w43973;
w43975 <= not w43922 and w43974;
w43976 <= not w43870 and not w43944;
w43977 <= pi0530 and not w43891;
w43978 <= not pi0241 and not w43890;
w43979 <= not w43940 and w43978;
w43980 <= not w43939 and not w43979;
w43981 <= not pi0490 and not w43980;
w43982 <= pi0241 and not w43890;
w43983 <= not w43938 and w43982;
w43984 <= not w43941 and not w43983;
w43985 <= pi0490 and not w43984;
w43986 <= not w43981 and not w43985;
w43987 <= not pi0530 and not w43986;
w43988 <= not pi0492 and not w43977;
w43989 <= not w43987 and w43988;
w43990 <= not w43976 and not w43989;
w43991 <= not w43871 and not w43946;
w43992 <= not pi0530 and not w43891;
w43993 <= pi0530 and not w43986;
w43994 <= pi0492 and not w43992;
w43995 <= not w43993 and w43994;
w43996 <= not w43991 and not w43995;
w43997 <= not w43990 and not w43996;
w43998 <= not pi0494 and w43997;
w43999 <= pi0494 and w43947;
w44000 <= pi0239 and not w43999;
w44001 <= not w43998 and w44000;
w44002 <= not w43894 and not w44001;
w44003 <= not pi0524 and not w44002;
w44004 <= pi0494 and w43997;
w44005 <= not pi0494 and w43947;
w44006 <= not pi0239 and not w44005;
w44007 <= not w44004 and w44006;
w44008 <= not w43896 and not w44007;
w44009 <= pi0524 and not w44008;
w44010 <= not w44003 and not w44009;
w44011 <= not pi0483 and w44010;
w44012 <= pi0483 and w43951;
w44013 <= not pi0242 and not w44012;
w44014 <= not w44011 and w44013;
w44015 <= not w43899 and not w44014;
w44016 <= not pi0573 and not w44015;
w44017 <= pi0483 and w44010;
w44018 <= not pi0483 and w43951;
w44019 <= pi0242 and not w44018;
w44020 <= not w44017 and w44019;
w44021 <= not w43901 and not w44020;
w44022 <= pi0573 and not w44021;
w44023 <= not w44016 and not w44022;
w44024 <= not pi0495 and w44023;
w44025 <= pi0495 and w43955;
w44026 <= not pi0235 and not w44025;
w44027 <= not w44024 and w44026;
w44028 <= not w43904 and not w44027;
w44029 <= not pi0575 and not w44028;
w44030 <= pi0495 and w44023;
w44031 <= not pi0495 and w43955;
w44032 <= pi0235 and not w44031;
w44033 <= not w44030 and w44032;
w44034 <= not w43906 and not w44033;
w44035 <= pi0575 and not w44034;
w44036 <= not w44029 and not w44035;
w44037 <= not pi0572 and w44036;
w44038 <= pi0572 and w43907;
w44039 <= not pi0244 and not w44038;
w44040 <= not w44037 and w44039;
w44041 <= not w43961 and not w44040;
w44042 <= not pi0493 and not w44041;
w44043 <= pi0572 and w44036;
w44044 <= not pi0572 and w43907;
w44045 <= pi0244 and not w44044;
w44046 <= not w44043 and w44045;
w44047 <= not w43963 and not w44046;
w44048 <= pi0493 and not w44047;
w44049 <= not w44042 and not w44048;
w44050 <= not pi0545 and w44049;
w44051 <= pi0545 and w43964;
w44052 <= not pi0245 and not w44051;
w44053 <= not w44050 and w44052;
w44054 <= not w43913 and not w44053;
w44055 <= not pi0525 and not w44054;
w44056 <= pi0545 and w44049;
w44057 <= not pi0545 and w43964;
w44058 <= pi0245 and not w44057;
w44059 <= not w44056 and w44058;
w44060 <= not w43915 and not w44059;
w44061 <= pi0525 and not w44060;
w44062 <= not w44055 and not w44061;
w44063 <= not pi0547 and w44062;
w44064 <= pi0547 and w43968;
w44065 <= not pi0247 and not w44064;
w44066 <= not w44063 and w44065;
w44067 <= not w43918 and not w44066;
w44068 <= not pi0527 and not w44067;
w44069 <= pi0547 and w44062;
w44070 <= not pi0547 and w43968;
w44071 <= pi0247 and not w44070;
w44072 <= not w44069 and w44071;
w44073 <= not w43920 and not w44072;
w44074 <= pi0527 and not w44073;
w44075 <= not w44068 and not w44074;
w44076 <= not pi0238 and w44075;
w44077 <= not pi0529 and not w44076;
w44078 <= not pi0491 and not w43975;
w44079 <= not w44077 and w44078;
w44080 <= pi0238 and w43921;
w44081 <= not pi0238 and w43972;
w44082 <= not pi0529 and not w44081;
w44083 <= not w44080 and w44082;
w44084 <= pi0238 and w44075;
w44085 <= pi0529 and not w44084;
w44086 <= pi0491 and not w44083;
w44087 <= not w44085 and w44086;
w44088 <= not w44079 and not w44087;
w44089 <= pi0233 and not w44088;
w44090 <= pi0485 and not w43466;
w44091 <= pi0240 and pi0551;
w44092 <= not pi0240 and not pi0551;
w44093 <= not w44091 and not w44092;
w44094 <= pi0249 and not pi0555;
w44095 <= not pi0249 and pi0555;
w44096 <= pi0241 and not pi0553;
w44097 <= not pi0241 and pi0553;
w44098 <= pi0248 and not pi0554;
w44099 <= not pi0248 and pi0554;
w44100 <= not pi0246 and pi0563;
w44101 <= pi0246 and not pi0563;
w44102 <= not pi0485 and not w42994;
w44103 <= not w44094 and not w44095;
w44104 <= not w44096 and not w44097;
w44105 <= not w44098 and not w44099;
w44106 <= not w44100 and not w44101;
w44107 <= w44105 and w44106;
w44108 <= w44103 and w44104;
w44109 <= not w44093 and w44108;
w44110 <= w44107 and w44109;
w44111 <= not w44090 and w44110;
w44112 <= not w44102 and w44111;
w44113 <= pi0550 and w44112;
w44114 <= not pi0239 and not w44113;
w44115 <= not pi0550 and w44112;
w44116 <= pi0239 and not w44115;
w44117 <= not w44114 and not w44116;
w44118 <= not pi0489 and w44117;
w44119 <= not pi0242 and not w44118;
w44120 <= pi0489 and w44117;
w44121 <= pi0242 and not w44120;
w44122 <= not w44119 and not w44121;
w44123 <= pi0549 and w44122;
w44124 <= pi0235 and not w44123;
w44125 <= not pi0549 and w44122;
w44126 <= not pi0235 and not w44125;
w44127 <= not w44124 and not w44126;
w44128 <= pi0486 and w44127;
w44129 <= pi0244 and not w44128;
w44130 <= not pi0486 and w44127;
w44131 <= not pi0244 and not w44130;
w44132 <= not w44129 and not w44131;
w44133 <= pi0245 and pi0580;
w44134 <= not pi0245 and not pi0580;
w44135 <= not w44133 and not w44134;
w44136 <= w44132 and not w44135;
w44137 <= pi0552 and w44136;
w44138 <= pi0247 and not w44137;
w44139 <= not pi0552 and w44136;
w44140 <= not pi0247 and not w44139;
w44141 <= not w44138 and not w44140;
w44142 <= pi0238 and w44141;
w44143 <= not pi0242 and not pi0556;
w44144 <= pi0242 and pi0556;
w44145 <= not w44143 and not w44144;
w44146 <= pi0246 and not pi0564;
w44147 <= pi0570 and not w43408;
w44148 <= not pi0246 and pi0564;
w44149 <= pi0249 and not pi0482;
w44150 <= not pi0249 and pi0482;
w44151 <= pi0241 and pi0562;
w44152 <= not pi0241 and not pi0562;
w44153 <= not w44151 and not w44152;
w44154 <= not pi0570 and not w43018;
w44155 <= not w44148 and not w44149;
w44156 <= not w44150 and w44155;
w44157 <= not w44153 and w44156;
w44158 <= not w44147 and w44157;
w44159 <= not w44154 and w44158;
w44160 <= pi0248 and not pi0565;
w44161 <= not pi0248 and pi0565;
w44162 <= not w44160 and not w44161;
w44163 <= pi0240 and pi0560;
w44164 <= not pi0240 and not pi0560;
w44165 <= not w44163 and not w44164;
w44166 <= not w44146 and w44162;
w44167 <= not w44165 and w44166;
w44168 <= w44159 and w44167;
w44169 <= not pi0240 and not w44168;
w44170 <= pi0560 and not w44146;
w44171 <= w44162 and w44170;
w44172 <= w44159 and w44171;
w44173 <= pi0240 and not w44172;
w44174 <= not w44169 and not w44173;
w44175 <= not pi0239 and pi0569;
w44176 <= pi0239 and not pi0569;
w44177 <= not w44175 and not w44176;
w44178 <= w44174 and not w44177;
w44179 <= not w44145 and w44178;
w44180 <= pi0235 and pi0531;
w44181 <= not pi0235 and not pi0531;
w44182 <= not w44180 and not w44181;
w44183 <= w44179 and not w44182;
w44184 <= pi0244 and pi0566;
w44185 <= not pi0244 and not pi0566;
w44186 <= not w44184 and not w44185;
w44187 <= w44183 and not w44186;
w44188 <= pi0568 and w44187;
w44189 <= pi0245 and not w44188;
w44190 <= not pi0568 and w44187;
w44191 <= not pi0245 and not w44190;
w44192 <= not w44189 and not w44191;
w44193 <= pi0247 and pi0532;
w44194 <= not pi0247 and not pi0532;
w44195 <= not w44193 and not w44194;
w44196 <= w44192 and not w44195;
w44197 <= not pi0238 and w44196;
w44198 <= pi0577 and not w44197;
w44199 <= not w44142 and w44198;
w44200 <= not w44119 and not w44143;
w44201 <= pi0489 and not w44178;
w44202 <= w44168 and w44176;
w44203 <= pi0569 and not w44116;
w44204 <= w44174 and w44203;
w44205 <= not w44117 and not w44202;
w44206 <= not w44204 and w44205;
w44207 <= not pi0489 and w44206;
w44208 <= not pi0556 and not w44201;
w44209 <= not w44207 and w44208;
w44210 <= not w44200 and not w44209;
w44211 <= not w44121 and not w44144;
w44212 <= not pi0489 and not w44178;
w44213 <= pi0489 and w44206;
w44214 <= pi0556 and not w44212;
w44215 <= not w44213 and w44214;
w44216 <= not w44211 and not w44215;
w44217 <= not w44210 and not w44216;
w44218 <= not pi0549 and w44217;
w44219 <= pi0549 and w44179;
w44220 <= not pi0235 and not w44219;
w44221 <= not w44218 and w44220;
w44222 <= not w44124 and not w44221;
w44223 <= not pi0531 and not w44222;
w44224 <= pi0549 and w44217;
w44225 <= not pi0549 and w44179;
w44226 <= pi0235 and not w44225;
w44227 <= not w44224 and w44226;
w44228 <= not w44126 and not w44227;
w44229 <= pi0531 and not w44228;
w44230 <= not w44223 and not w44229;
w44231 <= not pi0486 and w44230;
w44232 <= pi0486 and w44183;
w44233 <= not pi0244 and not w44232;
w44234 <= not w44231 and w44233;
w44235 <= not w44129 and not w44234;
w44236 <= not pi0566 and not w44235;
w44237 <= pi0486 and w44230;
w44238 <= not pi0486 and w44183;
w44239 <= pi0244 and not w44238;
w44240 <= not w44237 and w44239;
w44241 <= not w44131 and not w44240;
w44242 <= pi0566 and not w44241;
w44243 <= not w44236 and not w44242;
w44244 <= not pi0568 and w44243;
w44245 <= pi0568 and w44132;
w44246 <= not pi0245 and not w44245;
w44247 <= not w44244 and w44246;
w44248 <= not w44189 and not w44247;
w44249 <= not pi0580 and not w44248;
w44250 <= pi0568 and w44243;
w44251 <= not pi0568 and w44132;
w44252 <= pi0245 and not w44251;
w44253 <= not w44250 and w44252;
w44254 <= not w44191 and not w44253;
w44255 <= pi0580 and not w44254;
w44256 <= not w44249 and not w44255;
w44257 <= not pi0552 and w44256;
w44258 <= pi0552 and w44192;
w44259 <= not pi0247 and not w44258;
w44260 <= not w44257 and w44259;
w44261 <= not w44138 and not w44260;
w44262 <= not pi0532 and not w44261;
w44263 <= pi0552 and w44256;
w44264 <= not pi0552 and w44192;
w44265 <= pi0247 and not w44264;
w44266 <= not w44263 and w44265;
w44267 <= not w44140 and not w44266;
w44268 <= pi0532 and not w44267;
w44269 <= not w44262 and not w44268;
w44270 <= not pi0238 and w44269;
w44271 <= not pi0577 and not w44270;
w44272 <= not pi0498 and not w44199;
w44273 <= not w44271 and w44272;
w44274 <= not pi0238 and w44141;
w44275 <= pi0238 and w44196;
w44276 <= not pi0577 and not w44275;
w44277 <= not w44274 and w44276;
w44278 <= pi0238 and w44269;
w44279 <= pi0577 and not w44278;
w44280 <= pi0498 and not w44277;
w44281 <= not w44279 and w44280;
w44282 <= not w44273 and not w44281;
w44283 <= not pi0233 and not w44282;
w44284 <= not pi0237 and not w44283;
w44285 <= not w44089 and w44284;
w44286 <= not w43869 and not w44285;
w44287 <= not pi0806 and w42689;
w44288 <= not pi0332 and not pi0806;
w44289 <= pi0990 and w44288;
w44290 <= pi0600 and w44289;
w44291 <= not pi0332 and pi0594;
w44292 <= not w44290 and not w44291;
w44293 <= not w44287 and not w44292;
w44294 <= pi0605 and not pi0806;
w44295 <= w42672 and w44294;
w44296 <= not pi0595 and not w44295;
w44297 <= pi0595 and w44295;
w44298 <= not pi0332 and not w44296;
w44299 <= not w44297 and w44298;
w44300 <= not pi0332 and pi0596;
w44301 <= pi0595 and w42671;
w44302 <= w44289 and w44301;
w44303 <= not w44300 and not w44302;
w44304 <= pi0596 and w44302;
w44305 <= not w44303 and not w44304;
w44306 <= not pi0597 and not w44287;
w44307 <= pi0597 and w44287;
w44308 <= not pi0332 and not w44306;
w44309 <= not w44307 and w44308;
w44310 <= not pi0882 and w4989;
w44311 <= pi0947 and w44310;
w44312 <= pi0598 and not w44311;
w44313 <= pi0740 and pi0780;
w44314 <= w3755 and w44313;
w44315 <= not w44312 and not w44314;
w44316 <= not pi0332 and pi0599;
w44317 <= not w44304 and not w44316;
w44318 <= pi0599 and w44304;
w44319 <= not w44317 and not w44318;
w44320 <= not pi0332 and pi0600;
w44321 <= not w44289 and not w44320;
w44322 <= not w44290 and not w44321;
w44323 <= not pi0806 and not pi0989;
w44324 <= not pi0601 and pi0806;
w44325 <= not pi0332 and not w44323;
w44326 <= not w44324 and w44325;
w44327 <= not pi0230 and pi0602;
w44328 <= not pi0715 and not pi1160;
w44329 <= pi0715 and pi1160;
w44330 <= pi0790 and not w44328;
w44331 <= not w44329 and w44330;
w44332 <= pi0230 and w14207;
w44333 <= not w15419 and w44332;
w44334 <= not w16709 and not w16905;
w44335 <= not w44331 and w44334;
w44336 <= w44333 and w44335;
w44337 <= w16714 and w44336;
w44338 <= not w44327 and not w44337;
w44339 <= pi0871 and pi0966;
w44340 <= pi0872 and pi0966;
w44341 <= pi0832 and not pi1100;
w44342 <= not pi0980 and pi1038;
w44343 <= pi1060 and w44342;
w44344 <= pi0952 and not pi1061;
w44345 <= w44343 and w44344;
w44346 <= w44341 and w44345;
w44347 <= pi0832 and w44345;
w44348 <= not pi0603 and not w44347;
w44349 <= not pi0966 and not w44346;
w44350 <= not w44348 and w44349;
w44351 <= not w44339 and not w44340;
w44352 <= not w44350 and w44351;
w44353 <= pi0823 and w14220;
w44354 <= not pi0779 and w44353;
w44355 <= not pi0299 and pi0983;
w44356 <= pi0907 and w44355;
w44357 <= pi0604 and not w44356;
w44358 <= not w44353 and w44357;
w44359 <= not w44354 and not w44358;
w44360 <= not pi0605 and not w44288;
w44361 <= not pi0332 and not w44294;
w44362 <= not w44360 and w44361;
w44363 <= not pi0606 and not w44347;
w44364 <= not pi1104 and w44347;
w44365 <= not w44363 and not w44364;
w44366 <= not pi0966 and not w44365;
w44367 <= not pi0837 and pi0966;
w44368 <= not w44366 and not w44367;
w44369 <= not pi0607 and not w44347;
w44370 <= not pi1107 and w44347;
w44371 <= not pi0966 and not w44369;
w44372 <= not w44370 and w44371;
w44373 <= not pi0608 and not w44347;
w44374 <= not pi1116 and w44347;
w44375 <= not pi0966 and not w44373;
w44376 <= not w44374 and w44375;
w44377 <= not pi0609 and not w44347;
w44378 <= not pi1118 and w44347;
w44379 <= not pi0966 and not w44377;
w44380 <= not w44378 and w44379;
w44381 <= not pi0610 and not w44347;
w44382 <= not pi1113 and w44347;
w44383 <= not pi0966 and not w44381;
w44384 <= not w44382 and w44383;
w44385 <= not pi0611 and not w44347;
w44386 <= not pi1114 and w44347;
w44387 <= not pi0966 and not w44385;
w44388 <= not w44386 and w44387;
w44389 <= not pi0612 and not w44347;
w44390 <= not pi1111 and w44347;
w44391 <= not pi0966 and not w44389;
w44392 <= not w44390 and w44391;
w44393 <= not pi0613 and not w44347;
w44394 <= not pi1115 and w44347;
w44395 <= not pi0966 and not w44393;
w44396 <= not w44394 and w44395;
w44397 <= not pi0614 and not w44347;
w44398 <= not pi1102 and w44347;
w44399 <= not pi0966 and not w44397;
w44400 <= not w44398 and w44399;
w44401 <= not w44339 and not w44400;
w44402 <= pi0907 and w44310;
w44403 <= not pi0615 and not w44402;
w44404 <= pi0779 and pi0797;
w44405 <= w3758 and w44404;
w44406 <= not w44403 and not w44405;
w44407 <= not pi0616 and not w44347;
w44408 <= not pi1101 and w44347;
w44409 <= not pi0966 and not w44407;
w44410 <= not w44408 and w44409;
w44411 <= not w44340 and not w44410;
w44412 <= not pi0617 and not w44347;
w44413 <= not pi1105 and w44347;
w44414 <= not w44412 and not w44413;
w44415 <= not pi0966 and not w44414;
w44416 <= not pi0850 and pi0966;
w44417 <= not w44415 and not w44416;
w44418 <= not pi0618 and not w44347;
w44419 <= not pi1117 and w44347;
w44420 <= not pi0966 and not w44418;
w44421 <= not w44419 and w44420;
w44422 <= not pi0619 and not w44347;
w44423 <= not pi1122 and w44347;
w44424 <= not pi0966 and not w44422;
w44425 <= not w44423 and w44424;
w44426 <= not pi0620 and not w44347;
w44427 <= not pi1112 and w44347;
w44428 <= not pi0966 and not w44426;
w44429 <= not w44427 and w44428;
w44430 <= not pi0621 and not w44347;
w44431 <= not pi1108 and w44347;
w44432 <= not pi0966 and not w44430;
w44433 <= not w44431 and w44432;
w44434 <= not pi0622 and not w44347;
w44435 <= not pi1109 and w44347;
w44436 <= not pi0966 and not w44434;
w44437 <= not w44435 and w44436;
w44438 <= not pi0623 and not w44347;
w44439 <= not pi1106 and w44347;
w44440 <= not pi0966 and not w44438;
w44441 <= not w44439 and w44440;
w44442 <= pi0831 and w14730;
w44443 <= not pi0780 and w44442;
w44444 <= pi0947 and w44355;
w44445 <= pi0624 and not w44444;
w44446 <= not w44442 and w44445;
w44447 <= not w44443 and not w44446;
w44448 <= pi0832 and not pi0973;
w44449 <= not pi1054 and pi1066;
w44450 <= pi1088 and w44449;
w44451 <= w44448 and w44450;
w44452 <= not pi0953 and w44451;
w44453 <= not pi0625 and not w44452;
w44454 <= not pi1116 and w44452;
w44455 <= not pi0962 and not w44453;
w44456 <= not w44454 and w44455;
w44457 <= not pi0626 and not w44347;
w44458 <= not pi1121 and w44347;
w44459 <= not pi0966 and not w44457;
w44460 <= not w44458 and w44459;
w44461 <= not pi0627 and not w44452;
w44462 <= not pi1117 and w44452;
w44463 <= not pi0962 and not w44461;
w44464 <= not w44462 and w44463;
w44465 <= not pi0628 and not w44452;
w44466 <= not pi1119 and w44452;
w44467 <= not pi0962 and not w44465;
w44468 <= not w44466 and w44467;
w44469 <= not pi0629 and not w44347;
w44470 <= not pi1119 and w44347;
w44471 <= not pi0966 and not w44469;
w44472 <= not w44470 and w44471;
w44473 <= not pi0630 and not w44347;
w44474 <= not pi1120 and w44347;
w44475 <= not pi0966 and not w44473;
w44476 <= not w44474 and w44475;
w44477 <= not pi1113 and w44452;
w44478 <= pi0631 and not w44452;
w44479 <= not pi0962 and not w44477;
w44480 <= not w44478 and w44479;
w44481 <= not pi1115 and w44452;
w44482 <= pi0632 and not w44452;
w44483 <= not pi0962 and not w44481;
w44484 <= not w44482 and w44483;
w44485 <= not pi0633 and not w44347;
w44486 <= not pi1110 and w44347;
w44487 <= not pi0966 and not w44485;
w44488 <= not w44486 and w44487;
w44489 <= not pi0634 and not w44452;
w44490 <= not pi1110 and w44452;
w44491 <= not pi0962 and not w44489;
w44492 <= not w44490 and w44491;
w44493 <= not pi1112 and w44452;
w44494 <= pi0635 and not w44452;
w44495 <= not pi0962 and not w44493;
w44496 <= not w44494 and w44495;
w44497 <= not pi0636 and not w44347;
w44498 <= not pi1127 and w44347;
w44499 <= not pi0966 and not w44497;
w44500 <= not w44498 and w44499;
w44501 <= not pi0637 and not w44452;
w44502 <= not pi1105 and w44452;
w44503 <= not pi0962 and not w44501;
w44504 <= not w44502 and w44503;
w44505 <= not pi0638 and not w44452;
w44506 <= not pi1107 and w44452;
w44507 <= not pi0962 and not w44505;
w44508 <= not w44506 and w44507;
w44509 <= not pi0639 and not w44452;
w44510 <= not pi1109 and w44452;
w44511 <= not pi0962 and not w44509;
w44512 <= not w44510 and w44511;
w44513 <= not pi0640 and not w44347;
w44514 <= not pi1128 and w44347;
w44515 <= not pi0966 and not w44513;
w44516 <= not w44514 and w44515;
w44517 <= not pi0641 and not w44452;
w44518 <= not pi1121 and w44452;
w44519 <= not pi0962 and not w44517;
w44520 <= not w44518 and w44519;
w44521 <= not pi0642 and not w44347;
w44522 <= not pi1103 and w44347;
w44523 <= not pi0966 and not w44521;
w44524 <= not w44522 and w44523;
w44525 <= not pi0643 and not w44452;
w44526 <= not pi1104 and w44452;
w44527 <= not pi0962 and not w44525;
w44528 <= not w44526 and w44527;
w44529 <= not pi0644 and not w44347;
w44530 <= not pi1123 and w44347;
w44531 <= not pi0966 and not w44529;
w44532 <= not w44530 and w44531;
w44533 <= not pi0645 and not w44347;
w44534 <= not pi1125 and w44347;
w44535 <= not pi0966 and not w44533;
w44536 <= not w44534 and w44535;
w44537 <= not pi1114 and w44452;
w44538 <= pi0646 and not w44452;
w44539 <= not pi0962 and not w44537;
w44540 <= not w44538 and w44539;
w44541 <= not pi0647 and not w44452;
w44542 <= not pi1120 and w44452;
w44543 <= not pi0962 and not w44541;
w44544 <= not w44542 and w44543;
w44545 <= not pi0648 and not w44452;
w44546 <= not pi1122 and w44452;
w44547 <= not pi0962 and not w44545;
w44548 <= not w44546 and w44547;
w44549 <= not pi1126 and w44452;
w44550 <= pi0649 and not w44452;
w44551 <= not pi0962 and not w44549;
w44552 <= not w44550 and w44551;
w44553 <= not pi1127 and w44452;
w44554 <= pi0650 and not w44452;
w44555 <= not pi0962 and not w44553;
w44556 <= not w44554 and w44555;
w44557 <= not pi0651 and not w44347;
w44558 <= not pi1130 and w44347;
w44559 <= not pi0966 and not w44557;
w44560 <= not w44558 and w44559;
w44561 <= not pi0652 and not w44347;
w44562 <= not pi1131 and w44347;
w44563 <= not pi0966 and not w44561;
w44564 <= not w44562 and w44563;
w44565 <= not pi0653 and not w44347;
w44566 <= not pi1129 and w44347;
w44567 <= not pi0966 and not w44565;
w44568 <= not w44566 and w44567;
w44569 <= not pi1130 and w44452;
w44570 <= pi0654 and not w44452;
w44571 <= not pi0962 and not w44569;
w44572 <= not w44570 and w44571;
w44573 <= not pi1124 and w44452;
w44574 <= pi0655 and not w44452;
w44575 <= not pi0962 and not w44573;
w44576 <= not w44574 and w44575;
w44577 <= not pi0656 and not w44347;
w44578 <= not pi1126 and w44347;
w44579 <= not pi0966 and not w44577;
w44580 <= not w44578 and w44579;
w44581 <= not pi1131 and w44452;
w44582 <= pi0657 and not w44452;
w44583 <= not pi0962 and not w44581;
w44584 <= not w44582 and w44583;
w44585 <= not pi0658 and not w44347;
w44586 <= not pi1124 and w44347;
w44587 <= not pi0966 and not w44585;
w44588 <= not w44586 and w44587;
w44589 <= pi0266 and pi0992;
w44590 <= not pi0280 and w44589;
w44591 <= not pi0269 and w44590;
w44592 <= not pi0281 and w44591;
w44593 <= not pi0270 and not pi0277;
w44594 <= not pi0282 and w44593;
w44595 <= w44592 and w44594;
w44596 <= not pi0264 and w44595;
w44597 <= not pi0265 and w44596;
w44598 <= not pi0274 and w44597;
w44599 <= pi0274 and not w44597;
w44600 <= not w44598 and not w44599;
w44601 <= not pi0660 and not w44452;
w44602 <= not pi1118 and w44452;
w44603 <= not pi0962 and not w44601;
w44604 <= not w44602 and w44603;
w44605 <= not pi0661 and not w44452;
w44606 <= not pi1101 and w44452;
w44607 <= not pi0962 and not w44605;
w44608 <= not w44606 and w44607;
w44609 <= not pi0662 and not w44452;
w44610 <= not pi1102 and w44452;
w44611 <= not pi0962 and not w44609;
w44612 <= not w44610 and w44611;
w44613 <= not pi0223 and not pi0224;
w44614 <= not pi0199 and not pi0257;
w44615 <= pi0199 and not pi1065;
w44616 <= not w44613 and not w44614;
w44617 <= not w44615 and w44616;
w44618 <= not pi0592 and w5604;
w44619 <= pi0464 and w44618;
w44620 <= pi0588 and not w44619;
w44621 <= not pi0591 and pi0592;
w44622 <= pi0365 and w44621;
w44623 <= pi0334 and pi0591;
w44624 <= not pi0592 and w44623;
w44625 <= not w44622 and not w44624;
w44626 <= not pi0590 and not w44625;
w44627 <= pi0590 and not pi0591;
w44628 <= not pi0592 and w44627;
w44629 <= pi0323 and w44628;
w44630 <= not pi0588 and not w44629;
w44631 <= not w44626 and w44630;
w44632 <= w44613 and not w44620;
w44633 <= not w44631 and w44632;
w44634 <= not w44617 and not w44633;
w44635 <= w5206 and not w44634;
w44636 <= not pi1137 and not pi1138;
w44637 <= not pi1134 and w44636;
w44638 <= not pi0784 and not pi1136;
w44639 <= not pi0634 and pi1136;
w44640 <= pi1135 and not w44638;
w44641 <= not w44639 and w44640;
w44642 <= not pi0815 and not pi1136;
w44643 <= not pi0633 and pi1136;
w44644 <= not pi1135 and not w44642;
w44645 <= not w44643 and w44644;
w44646 <= not w44641 and not w44645;
w44647 <= w44637 and not w44646;
w44648 <= pi1135 and w44636;
w44649 <= pi1136 and not w44648;
w44650 <= not pi0766 and w44649;
w44651 <= not pi0855 and not pi1136;
w44652 <= not pi0700 and pi1135;
w44653 <= pi1135 and not pi1136;
w44654 <= pi1134 and w44636;
w44655 <= not w44653 and w44654;
w44656 <= not w44651 and not w44652;
w44657 <= w44655 and w44656;
w44658 <= not w44650 and w44657;
w44659 <= not w44647 and not w44658;
w44660 <= not w5206 and not w44659;
w44661 <= not w44635 and not w44660;
w44662 <= pi0429 and w44618;
w44663 <= pi0588 and not w44662;
w44664 <= not pi0590 and pi0591;
w44665 <= pi0404 and w44664;
w44666 <= not pi0590 and pi0592;
w44667 <= not pi0588 and not w44666;
w44668 <= not w44665 and w44667;
w44669 <= pi0380 and not pi0591;
w44670 <= pi0592 and not w44669;
w44671 <= not w44668 and not w44670;
w44672 <= pi0355 and w44628;
w44673 <= not w44671 and not w44672;
w44674 <= w44613 and not w44663;
w44675 <= not w44673 and w44674;
w44676 <= not pi0199 and not pi0292;
w44677 <= pi0199 and not pi1084;
w44678 <= not w44613 and not w44676;
w44679 <= not w44677 and w44678;
w44680 <= not w44675 and not w44679;
w44681 <= w5206 and not w44680;
w44682 <= not pi1135 and not pi1136;
w44683 <= pi0872 and w44682;
w44684 <= not pi0772 and not pi1135;
w44685 <= not pi0727 and pi1135;
w44686 <= pi1136 and not w44684;
w44687 <= not w44685 and w44686;
w44688 <= pi1134 and not w44683;
w44689 <= not w44687 and w44688;
w44690 <= not w5206 and w44636;
w44691 <= pi0614 and not pi1135;
w44692 <= pi0662 and pi1135;
w44693 <= pi1136 and not w44691;
w44694 <= not w44692 and w44693;
w44695 <= pi0811 and not pi1135;
w44696 <= pi0785 and pi1135;
w44697 <= not pi1136 and not w44695;
w44698 <= not w44696 and w44697;
w44699 <= not w44694 and not w44698;
w44700 <= not pi1134 and not w44699;
w44701 <= not w44689 and w44690;
w44702 <= not w44700 and w44701;
w44703 <= not w44681 and not w44702;
w44704 <= not pi0665 and not w44452;
w44705 <= not pi1108 and w44452;
w44706 <= not pi0962 and not w44704;
w44707 <= not w44705 and w44706;
w44708 <= not pi0607 and not pi1135;
w44709 <= not pi0638 and pi1135;
w44710 <= pi1136 and not w44708;
w44711 <= not w44709 and w44710;
w44712 <= not pi0790 and pi1135;
w44713 <= pi0799 and not pi1135;
w44714 <= not pi1136 and not w44712;
w44715 <= not w44713 and w44714;
w44716 <= not w44711 and not w44715;
w44717 <= w44637 and not w44716;
w44718 <= not pi0764 and w44649;
w44719 <= not pi0691 and pi1135;
w44720 <= not pi0873 and not pi1136;
w44721 <= not w44719 and not w44720;
w44722 <= w44655 and w44721;
w44723 <= not w44718 and w44722;
w44724 <= not w44717 and not w44723;
w44725 <= not w5206 and not w44724;
w44726 <= not pi0199 and not pi0297;
w44727 <= pi0199 and not pi1044;
w44728 <= not w44613 and not w44726;
w44729 <= not w44727 and w44728;
w44730 <= pi0443 and w44618;
w44731 <= pi0588 and not w44730;
w44732 <= pi0456 and w44664;
w44733 <= w44667 and not w44732;
w44734 <= pi0337 and not pi0591;
w44735 <= pi0592 and not w44734;
w44736 <= not w44733 and not w44735;
w44737 <= pi0441 and w44628;
w44738 <= not w44736 and not w44737;
w44739 <= w44613 and not w44731;
w44740 <= not w44738 and w44739;
w44741 <= not w44729 and not w44740;
w44742 <= w5206 and not w44741;
w44743 <= not w44725 and not w44742;
w44744 <= pi0444 and w44618;
w44745 <= pi0588 and not w44744;
w44746 <= pi0319 and w44664;
w44747 <= w44667 and not w44746;
w44748 <= pi0338 and not pi0591;
w44749 <= pi0592 and not w44748;
w44750 <= not w44747 and not w44749;
w44751 <= pi0458 and w44628;
w44752 <= not w44750 and not w44751;
w44753 <= w44613 and not w44745;
w44754 <= not w44752 and w44753;
w44755 <= not pi0199 and not pi0294;
w44756 <= pi0199 and not pi1072;
w44757 <= not w44613 and not w44755;
w44758 <= not w44756 and w44757;
w44759 <= not w44754 and not w44758;
w44760 <= w5206 and not w44759;
w44761 <= pi0871 and w44682;
w44762 <= not pi0763 and not pi1135;
w44763 <= not pi0699 and pi1135;
w44764 <= pi1136 and not w44762;
w44765 <= not w44763 and w44764;
w44766 <= pi1134 and not w44761;
w44767 <= not w44765 and w44766;
w44768 <= pi0792 and not pi1136;
w44769 <= pi0681 and pi1136;
w44770 <= pi1135 and not w44768;
w44771 <= not w44769 and w44770;
w44772 <= not pi0809 and not pi1136;
w44773 <= pi0642 and pi1136;
w44774 <= not pi1135 and not w44772;
w44775 <= not w44773 and w44774;
w44776 <= not w44771 and not w44775;
w44777 <= not pi1134 and not w44776;
w44778 <= w44690 and not w44767;
w44779 <= not w44777 and w44778;
w44780 <= not w44760 and not w44779;
w44781 <= not pi0603 and not pi1135;
w44782 <= not pi0680 and pi1135;
w44783 <= pi1136 and not w44781;
w44784 <= not w44782 and w44783;
w44785 <= not pi0981 and not pi1135;
w44786 <= not pi0778 and pi1135;
w44787 <= not pi1136 and not w44785;
w44788 <= not w44786 and w44787;
w44789 <= not w44784 and not w44788;
w44790 <= w44637 and not w44789;
w44791 <= not pi0759 and w44649;
w44792 <= not pi0696 and pi1135;
w44793 <= not pi0837 and not pi1136;
w44794 <= not w44792 and not w44793;
w44795 <= w44655 and w44794;
w44796 <= not w44791 and w44795;
w44797 <= not w44790 and not w44796;
w44798 <= not w5206 and not w44797;
w44799 <= not pi0199 and not pi0291;
w44800 <= pi0199 and not pi1049;
w44801 <= not w44613 and not w44799;
w44802 <= not w44800 and w44801;
w44803 <= pi0414 and w44618;
w44804 <= pi0588 and not w44803;
w44805 <= pi0390 and w44664;
w44806 <= w44667 and not w44805;
w44807 <= pi0363 and not pi0591;
w44808 <= pi0592 and not w44807;
w44809 <= not w44806 and not w44808;
w44810 <= pi0342 and w44628;
w44811 <= not w44809 and not w44810;
w44812 <= w44613 and not w44804;
w44813 <= not w44811 and w44812;
w44814 <= not w44802 and not w44813;
w44815 <= w5206 and not w44814;
w44816 <= not w44798 and not w44815;
w44817 <= not pi1125 and w44452;
w44818 <= pi0669 and not w44452;
w44819 <= not pi0962 and not w44817;
w44820 <= not w44818 and w44819;
w44821 <= not pi0199 and not pi0258;
w44822 <= pi0199 and not pi1062;
w44823 <= not w44613 and not w44821;
w44824 <= not w44822 and w44823;
w44825 <= pi0415 and w44618;
w44826 <= pi0588 and not w44825;
w44827 <= pi0364 and w44621;
w44828 <= pi0391 and pi0591;
w44829 <= not pi0592 and w44828;
w44830 <= not w44827 and not w44829;
w44831 <= not pi0590 and not w44830;
w44832 <= pi0343 and w44628;
w44833 <= not pi0588 and not w44832;
w44834 <= not w44831 and w44833;
w44835 <= w44613 and not w44826;
w44836 <= not w44834 and w44835;
w44837 <= not w44824 and not w44836;
w44838 <= w5206 and not w44837;
w44839 <= pi0723 and pi1135;
w44840 <= not pi0852 and not pi1136;
w44841 <= pi0745 and w44649;
w44842 <= not w44839 and not w44840;
w44843 <= w44655 and w44842;
w44844 <= not w44841 and w44843;
w44845 <= pi0695 and pi1135;
w44846 <= pi1136 and w44636;
w44847 <= not pi0612 and not pi1135;
w44848 <= not pi1134 and not w44845;
w44849 <= not w44847 and w44848;
w44850 <= w44846 and w44849;
w44851 <= not w44844 and not w44850;
w44852 <= not w5206 and not w44851;
w44853 <= not w44838 and not w44852;
w44854 <= not pi0199 and not pi0261;
w44855 <= pi0199 and not pi1040;
w44856 <= not w44613 and not w44854;
w44857 <= not w44855 and w44856;
w44858 <= pi0453 and w44618;
w44859 <= pi0588 and not w44858;
w44860 <= pi0447 and w44621;
w44861 <= pi0333 and pi0591;
w44862 <= not pi0592 and w44861;
w44863 <= not w44860 and not w44862;
w44864 <= not pi0590 and not w44863;
w44865 <= pi0327 and w44628;
w44866 <= not pi0588 and not w44865;
w44867 <= not w44864 and w44866;
w44868 <= w44613 and not w44859;
w44869 <= not w44867 and w44868;
w44870 <= not w44857 and not w44869;
w44871 <= w5206 and not w44870;
w44872 <= pi0724 and pi1135;
w44873 <= not pi0865 and not pi1136;
w44874 <= pi0741 and w44649;
w44875 <= not w44872 and not w44873;
w44876 <= w44655 and w44875;
w44877 <= not w44874 and w44876;
w44878 <= pi0646 and pi1135;
w44879 <= not pi0611 and not pi1135;
w44880 <= not pi1134 and not w44878;
w44881 <= not w44879 and w44880;
w44882 <= w44846 and w44881;
w44883 <= not w44877 and not w44882;
w44884 <= not w5206 and not w44883;
w44885 <= not w44871 and not w44884;
w44886 <= not pi0616 and not pi1135;
w44887 <= not pi0661 and pi1135;
w44888 <= pi1136 and not w44886;
w44889 <= not w44887 and w44888;
w44890 <= not pi0808 and not pi1135;
w44891 <= not pi0781 and pi1135;
w44892 <= not pi1136 and not w44890;
w44893 <= not w44891 and w44892;
w44894 <= not w44889 and not w44893;
w44895 <= w44637 and not w44894;
w44896 <= not pi0758 and w44649;
w44897 <= not pi0736 and pi1135;
w44898 <= not pi0850 and not pi1136;
w44899 <= not w44897 and not w44898;
w44900 <= w44655 and w44899;
w44901 <= not w44896 and w44900;
w44902 <= not w44895 and not w44901;
w44903 <= not w5206 and not w44902;
w44904 <= not pi0199 and not pi0290;
w44905 <= pi0199 and not pi1048;
w44906 <= not w44613 and not w44904;
w44907 <= not w44905 and w44906;
w44908 <= pi0422 and w44618;
w44909 <= pi0588 and not w44908;
w44910 <= pi0397 and w44664;
w44911 <= w44667 and not w44910;
w44912 <= pi0372 and not pi0591;
w44913 <= pi0592 and not w44912;
w44914 <= not w44911 and not w44913;
w44915 <= pi0320 and w44628;
w44916 <= not w44914 and not w44915;
w44917 <= w44613 and not w44909;
w44918 <= not w44916 and w44917;
w44919 <= not w44907 and not w44918;
w44920 <= w5206 and not w44919;
w44921 <= not w44903 and not w44920;
w44922 <= not pi0617 and not pi1135;
w44923 <= not pi0637 and pi1135;
w44924 <= pi1136 and not w44922;
w44925 <= not w44923 and w44924;
w44926 <= not pi0788 and pi1135;
w44927 <= pi0814 and not pi1135;
w44928 <= not pi1136 and not w44926;
w44929 <= not w44927 and w44928;
w44930 <= not w44925 and not w44929;
w44931 <= w44637 and not w44930;
w44932 <= not pi0749 and w44649;
w44933 <= not pi0706 and pi1135;
w44934 <= not pi0866 and not pi1136;
w44935 <= not w44933 and not w44934;
w44936 <= w44655 and w44935;
w44937 <= not w44932 and w44936;
w44938 <= not w44931 and not w44937;
w44939 <= not w5206 and not w44938;
w44940 <= not pi0199 and not pi0295;
w44941 <= pi0199 and not pi1053;
w44942 <= not w44613 and not w44940;
w44943 <= not w44941 and w44942;
w44944 <= pi0435 and w44618;
w44945 <= pi0588 and not w44944;
w44946 <= pi0411 and w44664;
w44947 <= w44667 and not w44946;
w44948 <= pi0387 and not pi0591;
w44949 <= pi0592 and not w44948;
w44950 <= not w44947 and not w44949;
w44951 <= pi0452 and w44628;
w44952 <= not w44950 and not w44951;
w44953 <= w44613 and not w44945;
w44954 <= not w44952 and w44953;
w44955 <= not w44943 and not w44954;
w44956 <= w5206 and not w44955;
w44957 <= not w44939 and not w44956;
w44958 <= not pi0199 and not pi0256;
w44959 <= pi0199 and not pi1070;
w44960 <= not w44613 and not w44958;
w44961 <= not w44959 and w44960;
w44962 <= pi0437 and w44618;
w44963 <= pi0588 and not w44962;
w44964 <= pi0336 and w44621;
w44965 <= pi0463 and pi0591;
w44966 <= not pi0592 and w44965;
w44967 <= not w44964 and not w44966;
w44968 <= not pi0590 and not w44967;
w44969 <= pi0362 and w44628;
w44970 <= not pi0588 and not w44969;
w44971 <= not w44968 and w44970;
w44972 <= w44613 and not w44963;
w44973 <= not w44971 and w44972;
w44974 <= not w44961 and not w44973;
w44975 <= w5206 and not w44974;
w44976 <= pi0859 and w44682;
w44977 <= not pi0743 and not pi1135;
w44978 <= not pi0735 and pi1135;
w44979 <= pi1136 and not w44977;
w44980 <= not w44978 and w44979;
w44981 <= pi1134 and not w44976;
w44982 <= not w44980 and w44981;
w44983 <= pi0622 and not pi1135;
w44984 <= pi0639 and pi1135;
w44985 <= pi1136 and not w44983;
w44986 <= not w44984 and w44985;
w44987 <= pi0804 and not pi1135;
w44988 <= pi0783 and pi1135;
w44989 <= not pi1136 and not w44987;
w44990 <= not w44988 and w44989;
w44991 <= not w44986 and not w44990;
w44992 <= not pi1134 and not w44991;
w44993 <= w44690 and not w44982;
w44994 <= not w44992 and w44993;
w44995 <= not w44975 and not w44994;
w44996 <= pi0876 and w44682;
w44997 <= not pi0748 and not pi1135;
w44998 <= not pi0730 and pi1135;
w44999 <= pi1136 and not w44997;
w45000 <= not w44998 and w44999;
w45001 <= not w44996 and not w45000;
w45002 <= w44654 and not w45001;
w45003 <= not pi0623 and w44649;
w45004 <= pi0789 and w44653;
w45005 <= not pi0710 and pi1135;
w45006 <= pi1136 and not w45005;
w45007 <= not pi0803 and not pi1135;
w45008 <= not w45004 and not w45007;
w45009 <= not w45006 and w45008;
w45010 <= w44637 and not w45003;
w45011 <= not w45009 and w45010;
w45012 <= not w45002 and not w45011;
w45013 <= not w5206 and not w45012;
w45014 <= not pi0199 and not pi0296;
w45015 <= pi0199 and not pi1037;
w45016 <= not w44613 and not w45014;
w45017 <= not w45015 and w45016;
w45018 <= pi0436 and w44618;
w45019 <= pi0588 and not w45018;
w45020 <= pi0412 and w44664;
w45021 <= w44667 and not w45020;
w45022 <= pi0388 and not pi0591;
w45023 <= pi0592 and not w45022;
w45024 <= not w45021 and not w45023;
w45025 <= pi0455 and w44628;
w45026 <= not w45024 and not w45025;
w45027 <= w44613 and not w45019;
w45028 <= not w45026 and w45027;
w45029 <= not w45017 and not w45028;
w45030 <= w5206 and not w45029;
w45031 <= not w45013 and not w45030;
w45032 <= not pi0606 and not pi1135;
w45033 <= not pi0643 and pi1135;
w45034 <= pi1136 and not w45032;
w45035 <= not w45033 and w45034;
w45036 <= not pi0787 and pi1135;
w45037 <= pi0812 and not pi1135;
w45038 <= not pi1136 and not w45036;
w45039 <= not w45037 and w45038;
w45040 <= not w45035 and not w45039;
w45041 <= w44637 and not w45040;
w45042 <= not pi0746 and w44649;
w45043 <= not pi0729 and pi1135;
w45044 <= not pi0881 and not pi1136;
w45045 <= not w45043 and not w45044;
w45046 <= w44655 and w45045;
w45047 <= not w45042 and w45046;
w45048 <= not w45041 and not w45047;
w45049 <= not w5206 and not w45048;
w45050 <= not pi0199 and not pi0293;
w45051 <= pi0199 and not pi1059;
w45052 <= not w44613 and not w45050;
w45053 <= not w45051 and w45052;
w45054 <= pi0434 and w44618;
w45055 <= pi0588 and not w45054;
w45056 <= pi0410 and w44664;
w45057 <= w44667 and not w45056;
w45058 <= pi0386 and not pi0591;
w45059 <= pi0592 and not w45058;
w45060 <= not w45057 and not w45059;
w45061 <= pi0361 and w44628;
w45062 <= not w45060 and not w45061;
w45063 <= w44613 and not w45055;
w45064 <= not w45062 and w45063;
w45065 <= not w45053 and not w45064;
w45066 <= w5206 and not w45065;
w45067 <= not w45049 and not w45066;
w45068 <= not pi0199 and not pi0259;
w45069 <= pi0199 and not pi1069;
w45070 <= not w44613 and not w45068;
w45071 <= not w45069 and w45070;
w45072 <= pi0416 and w44618;
w45073 <= pi0588 and not w45072;
w45074 <= pi0366 and w44621;
w45075 <= pi0335 and pi0591;
w45076 <= not pi0592 and w45075;
w45077 <= not w45074 and not w45076;
w45078 <= not pi0590 and not w45077;
w45079 <= pi0344 and w44628;
w45080 <= not pi0588 and not w45079;
w45081 <= not w45078 and w45080;
w45082 <= w44613 and not w45073;
w45083 <= not w45081 and w45082;
w45084 <= not w45071 and not w45083;
w45085 <= w5206 and not w45084;
w45086 <= pi0704 and pi1135;
w45087 <= not pi0870 and not pi1136;
w45088 <= pi0742 and w44649;
w45089 <= not w45086 and not w45087;
w45090 <= w44655 and w45089;
w45091 <= not w45088 and w45090;
w45092 <= pi0635 and pi1135;
w45093 <= not pi0620 and not pi1135;
w45094 <= not pi1134 and not w45092;
w45095 <= not w45093 and w45094;
w45096 <= w44846 and w45095;
w45097 <= not w45091 and not w45096;
w45098 <= not w5206 and not w45097;
w45099 <= not w45085 and not w45098;
w45100 <= not pi0199 and not pi0260;
w45101 <= pi0199 and not pi1067;
w45102 <= not w44613 and not w45100;
w45103 <= not w45101 and w45102;
w45104 <= pi0418 and w44618;
w45105 <= pi0588 and not w45104;
w45106 <= pi0368 and w44621;
w45107 <= pi0393 and pi0591;
w45108 <= not pi0592 and w45107;
w45109 <= not w45106 and not w45108;
w45110 <= not pi0590 and not w45109;
w45111 <= pi0346 and w44628;
w45112 <= not pi0588 and not w45111;
w45113 <= not w45110 and w45112;
w45114 <= w44613 and not w45105;
w45115 <= not w45113 and w45114;
w45116 <= not w45103 and not w45115;
w45117 <= w5206 and not w45116;
w45118 <= pi0688 and pi1135;
w45119 <= not pi0856 and not pi1136;
w45120 <= pi0760 and w44649;
w45121 <= not w45118 and not w45119;
w45122 <= w44655 and w45121;
w45123 <= not w45120 and w45122;
w45124 <= pi0632 and pi1135;
w45125 <= not pi0613 and not pi1135;
w45126 <= not pi1134 and not w45124;
w45127 <= not w45125 and w45126;
w45128 <= w44846 and w45127;
w45129 <= not w45123 and not w45128;
w45130 <= not w5206 and not w45129;
w45131 <= not w45117 and not w45130;
w45132 <= not pi0199 and not pi0255;
w45133 <= pi0199 and not pi1036;
w45134 <= not w44613 and not w45132;
w45135 <= not w45133 and w45134;
w45136 <= pi0438 and w44618;
w45137 <= pi0588 and not w45136;
w45138 <= pi0389 and w44621;
w45139 <= pi0413 and pi0591;
w45140 <= not pi0592 and w45139;
w45141 <= not w45138 and not w45140;
w45142 <= not pi0590 and not w45141;
w45143 <= pi0450 and w44628;
w45144 <= not pi0588 and not w45143;
w45145 <= not w45142 and w45144;
w45146 <= w44613 and not w45137;
w45147 <= not w45145 and w45146;
w45148 <= not w45135 and not w45147;
w45149 <= w5206 and not w45148;
w45150 <= not pi0791 and not pi1136;
w45151 <= not pi0665 and pi1136;
w45152 <= pi1135 and not w45150;
w45153 <= not w45151 and w45152;
w45154 <= not pi0810 and not pi1136;
w45155 <= not pi0621 and pi1136;
w45156 <= not pi1135 and not w45154;
w45157 <= not w45155 and w45156;
w45158 <= not w45153 and not w45157;
w45159 <= w44637 and not w45158;
w45160 <= not pi0739 and w44649;
w45161 <= not pi0874 and not pi1136;
w45162 <= not pi0690 and pi1135;
w45163 <= not w45161 and not w45162;
w45164 <= w44655 and w45163;
w45165 <= not w45160 and w45164;
w45166 <= not w45159 and not w45165;
w45167 <= not w5206 and not w45166;
w45168 <= not w45149 and not w45167;
w45169 <= not pi0680 and not w44452;
w45170 <= not pi1100 and w44452;
w45171 <= not pi0962 and not w45169;
w45172 <= not w45170 and w45171;
w45173 <= not pi0681 and not w44452;
w45174 <= not pi1103 and w44452;
w45175 <= not pi0962 and not w45173;
w45176 <= not w45174 and w45175;
w45177 <= not pi0199 and not pi0251;
w45178 <= pi0199 and not pi1039;
w45179 <= not w44613 and not w45177;
w45180 <= not w45178 and w45179;
w45181 <= pi0417 and w44618;
w45182 <= pi0588 and not w45181;
w45183 <= pi0367 and w44621;
w45184 <= pi0392 and pi0591;
w45185 <= not pi0592 and w45184;
w45186 <= not w45183 and not w45185;
w45187 <= not pi0590 and not w45186;
w45188 <= pi0345 and w44628;
w45189 <= not pi0588 and not w45188;
w45190 <= not w45187 and w45189;
w45191 <= w44613 and not w45182;
w45192 <= not w45190 and w45191;
w45193 <= not w45180 and not w45192;
w45194 <= w5206 and not w45193;
w45195 <= pi0686 and pi1135;
w45196 <= not pi0848 and not pi1136;
w45197 <= pi0757 and w44649;
w45198 <= not w45195 and not w45196;
w45199 <= w44655 and w45198;
w45200 <= not w45197 and w45199;
w45201 <= pi0631 and pi1135;
w45202 <= not pi0610 and not pi1135;
w45203 <= not pi1134 and not w45201;
w45204 <= not w45202 and w45203;
w45205 <= w44846 and w45204;
w45206 <= not w45200 and not w45205;
w45207 <= not w5206 and not w45206;
w45208 <= not w45194 and not w45207;
w45209 <= pi0953 and w44451;
w45210 <= not pi1130 and w45209;
w45211 <= pi0684 and not w45209;
w45212 <= not pi0962 and not w45210;
w45213 <= not w45211 and w45212;
w45214 <= pi0590 and not pi0592;
w45215 <= pi0357 and w45214;
w45216 <= pi0382 and w44666;
w45217 <= not w45215 and not w45216;
w45218 <= not pi0591 and not w45217;
w45219 <= pi0406 and not pi0592;
w45220 <= w44664 and w45219;
w45221 <= not w45218 and not w45220;
w45222 <= not pi0588 and not w45221;
w45223 <= not pi0591 and not pi0592;
w45224 <= pi0588 and not pi0590;
w45225 <= pi0430 and w45223;
w45226 <= w45224 and w45225;
w45227 <= not w45222 and not w45226;
w45228 <= w44613 and not w45227;
w45229 <= pi0199 and not pi1076;
w45230 <= not w44613 and not w45229;
w45231 <= not w40443 and w45230;
w45232 <= not w45228 and not w45231;
w45233 <= w5206 and not w45232;
w45234 <= pi0860 and w44682;
w45235 <= pi0744 and not pi1135;
w45236 <= pi0728 and pi1135;
w45237 <= pi1136 and not w45235;
w45238 <= not w45236 and w45237;
w45239 <= not w45234 and not w45238;
w45240 <= w44654 and not w45239;
w45241 <= pi1136 and not w44636;
w45242 <= not pi1134 and not w45241;
w45243 <= not pi0652 and not pi1135;
w45244 <= pi0657 and pi1135;
w45245 <= pi1136 and not w45243;
w45246 <= not w45244 and w45245;
w45247 <= pi0813 and w44636;
w45248 <= w44682 and w45247;
w45249 <= not w45246 and not w45248;
w45250 <= w45242 and not w45249;
w45251 <= not w45240 and not w45250;
w45252 <= not w5206 and not w45251;
w45253 <= not w45233 and not w45252;
w45254 <= not pi1113 and w45209;
w45255 <= pi0686 and not w45209;
w45256 <= not pi0962 and not w45254;
w45257 <= not w45255 and w45256;
w45258 <= not pi0687 and not w45209;
w45259 <= not pi1127 and w45209;
w45260 <= not pi0962 and not w45258;
w45261 <= not w45259 and w45260;
w45262 <= not pi1115 and w45209;
w45263 <= pi0688 and not w45209;
w45264 <= not pi0962 and not w45262;
w45265 <= not w45263 and w45264;
w45266 <= pi0351 and w45214;
w45267 <= pi0376 and w44666;
w45268 <= not w45266 and not w45267;
w45269 <= not pi0591 and not w45268;
w45270 <= pi0401 and not pi0592;
w45271 <= w44664 and w45270;
w45272 <= not w45269 and not w45271;
w45273 <= not pi0588 and not w45272;
w45274 <= pi0426 and w45223;
w45275 <= w45224 and w45274;
w45276 <= not w45273 and not w45275;
w45277 <= w44613 and not w45276;
w45278 <= pi0199 and not pi1079;
w45279 <= not pi0199 and w40412;
w45280 <= not w44613 and not w45278;
w45281 <= not w45279 and w45280;
w45282 <= not w45277 and not w45281;
w45283 <= w5206 and not w45282;
w45284 <= pi0798 and w44682;
w45285 <= not pi0658 and not pi1135;
w45286 <= pi0655 and pi1135;
w45287 <= pi1136 and not w45285;
w45288 <= not w45286 and w45287;
w45289 <= not w45284 and not w45288;
w45290 <= w44637 and not w45289;
w45291 <= pi0752 and w44649;
w45292 <= not pi0703 and pi1135;
w45293 <= not pi0843 and not pi1136;
w45294 <= not w45292 and not w45293;
w45295 <= w44655 and w45294;
w45296 <= not w45291 and w45295;
w45297 <= not w45290 and not w45296;
w45298 <= not w5206 and not w45297;
w45299 <= not w45283 and not w45298;
w45300 <= not pi0690 and not w45209;
w45301 <= not pi1108 and w45209;
w45302 <= not pi0962 and not w45300;
w45303 <= not w45301 and w45302;
w45304 <= not pi0691 and not w45209;
w45305 <= not pi1107 and w45209;
w45306 <= not pi0962 and not w45304;
w45307 <= not w45305 and w45306;
w45308 <= pi0352 and w45214;
w45309 <= pi0317 and w44666;
w45310 <= not w45308 and not w45309;
w45311 <= not pi0591 and not w45310;
w45312 <= pi0402 and not pi0592;
w45313 <= w44664 and w45312;
w45314 <= not w45311 and not w45313;
w45315 <= not pi0588 and not w45314;
w45316 <= pi0427 and w45223;
w45317 <= w45224 and w45316;
w45318 <= not w45315 and not w45317;
w45319 <= w44613 and not w45318;
w45320 <= pi0199 and not pi1078;
w45321 <= not pi0199 and w40424;
w45322 <= not w44613 and not w45320;
w45323 <= not w45321 and w45322;
w45324 <= not w45319 and not w45323;
w45325 <= w5206 and not w45324;
w45326 <= pi0844 and w44682;
w45327 <= not pi0726 and pi1135;
w45328 <= pi0770 and not pi1135;
w45329 <= pi1136 and not w45327;
w45330 <= not w45328 and w45329;
w45331 <= pi1134 and not w45326;
w45332 <= not w45330 and w45331;
w45333 <= pi0801 and w44682;
w45334 <= not pi0656 and not pi1135;
w45335 <= pi0649 and pi1135;
w45336 <= pi1136 and not w45334;
w45337 <= not w45335 and w45336;
w45338 <= not pi1134 and not w45333;
w45339 <= not w45337 and w45338;
w45340 <= w44690 and not w45332;
w45341 <= not w45339 and w45340;
w45342 <= not w45325 and not w45341;
w45343 <= not pi1129 and w44452;
w45344 <= pi0693 and not w44452;
w45345 <= not pi0962 and not w45343;
w45346 <= not w45344 and w45345;
w45347 <= not pi1128 and w45209;
w45348 <= pi0694 and not w45209;
w45349 <= not pi0962 and not w45347;
w45350 <= not w45348 and w45349;
w45351 <= not pi1111 and w44452;
w45352 <= pi0695 and not w44452;
w45353 <= not pi0962 and not w45351;
w45354 <= not w45352 and w45353;
w45355 <= not pi0696 and not w45209;
w45356 <= not pi1100 and w45209;
w45357 <= not pi0962 and not w45355;
w45358 <= not w45356 and w45357;
w45359 <= not pi1129 and w45209;
w45360 <= pi0697 and not w45209;
w45361 <= not pi0962 and not w45359;
w45362 <= not w45360 and w45361;
w45363 <= not pi1116 and w45209;
w45364 <= pi0698 and not w45209;
w45365 <= not pi0962 and not w45363;
w45366 <= not w45364 and w45365;
w45367 <= not pi0699 and not w45209;
w45368 <= not pi1103 and w45209;
w45369 <= not pi0962 and not w45367;
w45370 <= not w45368 and w45369;
w45371 <= not pi0700 and not w45209;
w45372 <= not pi1110 and w45209;
w45373 <= not pi0962 and not w45371;
w45374 <= not w45372 and w45373;
w45375 <= not pi1123 and w45209;
w45376 <= pi0701 and not w45209;
w45377 <= not pi0962 and not w45375;
w45378 <= not w45376 and w45377;
w45379 <= not pi1117 and w45209;
w45380 <= pi0702 and not w45209;
w45381 <= not pi0962 and not w45379;
w45382 <= not w45380 and w45381;
w45383 <= not pi0703 and not w45209;
w45384 <= not pi1124 and w45209;
w45385 <= not pi0962 and not w45383;
w45386 <= not w45384 and w45385;
w45387 <= not pi1112 and w45209;
w45388 <= pi0704 and not w45209;
w45389 <= not pi0962 and not w45387;
w45390 <= not w45388 and w45389;
w45391 <= not pi0705 and not w45209;
w45392 <= not pi1125 and w45209;
w45393 <= not pi0962 and not w45391;
w45394 <= not w45392 and w45393;
w45395 <= not pi0706 and not w45209;
w45396 <= not pi1105 and w45209;
w45397 <= not pi0962 and not w45395;
w45398 <= not w45396 and w45397;
w45399 <= pi0370 and w44621;
w45400 <= pi0395 and pi0591;
w45401 <= not pi0592 and w45400;
w45402 <= not w45399 and not w45401;
w45403 <= not pi0590 and not w45402;
w45404 <= pi0347 and w44628;
w45405 <= not w45403 and not w45404;
w45406 <= not pi0588 and w44613;
w45407 <= not w45405 and w45406;
w45408 <= pi0199 and not pi1055;
w45409 <= not pi0200 and not pi0304;
w45410 <= pi0200 and not pi1048;
w45411 <= not w45409 and not w45410;
w45412 <= not pi0199 and not w45411;
w45413 <= not w44613 and not w45408;
w45414 <= not w45412 and w45413;
w45415 <= w44613 and w44618;
w45416 <= pi0420 and pi0588;
w45417 <= w45415 and w45416;
w45418 <= not w45414 and not w45417;
w45419 <= not w45407 and w45418;
w45420 <= w5206 and not w45419;
w45421 <= not pi0627 and pi1135;
w45422 <= not pi0618 and not pi1135;
w45423 <= not pi1134 and not w45421;
w45424 <= not w45422 and w45423;
w45425 <= w44846 and w45424;
w45426 <= pi0702 and pi1135;
w45427 <= not pi0847 and not pi1136;
w45428 <= pi0753 and w44649;
w45429 <= not w45426 and not w45427;
w45430 <= w44655 and w45429;
w45431 <= not w45428 and w45430;
w45432 <= not w45425 and not w45431;
w45433 <= not w5206 and not w45432;
w45434 <= not w45420 and not w45433;
w45435 <= w44613 and w45223;
w45436 <= pi0459 and w45224;
w45437 <= w45435 and w45436;
w45438 <= w44613 and w44621;
w45439 <= pi0442 and w45438;
w45440 <= not pi0592 and w44613;
w45441 <= pi0328 and pi0591;
w45442 <= w45440 and w45441;
w45443 <= not w45439 and not w45442;
w45444 <= not pi0590 and not w45443;
w45445 <= pi0321 and w44613;
w45446 <= w44628 and w45445;
w45447 <= not w45444 and not w45446;
w45448 <= not pi0588 and not w45447;
w45449 <= pi0199 and not pi1058;
w45450 <= not pi0200 and not pi0305;
w45451 <= pi0200 and not pi1084;
w45452 <= not w45450 and not w45451;
w45453 <= not pi0199 and not w45452;
w45454 <= not w44613 and not w45449;
w45455 <= not w45453 and w45454;
w45456 <= w5206 and not w45437;
w45457 <= not w45455 and w45456;
w45458 <= not w45448 and w45457;
w45459 <= not pi0609 and not pi1135;
w45460 <= not pi0660 and pi1135;
w45461 <= not pi1134 and not w45459;
w45462 <= not w45460 and w45461;
w45463 <= w44846 and w45462;
w45464 <= w44636 and not w44653;
w45465 <= pi0709 and pi1135;
w45466 <= not pi0857 and not pi1136;
w45467 <= pi0754 and w44649;
w45468 <= pi1134 and not w45465;
w45469 <= not w45466 and w45468;
w45470 <= w45464 and w45469;
w45471 <= not w45467 and w45470;
w45472 <= not w5206 and not w45463;
w45473 <= not w45471 and w45472;
w45474 <= not w45458 and not w45473;
w45475 <= not pi1118 and w45209;
w45476 <= pi0709 and not w45209;
w45477 <= not pi0962 and not w45475;
w45478 <= not w45476 and w45477;
w45479 <= not pi0710 and not w44452;
w45480 <= not pi1106 and w44452;
w45481 <= not pi0962 and not w45479;
w45482 <= not w45480 and w45481;
w45483 <= pi0373 and w44621;
w45484 <= pi0398 and pi0591;
w45485 <= not pi0592 and w45484;
w45486 <= not w45483 and not w45485;
w45487 <= not pi0590 and not w45486;
w45488 <= pi0348 and w44628;
w45489 <= not w45487 and not w45488;
w45490 <= w45406 and not w45489;
w45491 <= pi0199 and not pi1087;
w45492 <= not pi0200 and not pi0306;
w45493 <= pi0200 and not pi1059;
w45494 <= not w45492 and not w45493;
w45495 <= not pi0199 and not w45494;
w45496 <= not w44613 and not w45491;
w45497 <= not w45495 and w45496;
w45498 <= pi0423 and pi0588;
w45499 <= w45415 and w45498;
w45500 <= not w45497 and not w45499;
w45501 <= not w45490 and w45500;
w45502 <= w5206 and not w45501;
w45503 <= not pi0647 and pi1135;
w45504 <= not pi0630 and not pi1135;
w45505 <= not pi1134 and not w45503;
w45506 <= not w45504 and w45505;
w45507 <= w44846 and w45506;
w45508 <= pi0725 and pi1135;
w45509 <= not pi0858 and not pi1136;
w45510 <= pi0755 and w44649;
w45511 <= not w45508 and not w45509;
w45512 <= w44655 and w45511;
w45513 <= not w45510 and w45512;
w45514 <= not w45507 and not w45513;
w45515 <= not w5206 and not w45514;
w45516 <= not w45502 and not w45515;
w45517 <= pi0701 and pi1135;
w45518 <= not pi0842 and not pi1136;
w45519 <= pi0751 and w44649;
w45520 <= pi1134 and not w45517;
w45521 <= not w45518 and w45520;
w45522 <= w45464 and w45521;
w45523 <= not w45519 and w45522;
w45524 <= not pi0715 and pi1135;
w45525 <= not pi0644 and not pi1135;
w45526 <= not pi1134 and not w45524;
w45527 <= not w45525 and w45526;
w45528 <= w44846 and w45527;
w45529 <= not w45523 and not w45528;
w45530 <= not w5206 and not w45529;
w45531 <= pi0199 and pi1035;
w45532 <= pi0298 and w8372;
w45533 <= pi1044 and w9007;
w45534 <= not w44613 and not w45531;
w45535 <= not w45532 and w45534;
w45536 <= not w45533 and w45535;
w45537 <= pi0425 and w45223;
w45538 <= w45224 and w45537;
w45539 <= pi0374 and w44621;
w45540 <= pi0400 and pi0591;
w45541 <= not pi0592 and w45540;
w45542 <= not w45539 and not w45541;
w45543 <= not pi0590 and not w45542;
w45544 <= pi0350 and w44628;
w45545 <= not w45543 and not w45544;
w45546 <= not pi0588 and not w45545;
w45547 <= w44613 and not w45538;
w45548 <= not w45546 and w45547;
w45549 <= w5206 and not w45536;
w45550 <= not w45548 and w45549;
w45551 <= not w45530 and not w45550;
w45552 <= pi0371 and w44621;
w45553 <= pi0396 and pi0591;
w45554 <= not pi0592 and w45553;
w45555 <= not w45552 and not w45554;
w45556 <= not pi0590 and not w45555;
w45557 <= pi0322 and w44628;
w45558 <= not w45556 and not w45557;
w45559 <= w45406 and not w45558;
w45560 <= pi0199 and not pi1051;
w45561 <= not pi0200 and not pi0309;
w45562 <= pi0200 and not pi1072;
w45563 <= not w45561 and not w45562;
w45564 <= not pi0199 and not w45563;
w45565 <= not w44613 and not w45560;
w45566 <= not w45564 and w45565;
w45567 <= pi0421 and pi0588;
w45568 <= w45415 and w45567;
w45569 <= not w45566 and not w45568;
w45570 <= not w45559 and w45569;
w45571 <= w5206 and not w45570;
w45572 <= not pi0628 and pi1135;
w45573 <= not pi0629 and not pi1135;
w45574 <= not pi1134 and not w45572;
w45575 <= not w45573 and w45574;
w45576 <= w44846 and w45575;
w45577 <= pi0734 and pi1135;
w45578 <= not pi0854 and not pi1136;
w45579 <= pi0756 and w44649;
w45580 <= not w45577 and not w45578;
w45581 <= w44655 and w45580;
w45582 <= not w45579 and w45581;
w45583 <= not w45576 and not w45582;
w45584 <= not w5206 and not w45583;
w45585 <= not w45571 and not w45584;
w45586 <= pi0461 and w45214;
w45587 <= pi0439 and w44666;
w45588 <= not w45586 and not w45587;
w45589 <= not pi0591 and not w45588;
w45590 <= pi0326 and not pi0592;
w45591 <= w44664 and w45590;
w45592 <= not w45589 and not w45591;
w45593 <= not pi0588 and not w45592;
w45594 <= pi0449 and w45223;
w45595 <= w45224 and w45594;
w45596 <= not w45593 and not w45595;
w45597 <= w44613 and not w45596;
w45598 <= pi0199 and not pi1057;
w45599 <= not w44613 and not w45598;
w45600 <= not w39902 and w45599;
w45601 <= not w45597 and not w45600;
w45602 <= w5206 and not w45601;
w45603 <= pi0867 and w44682;
w45604 <= pi0762 and not pi1135;
w45605 <= pi0697 and pi1135;
w45606 <= pi1136 and not w45604;
w45607 <= not w45605 and w45606;
w45608 <= not w45603 and not w45607;
w45609 <= w44654 and not w45608;
w45610 <= not pi0653 and not pi1135;
w45611 <= pi0693 and pi1135;
w45612 <= pi1136 and not w45610;
w45613 <= not w45611 and w45612;
w45614 <= pi0816 and w44636;
w45615 <= w44682 and w45614;
w45616 <= not w45613 and not w45615;
w45617 <= w45242 and not w45616;
w45618 <= not w45609 and not w45617;
w45619 <= not w5206 and not w45618;
w45620 <= not w45602 and not w45619;
w45621 <= not pi0715 and not w44452;
w45622 <= not pi1123 and w44452;
w45623 <= not pi0962 and not w45621;
w45624 <= not w45622 and w45623;
w45625 <= pi0454 and w45224;
w45626 <= w45435 and w45625;
w45627 <= pi0440 and w45438;
w45628 <= pi0329 and pi0591;
w45629 <= w45440 and w45628;
w45630 <= not w45627 and not w45629;
w45631 <= not pi0590 and not w45630;
w45632 <= pi0349 and w44613;
w45633 <= w44628 and w45632;
w45634 <= not w45631 and not w45633;
w45635 <= not pi0588 and not w45634;
w45636 <= pi0199 and not pi1043;
w45637 <= not pi0200 and not pi0307;
w45638 <= pi0200 and not pi1053;
w45639 <= not w45637 and not w45638;
w45640 <= not pi0199 and not w45639;
w45641 <= not w44613 and not w45636;
w45642 <= not w45640 and w45641;
w45643 <= w5206 and not w45626;
w45644 <= not w45642 and w45643;
w45645 <= not w45635 and w45644;
w45646 <= not pi0626 and not pi1135;
w45647 <= not pi0641 and pi1135;
w45648 <= not pi1134 and not w45646;
w45649 <= not w45647 and w45648;
w45650 <= w44846 and w45649;
w45651 <= pi0738 and pi1135;
w45652 <= not pi0845 and not pi1136;
w45653 <= pi0761 and w44649;
w45654 <= pi1134 and not w45651;
w45655 <= not w45652 and w45654;
w45656 <= w45464 and w45655;
w45657 <= not w45653 and w45656;
w45658 <= not w5206 and not w45650;
w45659 <= not w45657 and w45658;
w45660 <= not w45645 and not w45659;
w45661 <= pi0318 and pi0591;
w45662 <= not pi0592 and w45661;
w45663 <= not pi0591 and w6031;
w45664 <= not w45662 and not w45663;
w45665 <= not pi0590 and not w45664;
w45666 <= pi0462 and w44628;
w45667 <= not w45665 and not w45666;
w45668 <= w45406 and not w45667;
w45669 <= pi0199 and not pi1074;
w45670 <= not pi0199 and w40418;
w45671 <= not w44613 and not w45669;
w45672 <= not w45670 and w45671;
w45673 <= pi0448 and pi0588;
w45674 <= w45415 and w45673;
w45675 <= not w45672 and not w45674;
w45676 <= not w45668 and w45675;
w45677 <= w5206 and not w45676;
w45678 <= not pi0705 and pi1135;
w45679 <= pi0768 and w44649;
w45680 <= not pi0839 and not pi1136;
w45681 <= pi1134 and not w45678;
w45682 <= not w45680 and w45681;
w45683 <= w45464 and w45682;
w45684 <= not w45679 and w45683;
w45685 <= pi0800 and w44682;
w45686 <= not pi0645 and not pi1135;
w45687 <= pi0669 and pi1135;
w45688 <= pi1136 and not w45686;
w45689 <= not w45687 and w45688;
w45690 <= not w45685 and not w45689;
w45691 <= w44637 and not w45690;
w45692 <= not w45684 and not w45691;
w45693 <= not w5206 and not w45692;
w45694 <= not w45677 and not w45693;
w45695 <= pi0419 and w45224;
w45696 <= w45435 and w45695;
w45697 <= pi0369 and w45438;
w45698 <= pi0394 and pi0591;
w45699 <= w45440 and w45698;
w45700 <= not w45697 and not w45699;
w45701 <= not pi0590 and not w45700;
w45702 <= pi0315 and w44613;
w45703 <= w44628 and w45702;
w45704 <= not w45701 and not w45703;
w45705 <= not pi0588 and not w45704;
w45706 <= pi0199 and not pi1080;
w45707 <= not pi0200 and not pi0303;
w45708 <= pi0200 and not pi1049;
w45709 <= not w45707 and not w45708;
w45710 <= not pi0199 and not w45709;
w45711 <= not w44613 and not w45706;
w45712 <= not w45710 and w45711;
w45713 <= w5206 and not w45696;
w45714 <= not w45712 and w45713;
w45715 <= not w45705 and w45714;
w45716 <= not pi0608 and not pi1135;
w45717 <= not pi0625 and pi1135;
w45718 <= not pi1134 and not w45716;
w45719 <= not w45717 and w45718;
w45720 <= w44846 and w45719;
w45721 <= pi0698 and pi1135;
w45722 <= not pi0853 and not pi1136;
w45723 <= pi0767 and w44649;
w45724 <= pi1134 and not w45721;
w45725 <= not w45722 and w45724;
w45726 <= w45464 and w45725;
w45727 <= not w45723 and w45726;
w45728 <= not w5206 and not w45720;
w45729 <= not w45727 and w45728;
w45730 <= not w45715 and not w45729;
w45731 <= pi0378 and w44621;
w45732 <= pi0325 and pi0591;
w45733 <= not pi0592 and w45732;
w45734 <= not w45731 and not w45733;
w45735 <= not pi0590 and not w45734;
w45736 <= pi0353 and w44628;
w45737 <= not w45735 and not w45736;
w45738 <= w45406 and not w45737;
w45739 <= pi0199 and not pi1063;
w45740 <= not pi0199 and w40430;
w45741 <= not w44613 and not w45739;
w45742 <= not w45740 and w45741;
w45743 <= pi0451 and pi0588;
w45744 <= w45415 and w45743;
w45745 <= not w45742 and not w45744;
w45746 <= not w45738 and w45745;
w45747 <= w5206 and not w45746;
w45748 <= not pi0687 and pi1135;
w45749 <= pi0774 and w44649;
w45750 <= not pi0868 and not pi1136;
w45751 <= pi1134 and not w45748;
w45752 <= not w45750 and w45751;
w45753 <= w45464 and w45752;
w45754 <= not w45749 and w45753;
w45755 <= pi0807 and w44682;
w45756 <= not pi0636 and not pi1135;
w45757 <= pi0650 and pi1135;
w45758 <= pi1136 and not w45756;
w45759 <= not w45757 and w45758;
w45760 <= not w45755 and not w45759;
w45761 <= w44637 and not w45760;
w45762 <= not w45754 and not w45761;
w45763 <= not w5206 and not w45762;
w45764 <= not w45747 and not w45763;
w45765 <= pi0356 and w45214;
w45766 <= pi0381 and w44666;
w45767 <= not w45765 and not w45766;
w45768 <= not pi0591 and not w45767;
w45769 <= pi0405 and not pi0592;
w45770 <= w44664 and w45769;
w45771 <= not w45768 and not w45770;
w45772 <= not pi0588 and not w45771;
w45773 <= pi0445 and w45223;
w45774 <= w45224 and w45773;
w45775 <= not w45772 and not w45774;
w45776 <= w44613 and not w45775;
w45777 <= pi0199 and not pi1081;
w45778 <= not w44613 and not w45777;
w45779 <= not w40450 and w45778;
w45780 <= not w45776 and not w45779;
w45781 <= w5206 and not w45780;
w45782 <= pi0880 and w44682;
w45783 <= pi0750 and not pi1135;
w45784 <= pi0684 and pi1135;
w45785 <= pi1136 and not w45783;
w45786 <= not w45784 and w45785;
w45787 <= not w45782 and not w45786;
w45788 <= w44654 and not w45787;
w45789 <= not pi0651 and not pi1135;
w45790 <= pi0654 and pi1135;
w45791 <= pi1136 and not w45789;
w45792 <= not w45790 and w45791;
w45793 <= pi0794 and w44636;
w45794 <= w44682 and w45793;
w45795 <= not w45792 and not w45794;
w45796 <= w45242 and not w45795;
w45797 <= not w45788 and not w45796;
w45798 <= not w5206 and not w45797;
w45799 <= not w45781 and not w45798;
w45800 <= pi0721 and not pi0775;
w45801 <= pi0721 and pi0813;
w45802 <= not pi0773 and not pi0801;
w45803 <= pi0773 and pi0801;
w45804 <= not w45802 and not w45803;
w45805 <= not pi0771 and not pi0800;
w45806 <= pi0771 and pi0800;
w45807 <= not w45805 and not w45806;
w45808 <= not pi0769 and not pi0794;
w45809 <= pi0769 and pi0794;
w45810 <= not w45808 and not w45809;
w45811 <= not pi0765 and not pi0798;
w45812 <= pi0765 and pi0798;
w45813 <= not w45811 and not w45812;
w45814 <= pi0807 and not w45813;
w45815 <= pi0747 and w45814;
w45816 <= not pi0747 and not pi0807;
w45817 <= not w45813 and w45816;
w45818 <= not w45815 and not w45817;
w45819 <= not w45810 and not w45818;
w45820 <= not w45807 and w45819;
w45821 <= not w45804 and w45820;
w45822 <= w45801 and w45821;
w45823 <= not pi0775 and not pi0816;
w45824 <= pi0775 and pi0816;
w45825 <= not w45823 and not w45824;
w45826 <= w45822 and not w45825;
w45827 <= w45800 and not w45826;
w45828 <= pi0747 and pi0773;
w45829 <= pi0769 and w45828;
w45830 <= pi0721 and w45829;
w45831 <= not pi0721 and not w45829;
w45832 <= pi0775 and not w45830;
w45833 <= not w45831 and w45832;
w45834 <= not w45807 and w45814;
w45835 <= not pi0721 and not pi0813;
w45836 <= pi0794 and pi0801;
w45837 <= w45835 and w45836;
w45838 <= w45834 and w45837;
w45839 <= not w45822 and not w45838;
w45840 <= pi0816 and not w45839;
w45841 <= w45833 and not w45840;
w45842 <= pi0795 and not w45841;
w45843 <= not pi0945 and pi0988;
w45844 <= pi0731 and w45843;
w45845 <= not w45800 and not w45833;
w45846 <= w45844 and not w45845;
w45847 <= not w45842 and w45846;
w45848 <= not pi0731 and not pi0795;
w45849 <= pi0731 and pi0795;
w45850 <= not w45848 and not w45849;
w45851 <= w45826 and not w45850;
w45852 <= pi0721 and not w45844;
w45853 <= not w45851 and w45852;
w45854 <= not w45827 and not w45853;
w45855 <= not w45847 and w45854;
w45856 <= pi0379 and w44621;
w45857 <= pi0403 and pi0591;
w45858 <= not pi0592 and w45857;
w45859 <= not w45856 and not w45858;
w45860 <= not pi0590 and not w45859;
w45861 <= pi0354 and w44628;
w45862 <= not w45860 and not w45861;
w45863 <= w45406 and not w45862;
w45864 <= pi0199 and not pi1045;
w45865 <= not pi0199 and w40436;
w45866 <= not w44613 and not w45864;
w45867 <= not w45865 and w45866;
w45868 <= pi0428 and pi0588;
w45869 <= w45415 and w45868;
w45870 <= not w45867 and not w45869;
w45871 <= not w45863 and w45870;
w45872 <= w5206 and not w45871;
w45873 <= not pi0795 and not pi1134;
w45874 <= not pi0851 and pi1134;
w45875 <= not pi1136 and not w45873;
w45876 <= not w45874 and w45875;
w45877 <= not pi0640 and not pi1134;
w45878 <= pi0776 and pi1134;
w45879 <= pi1136 and not w45877;
w45880 <= not w45878 and w45879;
w45881 <= not w45876 and not w45880;
w45882 <= not pi1135 and not w45881;
w45883 <= pi0694 and pi1134;
w45884 <= pi0732 and not pi1134;
w45885 <= pi1135 and pi1136;
w45886 <= not w45883 and w45885;
w45887 <= not w45884 and w45886;
w45888 <= not w45882 and not w45887;
w45889 <= w44690 and not w45888;
w45890 <= not w45872 and not w45889;
w45891 <= not pi1111 and w45209;
w45892 <= pi0723 and not w45209;
w45893 <= not pi0962 and not w45891;
w45894 <= not w45892 and w45893;
w45895 <= not pi1114 and w45209;
w45896 <= pi0724 and not w45209;
w45897 <= not pi0962 and not w45895;
w45898 <= not w45896 and w45897;
w45899 <= not pi1120 and w45209;
w45900 <= pi0725 and not w45209;
w45901 <= not pi0962 and not w45899;
w45902 <= not w45900 and w45901;
w45903 <= not pi0726 and not w45209;
w45904 <= not pi1126 and w45209;
w45905 <= not pi0962 and not w45903;
w45906 <= not w45904 and w45905;
w45907 <= not pi0727 and not w45209;
w45908 <= not pi1102 and w45209;
w45909 <= not pi0962 and not w45907;
w45910 <= not w45908 and w45909;
w45911 <= not pi1131 and w45209;
w45912 <= pi0728 and not w45209;
w45913 <= not pi0962 and not w45911;
w45914 <= not w45912 and w45913;
w45915 <= not pi0729 and not w45209;
w45916 <= not pi1104 and w45209;
w45917 <= not pi0962 and not w45915;
w45918 <= not w45916 and w45917;
w45919 <= not pi0730 and not w45209;
w45920 <= not pi1106 and w45209;
w45921 <= not pi0962 and not w45919;
w45922 <= not w45920 and w45921;
w45923 <= not w45801 and not w45835;
w45924 <= w45821 and not w45923;
w45925 <= pi0795 and not w45825;
w45926 <= w45924 and w45925;
w45927 <= not w45828 and not w45926;
w45928 <= w45844 and not w45927;
w45929 <= pi0731 and not w45926;
w45930 <= not w45825 and not w45923;
w45931 <= not pi0795 and pi0801;
w45932 <= not w45810 and w45931;
w45933 <= w45930 and w45932;
w45934 <= w45834 and w45933;
w45935 <= w45828 and not w45934;
w45936 <= not pi0731 and not w45935;
w45937 <= w45843 and not w45936;
w45938 <= not w45929 and not w45937;
w45939 <= not w45928 and not w45938;
w45940 <= not pi1128 and w44452;
w45941 <= pi0732 and not w44452;
w45942 <= not pi0962 and not w45940;
w45943 <= not w45941 and w45942;
w45944 <= pi0424 and w45224;
w45945 <= w45435 and w45944;
w45946 <= pi0375 and w45438;
w45947 <= pi0399 and pi0591;
w45948 <= w45440 and w45947;
w45949 <= not w45946 and not w45948;
w45950 <= not pi0590 and not w45949;
w45951 <= pi0316 and w44613;
w45952 <= w44628 and w45951;
w45953 <= not w45950 and not w45952;
w45954 <= not pi0588 and not w45953;
w45955 <= pi0199 and not pi1047;
w45956 <= not pi0200 and not pi0308;
w45957 <= pi0200 and not pi1037;
w45958 <= not w45956 and not w45957;
w45959 <= not pi0199 and not w45958;
w45960 <= not w44613 and not w45955;
w45961 <= not w45959 and w45960;
w45962 <= w5206 and not w45945;
w45963 <= not w45961 and w45962;
w45964 <= not w45954 and w45963;
w45965 <= not pi0619 and not pi1135;
w45966 <= not pi0648 and pi1135;
w45967 <= not pi1134 and not w45965;
w45968 <= not w45966 and w45967;
w45969 <= w44846 and w45968;
w45970 <= pi0737 and pi1135;
w45971 <= not pi0838 and not pi1136;
w45972 <= pi0777 and w44649;
w45973 <= pi1134 and not w45970;
w45974 <= not w45971 and w45973;
w45975 <= w45464 and w45974;
w45976 <= not w45972 and w45975;
w45977 <= not w5206 and not w45969;
w45978 <= not w45976 and w45977;
w45979 <= not w45964 and not w45978;
w45980 <= not pi1119 and w45209;
w45981 <= pi0734 and not w45209;
w45982 <= not pi0962 and not w45980;
w45983 <= not w45981 and w45982;
w45984 <= not pi0735 and not w45209;
w45985 <= not pi1109 and w45209;
w45986 <= not pi0962 and not w45984;
w45987 <= not w45985 and w45986;
w45988 <= not pi0736 and not w45209;
w45989 <= not pi1101 and w45209;
w45990 <= not pi0962 and not w45988;
w45991 <= not w45989 and w45990;
w45992 <= not pi1122 and w45209;
w45993 <= pi0737 and not w45209;
w45994 <= not pi0962 and not w45992;
w45995 <= not w45993 and w45994;
w45996 <= not pi1121 and w45209;
w45997 <= pi0738 and not w45209;
w45998 <= not pi0962 and not w45996;
w45999 <= not w45997 and w45998;
w46000 <= not pi0952 and not pi1061;
w46001 <= w44343 and w46000;
w46002 <= pi0832 and w46001;
w46003 <= pi1108 and w46002;
w46004 <= pi0739 and not w46002;
w46005 <= not pi0966 and not w46003;
w46006 <= not w46004 and w46005;
w46007 <= not pi0741 and not w46002;
w46008 <= pi1114 and w46002;
w46009 <= not pi0966 and not w46007;
w46010 <= not w46008 and w46009;
w46011 <= not pi0742 and not w46002;
w46012 <= pi1112 and w46002;
w46013 <= not pi0966 and not w46011;
w46014 <= not w46012 and w46013;
w46015 <= pi1109 and w46002;
w46016 <= pi0743 and not w46002;
w46017 <= not pi0966 and not w46015;
w46018 <= not w46016 and w46017;
w46019 <= not pi0744 and not w46002;
w46020 <= pi1131 and w46002;
w46021 <= not pi0966 and not w46019;
w46022 <= not w46020 and w46021;
w46023 <= not pi0745 and not w46002;
w46024 <= pi1111 and w46002;
w46025 <= not pi0966 and not w46023;
w46026 <= not w46024 and w46025;
w46027 <= pi1104 and w46002;
w46028 <= pi0746 and not w46002;
w46029 <= not pi0966 and not w46027;
w46030 <= not w46028 and w46029;
w46031 <= pi0773 and w45843;
w46032 <= not pi0747 and not w46031;
w46033 <= w45828 and w45843;
w46034 <= not w45850 and w45930;
w46035 <= pi0801 and w45817;
w46036 <= not w45804 and not w46031;
w46037 <= w45814 and w46036;
w46038 <= not w46035 and not w46037;
w46039 <= not w45807 and not w45810;
w46040 <= w46034 and w46039;
w46041 <= not w46038 and w46040;
w46042 <= not w46032 and not w46033;
w46043 <= not w46041 and w46042;
w46044 <= pi1106 and w46002;
w46045 <= pi0748 and not w46002;
w46046 <= not pi0966 and not w46044;
w46047 <= not w46045 and w46046;
w46048 <= pi1105 and w46002;
w46049 <= pi0749 and not w46002;
w46050 <= not pi0966 and not w46048;
w46051 <= not w46049 and w46050;
w46052 <= not pi0750 and not w46002;
w46053 <= pi1130 and w46002;
w46054 <= not pi0966 and not w46052;
w46055 <= not w46053 and w46054;
w46056 <= not pi0751 and not w46002;
w46057 <= pi1123 and w46002;
w46058 <= not pi0966 and not w46056;
w46059 <= not w46057 and w46058;
w46060 <= not pi0752 and not w46002;
w46061 <= pi1124 and w46002;
w46062 <= not pi0966 and not w46060;
w46063 <= not w46061 and w46062;
w46064 <= not pi0753 and not w46002;
w46065 <= pi1117 and w46002;
w46066 <= not pi0966 and not w46064;
w46067 <= not w46065 and w46066;
w46068 <= not pi0754 and not w46002;
w46069 <= pi1118 and w46002;
w46070 <= not pi0966 and not w46068;
w46071 <= not w46069 and w46070;
w46072 <= not pi0755 and not w46002;
w46073 <= pi1120 and w46002;
w46074 <= not pi0966 and not w46072;
w46075 <= not w46073 and w46074;
w46076 <= not pi0756 and not w46002;
w46077 <= pi1119 and w46002;
w46078 <= not pi0966 and not w46076;
w46079 <= not w46077 and w46078;
w46080 <= not pi0757 and not w46002;
w46081 <= pi1113 and w46002;
w46082 <= not pi0966 and not w46080;
w46083 <= not w46081 and w46082;
w46084 <= pi1101 and w46002;
w46085 <= pi0758 and not w46002;
w46086 <= not pi0966 and not w46084;
w46087 <= not w46085 and w46086;
w46088 <= not pi0759 and not w46002;
w46089 <= w44341 and w46001;
w46090 <= not w46088 and not w46089;
w46091 <= not pi0966 and not w46090;
w46092 <= not pi0760 and not w46002;
w46093 <= pi1115 and w46002;
w46094 <= not pi0966 and not w46092;
w46095 <= not w46093 and w46094;
w46096 <= not pi0761 and not w46002;
w46097 <= pi1121 and w46002;
w46098 <= not pi0966 and not w46096;
w46099 <= not w46097 and w46098;
w46100 <= not pi0762 and not w46002;
w46101 <= pi1129 and w46002;
w46102 <= not pi0966 and not w46100;
w46103 <= not w46101 and w46102;
w46104 <= pi1103 and w46002;
w46105 <= pi0763 and not w46002;
w46106 <= not pi0966 and not w46104;
w46107 <= not w46105 and w46106;
w46108 <= pi1107 and w46002;
w46109 <= pi0764 and not w46002;
w46110 <= not pi0966 and not w46108;
w46111 <= not w46109 and w46110;
w46112 <= w45821 and w46034;
w46113 <= pi0765 and not w46112;
w46114 <= pi0945 and not w46113;
w46115 <= not w45822 and not w45835;
w46116 <= not pi0765 and not w45806;
w46117 <= not w45809 and w46116;
w46118 <= not w45815 and w46117;
w46119 <= w45802 and not w46118;
w46120 <= not w45803 and not w46119;
w46121 <= w45820 and not w46120;
w46122 <= not pi0721 and not w46121;
w46123 <= w45823 and not w46122;
w46124 <= not w46115 and w46123;
w46125 <= w45824 and w45924;
w46126 <= not pi0765 and not w46125;
w46127 <= not w46124 and w46126;
w46128 <= not pi0795 and not w46127;
w46129 <= not pi0731 and not w46128;
w46130 <= not pi0795 and w46129;
w46131 <= pi0765 and not w46130;
w46132 <= not w45929 and not w46129;
w46133 <= not w46131 and not w46132;
w46134 <= not pi0945 and not w46133;
w46135 <= not w46114 and not w46134;
w46136 <= pi1110 and w46002;
w46137 <= pi0766 and not w46002;
w46138 <= not pi0966 and not w46136;
w46139 <= not w46137 and w46138;
w46140 <= not pi0767 and not w46002;
w46141 <= pi1116 and w46002;
w46142 <= not pi0966 and not w46140;
w46143 <= not w46141 and w46142;
w46144 <= not pi0768 and not w46002;
w46145 <= pi1125 and w46002;
w46146 <= not pi0966 and not w46144;
w46147 <= not w46145 and w46146;
w46148 <= pi0794 and not w45804;
w46149 <= not w45807 and w46148;
w46150 <= w45930 and w46149;
w46151 <= not w45818 and w46150;
w46152 <= not pi0775 and w46151;
w46153 <= not w46125 and not w46152;
w46154 <= pi0795 and not w46153;
w46155 <= pi0775 and w45828;
w46156 <= pi0769 and not w46155;
w46157 <= not pi0769 and w46155;
w46158 <= not w46156 and not w46157;
w46159 <= w45844 and not w46158;
w46160 <= not w46154 and w46159;
w46161 <= not w45850 and w46151;
w46162 <= pi0769 and not w45844;
w46163 <= not w46161 and w46162;
w46164 <= not w46160 and not w46163;
w46165 <= not pi0770 and not w46002;
w46166 <= pi1126 and w46002;
w46167 <= not pi0966 and not w46165;
w46168 <= not w46166 and w46167;
w46169 <= not w45824 and not w46123;
w46170 <= w45848 and not w46169;
w46171 <= not w45825 and w45849;
w46172 <= not w46170 and not w46171;
w46173 <= w45924 and not w46172;
w46174 <= not pi0945 and pi0987;
w46175 <= not w46173 and w46174;
w46176 <= pi0771 and pi0945;
w46177 <= not w46112 and w46176;
w46178 <= not w46175 and not w46177;
w46179 <= pi1102 and w46002;
w46180 <= pi0772 and not w46002;
w46181 <= not pi0966 and not w46179;
w46182 <= not w46180 and w46181;
w46183 <= not pi0801 and w45820;
w46184 <= w46173 and w46183;
w46185 <= w45843 and not w46184;
w46186 <= pi0801 and not w46034;
w46187 <= w45821 and not w46186;
w46188 <= pi0773 and not w46187;
w46189 <= not w46185 and not w46188;
w46190 <= not w46031 and not w46189;
w46191 <= not pi0774 and not w46002;
w46192 <= pi1127 and w46002;
w46193 <= not pi0966 and not w46191;
w46194 <= not w46192 and w46193;
w46195 <= pi0775 and not w46112;
w46196 <= pi0731 and not pi0945;
w46197 <= pi0765 and pi0771;
w46198 <= w45828 and w46197;
w46199 <= pi0795 and pi0800;
w46200 <= pi0801 and not pi0816;
w46201 <= w46199 and w46200;
w46202 <= not w45923 and w46201;
w46203 <= w45819 and w46202;
w46204 <= w46198 and not w46203;
w46205 <= not pi0775 and not w46204;
w46206 <= w46196 and not w46205;
w46207 <= not w46195 and not w46206;
w46208 <= not w45926 and not w46198;
w46209 <= pi0775 and w46196;
w46210 <= not w46208 and w46209;
w46211 <= not w46207 and not w46210;
w46212 <= not pi0776 and not w46002;
w46213 <= pi1128 and w46002;
w46214 <= not pi0966 and not w46212;
w46215 <= not w46213 and w46214;
w46216 <= not pi0777 and not w46002;
w46217 <= pi1122 and w46002;
w46218 <= not pi0966 and not w46216;
w46219 <= not w46217 and w46218;
w46220 <= pi0832 and pi0956;
w46221 <= not pi1046 and not pi1083;
w46222 <= pi1085 and w46221;
w46223 <= w46220 and w46222;
w46224 <= not pi0968 and w46223;
w46225 <= pi0778 and not w46224;
w46226 <= pi1100 and w46224;
w46227 <= not w46225 and not w46226;
w46228 <= pi0779 and not w44402;
w46229 <= pi0780 and not w44311;
w46230 <= pi0781 and not w46224;
w46231 <= pi1101 and w46224;
w46232 <= not w46230 and not w46231;
w46233 <= not w39908 and not w44355;
w46234 <= not w44310 and w46233;
w46235 <= pi0783 and not w46224;
w46236 <= pi1109 and w46224;
w46237 <= not w46235 and not w46236;
w46238 <= pi0784 and not w46224;
w46239 <= pi1110 and w46224;
w46240 <= not w46238 and not w46239;
w46241 <= pi0785 and not w46224;
w46242 <= pi1102 and w46224;
w46243 <= not w46241 and not w46242;
w46244 <= pi0024 and not pi0954;
w46245 <= pi0786 and pi0954;
w46246 <= not w46244 and not w46245;
w46247 <= pi0787 and not w46224;
w46248 <= pi1104 and w46224;
w46249 <= not w46247 and not w46248;
w46250 <= pi0788 and not w46224;
w46251 <= pi1105 and w46224;
w46252 <= not w46250 and not w46251;
w46253 <= pi0789 and not w46224;
w46254 <= pi1106 and w46224;
w46255 <= not w46253 and not w46254;
w46256 <= pi0790 and not w46224;
w46257 <= pi1107 and w46224;
w46258 <= not w46256 and not w46257;
w46259 <= pi0791 and not w46224;
w46260 <= pi1108 and w46224;
w46261 <= not w46259 and not w46260;
w46262 <= pi0792 and not w46224;
w46263 <= pi1103 and w46224;
w46264 <= not w46262 and not w46263;
w46265 <= pi0968 and w46223;
w46266 <= pi0794 and not w46265;
w46267 <= pi1130 and w46265;
w46268 <= not w46266 and not w46267;
w46269 <= pi0795 and not w46265;
w46270 <= pi1128 and w46265;
w46271 <= not w46269 and not w46270;
w46272 <= pi0266 and not pi0269;
w46273 <= pi0278 and pi0279;
w46274 <= not pi0280 and w46273;
w46275 <= w46272 and w46274;
w46276 <= not pi0281 and w46275;
w46277 <= w44594 and w46276;
w46278 <= pi0264 and not w46277;
w46279 <= not pi0264 and w46277;
w46280 <= not w46278 and not w46279;
w46281 <= pi0798 and not w46265;
w46282 <= pi1124 and w46265;
w46283 <= not w46281 and not w46282;
w46284 <= pi0799 and not w46265;
w46285 <= not pi1107 and w46265;
w46286 <= not w46284 and not w46285;
w46287 <= pi0800 and not w46265;
w46288 <= pi1125 and w46265;
w46289 <= not w46287 and not w46288;
w46290 <= pi0801 and not w46265;
w46291 <= pi1126 and w46265;
w46292 <= not w46290 and not w46291;
w46293 <= pi0803 and not w46265;
w46294 <= not pi1106 and w46265;
w46295 <= not w46293 and not w46294;
w46296 <= pi0804 and not w46265;
w46297 <= pi1109 and w46265;
w46298 <= not w46296 and not w46297;
w46299 <= not pi0282 and w44592;
w46300 <= not pi0270 and w46299;
w46301 <= pi0270 and not w46299;
w46302 <= not w46300 and not w46301;
w46303 <= pi0807 and not w46265;
w46304 <= pi1127 and w46265;
w46305 <= not w46303 and not w46304;
w46306 <= pi0808 and not w46265;
w46307 <= pi1101 and w46265;
w46308 <= not w46306 and not w46307;
w46309 <= pi0809 and not w46265;
w46310 <= not pi1103 and w46265;
w46311 <= not w46309 and not w46310;
w46312 <= pi0810 and not w46265;
w46313 <= pi1108 and w46265;
w46314 <= not w46312 and not w46313;
w46315 <= pi0811 and not w46265;
w46316 <= pi1102 and w46265;
w46317 <= not w46315 and not w46316;
w46318 <= pi0812 and not w46265;
w46319 <= not pi1104 and w46265;
w46320 <= not w46318 and not w46319;
w46321 <= pi0813 and not w46265;
w46322 <= pi1131 and w46265;
w46323 <= not w46321 and not w46322;
w46324 <= pi0814 and not w46265;
w46325 <= not pi1105 and w46265;
w46326 <= not w46324 and not w46325;
w46327 <= pi0815 and not w46265;
w46328 <= pi1110 and w46265;
w46329 <= not w46327 and not w46328;
w46330 <= pi0816 and not w46265;
w46331 <= pi1129 and w46265;
w46332 <= not w46330 and not w46331;
w46333 <= pi0269 and not w44590;
w46334 <= not w44591 and not w46333;
w46335 <= w5206 and w11735;
w46336 <= not w11588 and not w46335;
w46337 <= pi0265 and not w44596;
w46338 <= not w44597 and not w46337;
w46339 <= pi0277 and not w46300;
w46340 <= not w44595 and not w46339;
w46341 <= not pi0811 and not pi0893;
w46342 <= not pi0982 and not w7637;
w46343 <= w5189 and w5206;
w46344 <= not w46342 and not w46343;
w46345 <= w495 and not w46344;
w46346 <= pi0123 and w167;
w46347 <= pi1131 and not w46346;
w46348 <= pi1127 and not w46346;
w46349 <= not w46347 and not w46348;
w46350 <= not pi0825 and w46346;
w46351 <= w46349 and not w46350;
w46352 <= pi1131 and w46348;
w46353 <= not w46351 and not w46352;
w46354 <= pi1124 and not pi1130;
w46355 <= not pi1124 and pi1130;
w46356 <= not w46354 and not w46355;
w46357 <= not pi1128 and not pi1129;
w46358 <= pi1128 and pi1129;
w46359 <= not w46357 and not w46358;
w46360 <= not pi1125 and not pi1126;
w46361 <= pi1125 and pi1126;
w46362 <= not w46360 and not w46361;
w46363 <= w46359 and not w46362;
w46364 <= not w46359 and w46362;
w46365 <= not w46363 and not w46364;
w46366 <= w46356 and w46365;
w46367 <= not w46356 and not w46365;
w46368 <= not w46366 and not w46367;
w46369 <= not w46353 and not w46368;
w46370 <= pi0825 and w46346;
w46371 <= w46349 and not w46370;
w46372 <= not w46352 and w46368;
w46373 <= not w46371 and w46372;
w46374 <= not w46369 and not w46373;
w46375 <= pi1123 and not w46346;
w46376 <= pi1122 and not w46346;
w46377 <= not w46375 and not w46376;
w46378 <= not pi0826 and w46346;
w46379 <= w46377 and not w46378;
w46380 <= pi1123 and w46376;
w46381 <= not w46379 and not w46380;
w46382 <= pi1118 and not pi1119;
w46383 <= not pi1118 and pi1119;
w46384 <= not w46382 and not w46383;
w46385 <= not pi1120 and not pi1121;
w46386 <= pi1120 and pi1121;
w46387 <= not w46385 and not w46386;
w46388 <= not pi1116 and not pi1117;
w46389 <= pi1116 and pi1117;
w46390 <= not w46388 and not w46389;
w46391 <= w46387 and not w46390;
w46392 <= not w46387 and w46390;
w46393 <= not w46391 and not w46392;
w46394 <= w46384 and w46393;
w46395 <= not w46384 and not w46393;
w46396 <= not w46394 and not w46395;
w46397 <= not w46381 and not w46396;
w46398 <= pi0826 and w46346;
w46399 <= w46377 and not w46398;
w46400 <= not w46380 and w46396;
w46401 <= not w46399 and w46400;
w46402 <= not w46397 and not w46401;
w46403 <= pi1100 and not w46346;
w46404 <= pi1107 and not w46346;
w46405 <= not w46403 and not w46404;
w46406 <= not pi0827 and w46346;
w46407 <= w46405 and not w46406;
w46408 <= pi1100 and w46404;
w46409 <= not w46407 and not w46408;
w46410 <= pi1103 and not pi1105;
w46411 <= not pi1103 and pi1105;
w46412 <= not w46410 and not w46411;
w46413 <= not pi1101 and not pi1102;
w46414 <= pi1101 and pi1102;
w46415 <= not w46413 and not w46414;
w46416 <= not pi1104 and not pi1106;
w46417 <= pi1104 and pi1106;
w46418 <= not w46416 and not w46417;
w46419 <= w46415 and not w46418;
w46420 <= not w46415 and w46418;
w46421 <= not w46419 and not w46420;
w46422 <= w46412 and w46421;
w46423 <= not w46412 and not w46421;
w46424 <= not w46422 and not w46423;
w46425 <= not w46409 and not w46424;
w46426 <= pi0827 and w46346;
w46427 <= w46405 and not w46426;
w46428 <= not w46408 and w46424;
w46429 <= not w46427 and w46428;
w46430 <= not w46425 and not w46429;
w46431 <= pi1115 and not w46346;
w46432 <= pi1114 and not w46346;
w46433 <= not w46431 and not w46432;
w46434 <= not pi0828 and w46346;
w46435 <= w46433 and not w46434;
w46436 <= pi1115 and w46432;
w46437 <= not w46435 and not w46436;
w46438 <= pi1110 and not pi1111;
w46439 <= not pi1110 and pi1111;
w46440 <= not w46438 and not w46439;
w46441 <= not pi1112 and not pi1113;
w46442 <= pi1112 and pi1113;
w46443 <= not w46441 and not w46442;
w46444 <= not pi1108 and not pi1109;
w46445 <= pi1108 and pi1109;
w46446 <= not w46444 and not w46445;
w46447 <= w46443 and not w46446;
w46448 <= not w46443 and w46446;
w46449 <= not w46447 and not w46448;
w46450 <= w46440 and w46449;
w46451 <= not w46440 and not w46449;
w46452 <= not w46450 and not w46451;
w46453 <= not w46437 and not w46452;
w46454 <= pi0828 and w46346;
w46455 <= w46433 and not w46454;
w46456 <= not w46436 and w46452;
w46457 <= not w46455 and w46456;
w46458 <= not w46453 and not w46457;
w46459 <= w493 and w5206;
w46460 <= pi0951 and not w46459;
w46461 <= pi1092 and not w46460;
w46462 <= pi0281 and not w46275;
w46463 <= not w46276 and not w46462;
w46464 <= not pi0832 and pi1091;
w46465 <= pi1162 and w46464;
w46466 <= w6437 and w46465;
w46467 <= pi0833 and not w489;
w46468 <= not w14450 and not w46467;
w46469 <= pi0946 and w489;
w46470 <= pi0282 and not w44592;
w46471 <= not w46299 and not w46470;
w46472 <= not pi0955 and pi1049;
w46473 <= pi0837 and pi0955;
w46474 <= not w46472 and not w46473;
w46475 <= not pi0955 and pi1047;
w46476 <= pi0838 and pi0955;
w46477 <= not w46475 and not w46476;
w46478 <= not pi0955 and pi1074;
w46479 <= pi0839 and pi0955;
w46480 <= not w46478 and not w46479;
w46481 <= pi0840 and not w489;
w46482 <= pi1196 and w489;
w46483 <= not w46481 and not w46482;
w46484 <= not pi0033 and w6542;
w46485 <= not pi0955 and pi1035;
w46486 <= pi0842 and pi0955;
w46487 <= not w46485 and not w46486;
w46488 <= not pi0955 and pi1079;
w46489 <= pi0843 and pi0955;
w46490 <= not w46488 and not w46489;
w46491 <= not pi0955 and pi1078;
w46492 <= pi0844 and pi0955;
w46493 <= not w46491 and not w46492;
w46494 <= not pi0955 and pi1043;
w46495 <= pi0845 and pi0955;
w46496 <= not w46494 and not w46495;
w46497 <= pi0846 and not w40465;
w46498 <= pi1134 and w40465;
w46499 <= not w46497 and not w46498;
w46500 <= not pi0955 and pi1055;
w46501 <= pi0847 and pi0955;
w46502 <= not w46500 and not w46501;
w46503 <= not pi0955 and pi1039;
w46504 <= pi0848 and pi0955;
w46505 <= not w46503 and not w46504;
w46506 <= pi0849 and not w489;
w46507 <= pi1198 and w489;
w46508 <= not w46506 and not w46507;
w46509 <= not pi0955 and pi1048;
w46510 <= pi0850 and pi0955;
w46511 <= not w46509 and not w46510;
w46512 <= not pi0955 and pi1045;
w46513 <= pi0851 and pi0955;
w46514 <= not w46512 and not w46513;
w46515 <= not pi0955 and pi1062;
w46516 <= pi0852 and pi0955;
w46517 <= not w46515 and not w46516;
w46518 <= not pi0955 and pi1080;
w46519 <= pi0853 and pi0955;
w46520 <= not w46518 and not w46519;
w46521 <= not pi0955 and pi1051;
w46522 <= pi0854 and pi0955;
w46523 <= not w46521 and not w46522;
w46524 <= not pi0955 and pi1065;
w46525 <= pi0855 and pi0955;
w46526 <= not w46524 and not w46525;
w46527 <= not pi0955 and pi1067;
w46528 <= pi0856 and pi0955;
w46529 <= not w46527 and not w46528;
w46530 <= not pi0955 and pi1058;
w46531 <= pi0857 and pi0955;
w46532 <= not w46530 and not w46531;
w46533 <= not pi0955 and pi1087;
w46534 <= pi0858 and pi0955;
w46535 <= not w46533 and not w46534;
w46536 <= not pi0955 and pi1070;
w46537 <= pi0859 and pi0955;
w46538 <= not w46536 and not w46537;
w46539 <= not pi0955 and pi1076;
w46540 <= pi0860 and pi0955;
w46541 <= not w46539 and not w46540;
w46542 <= pi1093 and pi1141;
w46543 <= pi0861 and not pi1093;
w46544 <= not w46542 and not w46543;
w46545 <= not pi0228 and not w46544;
w46546 <= not pi0123 and not pi1141;
w46547 <= pi0123 and not pi0861;
w46548 <= pi0228 and not w46546;
w46549 <= not w46547 and w46548;
w46550 <= not w46545 and not w46549;
w46551 <= pi0862 and not w40465;
w46552 <= pi1139 and w40465;
w46553 <= not w46551 and not w46552;
w46554 <= pi0863 and not w489;
w46555 <= pi1199 and w489;
w46556 <= not w46554 and not w46555;
w46557 <= pi0864 and not w489;
w46558 <= pi1197 and w489;
w46559 <= not w46557 and not w46558;
w46560 <= not pi0955 and pi1040;
w46561 <= pi0865 and pi0955;
w46562 <= not w46560 and not w46561;
w46563 <= not pi0955 and pi1053;
w46564 <= pi0866 and pi0955;
w46565 <= not w46563 and not w46564;
w46566 <= not pi0955 and pi1057;
w46567 <= pi0867 and pi0955;
w46568 <= not w46566 and not w46567;
w46569 <= not pi0955 and pi1063;
w46570 <= pi0868 and pi0955;
w46571 <= not w46569 and not w46570;
w46572 <= pi1093 and pi1140;
w46573 <= pi0869 and not pi1093;
w46574 <= not w46572 and not w46573;
w46575 <= not pi0228 and not w46574;
w46576 <= not pi0123 and not pi1140;
w46577 <= pi0123 and not pi0869;
w46578 <= pi0228 and not w46576;
w46579 <= not w46577 and w46578;
w46580 <= not w46575 and not w46579;
w46581 <= not pi0955 and pi1069;
w46582 <= pi0870 and pi0955;
w46583 <= not w46581 and not w46582;
w46584 <= not pi0955 and pi1072;
w46585 <= pi0871 and pi0955;
w46586 <= not w46584 and not w46585;
w46587 <= not pi0955 and pi1084;
w46588 <= pi0872 and pi0955;
w46589 <= not w46587 and not w46588;
w46590 <= not pi0955 and pi1044;
w46591 <= pi0873 and pi0955;
w46592 <= not w46590 and not w46591;
w46593 <= not pi0955 and pi1036;
w46594 <= pi0874 and pi0955;
w46595 <= not w46593 and not w46594;
w46596 <= pi1093 and not pi1136;
w46597 <= not pi0875 and not pi1093;
w46598 <= not w46596 and not w46597;
w46599 <= not pi0228 and not w46598;
w46600 <= not pi0123 and pi1136;
w46601 <= pi0123 and pi0875;
w46602 <= pi0228 and not w46600;
w46603 <= not w46601 and w46602;
w46604 <= not w46599 and not w46603;
w46605 <= not pi0955 and pi1037;
w46606 <= pi0876 and pi0955;
w46607 <= not w46605 and not w46606;
w46608 <= pi1093 and pi1138;
w46609 <= pi0877 and not pi1093;
w46610 <= not w46608 and not w46609;
w46611 <= not pi0228 and not w46610;
w46612 <= not pi0123 and not pi1138;
w46613 <= pi0123 and not pi0877;
w46614 <= pi0228 and not w46612;
w46615 <= not w46613 and w46614;
w46616 <= not w46611 and not w46615;
w46617 <= pi1093 and pi1137;
w46618 <= pi0878 and not pi1093;
w46619 <= not w46617 and not w46618;
w46620 <= not pi0228 and not w46619;
w46621 <= not pi0123 and not pi1137;
w46622 <= pi0123 and not pi0878;
w46623 <= pi0228 and not w46621;
w46624 <= not w46622 and w46623;
w46625 <= not w46620 and not w46624;
w46626 <= pi1093 and pi1135;
w46627 <= pi0879 and not pi1093;
w46628 <= not w46626 and not w46627;
w46629 <= not pi0228 and not w46628;
w46630 <= not pi0123 and not pi1135;
w46631 <= pi0123 and not pi0879;
w46632 <= pi0228 and not w46630;
w46633 <= not w46631 and w46632;
w46634 <= not w46629 and not w46633;
w46635 <= not pi0955 and pi1081;
w46636 <= pi0880 and pi0955;
w46637 <= not w46635 and not w46636;
w46638 <= not pi0955 and pi1059;
w46639 <= pi0881 and pi0955;
w46640 <= not w46638 and not w46639;
w46641 <= not pi0883 and w46346;
w46642 <= not w46404 and not w46641;
w46643 <= pi1124 and not w46346;
w46644 <= not pi0884 and w46346;
w46645 <= not w46643 and not w46644;
w46646 <= pi1125 and not w46346;
w46647 <= not pi0885 and w46346;
w46648 <= not w46646 and not w46647;
w46649 <= pi1109 and not w46346;
w46650 <= not pi0886 and w46346;
w46651 <= not w46649 and not w46650;
w46652 <= not pi0887 and w46346;
w46653 <= not w46403 and not w46652;
w46654 <= pi1120 and not w46346;
w46655 <= not pi0888 and w46346;
w46656 <= not w46654 and not w46655;
w46657 <= pi1103 and not w46346;
w46658 <= not pi0889 and w46346;
w46659 <= not w46657 and not w46658;
w46660 <= pi1126 and not w46346;
w46661 <= not pi0890 and w46346;
w46662 <= not w46660 and not w46661;
w46663 <= pi1116 and not w46346;
w46664 <= not pi0891 and w46346;
w46665 <= not w46663 and not w46664;
w46666 <= pi1101 and not w46346;
w46667 <= not pi0892 and w46346;
w46668 <= not w46666 and not w46667;
w46669 <= pi1119 and not w46346;
w46670 <= not pi0894 and w46346;
w46671 <= not w46669 and not w46670;
w46672 <= pi1113 and not w46346;
w46673 <= not pi0895 and w46346;
w46674 <= not w46672 and not w46673;
w46675 <= pi1118 and not w46346;
w46676 <= not pi0896 and w46346;
w46677 <= not w46675 and not w46676;
w46678 <= pi1129 and not w46346;
w46679 <= not pi0898 and w46346;
w46680 <= not w46678 and not w46679;
w46681 <= not pi0899 and w46346;
w46682 <= not w46431 and not w46681;
w46683 <= pi1110 and not w46346;
w46684 <= not pi0900 and w46346;
w46685 <= not w46683 and not w46684;
w46686 <= pi1111 and not w46346;
w46687 <= not pi0902 and w46346;
w46688 <= not w46686 and not w46687;
w46689 <= pi1121 and not w46346;
w46690 <= not pi0903 and w46346;
w46691 <= not w46689 and not w46690;
w46692 <= not pi0904 and w46346;
w46693 <= not w46348 and not w46692;
w46694 <= not pi0905 and w46346;
w46695 <= not w46347 and not w46694;
w46696 <= pi1128 and not w46346;
w46697 <= not pi0906 and w46346;
w46698 <= not w46696 and not w46697;
w46699 <= not pi0782 and not pi0907;
w46700 <= not pi0624 and not pi0979;
w46701 <= not pi0598 and pi0979;
w46702 <= pi0782 and not w46700;
w46703 <= not w46701 and w46702;
w46704 <= not pi0604 and not pi0979;
w46705 <= pi0615 and pi0979;
w46706 <= not w46704 and not w46705;
w46707 <= pi0782 and not w46706;
w46708 <= not w46699 and not w46703;
w46709 <= not w46707 and w46708;
w46710 <= not pi0908 and w46346;
w46711 <= not w46376 and not w46710;
w46712 <= pi1105 and not w46346;
w46713 <= not pi0909 and w46346;
w46714 <= not w46712 and not w46713;
w46715 <= pi1117 and not w46346;
w46716 <= not pi0910 and w46346;
w46717 <= not w46715 and not w46716;
w46718 <= pi1130 and not w46346;
w46719 <= not pi0911 and w46346;
w46720 <= not w46718 and not w46719;
w46721 <= not pi0912 and w46346;
w46722 <= not w46432 and not w46721;
w46723 <= pi1106 and not w46346;
w46724 <= not pi0913 and w46346;
w46725 <= not w46723 and not w46724;
w46726 <= pi0280 and not w44589;
w46727 <= not w44590 and not w46726;
w46728 <= pi1108 and not w46346;
w46729 <= not pi0915 and w46346;
w46730 <= not w46728 and not w46729;
w46731 <= not pi0916 and w46346;
w46732 <= not w46375 and not w46731;
w46733 <= pi1112 and not w46346;
w46734 <= not pi0917 and w46346;
w46735 <= not w46733 and not w46734;
w46736 <= pi1104 and not w46346;
w46737 <= not pi0918 and w46346;
w46738 <= not w46736 and not w46737;
w46739 <= pi1102 and not w46346;
w46740 <= not pi0919 and w46346;
w46741 <= not w46739 and not w46740;
w46742 <= pi1093 and pi1139;
w46743 <= pi0920 and not pi1093;
w46744 <= not w46742 and not w46743;
w46745 <= pi0921 and not pi1093;
w46746 <= not w46572 and not w46745;
w46747 <= not pi0922 and not pi1093;
w46748 <= pi1093 and not pi1152;
w46749 <= not w46747 and not w46748;
w46750 <= not pi0923 and not pi1093;
w46751 <= pi1093 and not pi1154;
w46752 <= not w46750 and not w46751;
w46753 <= not pi0300 and pi0301;
w46754 <= pi0311 and not pi0312;
w46755 <= w46753 and w46754;
w46756 <= not pi0925 and not pi1093;
w46757 <= pi1093 and not pi1155;
w46758 <= not w46756 and not w46757;
w46759 <= not pi0926 and not pi1093;
w46760 <= pi1093 and not pi1157;
w46761 <= not w46759 and not w46760;
w46762 <= not pi0927 and not pi1093;
w46763 <= pi1093 and not pi1145;
w46764 <= not w46762 and not w46763;
w46765 <= not pi0928 and not pi1093;
w46766 <= not w46596 and not w46765;
w46767 <= not pi0929 and not pi1093;
w46768 <= pi1093 and not pi1144;
w46769 <= not w46767 and not w46768;
w46770 <= not pi0930 and not pi1093;
w46771 <= pi1093 and not pi1134;
w46772 <= not w46770 and not w46771;
w46773 <= not pi0931 and not pi1093;
w46774 <= pi1093 and not pi1150;
w46775 <= not w46773 and not w46774;
w46776 <= pi0932 and not pi1093;
w46777 <= not w40454 and not w46776;
w46778 <= pi0933 and not pi1093;
w46779 <= not w46617 and not w46778;
w46780 <= not pi0934 and not pi1093;
w46781 <= pi1093 and not pi1147;
w46782 <= not w46780 and not w46781;
w46783 <= pi0935 and not pi1093;
w46784 <= not w46542 and not w46783;
w46785 <= not pi0936 and not pi1093;
w46786 <= pi1093 and not pi1149;
w46787 <= not w46785 and not w46786;
w46788 <= not pi0937 and not pi1093;
w46789 <= pi1093 and not pi1148;
w46790 <= not w46788 and not w46789;
w46791 <= pi0938 and not pi1093;
w46792 <= not w46626 and not w46791;
w46793 <= not pi0939 and not pi1093;
w46794 <= pi1093 and not pi1146;
w46795 <= not w46793 and not w46794;
w46796 <= pi0940 and not pi1093;
w46797 <= not w46608 and not w46796;
w46798 <= not pi0941 and not pi1093;
w46799 <= pi1093 and not pi1153;
w46800 <= not w46798 and not w46799;
w46801 <= not pi0942 and not pi1093;
w46802 <= pi1093 and not pi1156;
w46803 <= not w46801 and not w46802;
w46804 <= not pi0943 and not pi1093;
w46805 <= pi1093 and not pi1151;
w46806 <= not w46804 and not w46805;
w46807 <= pi1093 and pi1143;
w46808 <= pi0944 and not pi1093;
w46809 <= not w46807 and not w46808;
w46810 <= pi0230 and w489;
w46811 <= not pi0782 and pi0947;
w46812 <= not w46703 and not w46811;
w46813 <= not pi0266 and not pi0992;
w46814 <= not w44589 and not w46813;
w46815 <= not pi0313 and not pi0954;
w46816 <= pi0949 and pi0954;
w46817 <= not w46815 and not w46816;
w46818 <= not w5189 and w11834;
w46819 <= pi0957 and pi1092;
w46820 <= not pi0031 and not w46819;
w46821 <= not pi0782 and pi0960;
w46822 <= not pi0230 and pi0961;
w46823 <= not pi0782 and pi0963;
w46824 <= not pi0230 and pi0967;
w46825 <= not pi0230 and pi0969;
w46826 <= not pi0782 and pi0970;
w46827 <= not pi0230 and pi0971;
w46828 <= not pi0782 and pi0972;
w46829 <= not pi0230 and pi0974;
w46830 <= not pi0782 and pi0975;
w46831 <= not pi0230 and pi0977;
w46832 <= not pi0782 and pi0978;
w46833 <= not pi0598 and pi0615;
w46834 <= pi0824 and pi1092;
w46835 <= not pi0604 and not pi0624;
one <= '1';
po0000 <= pi0668;-- level 0
po0001 <= pi0672;-- level 0
po0002 <= pi0664;-- level 0
po0003 <= pi0667;-- level 0
po0004 <= pi0676;-- level 0
po0005 <= pi0673;-- level 0
po0006 <= pi0675;-- level 0
po0007 <= pi0666;-- level 0
po0008 <= pi0679;-- level 0
po0009 <= pi0674;-- level 0
po0010 <= pi0663;-- level 0
po0011 <= pi0670;-- level 0
po0012 <= pi0677;-- level 0
po0013 <= pi0682;-- level 0
po0014 <= pi0671;-- level 0
po0015 <= pi0678;-- level 0
po0016 <= pi0718;-- level 0
po0017 <= pi0707;-- level 0
po0018 <= pi0708;-- level 0
po0019 <= pi0713;-- level 0
po0020 <= pi0711;-- level 0
po0021 <= pi0716;-- level 0
po0022 <= pi0733;-- level 0
po0023 <= pi0712;-- level 0
po0024 <= pi0689;-- level 0
po0025 <= pi0717;-- level 0
po0026 <= pi0692;-- level 0
po0027 <= pi0719;-- level 0
po0028 <= pi0722;-- level 0
po0029 <= pi0714;-- level 0
po0030 <= pi0720;-- level 0
po0031 <= pi0685;-- level 0
po0032 <= pi0837;-- level 0
po0033 <= pi0850;-- level 0
po0034 <= pi0872;-- level 0
po0035 <= pi0871;-- level 0
po0036 <= pi0881;-- level 0
po0037 <= pi0866;-- level 0
po0038 <= pi0876;-- level 0
po0039 <= pi0873;-- level 0
po0040 <= pi0874;-- level 0
po0041 <= pi0859;-- level 0
po0042 <= pi0855;-- level 0
po0043 <= pi0852;-- level 0
po0044 <= pi0870;-- level 0
po0045 <= pi0848;-- level 0
po0046 <= pi0865;-- level 0
po0047 <= pi0856;-- level 0
po0048 <= pi0853;-- level 0
po0049 <= pi0847;-- level 0
po0050 <= pi0857;-- level 0
po0051 <= pi0854;-- level 0
po0052 <= pi0858;-- level 0
po0053 <= pi0845;-- level 0
po0054 <= pi0838;-- level 0
po0055 <= pi0842;-- level 0
po0056 <= pi0843;-- level 0
po0057 <= pi0839;-- level 0
po0058 <= pi0844;-- level 0
po0059 <= pi0868;-- level 0
po0060 <= pi0851;-- level 0
po0061 <= pi0867;-- level 0
po0062 <= pi0880;-- level 0
po0063 <= pi0860;-- level 0
po0064 <= pi1030;-- level 0
po0065 <= pi1034;-- level 0
po0066 <= pi1015;-- level 0
po0067 <= pi1020;-- level 0
po0068 <= pi1025;-- level 0
po0069 <= pi1005;-- level 0
po0070 <= pi0996;-- level 0
po0071 <= pi1012;-- level 0
po0072 <= pi0993;-- level 0
po0073 <= pi1016;-- level 0
po0074 <= pi1021;-- level 0
po0075 <= pi1010;-- level 0
po0076 <= pi1027;-- level 0
po0077 <= pi1018;-- level 0
po0078 <= pi1017;-- level 0
po0079 <= pi1024;-- level 0
po0080 <= pi1009;-- level 0
po0081 <= pi1032;-- level 0
po0082 <= pi1003;-- level 0
po0083 <= pi0997;-- level 0
po0084 <= pi1013;-- level 0
po0085 <= pi1011;-- level 0
po0086 <= pi1008;-- level 0
po0087 <= pi1019;-- level 0
po0088 <= pi1031;-- level 0
po0089 <= pi1022;-- level 0
po0090 <= pi1000;-- level 0
po0091 <= pi1023;-- level 0
po0092 <= pi1002;-- level 0
po0093 <= pi1026;-- level 0
po0094 <= pi1006;-- level 0
po0095 <= pi0998;-- level 0
po0096 <= pi0031;-- level 0
po0097 <= pi0080;-- level 0
po0098 <= pi0893;-- level 0
po0099 <= pi0467;-- level 0
po0100 <= pi0078;-- level 0
po0101 <= pi0112;-- level 0
po0102 <= pi0013;-- level 0
po0103 <= pi0025;-- level 0
po0104 <= pi0226;-- level 0
po0105 <= pi0127;-- level 0
po0106 <= pi0822;-- level 0
po0107 <= pi0808;-- level 0
po0108 <= pi0227;-- level 0
po0109 <= pi0477;-- level 0
po0110 <= pi0834;-- level 0
po0111 <= pi0229;-- level 0
po0112 <= pi0012;-- level 0
po0113 <= pi0011;-- level 0
po0114 <= pi0010;-- level 0
po0115 <= pi0009;-- level 0
po0116 <= pi0008;-- level 0
po0117 <= pi0007;-- level 0
po0118 <= pi0006;-- level 0
po0119 <= pi0005;-- level 0
po0120 <= pi0004;-- level 0
po0121 <= pi0003;-- level 0
po0122 <= pi0000;-- level 0
po0123 <= pi0002;-- level 0
po0124 <= pi0001;-- level 0
po0125 <= pi0310;-- level 0
po0126 <= pi0302;-- level 0
po0127 <= pi0475;-- level 0
po0128 <= pi0474;-- level 0
po0129 <= pi0466;-- level 0
po0130 <= pi0473;-- level 0
po0131 <= pi0471;-- level 0
po0132 <= pi0472;-- level 0
po0133 <= pi0470;-- level 0
po0134 <= pi0469;-- level 0
po0135 <= pi0465;-- level 0
po0136 <= pi1028;-- level 0
po0137 <= pi1033;-- level 0
po0138 <= pi0995;-- level 0
po0139 <= pi0994;-- level 0
po0140 <= pi0028;-- level 0
po0141 <= pi0027;-- level 0
po0142 <= pi0026;-- level 0
po0143 <= pi0029;-- level 0
po0144 <= pi0015;-- level 0
po0145 <= pi0014;-- level 0
po0146 <= pi0021;-- level 0
po0147 <= pi0020;-- level 0
po0148 <= pi0019;-- level 0
po0149 <= pi0018;-- level 0
po0150 <= pi0017;-- level 0
po0151 <= pi0016;-- level 0
po0152 <= pi1096;-- level 0
po0153 <= not w871;-- level 95
po0154 <= not w1105;-- level 78
po0155 <= w1276;-- level 80
po0156 <= w1506;-- level 83
po0157 <= not w1733;-- level 82
po0158 <= w1956;-- level 82
po0159 <= w2179;-- level 82
po0160 <= not w2410;-- level 83
po0161 <= w2633;-- level 82
po0162 <= w2856;-- level 82
po0163 <= not w3092;-- level 84
po0164 <= not w3327;-- level 84
po0165 <= w3682;-- level 83
po0166 <= one;-- level 0
po0167 <= w3866;-- level 69
po0168 <= pi0228;-- level 0
po0169 <= pi0022;-- level 0
po0170 <= not pi1090;-- level 0
po0171 <= w4134;-- level 68
po0172 <= w4257;-- level 68
po0173 <= w4387;-- level 69
po0174 <= w4483;-- level 69
po0175 <= w4579;-- level 69
po0176 <= w4675;-- level 69
po0177 <= w4771;-- level 69
po0178 <= w4863;-- level 69
po0179 <= pi1089;-- level 0
po0180 <= pi0023;-- level 0
po0181 <= w3866;-- level 69
po0182 <= w4918;-- level 69
po0183 <= not w4968;-- level 74
po0184 <= not w4973;-- level 4
po0185 <= not w4975;-- level 4
po0186 <= not w4977;-- level 4
po0187 <= not w4979;-- level 4
po0188 <= pi0037;-- level 0
po0189 <= not w6440;-- level 80
po0190 <= w6536;-- level 32
po0191 <= w7253;-- level 70
po0192 <= w7629;-- level 68
po0193 <= w7709;-- level 37
po0194 <= w7731;-- level 22
po0195 <= w4915;-- level 67
po0196 <= w7762;-- level 22
po0197 <= w7843;-- level 34
po0198 <= w7857;-- level 25
po0199 <= w8046;-- level 49
po0200 <= not w8291;-- level 60
po0201 <= not w8469;-- level 62
po0202 <= not w8544;-- level 46
po0203 <= w8548;-- level 23
po0204 <= w8568;-- level 23
po0205 <= w8613;-- level 29
po0206 <= w8619;-- level 9
po0207 <= w8638;-- level 23
po0208 <= w8664;-- level 28
po0209 <= w8672;-- level 12
po0210 <= w8823;-- level 62
po0211 <= w8835;-- level 23
po0212 <= w8855;-- level 23
po0213 <= w8869;-- level 25
po0214 <= w8877;-- level 25
po0215 <= w8887;-- level 27
po0216 <= w8890;-- level 21
po0217 <= w8896;-- level 27
po0218 <= w8905;-- level 25
po0219 <= w8910;-- level 20
po0220 <= w8915;-- level 26
po0221 <= w8921;-- level 23
po0222 <= w8931;-- level 18
po0223 <= w8935;-- level 29
po0224 <= w8952;-- level 19
po0225 <= w8957;-- level 11
po0226 <= w8965;-- level 29
po0227 <= w8978;-- level 18
po0228 <= w8998;-- level 24
po0229 <= w9020;-- level 21
po0230 <= w9035;-- level 31
po0231 <= w9047;-- level 31
po0232 <= w9062;-- level 26
po0233 <= w9072;-- level 27
po0234 <= w9225;-- level 46
po0235 <= w9235;-- level 25
po0236 <= w9237;-- level 2
po0237 <= not w9740;-- level 67
po0238 <= w10591;-- level 70
po0239 <= w10601;-- level 17
po0240 <= w10609;-- level 13
po0241 <= w10623;-- level 15
po0242 <= w10629;-- level 17
po0243 <= w10634;-- level 15
po0244 <= w10638;-- level 30
po0245 <= w10642;-- level 13
po0246 <= w10662;-- level 26
po0247 <= w10672;-- level 22
po0248 <= w10677;-- level 21
po0249 <= w10689;-- level 32
po0250 <= w10701;-- level 32
po0251 <= w10708;-- level 24
po0252 <= w10726;-- level 27
po0253 <= w10742;-- level 30
po0254 <= w10753;-- level 26
po0255 <= w10763;-- level 29
po0256 <= w10768;-- level 24
po0257 <= not w10845;-- level 50
po0258 <= w10862;-- level 22
po0259 <= not w10943;-- level 48
po0260 <= w10945;-- level 14
po0261 <= w10953;-- level 22
po0262 <= w10971;-- level 27
po0263 <= pi0117;-- level 0
po0264 <= w10981;-- level 25
po0265 <= w10983;-- level 14
po0266 <= w11001;-- level 28
po0267 <= w11003;-- level 20
po0268 <= w11014;-- level 23
po0269 <= w11020;-- level 23
po0270 <= not w11021;-- level 1
po0271 <= w11074;-- level 51
po0272 <= w11117;-- level 58
po0273 <= w11159;-- level 56
po0274 <= w11210;-- level 54
po0275 <= w11226;-- level 74
po0276 <= not w11531;-- level 65
po0277 <= not w11586;-- level 40
po0278 <= not w11989;-- level 52
po0279 <= not w12409;-- level 48
po0280 <= not w12417;-- level 48
po0281 <= w12471;-- level 37
po0282 <= not w12877;-- level 45
po0283 <= w13180;-- level 47
po0284 <= w13274;-- level 77
po0285 <= pi0131;-- level 0
po0286 <= w13299;-- level 75
po0287 <= w13434;-- level 43
po0288 <= w13442;-- level 38
po0289 <= not w13658;-- level 46
po0290 <= not w13719;-- level 40
po0291 <= not w13833;-- level 41
po0292 <= not w13952;-- level 45
po0293 <= not w14038;-- level 40
po0294 <= not w14051;-- level 27
po0295 <= w14136;-- level 58
po0296 <= w14190;-- level 58
po0297 <= w15628;-- level 113
po0298 <= w16153;-- level 111
po0299 <= w16928;-- level 113
po0300 <= w17454;-- level 113
po0301 <= w17973;-- level 114
po0302 <= w18461;-- level 99
po0303 <= not w18542;-- level 60
po0304 <= w18691;-- level 66
po0305 <= not w18755;-- level 65
po0306 <= w18814;-- level 65
po0307 <= w18870;-- level 65
po0308 <= w18948;-- level 64
po0309 <= not w19051;-- level 62
po0310 <= not w19132;-- level 65
po0311 <= w19184;-- level 65
po0312 <= w19224;-- level 67
po0313 <= w19254;-- level 66
po0314 <= w19311;-- level 66
po0315 <= w19367;-- level 65
po0316 <= w19423;-- level 65
po0317 <= w19482;-- level 65
po0318 <= not w19577;-- level 62
po0319 <= w19632;-- level 66
po0320 <= w19690;-- level 65
po0321 <= w19730;-- level 66
po0322 <= w19770;-- level 66
po0323 <= not w19867;-- level 62
po0324 <= w19910;-- level 65
po0325 <= not w19991;-- level 65
po0326 <= not w20072;-- level 65
po0327 <= not w20152;-- level 64
po0328 <= not w20233;-- level 65
po0329 <= not w20314;-- level 65
po0330 <= w20789;-- level 99
po0331 <= w21273;-- level 114
po0332 <= w21751;-- level 94
po0333 <= w22201;-- level 96
po0334 <= w22685;-- level 113
po0335 <= w23156;-- level 94
po0336 <= w23638;-- level 112
po0337 <= w24115;-- level 94
po0338 <= w24592;-- level 94
po0339 <= w25063;-- level 94
po0340 <= w25534;-- level 94
po0341 <= w26005;-- level 94
po0342 <= w26482;-- level 94
po0343 <= w26957;-- level 113
po0344 <= w27432;-- level 113
po0345 <= w27907;-- level 113
po0346 <= w28386;-- level 114
po0347 <= w28863;-- level 94
po0348 <= w29340;-- level 94
po0349 <= w29817;-- level 94
po0350 <= w30289;-- level 94
po0351 <= w30757;-- level 113
po0352 <= not w30807;-- level 56
po0353 <= not w30876;-- level 58
po0354 <= w30937;-- level 65
po0355 <= not w31573;-- level 94
po0356 <= not w31864;-- level 112
po0357 <= w32145;-- level 98
po0358 <= w32340;-- level 47
po0359 <= w32348;-- level 47
po0360 <= w32356;-- level 47
po0361 <= w32465;-- level 47
po0362 <= w32472;-- level 47
po0363 <= w32480;-- level 47
po0364 <= not w32972;-- level 107
po0365 <= not w33047;-- level 107
po0366 <= not w33207;-- level 107
po0367 <= w33333;-- level 53
po0368 <= not w33360;-- level 66
po0369 <= not w33381;-- level 66
po0370 <= not w33402;-- level 66
po0371 <= not w33423;-- level 66
po0372 <= not w33539;-- level 59
po0373 <= w33650;-- level 59
po0374 <= not w33669;-- level 106
po0375 <= w33676;-- level 47
po0376 <= not w33697;-- level 66
po0377 <= w33704;-- level 47
po0378 <= w33813;-- level 59
po0379 <= w34439;-- level 96
po0380 <= w35021;-- level 93
po0381 <= w35610;-- level 95
po0382 <= w35735;-- level 83
po0383 <= w35788;-- level 76
po0384 <= not w35819;-- level 31
po0385 <= not w35831;-- level 28
po0386 <= pi0232;-- level 0
po0387 <= w35914;-- level 41
po0388 <= pi0236;-- level 0
po0389 <= w35974;-- level 76
po0390 <= not w36386;-- level 25
po0391 <= not w36720;-- level 27
po0392 <= w36918;-- level 25
po0393 <= w36931;-- level 74
po0394 <= not w37193;-- level 25
po0395 <= not w37531;-- level 26
po0396 <= w37622;-- level 21
po0397 <= w38043;-- level 27
po0398 <= w38332;-- level 26
po0399 <= w38421;-- level 22
po0400 <= w38732;-- level 33
po0401 <= w38785;-- level 24
po0402 <= w39032;-- level 27
po0403 <= w39306;-- level 31
po0404 <= w39536;-- level 28
po0405 <= w39699;-- level 28
po0406 <= w39887;-- level 27
po0407 <= w39895;-- level 27
po0408 <= not w39905;-- level 5
po0409 <= w39947;-- level 37
po0410 <= w40183;-- level 33
po0411 <= w40409;-- level 31
po0412 <= w40415;-- level 5
po0413 <= w40421;-- level 5
po0414 <= w40427;-- level 5
po0415 <= w40433;-- level 5
po0416 <= w40439;-- level 5
po0417 <= not w40446;-- level 5
po0418 <= not w40453;-- level 5
po0419 <= not w40487;-- level 10
po0420 <= w40697;-- level 33
po0421 <= not w40742;-- level 14
po0422 <= not w40783;-- level 14
po0423 <= w40850;-- level 16
po0424 <= w41057;-- level 32
po0425 <= w41214;-- level 35
po0426 <= w41259;-- level 12
po0427 <= not w41303;-- level 12
po0428 <= w41352;-- level 17
po0429 <= w41453;-- level 35
po0430 <= not w41516;-- level 26
po0431 <= w41557;-- level 14
po0432 <= not w41631;-- level 35
po0433 <= not w41660;-- level 12
po0434 <= not w41703;-- level 14
po0435 <= w41772;-- level 18
po0436 <= w41831;-- level 14
po0437 <= w41875;-- level 13
po0438 <= w41914;-- level 12
po0439 <= w41953;-- level 12
po0440 <= w42012;-- level 33
po0441 <= not w42016;-- level 10
po0442 <= w42034;-- level 36
po0443 <= w42052;-- level 35
po0444 <= w42054;-- level 2
po0445 <= w42061;-- level 32
po0446 <= w42076;-- level 36
po0447 <= w42079;-- level 2
po0448 <= w42082;-- level 2
po0449 <= w42085;-- level 2
po0450 <= w42088;-- level 2
po0451 <= w42091;-- level 2
po0452 <= w42094;-- level 2
po0453 <= w42097;-- level 2
po0454 <= w42100;-- level 2
po0455 <= not w42103;-- level 2
po0456 <= w42111;-- level 26
po0457 <= not w42118;-- level 27
po0458 <= not w42122;-- level 28
po0459 <= w42144;-- level 10
po0460 <= not w42147;-- level 2
po0461 <= not w42150;-- level 2
po0462 <= not w42153;-- level 2
po0463 <= not w42156;-- level 2
po0464 <= not w42159;-- level 2
po0465 <= not w42162;-- level 2
po0466 <= not w42165;-- level 2
po0467 <= not w42192;-- level 13
po0468 <= w42196;-- level 28
po0469 <= w42199;-- level 26
po0470 <= w42206;-- level 24
po0471 <= w42218;-- level 24
po0472 <= not w42223;-- level 32
po0473 <= not w42226;-- level 32
po0474 <= not w42230;-- level 32
po0475 <= not w42235;-- level 32
po0476 <= not w42238;-- level 32
po0477 <= not w42241;-- level 32
po0478 <= not w42244;-- level 32
po0479 <= not w42247;-- level 32
po0480 <= not w42250;-- level 32
po0481 <= not w42253;-- level 32
po0482 <= not w42256;-- level 32
po0483 <= not w42259;-- level 32
po0484 <= not w42262;-- level 32
po0485 <= not w42265;-- level 32
po0486 <= not w42268;-- level 32
po0487 <= not w42276;-- level 32
po0488 <= not w42281;-- level 32
po0489 <= w42293;-- level 28
po0490 <= not w42296;-- level 32
po0491 <= not w42299;-- level 32
po0492 <= not w42302;-- level 32
po0493 <= not w42305;-- level 32
po0494 <= not w42308;-- level 32
po0495 <= not w42311;-- level 32
po0496 <= not w42314;-- level 32
po0497 <= w42320;-- level 32
po0498 <= w42323;-- level 32
po0499 <= not w42326;-- level 32
po0500 <= not w42329;-- level 32
po0501 <= not w42332;-- level 32
po0502 <= not w42335;-- level 32
po0503 <= not w42338;-- level 32
po0504 <= not w42341;-- level 32
po0505 <= not w42344;-- level 32
po0506 <= not w42347;-- level 32
po0507 <= not w42350;-- level 32
po0508 <= not w42353;-- level 32
po0509 <= not w42356;-- level 32
po0510 <= not w42359;-- level 32
po0511 <= not w42362;-- level 32
po0512 <= not w42365;-- level 32
po0513 <= not w42368;-- level 32
po0514 <= not w42371;-- level 32
po0515 <= not w42374;-- level 32
po0516 <= not w42377;-- level 32
po0517 <= not w42380;-- level 32
po0518 <= not w42383;-- level 32
po0519 <= not w42386;-- level 32
po0520 <= not w42389;-- level 32
po0521 <= not w42392;-- level 32
po0522 <= not w42395;-- level 32
po0523 <= not w42398;-- level 32
po0524 <= not w42401;-- level 32
po0525 <= not w42404;-- level 32
po0526 <= not w42407;-- level 32
po0527 <= not w42410;-- level 32
po0528 <= not w42413;-- level 32
po0529 <= not w42416;-- level 32
po0530 <= not w42419;-- level 32
po0531 <= not w42422;-- level 32
po0532 <= not w42425;-- level 32
po0533 <= not w42428;-- level 32
po0534 <= not w42431;-- level 32
po0535 <= not w42434;-- level 32
po0536 <= not w42437;-- level 32
po0537 <= not w42440;-- level 32
po0538 <= not w42443;-- level 32
po0539 <= not w42446;-- level 32
po0540 <= not w42449;-- level 32
po0541 <= not w42452;-- level 32
po0542 <= not w42455;-- level 32
po0543 <= not w42458;-- level 32
po0544 <= not w42461;-- level 32
po0545 <= not w42464;-- level 32
po0546 <= not w42467;-- level 32
po0547 <= not w42470;-- level 32
po0548 <= not w42473;-- level 32
po0549 <= not w42476;-- level 32
po0550 <= not w42479;-- level 32
po0551 <= not w42482;-- level 32
po0552 <= not w42485;-- level 32
po0553 <= not w42488;-- level 32
po0554 <= not w42491;-- level 32
po0555 <= not w42494;-- level 32
po0556 <= not w42497;-- level 32
po0557 <= not w42500;-- level 32
po0558 <= not w42503;-- level 32
po0559 <= not w42506;-- level 32
po0560 <= not w42509;-- level 32
po0561 <= not w42512;-- level 32
po0562 <= not w42515;-- level 32
po0563 <= not w42518;-- level 32
po0564 <= not w42521;-- level 32
po0565 <= not w42524;-- level 32
po0566 <= not w42527;-- level 32
po0567 <= not w42530;-- level 32
po0568 <= not w42533;-- level 32
po0569 <= not w42536;-- level 32
po0570 <= not w42539;-- level 32
po0571 <= not w42543;-- level 32
po0572 <= not w42546;-- level 32
po0573 <= not w42549;-- level 32
po0574 <= not w42552;-- level 32
po0575 <= not w42555;-- level 32
po0576 <= not w42558;-- level 32
po0577 <= not w42561;-- level 32
po0578 <= not w42564;-- level 32
po0579 <= not w42567;-- level 32
po0580 <= not w42570;-- level 32
po0581 <= not w42573;-- level 32
po0582 <= not w42576;-- level 32
po0583 <= not w42579;-- level 32
po0584 <= not w42582;-- level 32
po0585 <= not w42585;-- level 32
po0586 <= not w42588;-- level 32
po0587 <= not w42591;-- level 32
po0588 <= not w42594;-- level 32
po0589 <= not w42597;-- level 32
po0590 <= not w42600;-- level 32
po0591 <= not w42603;-- level 32
po0592 <= not w42606;-- level 32
po0593 <= not w42609;-- level 32
po0594 <= not w42612;-- level 32
po0595 <= not w42615;-- level 32
po0596 <= not w42618;-- level 32
po0597 <= not w42621;-- level 32
po0598 <= not w42624;-- level 32
po0599 <= not w42627;-- level 32
po0600 <= not w42630;-- level 32
po0601 <= not w42633;-- level 32
po0602 <= not w42636;-- level 32
po0603 <= not w42639;-- level 32
po0604 <= not w42642;-- level 32
po0605 <= not w42645;-- level 32
po0606 <= not w42648;-- level 32
po0607 <= not w42651;-- level 32
po0608 <= not w42654;-- level 32
po0609 <= not w42657;-- level 32
po0610 <= not w42660;-- level 32
po0611 <= not w42663;-- level 32
po0612 <= not w42666;-- level 32
po0613 <= not w42669;-- level 32
po0614 <= w42693;-- level 10
po0615 <= not w42696;-- level 32
po0616 <= not w42699;-- level 32
po0617 <= not w42702;-- level 32
po0618 <= not w42705;-- level 32
po0619 <= not w42708;-- level 32
po0620 <= not w42711;-- level 32
po0621 <= not w42714;-- level 32
po0622 <= w42739;-- level 10
po0623 <= w42757;-- level 12
po0624 <= w42787;-- level 28
po0625 <= not w42793;-- level 25
po0626 <= w42813;-- level 10
po0627 <= w42833;-- level 10
po0628 <= w42853;-- level 10
po0629 <= w42873;-- level 10
po0630 <= w42884;-- level 12
po0631 <= w42895;-- level 12
po0632 <= w42906;-- level 12
po0633 <= not w42918;-- level 15
po0634 <= not w42203;-- level 22
po0635 <= w42919;-- level 7
po0636 <= pi0583;-- level 0
po0637 <= w42057;-- level 29
po0638 <= not w42922;-- level 11
po0639 <= not w42925;-- level 11
po0640 <= not w42928;-- level 11
po0641 <= not w42931;-- level 11
po0642 <= not w42934;-- level 11
po0643 <= not w42937;-- level 11
po0644 <= not w42940;-- level 11
po0645 <= w42943;-- level 11
po0646 <= not w42946;-- level 11
po0647 <= not w42949;-- level 11
po0648 <= not w42952;-- level 11
po0649 <= not w42955;-- level 11
po0650 <= not w42958;-- level 11
po0651 <= w42961;-- level 11
po0652 <= not w42964;-- level 11
po0653 <= not w42967;-- level 11
po0654 <= w42970;-- level 11
po0655 <= not w42973;-- level 11
po0656 <= not w42976;-- level 11
po0657 <= not w42979;-- level 11
po0658 <= not w42982;-- level 11
po0659 <= not w42985;-- level 11
po0660 <= not w42988;-- level 11
po0661 <= not w42991;-- level 11
po0662 <= not w43000;-- level 12
po0663 <= not w43003;-- level 11
po0664 <= not w43006;-- level 11
po0665 <= not w43009;-- level 11
po0666 <= not w43012;-- level 11
po0667 <= not w43015;-- level 11
po0668 <= not w43021;-- level 11
po0669 <= not w43024;-- level 11
po0670 <= not w43027;-- level 11
po0671 <= not w43030;-- level 11
po0672 <= not w43033;-- level 11
po0673 <= not w43036;-- level 11
po0674 <= not w43039;-- level 11
po0675 <= not w43045;-- level 12
po0676 <= w43048;-- level 11
po0677 <= not w43051;-- level 11
po0678 <= not w43054;-- level 11
po0679 <= not w43057;-- level 11
po0680 <= not w43062;-- level 12
po0681 <= w43065;-- level 11
po0682 <= not w43068;-- level 11
po0683 <= not w43071;-- level 11
po0684 <= not w43074;-- level 11
po0685 <= not w43077;-- level 11
po0686 <= not w43080;-- level 11
po0687 <= not w43083;-- level 11
po0688 <= not w43086;-- level 11
po0689 <= not w43089;-- level 11
po0690 <= not w43092;-- level 11
po0691 <= w43095;-- level 11
po0692 <= not w43098;-- level 11
po0693 <= not w43101;-- level 11
po0694 <= not w43104;-- level 11
po0695 <= not w43107;-- level 11
po0696 <= not w43110;-- level 11
po0697 <= not w43113;-- level 11
po0698 <= not w43116;-- level 11
po0699 <= not w43119;-- level 11
po0700 <= not w43122;-- level 11
po0701 <= not w43127;-- level 12
po0702 <= not w43130;-- level 11
po0703 <= not w43133;-- level 11
po0704 <= not w43136;-- level 11
po0705 <= not w43139;-- level 11
po0706 <= not w43142;-- level 11
po0707 <= w43145;-- level 11
po0708 <= not w43148;-- level 11
po0709 <= not w43151;-- level 11
po0710 <= not w43154;-- level 11
po0711 <= not w43157;-- level 11
po0712 <= not w43160;-- level 11
po0713 <= not w43163;-- level 11
po0714 <= not w43168;-- level 12
po0715 <= not w43171;-- level 11
po0716 <= not w43174;-- level 11
po0717 <= not w43177;-- level 11
po0718 <= not w43180;-- level 11
po0719 <= not w43183;-- level 11
po0720 <= not w43186;-- level 11
po0721 <= not w43189;-- level 11
po0722 <= not w43192;-- level 11
po0723 <= not w43195;-- level 11
po0724 <= not w43306;-- level 33
po0725 <= not w43309;-- level 11
po0726 <= w43312;-- level 11
po0727 <= not w43317;-- level 12
po0728 <= not w43320;-- level 11
po0729 <= not w43323;-- level 11
po0730 <= not w43326;-- level 11
po0731 <= not w43329;-- level 11
po0732 <= not w43332;-- level 11
po0733 <= not w43335;-- level 11
po0734 <= not w43338;-- level 11
po0735 <= not w43341;-- level 11
po0736 <= not w43344;-- level 11
po0737 <= not w43347;-- level 11
po0738 <= not w43350;-- level 11
po0739 <= not w43353;-- level 11
po0740 <= w3841;-- level 3
po0741 <= not w43356;-- level 11
po0742 <= not w43359;-- level 11
po0743 <= not w43362;-- level 11
po0744 <= not w43369;-- level 8
po0745 <= w43374;-- level 5
po0746 <= w43395;-- level 13
po0747 <= not w43399;-- level 5
po0748 <= w43403;-- level 5
po0749 <= w43407;-- level 5
po0750 <= w44286;-- level 69
po0751 <= w44293;-- level 5
po0752 <= w44299;-- level 7
po0753 <= w44305;-- level 6
po0754 <= w44309;-- level 6
po0755 <= not w44315;-- level 8
po0756 <= w44319;-- level 7
po0757 <= w44322;-- level 4
po0758 <= w44326;-- level 3
po0759 <= not w44338;-- level 8
po0760 <= not w44352;-- level 7
po0761 <= not w44359;-- level 5
po0762 <= w44362;-- level 3
po0763 <= w44368;-- level 8
po0764 <= w44372;-- level 7
po0765 <= w44376;-- level 7
po0766 <= w44380;-- level 7
po0767 <= w44384;-- level 7
po0768 <= w44388;-- level 7
po0769 <= w44392;-- level 7
po0770 <= w44396;-- level 7
po0771 <= not w44401;-- level 8
po0772 <= not w44406;-- level 8
po0773 <= not w44411;-- level 8
po0774 <= w44417;-- level 8
po0775 <= w44421;-- level 7
po0776 <= w44425;-- level 7
po0777 <= w44429;-- level 7
po0778 <= w44433;-- level 7
po0779 <= w44437;-- level 7
po0780 <= w44441;-- level 7
po0781 <= not w44447;-- level 5
po0782 <= w44456;-- level 7
po0783 <= w44460;-- level 7
po0784 <= w44464;-- level 7
po0785 <= w44468;-- level 7
po0786 <= w44472;-- level 7
po0787 <= w44476;-- level 7
po0788 <= w44480;-- level 7
po0789 <= w44484;-- level 7
po0790 <= w44488;-- level 7
po0791 <= w44492;-- level 7
po0792 <= w44496;-- level 7
po0793 <= w44500;-- level 7
po0794 <= w44504;-- level 7
po0795 <= w44508;-- level 7
po0796 <= w44512;-- level 7
po0797 <= w44516;-- level 7
po0798 <= w44520;-- level 7
po0799 <= w44524;-- level 7
po0800 <= w44528;-- level 7
po0801 <= w44532;-- level 7
po0802 <= w44536;-- level 7
po0803 <= w44540;-- level 7
po0804 <= w44544;-- level 7
po0805 <= w44548;-- level 7
po0806 <= w44552;-- level 7
po0807 <= w44556;-- level 7
po0808 <= w44560;-- level 7
po0809 <= w44564;-- level 7
po0810 <= w44568;-- level 7
po0811 <= w44572;-- level 7
po0812 <= w44576;-- level 7
po0813 <= w44580;-- level 7
po0814 <= w44584;-- level 7
po0815 <= w44588;-- level 7
po0816 <= w44600;-- level 9
po0817 <= w44604;-- level 7
po0818 <= w44608;-- level 7
po0819 <= w44612;-- level 7
po0820 <= not w44661;-- level 9
po0821 <= not w44703;-- level 9
po0822 <= w44707;-- level 7
po0823 <= not w44743;-- level 9
po0824 <= not w44780;-- level 9
po0825 <= not w44816;-- level 9
po0826 <= w44820;-- level 7
po0827 <= not w44853;-- level 9
po0828 <= not w44885;-- level 9
po0829 <= not w44921;-- level 9
po0830 <= not w44957;-- level 9
po0831 <= not w44995;-- level 9
po0832 <= not w45031;-- level 9
po0833 <= not w45067;-- level 9
po0834 <= not w45099;-- level 9
po0835 <= not w45131;-- level 9
po0836 <= not w45168;-- level 9
po0837 <= w45172;-- level 7
po0838 <= w45176;-- level 7
po0839 <= not w45208;-- level 9
po0840 <= not w6468;-- level 4
po0841 <= w45213;-- level 7
po0842 <= not w45253;-- level 11
po0843 <= w45257;-- level 7
po0844 <= w45261;-- level 7
po0845 <= w45265;-- level 7
po0846 <= not w45299;-- level 11
po0847 <= w45303;-- level 7
po0848 <= w45307;-- level 7
po0849 <= not w45342;-- level 11
po0850 <= w45346;-- level 7
po0851 <= w45350;-- level 7
po0852 <= w45354;-- level 7
po0853 <= w45358;-- level 7
po0854 <= w45362;-- level 7
po0855 <= w45366;-- level 7
po0856 <= w45370;-- level 7
po0857 <= w45374;-- level 7
po0858 <= w45378;-- level 7
po0859 <= w45382;-- level 7
po0860 <= w45386;-- level 7
po0861 <= w45390;-- level 7
po0862 <= w45394;-- level 7
po0863 <= w45398;-- level 7
po0864 <= not w45434;-- level 9
po0865 <= w45474;-- level 9
po0866 <= w45478;-- level 7
po0867 <= w45482;-- level 7
po0868 <= not w45516;-- level 9
po0869 <= not w45551;-- level 9
po0870 <= not w45585;-- level 9
po0871 <= not w45620;-- level 11
po0872 <= w45624;-- level 7
po0873 <= w45660;-- level 9
po0874 <= not w45694;-- level 9
po0875 <= w45730;-- level 9
po0876 <= not w45764;-- level 9
po0877 <= not w45799;-- level 11
po0878 <= not w45855;-- level 15
po0879 <= not w45890;-- level 9
po0880 <= w45894;-- level 7
po0881 <= w45898;-- level 7
po0882 <= w45902;-- level 7
po0883 <= w45906;-- level 7
po0884 <= w45910;-- level 7
po0885 <= w45914;-- level 7
po0886 <= w45918;-- level 7
po0887 <= w45922;-- level 7
po0888 <= w45939;-- level 13
po0889 <= w45943;-- level 7
po0890 <= w45979;-- level 9
po0891 <= w45983;-- level 7
po0892 <= w45987;-- level 7
po0893 <= w45991;-- level 7
po0894 <= w45995;-- level 7
po0895 <= w45999;-- level 7
po0896 <= not w46006;-- level 7
po0897 <= w44347;-- level 4
po0898 <= not w46010;-- level 7
po0899 <= not w46014;-- level 7
po0900 <= not w46018;-- level 7
po0901 <= not w46022;-- level 7
po0902 <= not w46026;-- level 7
po0903 <= not w46030;-- level 7
po0904 <= w46043;-- level 7
po0905 <= not w46047;-- level 7
po0906 <= not w46051;-- level 7
po0907 <= not w46055;-- level 7
po0908 <= not w46059;-- level 7
po0909 <= not w46063;-- level 7
po0910 <= not w46067;-- level 7
po0911 <= not w46071;-- level 7
po0912 <= not w46075;-- level 7
po0913 <= not w46079;-- level 7
po0914 <= not w46083;-- level 7
po0915 <= not w46087;-- level 7
po0916 <= not w46091;-- level 7
po0917 <= not w46095;-- level 7
po0918 <= not w46099;-- level 7
po0919 <= not w46103;-- level 7
po0920 <= not w46107;-- level 7
po0921 <= not w46111;-- level 7
po0922 <= w46135;-- level 19
po0923 <= not w46139;-- level 7
po0924 <= not w46143;-- level 7
po0925 <= not w46147;-- level 7
po0926 <= not w46164;-- level 14
po0927 <= not w46168;-- level 7
po0928 <= not w46178;-- level 16
po0929 <= not w46182;-- level 7
po0930 <= w46190;-- level 18
po0931 <= not w46194;-- level 7
po0932 <= w46211;-- level 13
po0933 <= not w46215;-- level 7
po0934 <= not w46219;-- level 7
po0935 <= not w46227;-- level 6
po0936 <= not w46228;-- level 7
po0937 <= not w46229;-- level 7
po0938 <= not w46232;-- level 6
po0939 <= not w46234;-- level 6
po0940 <= not w46237;-- level 6
po0941 <= not w46240;-- level 6
po0942 <= not w46243;-- level 6
po0943 <= w46246;-- level 2
po0944 <= not w46249;-- level 6
po0945 <= not w46252;-- level 6
po0946 <= not w46255;-- level 6
po0947 <= not w46258;-- level 6
po0948 <= not w46261;-- level 6
po0949 <= not w46264;-- level 6
po0950 <= not w35951;-- level 6
po0951 <= not w46268;-- level 6
po0952 <= not w46271;-- level 6
po0953 <= w46280;-- level 7
po0954 <= w44452;-- level 4
po0955 <= not w46283;-- level 6
po0956 <= w46286;-- level 6
po0957 <= not w46289;-- level 6
po0958 <= not w46292;-- level 6
po0959 <= w44598;-- level 8
po0960 <= w46295;-- level 6
po0961 <= not w46298;-- level 6
po0962 <= w46302;-- level 7
po0963 <= w46173;-- level 14
po0964 <= not w46305;-- level 6
po0965 <= not w46308;-- level 6
po0966 <= w46311;-- level 6
po0967 <= not w46314;-- level 6
po0968 <= not w46317;-- level 6
po0969 <= w46320;-- level 6
po0970 <= not w46323;-- level 6
po0971 <= w46326;-- level 6
po0972 <= not w46329;-- level 6
po0973 <= not w46332;-- level 6
po0974 <= w46334;-- level 4
po0975 <= not w46336;-- level 5
po0976 <= w46338;-- level 8
po0977 <= w46340;-- level 8
po0978 <= w46112;-- level 9
po0979 <= w46341;-- level 1
po0980 <= w45209;-- level 4
po0981 <= w46345;-- level 5
po0982 <= w46374;-- level 9
po0983 <= w46402;-- level 9
po0984 <= w46430;-- level 9
po0985 <= w46458;-- level 9
po0986 <= w46461;-- level 5
po0987 <= w46463;-- level 5
po0988 <= w46002;-- level 4
po0989 <= w46466;-- level 3
po0990 <= not w46468;-- level 3
po0991 <= w46469;-- level 2
po0992 <= w46471;-- level 6
po0993 <= not w46474;-- level 2
po0994 <= not w46477;-- level 2
po0995 <= not w46480;-- level 2
po0996 <= not w46483;-- level 3
po0997 <= w46484;-- level 7
po0998 <= not w46487;-- level 2
po0999 <= not w46490;-- level 2
po1000 <= not w46493;-- level 2
po1001 <= not w46496;-- level 2
po1002 <= not w46499;-- level 4
po1003 <= not w46502;-- level 2
po1004 <= not w46505;-- level 2
po1005 <= not w46508;-- level 3
po1006 <= not w46511;-- level 2
po1007 <= not w46514;-- level 2
po1008 <= not w46517;-- level 2
po1009 <= not w46520;-- level 2
po1010 <= not w46523;-- level 2
po1011 <= not w46526;-- level 2
po1012 <= not w46529;-- level 2
po1013 <= not w46532;-- level 2
po1014 <= not w46535;-- level 2
po1015 <= not w46538;-- level 2
po1016 <= not w46541;-- level 2
po1017 <= not w46550;-- level 4
po1018 <= not w46553;-- level 4
po1019 <= not w46556;-- level 3
po1020 <= not w46559;-- level 3
po1021 <= not w46562;-- level 2
po1022 <= not w46565;-- level 2
po1023 <= not w46568;-- level 2
po1024 <= not w46571;-- level 2
po1025 <= not w46580;-- level 4
po1026 <= not w46583;-- level 2
po1027 <= not w46586;-- level 2
po1028 <= not w46589;-- level 2
po1029 <= not w46592;-- level 2
po1030 <= not w46595;-- level 2
po1031 <= w46604;-- level 4
po1032 <= not w46607;-- level 2
po1033 <= not w46616;-- level 4
po1034 <= not w46625;-- level 4
po1035 <= not w46634;-- level 4
po1036 <= not w46637;-- level 2
po1037 <= not w46640;-- level 2
po1038 <= not w4989;-- level 4
po1039 <= not w46642;-- level 5
po1040 <= not w46645;-- level 5
po1041 <= not w46648;-- level 5
po1042 <= not w46651;-- level 5
po1043 <= not w46653;-- level 5
po1044 <= not w46656;-- level 5
po1045 <= not w46659;-- level 5
po1046 <= not w46662;-- level 5
po1047 <= not w46665;-- level 5
po1048 <= not w46668;-- level 5
po1049 <= not w4000;-- level 2
po1050 <= not w46671;-- level 5
po1051 <= not w46674;-- level 5
po1052 <= not w46677;-- level 5
po1053 <= pi0067;-- level 0
po1054 <= not w46680;-- level 5
po1055 <= not w46682;-- level 5
po1056 <= not w46685;-- level 5
po1057 <= not w3837;-- level 5
po1058 <= not w46688;-- level 5
po1059 <= not w46691;-- level 5
po1060 <= not w46693;-- level 5
po1061 <= not w46695;-- level 5
po1062 <= not w46698;-- level 5
po1063 <= w46709;-- level 5
po1064 <= not w46711;-- level 5
po1065 <= not w46714;-- level 5
po1066 <= not w46717;-- level 5
po1067 <= not w46720;-- level 5
po1068 <= not w46722;-- level 5
po1069 <= not w46725;-- level 5
po1070 <= w46727;-- level 3
po1071 <= not w46730;-- level 5
po1072 <= not w46732;-- level 5
po1073 <= not w46735;-- level 5
po1074 <= not w46738;-- level 5
po1075 <= not w46741;-- level 5
po1076 <= not w46744;-- level 2
po1077 <= not w46746;-- level 2
po1078 <= w46749;-- level 2
po1079 <= w46752;-- level 2
po1080 <= w46755;-- level 2
po1081 <= w46758;-- level 2
po1082 <= w46761;-- level 2
po1083 <= w46764;-- level 2
po1084 <= w46766;-- level 2
po1085 <= w46769;-- level 2
po1086 <= w46772;-- level 2
po1087 <= w46775;-- level 2
po1088 <= not w46777;-- level 2
po1089 <= not w46779;-- level 2
po1090 <= w46782;-- level 2
po1091 <= not w46784;-- level 2
po1092 <= w46787;-- level 2
po1093 <= w46790;-- level 2
po1094 <= not w46792;-- level 2
po1095 <= w46795;-- level 2
po1096 <= not w46797;-- level 2
po1097 <= w46800;-- level 2
po1098 <= w46803;-- level 2
po1099 <= w46806;-- level 2
po1100 <= not w46809;-- level 2
po1101 <= not w3759;-- level 4
po1102 <= w46810;-- level 2
po1103 <= not w46812;-- level 4
po1104 <= w46814;-- level 2
po1105 <= not w46817;-- level 2
po1106 <= w14451;-- level 3
po1107 <= w46818;-- level 2
po1108 <= pi1134;-- level 0
po1109 <= pi0964;-- level 0
po1110 <= not pi0954;-- level 0
po1111 <= pi0965;-- level 0
po1112 <= not w46820;-- level 2
po1113 <= pi0991;-- level 0
po1114 <= pi0985;-- level 0
po1115 <= w46821;-- level 1
po1116 <= w46822;-- level 1
po1117 <= pi1014;-- level 0
po1118 <= w46823;-- level 1
po1119 <= pi1029;-- level 0
po1120 <= pi1004;-- level 0
po1121 <= pi1007;-- level 0
po1122 <= w46824;-- level 1
po1123 <= pi1135;-- level 0
po1124 <= w46825;-- level 1
po1125 <= w46826;-- level 1
po1126 <= w46827;-- level 1
po1127 <= w46828;-- level 1
po1128 <= w46829;-- level 1
po1129 <= w46830;-- level 1
po1130 <= not pi0278;-- level 0
po1131 <= w46831;-- level 1
po1132 <= w46832;-- level 1
po1133 <= not w46833;-- level 1
po1134 <= pi1064;-- level 0
po1135 <= w46834;-- level 1
po1136 <= pi0299;-- level 0
po1137 <= not w46835;-- level 1
po1138 <= pi1075;-- level 0
po1139 <= pi1052;-- level 0
po1140 <= pi0771;-- level 0
po1141 <= pi0765;-- level 0
po1142 <= pi0605;-- level 0
po1143 <= pi0601;-- level 0
po1144 <= pi0278;-- level 0
po1145 <= pi0279;-- level 0
po1146 <= not pi0915;-- level 0
po1147 <= not pi0825;-- level 0
po1148 <= not pi0826;-- level 0
po1149 <= not pi0913;-- level 0
po1150 <= not pi0894;-- level 0
po1151 <= not pi0905;-- level 0
po1152 <= pi1095;-- level 0
po1153 <= not pi0890;-- level 0
po1154 <= pi1094;-- level 0
po1155 <= not pi0906;-- level 0
po1156 <= not pi0896;-- level 0
po1157 <= not pi0909;-- level 0
po1158 <= not pi0911;-- level 0
po1159 <= not pi0908;-- level 0
po1160 <= not pi0891;-- level 0
po1161 <= not pi0902;-- level 0
po1162 <= not pi0903;-- level 0
po1163 <= not pi0883;-- level 0
po1164 <= not pi0888;-- level 0
po1165 <= not pi0919;-- level 0
po1166 <= not pi0886;-- level 0
po1167 <= not pi0912;-- level 0
po1168 <= not pi0895;-- level 0
po1169 <= not pi0916;-- level 0
po1170 <= not pi0889;-- level 0
po1171 <= not pi0900;-- level 0
po1172 <= not pi0885;-- level 0
po1173 <= not pi0904;-- level 0
po1174 <= not pi0899;-- level 0
po1175 <= not pi0918;-- level 0
po1176 <= not pi0898;-- level 0
po1177 <= not pi0917;-- level 0
po1178 <= not pi0827;-- level 0
po1179 <= not pi0887;-- level 0
po1180 <= not pi0884;-- level 0
po1181 <= not pi0910;-- level 0
po1182 <= not pi0828;-- level 0
po1183 <= not pi0892;-- level 0
po1184 <= pi1187;-- level 0
po1185 <= pi1172;-- level 0
po1186 <= pi1170;-- level 0
po1187 <= pi1138;-- level 0
po1188 <= pi1177;-- level 0
po1189 <= pi1178;-- level 0
po1190 <= pi0863;-- level 0
po1191 <= pi1203;-- level 0
po1192 <= pi1185;-- level 0
po1193 <= pi1171;-- level 0
po1194 <= pi1192;-- level 0
po1195 <= pi1137;-- level 0
po1196 <= pi1186;-- level 0
po1197 <= pi1165;-- level 0
po1198 <= pi1164;-- level 0
po1199 <= pi1098;-- level 0
po1200 <= pi1183;-- level 0
po1201 <= pi0230;-- level 0
po1202 <= pi1169;-- level 0
po1203 <= pi1136;-- level 0
po1204 <= pi1181;-- level 0
po1205 <= pi0849;-- level 0
po1206 <= pi1193;-- level 0
po1207 <= pi1182;-- level 0
po1208 <= pi1168;-- level 0
po1209 <= pi1175;-- level 0
po1210 <= pi1191;-- level 0
po1211 <= pi1099;-- level 0
po1212 <= pi1174;-- level 0
po1213 <= pi1179;-- level 0
po1214 <= pi1202;-- level 0
po1215 <= pi1176;-- level 0
po1216 <= pi1173;-- level 0
po1217 <= pi1201;-- level 0
po1218 <= pi1167;-- level 0
po1219 <= pi0840;-- level 0
po1220 <= pi1189;-- level 0
po1221 <= pi1195;-- level 0
po1222 <= pi0864;-- level 0
po1223 <= pi1190;-- level 0
po1224 <= pi1188;-- level 0
po1225 <= pi1180;-- level 0
po1226 <= pi1194;-- level 0
po1227 <= pi1097;-- level 0
po1228 <= pi1166;-- level 0
po1229 <= pi1200;-- level 0
po1230 <= pi1184;-- level 0
end Behavioral;
