library ieee;
use ieee.std_logic_1164.all;

entity top is
 port(count: in std_logic_vector(7 downto 0);
 selectp1: out std_logic_vector(127 downto 0);
 selectp2: out std_logic_vector(127 downto 0));
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303: std_logic;

begin

w0 <= not count(4) and not count(5);
w1 <= not count(6) and count(7);
w2 <= w0 and w1;
w3 <= not count(0) and not count(2);
w4 <= not count(1) and not count(3);
w5 <= w3 and w4;
w6 <= w2 and w5;
w7 <= count(0) and not count(2);
w8 <= w4 and w7;
w9 <= w2 and w8;
w10 <= count(1) and not count(3);
w11 <= w3 and w10;
w12 <= w2 and w11;
w13 <= w7 and w10;
w14 <= w2 and w13;
w15 <= not count(0) and count(2);
w16 <= w4 and w15;
w17 <= w2 and w16;
w18 <= count(0) and count(2);
w19 <= w4 and w18;
w20 <= w2 and w19;
w21 <= w10 and w15;
w22 <= w2 and w21;
w23 <= w10 and w18;
w24 <= w2 and w23;
w25 <= not count(1) and count(3);
w26 <= w3 and w25;
w27 <= w2 and w26;
w28 <= w7 and w25;
w29 <= w2 and w28;
w30 <= count(1) and count(3);
w31 <= w3 and w30;
w32 <= w2 and w31;
w33 <= w7 and w30;
w34 <= w2 and w33;
w35 <= w15 and w25;
w36 <= w2 and w35;
w37 <= w18 and w25;
w38 <= w2 and w37;
w39 <= w15 and w30;
w40 <= w2 and w39;
w41 <= w18 and w30;
w42 <= w2 and w41;
w43 <= count(4) and not count(5);
w44 <= w1 and w43;
w45 <= w5 and w44;
w46 <= w8 and w44;
w47 <= w11 and w44;
w48 <= w13 and w44;
w49 <= w16 and w44;
w50 <= w19 and w44;
w51 <= w21 and w44;
w52 <= w23 and w44;
w53 <= w26 and w44;
w54 <= w28 and w44;
w55 <= w31 and w44;
w56 <= w33 and w44;
w57 <= w35 and w44;
w58 <= w37 and w44;
w59 <= w39 and w44;
w60 <= w41 and w44;
w61 <= not count(4) and count(5);
w62 <= w1 and w61;
w63 <= w5 and w62;
w64 <= w8 and w62;
w65 <= w11 and w62;
w66 <= w13 and w62;
w67 <= w16 and w62;
w68 <= w19 and w62;
w69 <= w21 and w62;
w70 <= w23 and w62;
w71 <= w26 and w62;
w72 <= w28 and w62;
w73 <= w31 and w62;
w74 <= w33 and w62;
w75 <= w35 and w62;
w76 <= w37 and w62;
w77 <= w39 and w62;
w78 <= w41 and w62;
w79 <= count(4) and count(5);
w80 <= w1 and w79;
w81 <= w5 and w80;
w82 <= w8 and w80;
w83 <= w11 and w80;
w84 <= w13 and w80;
w85 <= w16 and w80;
w86 <= w19 and w80;
w87 <= w21 and w80;
w88 <= w23 and w80;
w89 <= w26 and w80;
w90 <= w28 and w80;
w91 <= w31 and w80;
w92 <= w33 and w80;
w93 <= w35 and w80;
w94 <= w37 and w80;
w95 <= w39 and w80;
w96 <= w41 and w80;
w97 <= count(6) and count(7);
w98 <= w0 and w97;
w99 <= w5 and w98;
w100 <= w8 and w98;
w101 <= w11 and w98;
w102 <= w13 and w98;
w103 <= w16 and w98;
w104 <= w19 and w98;
w105 <= w21 and w98;
w106 <= w23 and w98;
w107 <= w26 and w98;
w108 <= w28 and w98;
w109 <= w31 and w98;
w110 <= w33 and w98;
w111 <= w35 and w98;
w112 <= w37 and w98;
w113 <= w39 and w98;
w114 <= w41 and w98;
w115 <= w43 and w97;
w116 <= w5 and w115;
w117 <= w8 and w115;
w118 <= w11 and w115;
w119 <= w13 and w115;
w120 <= w16 and w115;
w121 <= w19 and w115;
w122 <= w21 and w115;
w123 <= w23 and w115;
w124 <= w26 and w115;
w125 <= w28 and w115;
w126 <= w31 and w115;
w127 <= w33 and w115;
w128 <= w35 and w115;
w129 <= w37 and w115;
w130 <= w39 and w115;
w131 <= w41 and w115;
w132 <= w61 and w97;
w133 <= w5 and w132;
w134 <= w8 and w132;
w135 <= w11 and w132;
w136 <= w13 and w132;
w137 <= w16 and w132;
w138 <= w19 and w132;
w139 <= w21 and w132;
w140 <= w23 and w132;
w141 <= w26 and w132;
w142 <= w28 and w132;
w143 <= w31 and w132;
w144 <= w33 and w132;
w145 <= w35 and w132;
w146 <= w37 and w132;
w147 <= w39 and w132;
w148 <= w41 and w132;
w149 <= w79 and w97;
w150 <= w5 and w149;
w151 <= w8 and w149;
w152 <= w11 and w149;
w153 <= w13 and w149;
w154 <= w16 and w149;
w155 <= w19 and w149;
w156 <= w21 and w149;
w157 <= w23 and w149;
w158 <= w26 and w149;
w159 <= w28 and w149;
w160 <= w31 and w149;
w161 <= w33 and w149;
w162 <= w35 and w149;
w163 <= w37 and w149;
w164 <= w39 and w149;
w165 <= w41 and w149;
w166 <= not count(6) and not count(7);
w167 <= w0 and w166;
w168 <= w5 and w167;
w169 <= w8 and w167;
w170 <= w11 and w167;
w171 <= w13 and w167;
w172 <= w16 and w167;
w173 <= w19 and w167;
w174 <= w21 and w167;
w175 <= w23 and w167;
w176 <= w26 and w167;
w177 <= w28 and w167;
w178 <= w31 and w167;
w179 <= w33 and w167;
w180 <= w35 and w167;
w181 <= w37 and w167;
w182 <= w39 and w167;
w183 <= w41 and w167;
w184 <= w43 and w166;
w185 <= w5 and w184;
w186 <= w8 and w184;
w187 <= w11 and w184;
w188 <= w13 and w184;
w189 <= w16 and w184;
w190 <= w19 and w184;
w191 <= w21 and w184;
w192 <= w23 and w184;
w193 <= w26 and w184;
w194 <= w28 and w184;
w195 <= w31 and w184;
w196 <= w33 and w184;
w197 <= w35 and w184;
w198 <= w37 and w184;
w199 <= w39 and w184;
w200 <= w41 and w184;
w201 <= w61 and w166;
w202 <= w5 and w201;
w203 <= w8 and w201;
w204 <= w11 and w201;
w205 <= w13 and w201;
w206 <= w16 and w201;
w207 <= w19 and w201;
w208 <= w21 and w201;
w209 <= w23 and w201;
w210 <= w26 and w201;
w211 <= w28 and w201;
w212 <= w31 and w201;
w213 <= w33 and w201;
w214 <= w35 and w201;
w215 <= w37 and w201;
w216 <= w39 and w201;
w217 <= w41 and w201;
w218 <= w79 and w166;
w219 <= w5 and w218;
w220 <= w8 and w218;
w221 <= w11 and w218;
w222 <= w13 and w218;
w223 <= w16 and w218;
w224 <= w19 and w218;
w225 <= w21 and w218;
w226 <= w23 and w218;
w227 <= w26 and w218;
w228 <= w28 and w218;
w229 <= w31 and w218;
w230 <= w33 and w218;
w231 <= w35 and w218;
w232 <= w37 and w218;
w233 <= w39 and w218;
w234 <= w41 and w218;
w235 <= count(6) and not count(7);
w236 <= w0 and w235;
w237 <= w5 and w236;
w238 <= w8 and w236;
w239 <= w11 and w236;
w240 <= w13 and w236;
w241 <= w16 and w236;
w242 <= w19 and w236;
w243 <= w21 and w236;
w244 <= w23 and w236;
w245 <= w26 and w236;
w246 <= w28 and w236;
w247 <= w31 and w236;
w248 <= w33 and w236;
w249 <= w35 and w236;
w250 <= w37 and w236;
w251 <= w39 and w236;
w252 <= w41 and w236;
w253 <= w43 and w235;
w254 <= w5 and w253;
w255 <= w8 and w253;
w256 <= w11 and w253;
w257 <= w13 and w253;
w258 <= w16 and w253;
w259 <= w19 and w253;
w260 <= w21 and w253;
w261 <= w23 and w253;
w262 <= w26 and w253;
w263 <= w28 and w253;
w264 <= w31 and w253;
w265 <= w33 and w253;
w266 <= w35 and w253;
w267 <= w37 and w253;
w268 <= w39 and w253;
w269 <= w41 and w253;
w270 <= w61 and w235;
w271 <= w5 and w270;
w272 <= w8 and w270;
w273 <= w11 and w270;
w274 <= w13 and w270;
w275 <= w16 and w270;
w276 <= w19 and w270;
w277 <= w21 and w270;
w278 <= w23 and w270;
w279 <= w26 and w270;
w280 <= w28 and w270;
w281 <= w31 and w270;
w282 <= w33 and w270;
w283 <= w35 and w270;
w284 <= w37 and w270;
w285 <= w39 and w270;
w286 <= w41 and w270;
w287 <= w79 and w235;
w288 <= w5 and w287;
w289 <= w8 and w287;
w290 <= w11 and w287;
w291 <= w13 and w287;
w292 <= w16 and w287;
w293 <= w19 and w287;
w294 <= w21 and w287;
w295 <= w23 and w287;
w296 <= w26 and w287;
w297 <= w28 and w287;
w298 <= w31 and w287;
w299 <= w33 and w287;
w300 <= w35 and w287;
w301 <= w37 and w287;
w302 <= w39 and w287;
w303 <= w41 and w287;
one <= '1';
selectp1(0) <= w6;-- level 3
selectp1(1) <= w9;-- level 3
selectp1(2) <= w12;-- level 3
selectp1(3) <= w14;-- level 3
selectp1(4) <= w17;-- level 3
selectp1(5) <= w20;-- level 3
selectp1(6) <= w22;-- level 3
selectp1(7) <= w24;-- level 3
selectp1(8) <= w27;-- level 3
selectp1(9) <= w29;-- level 3
selectp1(10) <= w32;-- level 3
selectp1(11) <= w34;-- level 3
selectp1(12) <= w36;-- level 3
selectp1(13) <= w38;-- level 3
selectp1(14) <= w40;-- level 3
selectp1(15) <= w42;-- level 3
selectp1(16) <= w45;-- level 3
selectp1(17) <= w46;-- level 3
selectp1(18) <= w47;-- level 3
selectp1(19) <= w48;-- level 3
selectp1(20) <= w49;-- level 3
selectp1(21) <= w50;-- level 3
selectp1(22) <= w51;-- level 3
selectp1(23) <= w52;-- level 3
selectp1(24) <= w53;-- level 3
selectp1(25) <= w54;-- level 3
selectp1(26) <= w55;-- level 3
selectp1(27) <= w56;-- level 3
selectp1(28) <= w57;-- level 3
selectp1(29) <= w58;-- level 3
selectp1(30) <= w59;-- level 3
selectp1(31) <= w60;-- level 3
selectp1(32) <= w63;-- level 3
selectp1(33) <= w64;-- level 3
selectp1(34) <= w65;-- level 3
selectp1(35) <= w66;-- level 3
selectp1(36) <= w67;-- level 3
selectp1(37) <= w68;-- level 3
selectp1(38) <= w69;-- level 3
selectp1(39) <= w70;-- level 3
selectp1(40) <= w71;-- level 3
selectp1(41) <= w72;-- level 3
selectp1(42) <= w73;-- level 3
selectp1(43) <= w74;-- level 3
selectp1(44) <= w75;-- level 3
selectp1(45) <= w76;-- level 3
selectp1(46) <= w77;-- level 3
selectp1(47) <= w78;-- level 3
selectp1(48) <= w81;-- level 3
selectp1(49) <= w82;-- level 3
selectp1(50) <= w83;-- level 3
selectp1(51) <= w84;-- level 3
selectp1(52) <= w85;-- level 3
selectp1(53) <= w86;-- level 3
selectp1(54) <= w87;-- level 3
selectp1(55) <= w88;-- level 3
selectp1(56) <= w89;-- level 3
selectp1(57) <= w90;-- level 3
selectp1(58) <= w91;-- level 3
selectp1(59) <= w92;-- level 3
selectp1(60) <= w93;-- level 3
selectp1(61) <= w94;-- level 3
selectp1(62) <= w95;-- level 3
selectp1(63) <= w96;-- level 3
selectp1(64) <= w99;-- level 3
selectp1(65) <= w100;-- level 3
selectp1(66) <= w101;-- level 3
selectp1(67) <= w102;-- level 3
selectp1(68) <= w103;-- level 3
selectp1(69) <= w104;-- level 3
selectp1(70) <= w105;-- level 3
selectp1(71) <= w106;-- level 3
selectp1(72) <= w107;-- level 3
selectp1(73) <= w108;-- level 3
selectp1(74) <= w109;-- level 3
selectp1(75) <= w110;-- level 3
selectp1(76) <= w111;-- level 3
selectp1(77) <= w112;-- level 3
selectp1(78) <= w113;-- level 3
selectp1(79) <= w114;-- level 3
selectp1(80) <= w116;-- level 3
selectp1(81) <= w117;-- level 3
selectp1(82) <= w118;-- level 3
selectp1(83) <= w119;-- level 3
selectp1(84) <= w120;-- level 3
selectp1(85) <= w121;-- level 3
selectp1(86) <= w122;-- level 3
selectp1(87) <= w123;-- level 3
selectp1(88) <= w124;-- level 3
selectp1(89) <= w125;-- level 3
selectp1(90) <= w126;-- level 3
selectp1(91) <= w127;-- level 3
selectp1(92) <= w128;-- level 3
selectp1(93) <= w129;-- level 3
selectp1(94) <= w130;-- level 3
selectp1(95) <= w131;-- level 3
selectp1(96) <= w133;-- level 3
selectp1(97) <= w134;-- level 3
selectp1(98) <= w135;-- level 3
selectp1(99) <= w136;-- level 3
selectp1(100) <= w137;-- level 3
selectp1(101) <= w138;-- level 3
selectp1(102) <= w139;-- level 3
selectp1(103) <= w140;-- level 3
selectp1(104) <= w141;-- level 3
selectp1(105) <= w142;-- level 3
selectp1(106) <= w143;-- level 3
selectp1(107) <= w144;-- level 3
selectp1(108) <= w145;-- level 3
selectp1(109) <= w146;-- level 3
selectp1(110) <= w147;-- level 3
selectp1(111) <= w148;-- level 3
selectp1(112) <= w150;-- level 3
selectp1(113) <= w151;-- level 3
selectp1(114) <= w152;-- level 3
selectp1(115) <= w153;-- level 3
selectp1(116) <= w154;-- level 3
selectp1(117) <= w155;-- level 3
selectp1(118) <= w156;-- level 3
selectp1(119) <= w157;-- level 3
selectp1(120) <= w158;-- level 3
selectp1(121) <= w159;-- level 3
selectp1(122) <= w160;-- level 3
selectp1(123) <= w161;-- level 3
selectp1(124) <= w162;-- level 3
selectp1(125) <= w163;-- level 3
selectp1(126) <= w164;-- level 3
selectp1(127) <= w165;-- level 3
selectp2(0) <= w168;-- level 3
selectp2(1) <= w169;-- level 3
selectp2(2) <= w170;-- level 3
selectp2(3) <= w171;-- level 3
selectp2(4) <= w172;-- level 3
selectp2(5) <= w173;-- level 3
selectp2(6) <= w174;-- level 3
selectp2(7) <= w175;-- level 3
selectp2(8) <= w176;-- level 3
selectp2(9) <= w177;-- level 3
selectp2(10) <= w178;-- level 3
selectp2(11) <= w179;-- level 3
selectp2(12) <= w180;-- level 3
selectp2(13) <= w181;-- level 3
selectp2(14) <= w182;-- level 3
selectp2(15) <= w183;-- level 3
selectp2(16) <= w185;-- level 3
selectp2(17) <= w186;-- level 3
selectp2(18) <= w187;-- level 3
selectp2(19) <= w188;-- level 3
selectp2(20) <= w189;-- level 3
selectp2(21) <= w190;-- level 3
selectp2(22) <= w191;-- level 3
selectp2(23) <= w192;-- level 3
selectp2(24) <= w193;-- level 3
selectp2(25) <= w194;-- level 3
selectp2(26) <= w195;-- level 3
selectp2(27) <= w196;-- level 3
selectp2(28) <= w197;-- level 3
selectp2(29) <= w198;-- level 3
selectp2(30) <= w199;-- level 3
selectp2(31) <= w200;-- level 3
selectp2(32) <= w202;-- level 3
selectp2(33) <= w203;-- level 3
selectp2(34) <= w204;-- level 3
selectp2(35) <= w205;-- level 3
selectp2(36) <= w206;-- level 3
selectp2(37) <= w207;-- level 3
selectp2(38) <= w208;-- level 3
selectp2(39) <= w209;-- level 3
selectp2(40) <= w210;-- level 3
selectp2(41) <= w211;-- level 3
selectp2(42) <= w212;-- level 3
selectp2(43) <= w213;-- level 3
selectp2(44) <= w214;-- level 3
selectp2(45) <= w215;-- level 3
selectp2(46) <= w216;-- level 3
selectp2(47) <= w217;-- level 3
selectp2(48) <= w219;-- level 3
selectp2(49) <= w220;-- level 3
selectp2(50) <= w221;-- level 3
selectp2(51) <= w222;-- level 3
selectp2(52) <= w223;-- level 3
selectp2(53) <= w224;-- level 3
selectp2(54) <= w225;-- level 3
selectp2(55) <= w226;-- level 3
selectp2(56) <= w227;-- level 3
selectp2(57) <= w228;-- level 3
selectp2(58) <= w229;-- level 3
selectp2(59) <= w230;-- level 3
selectp2(60) <= w231;-- level 3
selectp2(61) <= w232;-- level 3
selectp2(62) <= w233;-- level 3
selectp2(63) <= w234;-- level 3
selectp2(64) <= w237;-- level 3
selectp2(65) <= w238;-- level 3
selectp2(66) <= w239;-- level 3
selectp2(67) <= w240;-- level 3
selectp2(68) <= w241;-- level 3
selectp2(69) <= w242;-- level 3
selectp2(70) <= w243;-- level 3
selectp2(71) <= w244;-- level 3
selectp2(72) <= w245;-- level 3
selectp2(73) <= w246;-- level 3
selectp2(74) <= w247;-- level 3
selectp2(75) <= w248;-- level 3
selectp2(76) <= w249;-- level 3
selectp2(77) <= w250;-- level 3
selectp2(78) <= w251;-- level 3
selectp2(79) <= w252;-- level 3
selectp2(80) <= w254;-- level 3
selectp2(81) <= w255;-- level 3
selectp2(82) <= w256;-- level 3
selectp2(83) <= w257;-- level 3
selectp2(84) <= w258;-- level 3
selectp2(85) <= w259;-- level 3
selectp2(86) <= w260;-- level 3
selectp2(87) <= w261;-- level 3
selectp2(88) <= w262;-- level 3
selectp2(89) <= w263;-- level 3
selectp2(90) <= w264;-- level 3
selectp2(91) <= w265;-- level 3
selectp2(92) <= w266;-- level 3
selectp2(93) <= w267;-- level 3
selectp2(94) <= w268;-- level 3
selectp2(95) <= w269;-- level 3
selectp2(96) <= w271;-- level 3
selectp2(97) <= w272;-- level 3
selectp2(98) <= w273;-- level 3
selectp2(99) <= w274;-- level 3
selectp2(100) <= w275;-- level 3
selectp2(101) <= w276;-- level 3
selectp2(102) <= w277;-- level 3
selectp2(103) <= w278;-- level 3
selectp2(104) <= w279;-- level 3
selectp2(105) <= w280;-- level 3
selectp2(106) <= w281;-- level 3
selectp2(107) <= w282;-- level 3
selectp2(108) <= w283;-- level 3
selectp2(109) <= w284;-- level 3
selectp2(110) <= w285;-- level 3
selectp2(111) <= w286;-- level 3
selectp2(112) <= w288;-- level 3
selectp2(113) <= w289;-- level 3
selectp2(114) <= w290;-- level 3
selectp2(115) <= w291;-- level 3
selectp2(116) <= w292;-- level 3
selectp2(117) <= w293;-- level 3
selectp2(118) <= w294;-- level 3
selectp2(119) <= w295;-- level 3
selectp2(120) <= w296;-- level 3
selectp2(121) <= w297;-- level 3
selectp2(122) <= w298;-- level 3
selectp2(123) <= w299;-- level 3
selectp2(124) <= w300;-- level 3
selectp2(125) <= w301;-- level 3
selectp2(126) <= w302;-- level 3
selectp2(127) <= w303;-- level 3
end Behavioral;
