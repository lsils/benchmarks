module top ( 
    \dest_x[0] , \dest_x[1] , \dest_x[2] , \dest_x[3] , \dest_x[4] ,
    \dest_x[5] , \dest_x[6] , \dest_x[7] , \dest_x[8] , \dest_x[9] ,
    \dest_x[10] , \dest_x[11] , \dest_x[12] , \dest_x[13] , \dest_x[14] ,
    \dest_x[15] , \dest_x[16] , \dest_x[17] , \dest_x[18] , \dest_x[19] ,
    \dest_x[20] , \dest_x[21] , \dest_x[22] , \dest_x[23] , \dest_x[24] ,
    \dest_x[25] , \dest_x[26] , \dest_x[27] , \dest_x[28] , \dest_x[29] ,
    \dest_y[0] , \dest_y[1] , \dest_y[2] , \dest_y[3] , \dest_y[4] ,
    \dest_y[5] , \dest_y[6] , \dest_y[7] , \dest_y[8] , \dest_y[9] ,
    \dest_y[10] , \dest_y[11] , \dest_y[12] , \dest_y[13] , \dest_y[14] ,
    \dest_y[15] , \dest_y[16] , \dest_y[17] , \dest_y[18] , \dest_y[19] ,
    \dest_y[20] , \dest_y[21] , \dest_y[22] , \dest_y[23] , \dest_y[24] ,
    \dest_y[25] , \dest_y[26] , \dest_y[27] , \dest_y[28] , \dest_y[29] ,
    \outport[0] , \outport[1] , \outport[2] , \outport[3] , \outport[4] ,
    \outport[5] , \outport[6] , \outport[7] , \outport[8] , \outport[9] ,
    \outport[10] , \outport[11] , \outport[12] , \outport[13] ,
    \outport[14] , \outport[15] , \outport[16] , \outport[17] ,
    \outport[18] , \outport[19] , \outport[20] , \outport[21] ,
    \outport[22] , \outport[23] , \outport[24] , \outport[25] ,
    \outport[26] , \outport[27] , \outport[28] , \outport[29]   );
  input  \dest_x[0] , \dest_x[1] , \dest_x[2] , \dest_x[3] , \dest_x[4] ,
    \dest_x[5] , \dest_x[6] , \dest_x[7] , \dest_x[8] , \dest_x[9] ,
    \dest_x[10] , \dest_x[11] , \dest_x[12] , \dest_x[13] , \dest_x[14] ,
    \dest_x[15] , \dest_x[16] , \dest_x[17] , \dest_x[18] , \dest_x[19] ,
    \dest_x[20] , \dest_x[21] , \dest_x[22] , \dest_x[23] , \dest_x[24] ,
    \dest_x[25] , \dest_x[26] , \dest_x[27] , \dest_x[28] , \dest_x[29] ,
    \dest_y[0] , \dest_y[1] , \dest_y[2] , \dest_y[3] , \dest_y[4] ,
    \dest_y[5] , \dest_y[6] , \dest_y[7] , \dest_y[8] , \dest_y[9] ,
    \dest_y[10] , \dest_y[11] , \dest_y[12] , \dest_y[13] , \dest_y[14] ,
    \dest_y[15] , \dest_y[16] , \dest_y[17] , \dest_y[18] , \dest_y[19] ,
    \dest_y[20] , \dest_y[21] , \dest_y[22] , \dest_y[23] , \dest_y[24] ,
    \dest_y[25] , \dest_y[26] , \dest_y[27] , \dest_y[28] , \dest_y[29] ;
  output \outport[0] , \outport[1] , \outport[2] , \outport[3] , \outport[4] ,
    \outport[5] , \outport[6] , \outport[7] , \outport[8] , \outport[9] ,
    \outport[10] , \outport[11] , \outport[12] , \outport[13] ,
    \outport[14] , \outport[15] , \outport[16] , \outport[17] ,
    \outport[18] , \outport[19] , \outport[20] , \outport[21] ,
    \outport[22] , \outport[23] , \outport[24] , \outport[25] ,
    \outport[26] , \outport[27] , \outport[28] , \outport[29] ;
  wire n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
    n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n345, n346,
    n347;
  assign n92 = ~\dest_x[9]  & ~\dest_x[10] ;
  assign n93 = \dest_x[9]  & \dest_x[10] ;
  assign n94 = ~n92 & ~n93;
  assign n95 = \dest_x[11]  & ~n92;
  assign n96 = ~\dest_x[11]  & n92;
  assign n97 = ~n95 & ~n96;
  assign n98 = ~\dest_x[12]  & ~n95;
  assign n99 = \dest_x[12]  & n95;
  assign n100 = ~n98 & ~n99;
  assign n101 = ~\dest_x[13]  & n98;
  assign n102 = \dest_x[13]  & ~n98;
  assign n103 = ~n101 & ~n102;
  assign n104 = \dest_x[14]  & ~n101;
  assign n105 = ~\dest_x[14]  & n101;
  assign n106 = ~n104 & ~n105;
  assign n107 = \dest_x[15]  & ~n104;
  assign n108 = ~\dest_x[15]  & n104;
  assign n109 = ~n107 & ~n108;
  assign n110 = \dest_x[15]  & n104;
  assign n111 = ~\dest_x[16]  & ~n110;
  assign n112 = \dest_x[16]  & n110;
  assign n113 = ~n111 & ~n112;
  assign n114 = \dest_x[17]  & ~n111;
  assign n115 = ~\dest_x[17]  & n111;
  assign n116 = ~n114 & ~n115;
  assign n117 = ~\dest_x[18]  & ~n114;
  assign n118 = \dest_x[18]  & n114;
  assign n119 = ~n117 & ~n118;
  assign n120 = \dest_x[19]  & ~n117;
  assign n121 = ~\dest_x[19]  & n117;
  assign n122 = ~n120 & ~n121;
  assign n123 = \dest_x[20]  & ~n120;
  assign n124 = ~\dest_x[20]  & n120;
  assign n125 = ~n123 & ~n124;
  assign n126 = \dest_x[20]  & n120;
  assign n127 = ~\dest_x[21]  & ~n126;
  assign n128 = \dest_x[21]  & n126;
  assign n129 = ~n127 & ~n128;
  assign n130 = ~\dest_x[22]  & n127;
  assign n131 = \dest_x[22]  & ~n127;
  assign n132 = ~n130 & ~n131;
  assign n133 = \dest_x[23]  & ~n130;
  assign n134 = ~\dest_x[23]  & n130;
  assign n135 = ~n133 & ~n134;
  assign n136 = \dest_x[24]  & ~n133;
  assign n137 = ~\dest_x[24]  & n133;
  assign n138 = ~n136 & ~n137;
  assign n139 = \dest_x[24]  & n133;
  assign n140 = \dest_x[25]  & ~n139;
  assign n141 = ~\dest_x[25]  & n139;
  assign n142 = ~n140 & ~n141;
  assign n143 = \dest_x[25]  & n139;
  assign n144 = ~\dest_x[26]  & ~n143;
  assign n145 = \dest_x[26]  & n143;
  assign n146 = ~n144 & ~n145;
  assign n147 = \dest_x[27]  & ~n144;
  assign n148 = ~\dest_x[27]  & n144;
  assign n149 = ~n147 & ~n148;
  assign n150 = \dest_x[28]  & ~n147;
  assign n151 = ~\dest_x[28]  & n147;
  assign n152 = ~n150 & ~n151;
  assign n153 = \dest_x[28]  & n147;
  assign n154 = ~\dest_x[29]  & n153;
  assign n155 = \dest_x[29]  & ~n153;
  assign n156 = ~n154 & ~n155;
  assign n157 = ~\dest_x[9]  & ~n156;
  assign n158 = ~n152 & n157;
  assign n159 = n149 & n158;
  assign n160 = ~n146 & n159;
  assign n161 = ~n142 & n160;
  assign n162 = ~n138 & n161;
  assign n163 = n135 & n162;
  assign n164 = ~n132 & n163;
  assign n165 = ~n129 & n164;
  assign n166 = ~n125 & n165;
  assign n167 = n122 & n166;
  assign n168 = ~n119 & n167;
  assign n169 = n116 & n168;
  assign n170 = ~n113 & n169;
  assign n171 = ~n109 & n170;
  assign n172 = n106 & n171;
  assign n173 = ~n103 & n172;
  assign n174 = ~n100 & n173;
  assign n175 = n97 & n174;
  assign n176 = ~n94 & n175;
  assign n177 = \dest_x[8]  & n176;
  assign n178 = \dest_x[7]  & n177;
  assign n179 = \dest_x[6]  & n178;
  assign n180 = \dest_x[5]  & n179;
  assign n181 = \dest_x[4]  & n180;
  assign n182 = \dest_x[3]  & n181;
  assign n183 = \dest_x[2]  & n182;
  assign n184 = \dest_x[1]  & n183;
  assign n185 = \dest_x[0]  & n184;
  assign n186 = \dest_x[29]  & n153;
  assign n187 = ~n185 & ~n186;
  assign n188 = ~\dest_x[1]  & ~\dest_x[2] ;
  assign n189 = ~\dest_x[3]  & n188;
  assign n190 = ~\dest_x[4]  & n189;
  assign n191 = ~\dest_x[5]  & n190;
  assign n192 = ~\dest_x[6]  & n191;
  assign n193 = ~\dest_x[7]  & n192;
  assign n194 = ~\dest_x[8]  & n193;
  assign n195 = n94 & n194;
  assign n196 = ~n97 & n195;
  assign n197 = n100 & n196;
  assign n198 = n103 & n197;
  assign n199 = ~n106 & n198;
  assign n200 = n109 & n199;
  assign n201 = n113 & n200;
  assign n202 = ~n116 & n201;
  assign n203 = n119 & n202;
  assign n204 = ~n122 & n203;
  assign n205 = n125 & n204;
  assign n206 = n129 & n205;
  assign n207 = n132 & n206;
  assign n208 = ~n135 & n207;
  assign n209 = n138 & n208;
  assign n210 = n142 & n209;
  assign n211 = n146 & n210;
  assign n212 = ~n149 & n211;
  assign n213 = n152 & n212;
  assign n214 = \dest_x[9]  & n213;
  assign n215 = n186 & ~n214;
  assign \outport[0]  = n187 | n215;
  assign n217 = ~\dest_y[9]  & ~\dest_y[10] ;
  assign n218 = \dest_y[11]  & ~n217;
  assign n219 = ~\dest_y[12]  & ~n218;
  assign n220 = ~\dest_y[13]  & n219;
  assign n221 = \dest_y[14]  & ~n220;
  assign n222 = \dest_y[15]  & n221;
  assign n223 = ~\dest_y[16]  & ~n222;
  assign n224 = \dest_y[17]  & ~n223;
  assign n225 = ~\dest_y[18]  & ~n224;
  assign n226 = \dest_y[19]  & ~n225;
  assign n227 = \dest_y[20]  & n226;
  assign n228 = ~\dest_y[21]  & ~n227;
  assign n229 = ~\dest_y[22]  & n228;
  assign n230 = \dest_y[23]  & ~n229;
  assign n231 = \dest_y[24]  & n230;
  assign n232 = \dest_y[25]  & n231;
  assign n233 = ~\dest_y[26]  & ~n232;
  assign n234 = \dest_y[27]  & ~n233;
  assign n235 = \dest_y[28]  & n234;
  assign n236 = \dest_y[29]  & n235;
  assign n237 = \dest_x[0]  & ~n236;
  assign n238 = ~\dest_x[0]  & ~\dest_y[0] ;
  assign n239 = n236 & ~n238;
  assign n240 = \dest_y[9]  & \dest_y[10] ;
  assign n241 = ~n217 & ~n240;
  assign n242 = ~\dest_y[11]  & n217;
  assign n243 = ~n218 & ~n242;
  assign n244 = \dest_y[12]  & n218;
  assign n245 = ~n219 & ~n244;
  assign n246 = \dest_y[13]  & ~n219;
  assign n247 = ~n220 & ~n246;
  assign n248 = ~\dest_y[14]  & n220;
  assign n249 = ~n221 & ~n248;
  assign n250 = \dest_y[15]  & ~n221;
  assign n251 = ~\dest_y[15]  & n221;
  assign n252 = ~n250 & ~n251;
  assign n253 = \dest_y[16]  & n222;
  assign n254 = ~n223 & ~n253;
  assign n255 = ~\dest_y[17]  & n223;
  assign n256 = ~n224 & ~n255;
  assign n257 = \dest_y[18]  & n224;
  assign n258 = ~n225 & ~n257;
  assign n259 = ~\dest_y[19]  & n225;
  assign n260 = ~n226 & ~n259;
  assign n261 = \dest_y[20]  & ~n226;
  assign n262 = ~\dest_y[20]  & n226;
  assign n263 = ~n261 & ~n262;
  assign n264 = \dest_y[21]  & n227;
  assign n265 = ~n228 & ~n264;
  assign n266 = \dest_y[22]  & ~n228;
  assign n267 = ~n229 & ~n266;
  assign n268 = ~\dest_y[23]  & n229;
  assign n269 = ~n230 & ~n268;
  assign n270 = \dest_y[24]  & ~n230;
  assign n271 = ~\dest_y[24]  & n230;
  assign n272 = ~n270 & ~n271;
  assign n273 = \dest_y[25]  & ~n231;
  assign n274 = ~\dest_y[25]  & n231;
  assign n275 = ~n273 & ~n274;
  assign n276 = \dest_y[26]  & n232;
  assign n277 = ~n233 & ~n276;
  assign n278 = ~\dest_y[27]  & n233;
  assign n279 = ~n234 & ~n278;
  assign n280 = \dest_y[28]  & ~n234;
  assign n281 = ~\dest_y[28]  & n234;
  assign n282 = ~n280 & ~n281;
  assign n283 = \dest_y[0]  & ~\dest_y[9] ;
  assign n284 = \dest_y[29]  & n283;
  assign n285 = ~n282 & n284;
  assign n286 = n279 & n285;
  assign n287 = ~n277 & n286;
  assign n288 = ~n275 & n287;
  assign n289 = ~n272 & n288;
  assign n290 = n269 & n289;
  assign n291 = ~n267 & n290;
  assign n292 = ~n265 & n291;
  assign n293 = ~n263 & n292;
  assign n294 = n260 & n293;
  assign n295 = ~n258 & n294;
  assign n296 = n256 & n295;
  assign n297 = ~n254 & n296;
  assign n298 = ~n252 & n297;
  assign n299 = n249 & n298;
  assign n300 = ~n247 & n299;
  assign n301 = ~n245 & n300;
  assign n302 = n243 & n301;
  assign n303 = ~n241 & n302;
  assign n304 = \dest_y[8]  & n303;
  assign n305 = \dest_y[7]  & n304;
  assign n306 = \dest_y[6]  & n305;
  assign n307 = \dest_y[5]  & n306;
  assign n308 = \dest_y[4]  & n307;
  assign n309 = \dest_y[3]  & n308;
  assign n310 = \dest_y[2]  & n309;
  assign n311 = \dest_y[1]  & n310;
  assign n312 = ~\dest_y[1]  & ~\dest_y[2] ;
  assign n313 = ~\dest_y[3]  & n312;
  assign n314 = ~\dest_y[4]  & n313;
  assign n315 = ~\dest_y[5]  & n314;
  assign n316 = ~\dest_y[6]  & n315;
  assign n317 = ~\dest_y[7]  & n316;
  assign n318 = ~\dest_y[8]  & n317;
  assign n319 = n241 & n318;
  assign n320 = ~n243 & n319;
  assign n321 = n245 & n320;
  assign n322 = n247 & n321;
  assign n323 = ~n249 & n322;
  assign n324 = n252 & n323;
  assign n325 = n254 & n324;
  assign n326 = ~n256 & n325;
  assign n327 = n258 & n326;
  assign n328 = ~n260 & n327;
  assign n329 = n263 & n328;
  assign n330 = n265 & n329;
  assign n331 = n267 & n330;
  assign n332 = ~n269 & n331;
  assign n333 = n272 & n332;
  assign n334 = n275 & n333;
  assign n335 = n277 & n334;
  assign n336 = ~n279 & n335;
  assign n337 = n282 & n336;
  assign n338 = \dest_y[9]  & n337;
  assign n339 = n236 & ~n338;
  assign n340 = ~n311 & ~n339;
  assign n341 = ~n239 & n340;
  assign n342 = ~n187 & ~n341;
  assign n343 = ~n237 & n342;
  assign \outport[1]  = ~n215 & ~n343;
  assign n345 = \dest_x[0]  & n236;
  assign n346 = \dest_y[0]  & n345;
  assign n347 = ~n339 & ~n346;
  assign \outport[2]  = ~\outport[0]  & ~n347;
  assign \outport[3]  = 1'b0;
  assign \outport[4]  = 1'b0;
  assign \outport[5]  = 1'b0;
  assign \outport[6]  = 1'b0;
  assign \outport[7]  = 1'b0;
  assign \outport[8]  = 1'b0;
  assign \outport[9]  = 1'b0;
  assign \outport[10]  = 1'b0;
  assign \outport[11]  = 1'b0;
  assign \outport[12]  = 1'b0;
  assign \outport[13]  = 1'b0;
  assign \outport[14]  = 1'b0;
  assign \outport[15]  = 1'b0;
  assign \outport[16]  = 1'b0;
  assign \outport[17]  = 1'b0;
  assign \outport[18]  = 1'b0;
  assign \outport[19]  = 1'b0;
  assign \outport[20]  = 1'b0;
  assign \outport[21]  = 1'b0;
  assign \outport[22]  = 1'b0;
  assign \outport[23]  = 1'b0;
  assign \outport[24]  = 1'b0;
  assign \outport[25]  = 1'b0;
  assign \outport[26]  = 1'b0;
  assign \outport[27]  = 1'b0;
  assign \outport[28]  = 1'b0;
  assign \outport[29]  = 1'b0;
endmodule


