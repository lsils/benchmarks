library ieee;
use ieee.std_logic_1164.all;

entity top is
port (a, b: in std_logic_vector(63 downto 0);
      quotient, remainder: out std_logic_vector(63 downto 0));
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200, w19201, w19202, w19203, w19204, w19205, w19206, w19207, w19208, w19209, w19210, w19211, w19212, w19213, w19214, w19215, w19216, w19217, w19218, w19219, w19220, w19221, w19222, w19223, w19224, w19225, w19226, w19227, w19228, w19229, w19230, w19231, w19232, w19233, w19234, w19235, w19236, w19237, w19238, w19239, w19240, w19241, w19242, w19243, w19244, w19245, w19246, w19247, w19248, w19249, w19250, w19251, w19252, w19253, w19254, w19255, w19256, w19257, w19258, w19259, w19260, w19261, w19262, w19263, w19264, w19265, w19266, w19267, w19268, w19269, w19270, w19271, w19272, w19273, w19274, w19275, w19276, w19277, w19278, w19279, w19280, w19281, w19282, w19283, w19284, w19285, w19286, w19287, w19288, w19289, w19290, w19291, w19292, w19293, w19294, w19295, w19296, w19297, w19298, w19299, w19300, w19301, w19302, w19303, w19304, w19305, w19306, w19307, w19308, w19309, w19310, w19311, w19312, w19313, w19314, w19315, w19316, w19317, w19318, w19319, w19320, w19321, w19322, w19323, w19324, w19325, w19326, w19327, w19328, w19329, w19330, w19331, w19332, w19333, w19334, w19335, w19336, w19337, w19338, w19339, w19340, w19341, w19342, w19343, w19344, w19345, w19346, w19347, w19348, w19349, w19350, w19351, w19352, w19353, w19354, w19355, w19356, w19357, w19358, w19359, w19360, w19361, w19362, w19363, w19364, w19365, w19366, w19367, w19368, w19369, w19370, w19371, w19372, w19373, w19374, w19375, w19376, w19377, w19378, w19379, w19380, w19381, w19382, w19383, w19384, w19385, w19386, w19387, w19388, w19389, w19390, w19391, w19392, w19393, w19394, w19395, w19396, w19397, w19398, w19399, w19400, w19401, w19402, w19403, w19404, w19405, w19406, w19407, w19408, w19409, w19410, w19411, w19412, w19413, w19414, w19415, w19416, w19417, w19418, w19419, w19420, w19421, w19422, w19423, w19424, w19425, w19426, w19427, w19428, w19429, w19430, w19431, w19432, w19433, w19434, w19435, w19436, w19437, w19438, w19439, w19440, w19441, w19442, w19443, w19444, w19445, w19446, w19447, w19448, w19449, w19450, w19451, w19452, w19453, w19454, w19455, w19456, w19457, w19458, w19459, w19460, w19461, w19462, w19463, w19464, w19465, w19466, w19467, w19468, w19469, w19470, w19471, w19472, w19473, w19474, w19475, w19476, w19477, w19478, w19479, w19480, w19481, w19482, w19483, w19484, w19485, w19486, w19487, w19488, w19489, w19490, w19491, w19492, w19493, w19494, w19495, w19496, w19497, w19498, w19499, w19500, w19501, w19502, w19503, w19504, w19505, w19506, w19507, w19508, w19509, w19510, w19511, w19512, w19513, w19514, w19515, w19516, w19517, w19518, w19519, w19520, w19521, w19522, w19523, w19524, w19525, w19526, w19527, w19528, w19529, w19530, w19531, w19532, w19533, w19534, w19535, w19536, w19537, w19538, w19539, w19540, w19541, w19542, w19543, w19544, w19545, w19546, w19547, w19548, w19549, w19550, w19551, w19552, w19553, w19554, w19555, w19556, w19557, w19558, w19559, w19560, w19561, w19562, w19563, w19564, w19565, w19566, w19567, w19568, w19569, w19570, w19571, w19572, w19573, w19574, w19575, w19576, w19577, w19578, w19579, w19580, w19581, w19582, w19583, w19584, w19585, w19586, w19587, w19588, w19589, w19590, w19591, w19592, w19593, w19594, w19595, w19596, w19597, w19598, w19599, w19600, w19601, w19602, w19603, w19604, w19605, w19606, w19607, w19608, w19609, w19610, w19611, w19612, w19613, w19614, w19615, w19616, w19617, w19618, w19619, w19620, w19621, w19622, w19623, w19624, w19625, w19626, w19627, w19628, w19629, w19630, w19631, w19632, w19633, w19634, w19635, w19636, w19637, w19638, w19639, w19640, w19641, w19642, w19643, w19644, w19645, w19646, w19647, w19648, w19649, w19650, w19651, w19652, w19653, w19654, w19655, w19656, w19657, w19658, w19659, w19660, w19661, w19662, w19663, w19664, w19665, w19666, w19667, w19668, w19669, w19670, w19671, w19672, w19673, w19674, w19675, w19676, w19677, w19678, w19679, w19680, w19681, w19682, w19683, w19684, w19685, w19686, w19687, w19688, w19689, w19690, w19691, w19692, w19693, w19694, w19695, w19696, w19697, w19698, w19699, w19700, w19701, w19702, w19703, w19704, w19705, w19706, w19707, w19708, w19709, w19710, w19711, w19712, w19713, w19714, w19715, w19716, w19717, w19718, w19719, w19720, w19721, w19722, w19723, w19724, w19725, w19726, w19727, w19728, w19729, w19730, w19731, w19732, w19733, w19734, w19735, w19736, w19737, w19738, w19739, w19740, w19741, w19742, w19743, w19744, w19745, w19746, w19747, w19748, w19749, w19750, w19751, w19752, w19753, w19754, w19755, w19756, w19757, w19758, w19759, w19760, w19761, w19762, w19763, w19764, w19765, w19766, w19767, w19768, w19769, w19770, w19771, w19772, w19773, w19774, w19775, w19776, w19777, w19778, w19779, w19780, w19781, w19782, w19783, w19784, w19785, w19786, w19787, w19788, w19789, w19790, w19791, w19792, w19793, w19794, w19795, w19796, w19797, w19798, w19799, w19800, w19801, w19802, w19803, w19804, w19805, w19806, w19807, w19808, w19809, w19810, w19811, w19812, w19813, w19814, w19815, w19816, w19817, w19818, w19819, w19820, w19821, w19822, w19823, w19824, w19825, w19826, w19827, w19828, w19829, w19830, w19831, w19832, w19833, w19834, w19835, w19836, w19837, w19838, w19839, w19840, w19841, w19842, w19843, w19844, w19845, w19846, w19847, w19848, w19849, w19850, w19851, w19852, w19853, w19854, w19855, w19856, w19857, w19858, w19859, w19860, w19861, w19862, w19863, w19864, w19865, w19866, w19867, w19868, w19869, w19870, w19871, w19872, w19873, w19874, w19875, w19876, w19877, w19878, w19879, w19880, w19881, w19882, w19883, w19884, w19885, w19886, w19887, w19888, w19889, w19890, w19891, w19892, w19893, w19894, w19895, w19896, w19897, w19898, w19899, w19900, w19901, w19902, w19903, w19904, w19905, w19906, w19907, w19908, w19909, w19910, w19911, w19912, w19913, w19914, w19915, w19916, w19917, w19918, w19919, w19920, w19921, w19922, w19923, w19924, w19925, w19926, w19927, w19928, w19929, w19930, w19931, w19932, w19933, w19934, w19935, w19936, w19937, w19938, w19939, w19940, w19941, w19942, w19943, w19944, w19945, w19946, w19947, w19948, w19949, w19950, w19951, w19952, w19953, w19954, w19955, w19956, w19957, w19958, w19959, w19960, w19961, w19962, w19963, w19964, w19965, w19966, w19967, w19968, w19969, w19970, w19971, w19972, w19973, w19974, w19975, w19976, w19977, w19978, w19979, w19980, w19981, w19982, w19983, w19984, w19985, w19986, w19987, w19988, w19989, w19990, w19991, w19992, w19993, w19994, w19995, w19996, w19997, w19998, w19999, w20000, w20001, w20002, w20003, w20004, w20005, w20006, w20007, w20008, w20009, w20010, w20011, w20012, w20013, w20014, w20015, w20016, w20017, w20018, w20019, w20020, w20021, w20022, w20023, w20024, w20025, w20026, w20027, w20028, w20029, w20030, w20031, w20032, w20033, w20034, w20035, w20036, w20037, w20038, w20039, w20040, w20041, w20042, w20043, w20044, w20045, w20046, w20047, w20048, w20049, w20050, w20051, w20052, w20053, w20054, w20055, w20056, w20057, w20058, w20059, w20060, w20061, w20062, w20063, w20064, w20065, w20066, w20067, w20068, w20069, w20070, w20071, w20072, w20073, w20074, w20075, w20076, w20077, w20078, w20079, w20080, w20081, w20082, w20083, w20084, w20085, w20086, w20087, w20088, w20089, w20090, w20091, w20092, w20093, w20094, w20095, w20096, w20097, w20098, w20099, w20100, w20101, w20102, w20103, w20104, w20105, w20106, w20107, w20108, w20109, w20110, w20111, w20112, w20113, w20114, w20115, w20116, w20117, w20118, w20119, w20120, w20121, w20122, w20123, w20124, w20125, w20126, w20127, w20128, w20129, w20130, w20131, w20132, w20133, w20134, w20135, w20136, w20137, w20138, w20139, w20140, w20141, w20142, w20143, w20144, w20145, w20146, w20147, w20148, w20149, w20150, w20151, w20152, w20153, w20154, w20155, w20156, w20157, w20158, w20159, w20160, w20161, w20162, w20163, w20164, w20165, w20166, w20167, w20168, w20169, w20170, w20171, w20172, w20173, w20174, w20175, w20176, w20177, w20178, w20179, w20180, w20181, w20182, w20183, w20184, w20185, w20186, w20187, w20188, w20189, w20190, w20191, w20192, w20193, w20194, w20195, w20196, w20197, w20198, w20199, w20200, w20201, w20202, w20203, w20204, w20205, w20206, w20207, w20208, w20209, w20210, w20211, w20212, w20213, w20214, w20215, w20216, w20217, w20218, w20219, w20220, w20221, w20222, w20223, w20224, w20225, w20226, w20227, w20228, w20229, w20230, w20231, w20232, w20233, w20234, w20235, w20236, w20237, w20238, w20239, w20240, w20241, w20242, w20243, w20244, w20245, w20246, w20247, w20248, w20249, w20250, w20251, w20252, w20253, w20254, w20255, w20256, w20257, w20258, w20259, w20260, w20261, w20262, w20263, w20264, w20265, w20266, w20267, w20268, w20269, w20270, w20271, w20272, w20273, w20274, w20275, w20276, w20277, w20278, w20279, w20280, w20281, w20282, w20283, w20284, w20285, w20286, w20287, w20288, w20289, w20290, w20291, w20292, w20293, w20294, w20295, w20296, w20297, w20298, w20299, w20300, w20301, w20302, w20303, w20304, w20305, w20306, w20307, w20308, w20309, w20310, w20311, w20312, w20313, w20314, w20315, w20316, w20317, w20318, w20319, w20320, w20321, w20322, w20323, w20324, w20325, w20326, w20327, w20328, w20329, w20330, w20331, w20332, w20333, w20334, w20335, w20336, w20337, w20338, w20339, w20340, w20341, w20342, w20343, w20344, w20345, w20346, w20347, w20348, w20349, w20350, w20351, w20352, w20353, w20354, w20355, w20356, w20357, w20358, w20359, w20360, w20361, w20362, w20363, w20364, w20365, w20366, w20367, w20368, w20369, w20370, w20371, w20372, w20373, w20374, w20375, w20376, w20377, w20378, w20379, w20380, w20381, w20382, w20383, w20384, w20385, w20386, w20387, w20388, w20389, w20390, w20391, w20392, w20393, w20394, w20395, w20396, w20397, w20398, w20399, w20400, w20401, w20402, w20403, w20404, w20405, w20406, w20407, w20408, w20409, w20410, w20411, w20412, w20413, w20414, w20415, w20416, w20417, w20418, w20419, w20420, w20421, w20422, w20423, w20424, w20425, w20426, w20427, w20428, w20429, w20430, w20431, w20432, w20433, w20434, w20435, w20436, w20437, w20438, w20439, w20440, w20441, w20442, w20443, w20444, w20445, w20446, w20447, w20448, w20449, w20450, w20451, w20452, w20453, w20454, w20455, w20456, w20457, w20458, w20459, w20460, w20461, w20462, w20463, w20464, w20465, w20466, w20467, w20468, w20469, w20470, w20471, w20472, w20473, w20474, w20475, w20476, w20477, w20478, w20479, w20480, w20481, w20482, w20483, w20484, w20485, w20486, w20487, w20488, w20489, w20490, w20491, w20492, w20493, w20494, w20495, w20496, w20497, w20498, w20499, w20500, w20501, w20502, w20503, w20504, w20505, w20506, w20507, w20508, w20509, w20510, w20511, w20512, w20513, w20514, w20515, w20516, w20517, w20518, w20519, w20520, w20521, w20522, w20523, w20524, w20525, w20526, w20527, w20528, w20529, w20530, w20531, w20532, w20533, w20534, w20535, w20536, w20537, w20538, w20539, w20540, w20541, w20542, w20543, w20544, w20545, w20546, w20547, w20548, w20549, w20550, w20551, w20552, w20553, w20554, w20555, w20556, w20557, w20558, w20559, w20560, w20561, w20562, w20563, w20564, w20565, w20566, w20567, w20568, w20569, w20570, w20571, w20572, w20573, w20574, w20575, w20576, w20577, w20578, w20579, w20580, w20581, w20582, w20583, w20584, w20585, w20586, w20587, w20588, w20589, w20590, w20591, w20592, w20593, w20594, w20595, w20596, w20597, w20598, w20599, w20600, w20601, w20602, w20603, w20604, w20605, w20606, w20607, w20608, w20609, w20610, w20611, w20612, w20613, w20614, w20615, w20616, w20617, w20618, w20619, w20620, w20621, w20622, w20623, w20624, w20625, w20626, w20627, w20628, w20629, w20630, w20631, w20632, w20633, w20634, w20635, w20636, w20637, w20638, w20639, w20640, w20641, w20642, w20643, w20644, w20645, w20646, w20647, w20648, w20649, w20650, w20651, w20652, w20653, w20654, w20655, w20656, w20657, w20658, w20659, w20660, w20661, w20662, w20663, w20664, w20665, w20666, w20667, w20668, w20669, w20670, w20671, w20672, w20673, w20674, w20675, w20676, w20677, w20678, w20679, w20680, w20681, w20682, w20683, w20684, w20685, w20686, w20687, w20688, w20689, w20690, w20691, w20692, w20693, w20694, w20695, w20696, w20697, w20698, w20699, w20700, w20701, w20702, w20703, w20704, w20705, w20706, w20707, w20708, w20709, w20710, w20711, w20712, w20713, w20714, w20715, w20716, w20717, w20718, w20719, w20720, w20721, w20722, w20723, w20724, w20725, w20726, w20727, w20728, w20729, w20730, w20731, w20732, w20733, w20734, w20735, w20736, w20737, w20738, w20739, w20740, w20741, w20742, w20743, w20744, w20745, w20746, w20747, w20748, w20749, w20750, w20751, w20752, w20753, w20754, w20755, w20756, w20757, w20758, w20759, w20760, w20761, w20762, w20763, w20764, w20765, w20766, w20767, w20768, w20769, w20770, w20771, w20772, w20773, w20774, w20775, w20776, w20777, w20778, w20779, w20780, w20781, w20782, w20783, w20784, w20785, w20786, w20787, w20788, w20789, w20790, w20791, w20792, w20793, w20794, w20795, w20796, w20797, w20798, w20799, w20800, w20801, w20802, w20803, w20804, w20805, w20806, w20807, w20808, w20809, w20810, w20811, w20812, w20813, w20814, w20815, w20816, w20817, w20818, w20819, w20820, w20821, w20822, w20823, w20824, w20825, w20826, w20827, w20828, w20829, w20830, w20831, w20832, w20833, w20834, w20835, w20836, w20837, w20838, w20839, w20840, w20841, w20842, w20843, w20844, w20845, w20846, w20847, w20848, w20849, w20850, w20851, w20852, w20853, w20854, w20855, w20856, w20857, w20858, w20859, w20860, w20861, w20862, w20863, w20864, w20865, w20866, w20867, w20868, w20869, w20870, w20871, w20872, w20873, w20874, w20875, w20876, w20877, w20878, w20879, w20880, w20881, w20882, w20883, w20884, w20885, w20886, w20887, w20888, w20889, w20890, w20891, w20892, w20893, w20894, w20895, w20896, w20897, w20898, w20899, w20900, w20901, w20902, w20903, w20904, w20905, w20906, w20907, w20908, w20909, w20910, w20911, w20912, w20913, w20914, w20915, w20916, w20917, w20918, w20919, w20920, w20921, w20922, w20923, w20924, w20925, w20926, w20927, w20928, w20929, w20930, w20931, w20932, w20933, w20934, w20935, w20936, w20937, w20938, w20939, w20940, w20941, w20942, w20943, w20944, w20945, w20946, w20947, w20948, w20949, w20950, w20951, w20952, w20953, w20954, w20955, w20956, w20957, w20958, w20959, w20960, w20961, w20962, w20963, w20964, w20965, w20966, w20967, w20968, w20969, w20970, w20971, w20972, w20973, w20974, w20975, w20976, w20977, w20978, w20979, w20980, w20981, w20982, w20983, w20984, w20985, w20986, w20987, w20988, w20989, w20990, w20991, w20992, w20993, w20994, w20995, w20996, w20997, w20998, w20999, w21000, w21001, w21002, w21003, w21004, w21005, w21006, w21007, w21008, w21009, w21010, w21011, w21012, w21013, w21014, w21015, w21016, w21017, w21018, w21019, w21020, w21021, w21022, w21023, w21024, w21025, w21026, w21027, w21028, w21029, w21030, w21031, w21032, w21033, w21034, w21035, w21036, w21037, w21038, w21039, w21040, w21041, w21042, w21043, w21044, w21045, w21046, w21047, w21048, w21049, w21050, w21051, w21052, w21053, w21054, w21055, w21056, w21057, w21058, w21059, w21060, w21061, w21062, w21063, w21064, w21065, w21066, w21067, w21068, w21069, w21070, w21071, w21072, w21073, w21074, w21075, w21076, w21077, w21078, w21079, w21080, w21081, w21082, w21083, w21084, w21085, w21086, w21087, w21088, w21089, w21090, w21091, w21092, w21093, w21094, w21095, w21096, w21097, w21098, w21099, w21100, w21101, w21102, w21103, w21104, w21105, w21106, w21107, w21108, w21109, w21110, w21111, w21112, w21113, w21114, w21115, w21116, w21117, w21118, w21119, w21120, w21121, w21122, w21123, w21124, w21125, w21126, w21127, w21128, w21129, w21130, w21131, w21132, w21133, w21134, w21135, w21136, w21137, w21138, w21139, w21140, w21141, w21142, w21143, w21144, w21145, w21146, w21147, w21148, w21149, w21150, w21151, w21152, w21153, w21154, w21155, w21156, w21157, w21158, w21159, w21160, w21161, w21162, w21163, w21164, w21165, w21166, w21167, w21168, w21169, w21170, w21171, w21172, w21173, w21174, w21175, w21176, w21177, w21178, w21179, w21180, w21181, w21182, w21183, w21184, w21185, w21186, w21187, w21188, w21189, w21190, w21191, w21192, w21193, w21194, w21195, w21196, w21197, w21198, w21199, w21200, w21201, w21202, w21203, w21204, w21205, w21206, w21207, w21208, w21209, w21210, w21211, w21212, w21213, w21214, w21215, w21216, w21217, w21218, w21219, w21220, w21221, w21222, w21223, w21224, w21225, w21226, w21227, w21228, w21229, w21230, w21231, w21232, w21233, w21234, w21235, w21236, w21237, w21238, w21239, w21240, w21241, w21242, w21243, w21244, w21245, w21246, w21247, w21248, w21249, w21250, w21251, w21252, w21253, w21254, w21255, w21256, w21257, w21258, w21259, w21260, w21261, w21262, w21263, w21264, w21265, w21266, w21267, w21268, w21269, w21270, w21271, w21272, w21273, w21274, w21275, w21276, w21277, w21278, w21279, w21280, w21281, w21282, w21283, w21284, w21285, w21286, w21287, w21288, w21289, w21290, w21291, w21292, w21293, w21294, w21295, w21296, w21297, w21298, w21299, w21300, w21301, w21302, w21303, w21304, w21305, w21306, w21307, w21308, w21309, w21310, w21311, w21312, w21313, w21314, w21315, w21316, w21317, w21318, w21319, w21320, w21321, w21322, w21323, w21324, w21325, w21326, w21327, w21328, w21329, w21330, w21331, w21332, w21333, w21334, w21335, w21336, w21337, w21338, w21339, w21340, w21341, w21342, w21343, w21344, w21345, w21346, w21347, w21348, w21349, w21350, w21351, w21352, w21353, w21354, w21355, w21356, w21357, w21358, w21359, w21360, w21361, w21362, w21363, w21364, w21365, w21366, w21367, w21368, w21369, w21370, w21371, w21372, w21373, w21374, w21375, w21376, w21377, w21378, w21379, w21380, w21381, w21382, w21383, w21384, w21385, w21386, w21387, w21388, w21389, w21390, w21391, w21392, w21393, w21394, w21395, w21396, w21397, w21398, w21399, w21400, w21401, w21402, w21403, w21404, w21405, w21406, w21407, w21408, w21409, w21410, w21411, w21412, w21413, w21414, w21415, w21416, w21417, w21418, w21419, w21420, w21421, w21422, w21423, w21424, w21425, w21426, w21427, w21428, w21429, w21430, w21431, w21432, w21433, w21434, w21435, w21436, w21437, w21438, w21439, w21440, w21441, w21442, w21443, w21444, w21445, w21446, w21447, w21448, w21449, w21450, w21451, w21452, w21453, w21454, w21455, w21456, w21457, w21458, w21459, w21460, w21461, w21462, w21463, w21464, w21465, w21466, w21467, w21468, w21469, w21470, w21471, w21472, w21473, w21474, w21475, w21476, w21477, w21478, w21479, w21480, w21481, w21482, w21483, w21484, w21485, w21486, w21487, w21488, w21489, w21490, w21491, w21492, w21493, w21494, w21495, w21496, w21497, w21498, w21499, w21500, w21501, w21502, w21503, w21504, w21505, w21506, w21507, w21508, w21509, w21510, w21511, w21512, w21513, w21514, w21515, w21516, w21517, w21518, w21519, w21520, w21521, w21522, w21523, w21524, w21525, w21526, w21527, w21528, w21529, w21530, w21531, w21532, w21533, w21534, w21535, w21536, w21537, w21538, w21539, w21540, w21541, w21542, w21543, w21544, w21545, w21546, w21547, w21548, w21549, w21550, w21551, w21552, w21553, w21554, w21555, w21556, w21557, w21558, w21559, w21560, w21561, w21562, w21563, w21564, w21565, w21566, w21567, w21568, w21569, w21570, w21571, w21572, w21573, w21574, w21575, w21576, w21577, w21578, w21579, w21580, w21581, w21582, w21583, w21584, w21585, w21586, w21587, w21588, w21589, w21590, w21591, w21592, w21593, w21594, w21595, w21596, w21597, w21598, w21599, w21600, w21601, w21602, w21603, w21604, w21605, w21606, w21607, w21608, w21609, w21610, w21611, w21612, w21613, w21614, w21615, w21616, w21617, w21618, w21619, w21620, w21621, w21622, w21623, w21624, w21625, w21626, w21627, w21628, w21629, w21630, w21631, w21632, w21633, w21634, w21635, w21636, w21637, w21638, w21639, w21640, w21641, w21642, w21643, w21644, w21645, w21646, w21647, w21648, w21649, w21650, w21651, w21652, w21653, w21654, w21655, w21656, w21657, w21658, w21659, w21660, w21661, w21662, w21663, w21664, w21665, w21666, w21667, w21668, w21669, w21670, w21671, w21672, w21673, w21674, w21675, w21676, w21677, w21678, w21679, w21680, w21681, w21682, w21683, w21684, w21685, w21686, w21687, w21688, w21689, w21690, w21691, w21692, w21693, w21694, w21695, w21696, w21697, w21698, w21699, w21700, w21701, w21702, w21703, w21704, w21705, w21706, w21707, w21708, w21709, w21710, w21711, w21712, w21713, w21714, w21715, w21716, w21717, w21718, w21719, w21720, w21721, w21722, w21723, w21724, w21725, w21726, w21727, w21728, w21729, w21730, w21731, w21732, w21733, w21734, w21735, w21736, w21737, w21738, w21739, w21740, w21741, w21742, w21743, w21744, w21745, w21746, w21747, w21748, w21749, w21750, w21751, w21752, w21753, w21754, w21755, w21756, w21757, w21758, w21759, w21760, w21761, w21762, w21763, w21764, w21765, w21766, w21767, w21768, w21769, w21770, w21771, w21772, w21773, w21774, w21775, w21776, w21777, w21778, w21779, w21780, w21781, w21782, w21783, w21784, w21785, w21786, w21787, w21788, w21789, w21790, w21791, w21792, w21793, w21794, w21795, w21796, w21797, w21798, w21799, w21800, w21801, w21802, w21803, w21804, w21805, w21806, w21807, w21808, w21809, w21810, w21811, w21812, w21813, w21814, w21815, w21816, w21817, w21818, w21819, w21820, w21821, w21822, w21823, w21824, w21825, w21826, w21827, w21828, w21829, w21830, w21831, w21832, w21833, w21834, w21835, w21836, w21837, w21838, w21839, w21840, w21841, w21842, w21843, w21844, w21845, w21846, w21847, w21848, w21849, w21850, w21851, w21852, w21853, w21854, w21855, w21856, w21857, w21858, w21859, w21860, w21861, w21862, w21863, w21864, w21865, w21866, w21867, w21868, w21869, w21870, w21871, w21872, w21873, w21874, w21875, w21876, w21877, w21878, w21879, w21880, w21881, w21882, w21883, w21884, w21885, w21886, w21887, w21888, w21889, w21890, w21891, w21892, w21893, w21894, w21895, w21896, w21897, w21898, w21899, w21900, w21901, w21902, w21903, w21904, w21905, w21906, w21907, w21908, w21909, w21910, w21911, w21912, w21913, w21914, w21915, w21916, w21917, w21918, w21919, w21920, w21921, w21922, w21923, w21924, w21925, w21926, w21927, w21928, w21929, w21930, w21931, w21932, w21933, w21934, w21935, w21936, w21937, w21938, w21939, w21940, w21941, w21942, w21943, w21944, w21945, w21946, w21947, w21948, w21949, w21950, w21951, w21952, w21953, w21954, w21955, w21956, w21957, w21958, w21959, w21960, w21961, w21962, w21963, w21964, w21965, w21966, w21967, w21968, w21969, w21970, w21971, w21972, w21973, w21974, w21975, w21976, w21977, w21978, w21979, w21980, w21981, w21982, w21983, w21984, w21985, w21986, w21987, w21988, w21989, w21990, w21991, w21992, w21993, w21994, w21995, w21996, w21997, w21998, w21999, w22000, w22001, w22002, w22003, w22004, w22005, w22006, w22007, w22008, w22009, w22010, w22011, w22012, w22013, w22014, w22015, w22016, w22017, w22018, w22019, w22020, w22021, w22022, w22023, w22024, w22025, w22026, w22027, w22028, w22029, w22030, w22031, w22032, w22033, w22034, w22035, w22036, w22037, w22038, w22039, w22040, w22041, w22042, w22043, w22044, w22045, w22046, w22047, w22048, w22049, w22050, w22051, w22052, w22053, w22054, w22055, w22056, w22057, w22058, w22059, w22060, w22061, w22062, w22063, w22064, w22065, w22066, w22067, w22068, w22069, w22070, w22071, w22072, w22073, w22074, w22075, w22076, w22077, w22078, w22079, w22080, w22081, w22082, w22083, w22084, w22085, w22086, w22087, w22088, w22089, w22090, w22091, w22092, w22093, w22094, w22095, w22096, w22097, w22098, w22099, w22100, w22101, w22102, w22103, w22104, w22105, w22106, w22107, w22108, w22109, w22110, w22111, w22112, w22113, w22114, w22115, w22116, w22117, w22118, w22119, w22120, w22121, w22122, w22123, w22124, w22125, w22126, w22127, w22128, w22129, w22130, w22131, w22132, w22133, w22134, w22135, w22136, w22137, w22138, w22139, w22140, w22141, w22142, w22143, w22144, w22145, w22146, w22147, w22148, w22149, w22150, w22151, w22152, w22153, w22154, w22155, w22156, w22157, w22158, w22159, w22160, w22161, w22162, w22163, w22164, w22165, w22166, w22167, w22168, w22169, w22170, w22171, w22172, w22173, w22174, w22175, w22176, w22177, w22178, w22179, w22180, w22181, w22182, w22183, w22184, w22185, w22186, w22187, w22188, w22189, w22190, w22191, w22192, w22193, w22194, w22195, w22196, w22197, w22198, w22199, w22200, w22201, w22202, w22203, w22204, w22205, w22206, w22207, w22208, w22209, w22210, w22211, w22212, w22213, w22214, w22215, w22216, w22217, w22218, w22219, w22220, w22221, w22222, w22223, w22224, w22225, w22226, w22227, w22228, w22229, w22230, w22231, w22232, w22233, w22234, w22235, w22236, w22237, w22238, w22239, w22240, w22241, w22242, w22243, w22244, w22245, w22246, w22247, w22248, w22249, w22250, w22251, w22252, w22253, w22254, w22255, w22256, w22257, w22258, w22259, w22260, w22261, w22262, w22263, w22264, w22265, w22266, w22267, w22268, w22269, w22270, w22271, w22272, w22273, w22274, w22275, w22276, w22277, w22278, w22279, w22280, w22281, w22282, w22283, w22284, w22285, w22286, w22287, w22288, w22289, w22290, w22291, w22292, w22293, w22294, w22295, w22296, w22297, w22298, w22299, w22300, w22301, w22302, w22303, w22304, w22305, w22306, w22307, w22308, w22309, w22310, w22311, w22312, w22313, w22314, w22315, w22316, w22317, w22318, w22319, w22320, w22321, w22322, w22323, w22324, w22325, w22326, w22327, w22328, w22329, w22330, w22331, w22332, w22333, w22334, w22335, w22336, w22337, w22338, w22339, w22340, w22341, w22342, w22343, w22344, w22345, w22346, w22347, w22348, w22349, w22350, w22351, w22352, w22353, w22354, w22355, w22356, w22357, w22358, w22359, w22360, w22361, w22362, w22363, w22364, w22365, w22366, w22367, w22368, w22369, w22370, w22371, w22372, w22373, w22374, w22375, w22376, w22377, w22378, w22379, w22380, w22381, w22382, w22383, w22384, w22385, w22386, w22387, w22388, w22389, w22390, w22391, w22392, w22393, w22394, w22395, w22396, w22397, w22398, w22399, w22400, w22401, w22402, w22403, w22404, w22405, w22406, w22407, w22408, w22409, w22410, w22411, w22412, w22413, w22414, w22415, w22416, w22417, w22418, w22419, w22420, w22421, w22422, w22423, w22424, w22425, w22426, w22427, w22428, w22429, w22430, w22431, w22432, w22433, w22434, w22435, w22436, w22437, w22438, w22439, w22440, w22441, w22442, w22443, w22444, w22445, w22446, w22447, w22448, w22449, w22450, w22451, w22452, w22453, w22454, w22455, w22456, w22457, w22458, w22459, w22460, w22461, w22462, w22463, w22464, w22465, w22466, w22467, w22468, w22469, w22470, w22471, w22472, w22473, w22474, w22475, w22476, w22477, w22478, w22479, w22480, w22481, w22482, w22483, w22484, w22485, w22486, w22487, w22488, w22489, w22490, w22491, w22492, w22493, w22494, w22495, w22496, w22497, w22498, w22499, w22500, w22501, w22502, w22503, w22504, w22505, w22506, w22507, w22508, w22509, w22510, w22511, w22512, w22513, w22514, w22515, w22516, w22517, w22518, w22519, w22520, w22521, w22522, w22523, w22524, w22525, w22526, w22527, w22528, w22529, w22530, w22531, w22532, w22533, w22534, w22535, w22536, w22537, w22538, w22539, w22540, w22541, w22542, w22543, w22544, w22545, w22546, w22547, w22548, w22549, w22550, w22551, w22552, w22553, w22554, w22555, w22556, w22557, w22558, w22559, w22560, w22561, w22562, w22563, w22564, w22565, w22566, w22567, w22568, w22569, w22570, w22571, w22572, w22573, w22574, w22575, w22576, w22577, w22578, w22579, w22580, w22581, w22582, w22583, w22584, w22585, w22586, w22587, w22588, w22589, w22590, w22591, w22592, w22593, w22594, w22595, w22596, w22597, w22598, w22599, w22600, w22601, w22602, w22603, w22604, w22605, w22606, w22607, w22608, w22609, w22610, w22611, w22612, w22613, w22614, w22615, w22616, w22617, w22618, w22619, w22620, w22621, w22622, w22623, w22624, w22625, w22626, w22627, w22628, w22629, w22630, w22631, w22632, w22633, w22634, w22635, w22636, w22637, w22638, w22639, w22640, w22641, w22642, w22643, w22644, w22645, w22646, w22647, w22648, w22649, w22650, w22651, w22652, w22653, w22654, w22655, w22656, w22657, w22658, w22659, w22660, w22661, w22662, w22663, w22664, w22665, w22666, w22667, w22668, w22669, w22670, w22671, w22672, w22673, w22674, w22675, w22676, w22677, w22678, w22679, w22680, w22681, w22682, w22683, w22684, w22685, w22686, w22687, w22688, w22689, w22690, w22691, w22692, w22693, w22694, w22695, w22696, w22697, w22698, w22699, w22700, w22701, w22702, w22703, w22704, w22705, w22706, w22707, w22708, w22709, w22710, w22711, w22712, w22713, w22714, w22715, w22716, w22717, w22718, w22719, w22720, w22721, w22722, w22723, w22724, w22725, w22726, w22727, w22728, w22729, w22730, w22731, w22732, w22733, w22734, w22735, w22736, w22737, w22738, w22739, w22740, w22741, w22742, w22743, w22744, w22745, w22746, w22747, w22748, w22749, w22750, w22751, w22752, w22753, w22754, w22755, w22756, w22757, w22758, w22759, w22760, w22761, w22762, w22763, w22764, w22765, w22766, w22767, w22768, w22769, w22770, w22771, w22772, w22773, w22774, w22775, w22776, w22777, w22778, w22779, w22780, w22781, w22782, w22783, w22784, w22785, w22786, w22787, w22788, w22789, w22790, w22791, w22792, w22793, w22794, w22795, w22796, w22797, w22798, w22799, w22800, w22801, w22802, w22803, w22804, w22805, w22806, w22807, w22808, w22809, w22810, w22811, w22812, w22813, w22814, w22815, w22816, w22817, w22818, w22819, w22820, w22821, w22822, w22823, w22824, w22825, w22826, w22827, w22828, w22829, w22830, w22831, w22832, w22833, w22834, w22835, w22836, w22837, w22838, w22839, w22840, w22841, w22842, w22843, w22844, w22845, w22846, w22847, w22848, w22849, w22850, w22851, w22852, w22853, w22854, w22855, w22856, w22857, w22858, w22859, w22860, w22861, w22862, w22863, w22864, w22865, w22866, w22867, w22868, w22869, w22870, w22871, w22872, w22873, w22874, w22875, w22876, w22877, w22878, w22879, w22880, w22881, w22882, w22883, w22884, w22885, w22886, w22887, w22888, w22889, w22890, w22891, w22892, w22893, w22894, w22895, w22896, w22897, w22898, w22899, w22900, w22901, w22902, w22903, w22904, w22905, w22906, w22907, w22908, w22909, w22910, w22911, w22912, w22913, w22914, w22915, w22916, w22917, w22918, w22919, w22920, w22921, w22922, w22923, w22924, w22925, w22926, w22927, w22928, w22929, w22930, w22931, w22932, w22933, w22934, w22935, w22936, w22937, w22938, w22939, w22940, w22941, w22942, w22943, w22944, w22945, w22946, w22947, w22948, w22949, w22950, w22951, w22952, w22953, w22954, w22955, w22956, w22957, w22958, w22959, w22960, w22961, w22962, w22963, w22964, w22965, w22966, w22967, w22968, w22969, w22970, w22971, w22972, w22973, w22974, w22975, w22976, w22977, w22978, w22979, w22980, w22981, w22982, w22983, w22984, w22985, w22986, w22987, w22988, w22989, w22990, w22991, w22992, w22993, w22994, w22995, w22996, w22997, w22998, w22999, w23000, w23001, w23002, w23003, w23004, w23005, w23006, w23007, w23008, w23009, w23010, w23011, w23012, w23013, w23014, w23015, w23016, w23017, w23018, w23019, w23020, w23021, w23022, w23023, w23024, w23025, w23026, w23027, w23028, w23029, w23030, w23031, w23032, w23033, w23034, w23035, w23036, w23037, w23038, w23039, w23040, w23041, w23042, w23043, w23044, w23045, w23046, w23047, w23048, w23049, w23050, w23051, w23052, w23053, w23054, w23055, w23056, w23057, w23058, w23059, w23060, w23061, w23062, w23063, w23064, w23065, w23066, w23067, w23068, w23069, w23070, w23071, w23072, w23073, w23074, w23075, w23076, w23077, w23078, w23079, w23080, w23081, w23082, w23083, w23084, w23085, w23086, w23087, w23088, w23089, w23090, w23091, w23092, w23093, w23094, w23095, w23096, w23097, w23098, w23099, w23100, w23101, w23102, w23103, w23104, w23105, w23106, w23107, w23108, w23109, w23110, w23111, w23112, w23113, w23114, w23115, w23116, w23117, w23118, w23119, w23120, w23121, w23122, w23123, w23124, w23125, w23126, w23127, w23128, w23129, w23130, w23131, w23132, w23133, w23134, w23135, w23136, w23137, w23138, w23139, w23140, w23141, w23142, w23143, w23144, w23145, w23146, w23147, w23148, w23149, w23150, w23151, w23152, w23153, w23154, w23155, w23156, w23157, w23158, w23159, w23160, w23161, w23162, w23163, w23164, w23165, w23166, w23167, w23168, w23169, w23170, w23171, w23172, w23173, w23174, w23175, w23176, w23177, w23178, w23179, w23180, w23181, w23182, w23183, w23184, w23185, w23186, w23187, w23188, w23189, w23190, w23191, w23192, w23193, w23194, w23195, w23196, w23197, w23198, w23199, w23200, w23201, w23202, w23203, w23204, w23205, w23206, w23207, w23208, w23209, w23210, w23211, w23212, w23213, w23214, w23215, w23216, w23217, w23218, w23219, w23220, w23221, w23222, w23223, w23224, w23225, w23226, w23227, w23228, w23229, w23230, w23231, w23232, w23233, w23234, w23235, w23236, w23237, w23238, w23239, w23240, w23241, w23242, w23243, w23244, w23245, w23246, w23247, w23248, w23249, w23250, w23251, w23252, w23253, w23254, w23255, w23256, w23257, w23258, w23259, w23260, w23261, w23262, w23263, w23264, w23265, w23266, w23267, w23268, w23269, w23270, w23271, w23272, w23273, w23274, w23275, w23276, w23277, w23278, w23279, w23280, w23281, w23282, w23283, w23284, w23285, w23286, w23287, w23288, w23289, w23290, w23291, w23292, w23293, w23294, w23295, w23296, w23297, w23298, w23299, w23300, w23301, w23302, w23303, w23304, w23305, w23306, w23307, w23308, w23309, w23310, w23311, w23312, w23313, w23314, w23315, w23316, w23317, w23318, w23319, w23320, w23321, w23322, w23323, w23324, w23325, w23326, w23327, w23328, w23329, w23330, w23331, w23332, w23333, w23334, w23335, w23336, w23337, w23338, w23339, w23340, w23341, w23342, w23343, w23344, w23345, w23346, w23347, w23348, w23349, w23350, w23351, w23352, w23353, w23354, w23355, w23356, w23357, w23358, w23359, w23360, w23361, w23362, w23363, w23364, w23365, w23366, w23367, w23368, w23369, w23370, w23371, w23372, w23373, w23374, w23375, w23376, w23377, w23378, w23379, w23380, w23381, w23382, w23383, w23384, w23385, w23386, w23387, w23388, w23389, w23390, w23391, w23392, w23393, w23394, w23395, w23396, w23397, w23398, w23399, w23400, w23401, w23402, w23403, w23404, w23405, w23406, w23407, w23408, w23409, w23410, w23411, w23412, w23413, w23414, w23415, w23416, w23417, w23418, w23419, w23420, w23421, w23422, w23423, w23424, w23425, w23426, w23427, w23428, w23429, w23430, w23431, w23432, w23433, w23434, w23435, w23436, w23437, w23438, w23439, w23440, w23441, w23442, w23443, w23444, w23445, w23446, w23447, w23448, w23449, w23450, w23451, w23452, w23453, w23454, w23455, w23456, w23457, w23458, w23459, w23460, w23461, w23462, w23463, w23464, w23465, w23466, w23467, w23468, w23469, w23470, w23471, w23472, w23473, w23474, w23475, w23476, w23477, w23478, w23479, w23480, w23481, w23482, w23483, w23484, w23485, w23486, w23487, w23488, w23489, w23490, w23491, w23492, w23493, w23494, w23495, w23496, w23497, w23498, w23499, w23500, w23501, w23502, w23503, w23504, w23505, w23506, w23507, w23508, w23509, w23510, w23511, w23512, w23513, w23514, w23515, w23516, w23517, w23518, w23519, w23520, w23521, w23522, w23523, w23524, w23525, w23526, w23527, w23528, w23529, w23530, w23531, w23532, w23533, w23534, w23535, w23536, w23537, w23538, w23539, w23540, w23541, w23542, w23543, w23544, w23545, w23546, w23547, w23548, w23549, w23550, w23551, w23552, w23553, w23554, w23555, w23556, w23557, w23558, w23559, w23560, w23561, w23562, w23563, w23564, w23565, w23566, w23567, w23568, w23569, w23570, w23571, w23572, w23573, w23574, w23575, w23576, w23577, w23578, w23579, w23580, w23581, w23582, w23583, w23584, w23585, w23586, w23587, w23588, w23589, w23590, w23591, w23592, w23593, w23594, w23595, w23596, w23597, w23598, w23599, w23600, w23601, w23602, w23603, w23604, w23605, w23606, w23607, w23608, w23609, w23610, w23611, w23612, w23613, w23614, w23615, w23616, w23617, w23618, w23619, w23620, w23621, w23622, w23623, w23624, w23625, w23626, w23627, w23628, w23629, w23630, w23631, w23632, w23633, w23634, w23635, w23636, w23637, w23638, w23639, w23640, w23641, w23642, w23643, w23644, w23645, w23646, w23647, w23648, w23649, w23650, w23651, w23652, w23653, w23654, w23655, w23656, w23657, w23658, w23659, w23660, w23661, w23662, w23663, w23664, w23665, w23666, w23667, w23668, w23669, w23670, w23671, w23672, w23673, w23674, w23675, w23676, w23677, w23678, w23679, w23680, w23681, w23682, w23683, w23684, w23685, w23686, w23687, w23688, w23689, w23690, w23691, w23692, w23693, w23694, w23695, w23696, w23697, w23698, w23699, w23700, w23701, w23702, w23703, w23704, w23705, w23706, w23707, w23708, w23709, w23710, w23711, w23712, w23713, w23714, w23715, w23716, w23717, w23718, w23719, w23720, w23721, w23722, w23723, w23724, w23725, w23726, w23727, w23728, w23729, w23730, w23731, w23732, w23733, w23734, w23735, w23736, w23737, w23738, w23739, w23740, w23741, w23742, w23743, w23744, w23745, w23746, w23747, w23748, w23749, w23750, w23751, w23752, w23753, w23754, w23755, w23756, w23757, w23758, w23759, w23760, w23761, w23762, w23763, w23764, w23765, w23766, w23767, w23768, w23769, w23770, w23771, w23772, w23773, w23774, w23775, w23776, w23777, w23778, w23779, w23780, w23781, w23782, w23783, w23784, w23785, w23786, w23787, w23788, w23789, w23790, w23791, w23792, w23793, w23794, w23795, w23796, w23797, w23798, w23799, w23800, w23801, w23802, w23803, w23804, w23805, w23806, w23807, w23808, w23809, w23810, w23811, w23812, w23813, w23814, w23815, w23816, w23817, w23818, w23819, w23820, w23821, w23822, w23823, w23824, w23825, w23826, w23827, w23828, w23829, w23830, w23831, w23832, w23833, w23834, w23835, w23836, w23837, w23838, w23839, w23840, w23841, w23842, w23843, w23844, w23845, w23846, w23847, w23848, w23849, w23850, w23851, w23852, w23853, w23854, w23855, w23856, w23857, w23858, w23859, w23860, w23861, w23862, w23863, w23864, w23865, w23866, w23867, w23868, w23869, w23870, w23871, w23872, w23873, w23874, w23875, w23876, w23877, w23878, w23879, w23880, w23881, w23882, w23883, w23884, w23885, w23886, w23887, w23888, w23889, w23890, w23891, w23892, w23893, w23894, w23895, w23896, w23897, w23898, w23899, w23900, w23901, w23902, w23903, w23904, w23905, w23906, w23907, w23908, w23909, w23910, w23911, w23912, w23913, w23914, w23915, w23916, w23917, w23918, w23919, w23920, w23921, w23922, w23923, w23924, w23925, w23926, w23927, w23928, w23929, w23930, w23931, w23932, w23933, w23934, w23935, w23936, w23937, w23938, w23939, w23940, w23941, w23942, w23943, w23944, w23945, w23946, w23947, w23948, w23949, w23950, w23951, w23952, w23953, w23954, w23955, w23956, w23957, w23958, w23959, w23960, w23961, w23962, w23963, w23964, w23965, w23966, w23967, w23968, w23969, w23970, w23971, w23972, w23973, w23974, w23975, w23976, w23977, w23978, w23979, w23980, w23981, w23982, w23983, w23984, w23985, w23986, w23987, w23988, w23989, w23990, w23991, w23992, w23993, w23994, w23995, w23996, w23997, w23998, w23999, w24000, w24001, w24002, w24003, w24004, w24005, w24006, w24007, w24008, w24009, w24010, w24011, w24012, w24013, w24014, w24015, w24016, w24017, w24018, w24019, w24020, w24021, w24022, w24023, w24024, w24025, w24026, w24027, w24028, w24029, w24030, w24031, w24032, w24033, w24034, w24035, w24036, w24037, w24038, w24039, w24040, w24041, w24042, w24043, w24044, w24045, w24046, w24047, w24048, w24049, w24050, w24051, w24052, w24053, w24054, w24055, w24056, w24057, w24058, w24059, w24060, w24061, w24062, w24063, w24064, w24065, w24066, w24067, w24068, w24069, w24070, w24071, w24072, w24073, w24074, w24075, w24076, w24077, w24078, w24079, w24080, w24081, w24082, w24083, w24084, w24085, w24086, w24087, w24088, w24089, w24090, w24091, w24092, w24093, w24094, w24095, w24096, w24097, w24098, w24099, w24100, w24101, w24102, w24103, w24104, w24105, w24106, w24107, w24108, w24109, w24110, w24111, w24112, w24113, w24114, w24115, w24116, w24117, w24118, w24119, w24120, w24121, w24122, w24123, w24124, w24125, w24126, w24127, w24128, w24129, w24130, w24131, w24132, w24133, w24134, w24135, w24136, w24137, w24138, w24139, w24140, w24141, w24142, w24143, w24144, w24145, w24146, w24147, w24148, w24149, w24150, w24151, w24152, w24153, w24154, w24155, w24156, w24157, w24158, w24159, w24160, w24161, w24162, w24163, w24164, w24165, w24166, w24167, w24168, w24169, w24170, w24171, w24172, w24173, w24174, w24175, w24176, w24177, w24178, w24179, w24180, w24181, w24182, w24183, w24184, w24185, w24186, w24187, w24188, w24189, w24190, w24191, w24192, w24193, w24194, w24195, w24196, w24197, w24198, w24199, w24200, w24201, w24202, w24203, w24204, w24205, w24206, w24207, w24208, w24209, w24210, w24211, w24212, w24213, w24214, w24215, w24216, w24217, w24218, w24219, w24220, w24221, w24222, w24223, w24224, w24225, w24226, w24227, w24228, w24229, w24230, w24231, w24232, w24233, w24234, w24235, w24236, w24237, w24238, w24239, w24240, w24241, w24242, w24243, w24244, w24245, w24246, w24247, w24248, w24249, w24250, w24251, w24252, w24253, w24254, w24255, w24256, w24257, w24258, w24259, w24260, w24261, w24262, w24263, w24264, w24265, w24266, w24267, w24268, w24269, w24270, w24271, w24272, w24273, w24274, w24275, w24276, w24277, w24278, w24279, w24280, w24281, w24282, w24283, w24284, w24285, w24286, w24287, w24288, w24289, w24290, w24291, w24292, w24293, w24294, w24295, w24296, w24297, w24298, w24299, w24300, w24301, w24302, w24303, w24304, w24305, w24306, w24307, w24308, w24309, w24310, w24311, w24312, w24313, w24314, w24315, w24316, w24317, w24318, w24319, w24320, w24321, w24322, w24323, w24324, w24325, w24326, w24327, w24328, w24329, w24330, w24331, w24332, w24333, w24334, w24335, w24336, w24337, w24338, w24339, w24340, w24341, w24342, w24343, w24344, w24345, w24346, w24347, w24348, w24349, w24350, w24351, w24352, w24353, w24354, w24355, w24356, w24357, w24358, w24359, w24360, w24361, w24362, w24363, w24364, w24365, w24366, w24367, w24368, w24369, w24370, w24371, w24372, w24373, w24374, w24375, w24376, w24377, w24378, w24379, w24380, w24381, w24382, w24383, w24384, w24385, w24386, w24387, w24388, w24389, w24390, w24391, w24392, w24393, w24394, w24395, w24396, w24397, w24398, w24399, w24400, w24401, w24402, w24403, w24404, w24405, w24406, w24407, w24408, w24409, w24410, w24411, w24412, w24413, w24414, w24415, w24416, w24417, w24418, w24419, w24420, w24421, w24422, w24423, w24424, w24425, w24426, w24427, w24428, w24429, w24430, w24431, w24432, w24433, w24434, w24435, w24436, w24437, w24438, w24439, w24440, w24441, w24442, w24443, w24444, w24445, w24446, w24447, w24448, w24449, w24450, w24451, w24452, w24453, w24454, w24455, w24456, w24457, w24458, w24459, w24460, w24461, w24462, w24463, w24464, w24465, w24466, w24467, w24468, w24469, w24470, w24471, w24472, w24473, w24474, w24475, w24476, w24477, w24478, w24479, w24480, w24481, w24482, w24483, w24484, w24485, w24486, w24487, w24488, w24489, w24490, w24491, w24492, w24493, w24494, w24495, w24496, w24497, w24498, w24499, w24500, w24501, w24502, w24503, w24504, w24505, w24506, w24507, w24508, w24509, w24510, w24511, w24512, w24513, w24514, w24515, w24516, w24517, w24518, w24519, w24520, w24521, w24522, w24523, w24524, w24525, w24526, w24527, w24528, w24529, w24530, w24531, w24532, w24533, w24534, w24535, w24536, w24537, w24538, w24539, w24540, w24541, w24542, w24543, w24544, w24545, w24546, w24547, w24548, w24549, w24550, w24551, w24552, w24553, w24554, w24555, w24556, w24557, w24558, w24559, w24560, w24561, w24562, w24563, w24564, w24565, w24566, w24567, w24568, w24569, w24570, w24571, w24572, w24573, w24574, w24575, w24576, w24577, w24578, w24579, w24580, w24581, w24582, w24583, w24584, w24585, w24586, w24587, w24588, w24589, w24590, w24591, w24592, w24593, w24594, w24595, w24596, w24597, w24598, w24599, w24600, w24601, w24602, w24603, w24604, w24605, w24606, w24607, w24608, w24609, w24610, w24611, w24612, w24613, w24614, w24615, w24616, w24617, w24618, w24619, w24620, w24621, w24622, w24623, w24624, w24625, w24626, w24627, w24628, w24629, w24630, w24631, w24632, w24633, w24634, w24635, w24636, w24637, w24638, w24639, w24640, w24641, w24642, w24643, w24644, w24645, w24646, w24647, w24648, w24649, w24650, w24651, w24652, w24653, w24654, w24655, w24656, w24657, w24658, w24659, w24660, w24661, w24662, w24663, w24664, w24665, w24666, w24667, w24668, w24669, w24670, w24671, w24672, w24673, w24674, w24675, w24676, w24677, w24678, w24679, w24680, w24681, w24682, w24683, w24684, w24685, w24686, w24687, w24688, w24689, w24690, w24691, w24692, w24693, w24694, w24695, w24696, w24697, w24698, w24699, w24700, w24701, w24702, w24703, w24704, w24705, w24706, w24707, w24708, w24709, w24710, w24711, w24712, w24713, w24714, w24715, w24716, w24717, w24718, w24719, w24720, w24721, w24722, w24723, w24724, w24725, w24726, w24727, w24728, w24729, w24730, w24731, w24732, w24733, w24734, w24735, w24736, w24737, w24738, w24739, w24740, w24741, w24742, w24743, w24744, w24745, w24746, w24747, w24748, w24749, w24750, w24751, w24752, w24753, w24754, w24755, w24756, w24757, w24758, w24759, w24760, w24761, w24762, w24763, w24764, w24765, w24766, w24767, w24768, w24769, w24770, w24771, w24772, w24773, w24774, w24775, w24776, w24777, w24778, w24779, w24780, w24781, w24782, w24783, w24784, w24785, w24786, w24787, w24788, w24789, w24790, w24791, w24792, w24793, w24794, w24795, w24796, w24797, w24798, w24799, w24800, w24801, w24802, w24803, w24804, w24805, w24806, w24807, w24808, w24809, w24810, w24811, w24812, w24813, w24814, w24815, w24816, w24817, w24818, w24819, w24820, w24821, w24822, w24823, w24824, w24825, w24826, w24827, w24828, w24829, w24830, w24831, w24832, w24833, w24834, w24835, w24836, w24837, w24838, w24839, w24840, w24841, w24842, w24843, w24844, w24845, w24846, w24847, w24848, w24849, w24850, w24851, w24852, w24853, w24854, w24855, w24856, w24857, w24858, w24859, w24860, w24861, w24862, w24863, w24864, w24865, w24866, w24867, w24868, w24869, w24870, w24871, w24872, w24873, w24874, w24875, w24876, w24877, w24878, w24879, w24880, w24881, w24882, w24883, w24884, w24885, w24886, w24887, w24888, w24889, w24890, w24891, w24892, w24893, w24894, w24895, w24896, w24897, w24898, w24899, w24900, w24901, w24902, w24903, w24904, w24905, w24906, w24907, w24908, w24909, w24910, w24911, w24912, w24913, w24914, w24915, w24916, w24917, w24918, w24919, w24920, w24921, w24922, w24923, w24924, w24925, w24926, w24927, w24928, w24929, w24930, w24931, w24932, w24933, w24934, w24935, w24936, w24937, w24938, w24939, w24940, w24941, w24942, w24943, w24944, w24945, w24946, w24947, w24948, w24949, w24950, w24951, w24952, w24953, w24954, w24955, w24956, w24957, w24958, w24959, w24960, w24961, w24962, w24963, w24964, w24965, w24966, w24967, w24968, w24969, w24970, w24971, w24972, w24973, w24974, w24975, w24976, w24977, w24978, w24979, w24980, w24981, w24982, w24983, w24984, w24985, w24986, w24987, w24988, w24989, w24990, w24991, w24992, w24993, w24994, w24995, w24996, w24997, w24998, w24999, w25000, w25001, w25002, w25003, w25004, w25005, w25006, w25007, w25008, w25009, w25010, w25011, w25012, w25013, w25014, w25015, w25016, w25017, w25018, w25019, w25020, w25021, w25022, w25023, w25024, w25025, w25026, w25027, w25028, w25029, w25030, w25031, w25032, w25033, w25034, w25035, w25036, w25037, w25038, w25039, w25040, w25041, w25042, w25043, w25044, w25045, w25046, w25047, w25048, w25049, w25050, w25051, w25052, w25053, w25054, w25055, w25056, w25057, w25058, w25059, w25060, w25061, w25062, w25063, w25064, w25065, w25066, w25067, w25068, w25069, w25070, w25071, w25072, w25073, w25074, w25075, w25076, w25077, w25078, w25079, w25080, w25081, w25082, w25083, w25084, w25085, w25086, w25087, w25088, w25089, w25090, w25091, w25092, w25093, w25094, w25095, w25096, w25097, w25098, w25099, w25100, w25101, w25102, w25103, w25104, w25105, w25106, w25107, w25108, w25109, w25110, w25111, w25112, w25113, w25114, w25115, w25116, w25117, w25118, w25119, w25120, w25121, w25122, w25123, w25124, w25125, w25126, w25127, w25128, w25129, w25130, w25131, w25132, w25133, w25134, w25135, w25136, w25137, w25138, w25139, w25140, w25141, w25142, w25143, w25144, w25145, w25146, w25147, w25148, w25149, w25150, w25151, w25152, w25153, w25154, w25155, w25156, w25157, w25158, w25159, w25160, w25161, w25162, w25163, w25164, w25165, w25166, w25167, w25168, w25169, w25170, w25171, w25172, w25173, w25174, w25175, w25176, w25177, w25178, w25179, w25180, w25181, w25182, w25183, w25184, w25185, w25186, w25187, w25188, w25189, w25190, w25191, w25192, w25193, w25194, w25195, w25196, w25197, w25198, w25199, w25200, w25201, w25202, w25203, w25204, w25205, w25206, w25207, w25208, w25209, w25210, w25211, w25212, w25213, w25214, w25215, w25216, w25217, w25218, w25219, w25220, w25221, w25222, w25223, w25224, w25225, w25226, w25227, w25228, w25229, w25230, w25231, w25232, w25233, w25234, w25235, w25236, w25237, w25238, w25239, w25240, w25241, w25242, w25243, w25244, w25245, w25246, w25247, w25248, w25249, w25250, w25251, w25252, w25253, w25254, w25255, w25256, w25257, w25258, w25259, w25260, w25261, w25262, w25263, w25264, w25265, w25266, w25267, w25268, w25269, w25270, w25271, w25272, w25273, w25274, w25275, w25276, w25277, w25278, w25279, w25280, w25281, w25282, w25283, w25284, w25285, w25286, w25287, w25288, w25289, w25290, w25291, w25292, w25293, w25294, w25295, w25296, w25297, w25298, w25299, w25300, w25301, w25302, w25303, w25304, w25305, w25306, w25307, w25308, w25309, w25310, w25311, w25312, w25313, w25314, w25315, w25316, w25317, w25318, w25319, w25320, w25321, w25322, w25323, w25324, w25325, w25326, w25327, w25328, w25329, w25330, w25331, w25332, w25333, w25334, w25335, w25336, w25337, w25338, w25339, w25340, w25341, w25342, w25343, w25344, w25345, w25346, w25347, w25348, w25349, w25350, w25351, w25352, w25353, w25354, w25355, w25356, w25357, w25358, w25359, w25360, w25361, w25362, w25363, w25364, w25365, w25366, w25367, w25368, w25369, w25370, w25371, w25372, w25373, w25374, w25375, w25376, w25377, w25378, w25379, w25380, w25381, w25382, w25383, w25384, w25385, w25386, w25387, w25388, w25389, w25390, w25391, w25392, w25393, w25394, w25395, w25396, w25397, w25398, w25399, w25400, w25401, w25402, w25403, w25404, w25405, w25406, w25407, w25408, w25409, w25410, w25411, w25412, w25413, w25414, w25415, w25416, w25417, w25418, w25419, w25420, w25421, w25422, w25423, w25424, w25425, w25426, w25427, w25428, w25429, w25430, w25431, w25432, w25433, w25434, w25435, w25436, w25437, w25438, w25439, w25440, w25441, w25442, w25443, w25444, w25445, w25446, w25447, w25448, w25449, w25450, w25451, w25452, w25453, w25454, w25455, w25456, w25457, w25458, w25459, w25460, w25461, w25462, w25463, w25464, w25465, w25466, w25467, w25468, w25469, w25470, w25471, w25472, w25473, w25474, w25475, w25476, w25477, w25478, w25479, w25480, w25481, w25482, w25483, w25484, w25485, w25486, w25487, w25488, w25489, w25490, w25491, w25492, w25493, w25494, w25495, w25496, w25497, w25498, w25499, w25500, w25501, w25502, w25503, w25504, w25505, w25506, w25507, w25508, w25509, w25510, w25511, w25512, w25513, w25514, w25515, w25516, w25517, w25518, w25519, w25520, w25521, w25522, w25523, w25524, w25525, w25526, w25527, w25528, w25529, w25530, w25531, w25532, w25533, w25534, w25535, w25536, w25537, w25538, w25539, w25540, w25541, w25542, w25543, w25544, w25545, w25546, w25547, w25548, w25549, w25550, w25551, w25552, w25553, w25554, w25555, w25556, w25557, w25558, w25559, w25560, w25561, w25562, w25563, w25564, w25565, w25566, w25567, w25568, w25569, w25570, w25571, w25572, w25573, w25574, w25575, w25576, w25577, w25578, w25579, w25580, w25581, w25582, w25583, w25584, w25585, w25586, w25587, w25588, w25589, w25590, w25591, w25592, w25593, w25594, w25595, w25596, w25597, w25598, w25599, w25600, w25601, w25602, w25603, w25604, w25605, w25606, w25607, w25608, w25609, w25610, w25611, w25612, w25613, w25614, w25615, w25616, w25617, w25618, w25619, w25620, w25621, w25622, w25623, w25624, w25625, w25626, w25627, w25628, w25629, w25630, w25631, w25632, w25633, w25634, w25635, w25636, w25637, w25638, w25639, w25640, w25641, w25642, w25643, w25644, w25645, w25646, w25647, w25648, w25649, w25650, w25651, w25652, w25653, w25654, w25655, w25656, w25657, w25658, w25659, w25660, w25661, w25662, w25663, w25664, w25665, w25666, w25667, w25668, w25669, w25670, w25671, w25672, w25673, w25674, w25675, w25676, w25677, w25678, w25679, w25680, w25681, w25682, w25683, w25684, w25685, w25686, w25687, w25688, w25689, w25690, w25691, w25692, w25693, w25694, w25695, w25696, w25697, w25698, w25699, w25700, w25701, w25702, w25703, w25704, w25705, w25706, w25707, w25708, w25709, w25710, w25711, w25712, w25713, w25714, w25715, w25716, w25717, w25718, w25719, w25720, w25721, w25722, w25723, w25724, w25725, w25726, w25727, w25728, w25729, w25730, w25731, w25732, w25733, w25734, w25735, w25736, w25737, w25738, w25739, w25740, w25741, w25742, w25743, w25744, w25745, w25746, w25747, w25748, w25749, w25750, w25751, w25752, w25753, w25754, w25755, w25756, w25757, w25758, w25759, w25760, w25761, w25762, w25763, w25764, w25765, w25766, w25767, w25768, w25769, w25770, w25771, w25772, w25773, w25774, w25775, w25776, w25777, w25778, w25779, w25780, w25781, w25782, w25783, w25784, w25785, w25786, w25787, w25788, w25789, w25790, w25791, w25792, w25793, w25794, w25795, w25796, w25797, w25798, w25799, w25800, w25801, w25802, w25803, w25804, w25805, w25806, w25807, w25808, w25809, w25810, w25811, w25812, w25813, w25814, w25815, w25816, w25817, w25818, w25819, w25820, w25821, w25822, w25823, w25824, w25825, w25826, w25827, w25828, w25829, w25830, w25831, w25832, w25833, w25834, w25835, w25836, w25837, w25838, w25839, w25840, w25841, w25842, w25843, w25844, w25845, w25846, w25847, w25848, w25849, w25850, w25851, w25852, w25853, w25854, w25855, w25856, w25857, w25858, w25859, w25860, w25861, w25862, w25863, w25864, w25865, w25866, w25867, w25868, w25869, w25870, w25871, w25872, w25873, w25874, w25875, w25876, w25877, w25878, w25879, w25880, w25881, w25882, w25883, w25884, w25885, w25886, w25887, w25888, w25889, w25890, w25891, w25892, w25893, w25894, w25895, w25896, w25897, w25898, w25899, w25900, w25901, w25902, w25903, w25904, w25905, w25906, w25907, w25908, w25909, w25910, w25911, w25912, w25913, w25914, w25915, w25916, w25917, w25918, w25919, w25920, w25921, w25922, w25923, w25924, w25925, w25926, w25927, w25928, w25929, w25930, w25931, w25932, w25933, w25934, w25935, w25936, w25937, w25938, w25939, w25940, w25941, w25942, w25943, w25944, w25945, w25946, w25947, w25948, w25949, w25950, w25951, w25952, w25953, w25954, w25955, w25956, w25957, w25958, w25959, w25960, w25961, w25962, w25963, w25964, w25965, w25966, w25967, w25968, w25969, w25970, w25971, w25972, w25973, w25974, w25975, w25976, w25977, w25978, w25979, w25980, w25981, w25982, w25983, w25984, w25985, w25986, w25987, w25988, w25989, w25990, w25991, w25992, w25993, w25994, w25995, w25996, w25997, w25998, w25999, w26000, w26001, w26002, w26003, w26004, w26005, w26006, w26007, w26008, w26009, w26010, w26011, w26012, w26013, w26014, w26015, w26016, w26017, w26018, w26019, w26020, w26021, w26022, w26023, w26024, w26025, w26026, w26027, w26028, w26029, w26030, w26031, w26032, w26033, w26034, w26035, w26036, w26037, w26038, w26039, w26040, w26041, w26042, w26043, w26044, w26045, w26046, w26047, w26048, w26049, w26050, w26051, w26052, w26053, w26054, w26055, w26056, w26057, w26058, w26059, w26060, w26061, w26062, w26063, w26064, w26065, w26066, w26067, w26068, w26069, w26070, w26071, w26072, w26073, w26074, w26075, w26076, w26077, w26078, w26079, w26080, w26081, w26082, w26083, w26084, w26085, w26086, w26087, w26088, w26089, w26090, w26091, w26092, w26093, w26094, w26095, w26096, w26097, w26098, w26099, w26100, w26101, w26102, w26103, w26104, w26105, w26106, w26107, w26108, w26109, w26110, w26111, w26112, w26113, w26114, w26115, w26116, w26117, w26118, w26119, w26120, w26121, w26122, w26123, w26124, w26125, w26126, w26127, w26128, w26129, w26130, w26131, w26132, w26133, w26134, w26135, w26136, w26137, w26138, w26139, w26140, w26141, w26142, w26143, w26144, w26145, w26146, w26147, w26148, w26149, w26150, w26151, w26152, w26153, w26154, w26155, w26156, w26157, w26158, w26159, w26160, w26161, w26162, w26163, w26164, w26165, w26166, w26167, w26168, w26169, w26170, w26171, w26172, w26173, w26174, w26175, w26176, w26177, w26178, w26179, w26180, w26181, w26182, w26183, w26184, w26185, w26186, w26187, w26188, w26189, w26190, w26191, w26192, w26193, w26194, w26195, w26196, w26197, w26198, w26199, w26200, w26201, w26202, w26203, w26204, w26205, w26206, w26207, w26208, w26209, w26210, w26211, w26212, w26213, w26214, w26215, w26216, w26217, w26218, w26219, w26220, w26221, w26222, w26223, w26224, w26225, w26226, w26227, w26228, w26229, w26230, w26231, w26232, w26233, w26234, w26235, w26236, w26237, w26238, w26239, w26240, w26241, w26242, w26243, w26244, w26245, w26246, w26247, w26248, w26249, w26250, w26251, w26252, w26253, w26254, w26255, w26256, w26257, w26258, w26259, w26260, w26261, w26262, w26263, w26264, w26265, w26266, w26267, w26268, w26269, w26270, w26271, w26272, w26273, w26274, w26275, w26276, w26277, w26278, w26279, w26280, w26281, w26282, w26283, w26284, w26285, w26286, w26287, w26288, w26289, w26290, w26291, w26292, w26293, w26294, w26295, w26296, w26297, w26298, w26299, w26300, w26301, w26302, w26303, w26304, w26305, w26306, w26307, w26308, w26309, w26310, w26311, w26312, w26313, w26314, w26315, w26316, w26317, w26318, w26319, w26320, w26321, w26322, w26323, w26324, w26325, w26326, w26327, w26328, w26329, w26330, w26331, w26332, w26333, w26334, w26335, w26336, w26337, w26338, w26339, w26340, w26341, w26342, w26343, w26344, w26345, w26346, w26347, w26348, w26349, w26350, w26351, w26352, w26353, w26354, w26355, w26356, w26357, w26358, w26359, w26360, w26361, w26362, w26363, w26364, w26365, w26366, w26367, w26368, w26369, w26370, w26371, w26372, w26373, w26374, w26375, w26376, w26377, w26378, w26379, w26380, w26381, w26382, w26383, w26384, w26385, w26386, w26387, w26388, w26389, w26390, w26391, w26392, w26393, w26394, w26395, w26396, w26397, w26398, w26399, w26400, w26401, w26402, w26403, w26404, w26405, w26406, w26407, w26408, w26409, w26410, w26411, w26412, w26413, w26414, w26415, w26416, w26417, w26418, w26419, w26420, w26421, w26422, w26423, w26424, w26425, w26426, w26427, w26428, w26429, w26430, w26431, w26432, w26433, w26434, w26435, w26436, w26437, w26438, w26439, w26440, w26441, w26442, w26443, w26444, w26445, w26446, w26447, w26448, w26449, w26450, w26451, w26452, w26453, w26454, w26455, w26456, w26457, w26458, w26459, w26460, w26461, w26462, w26463, w26464, w26465, w26466, w26467, w26468, w26469, w26470, w26471, w26472, w26473, w26474, w26475, w26476, w26477, w26478, w26479, w26480, w26481, w26482, w26483, w26484, w26485, w26486, w26487, w26488, w26489, w26490, w26491, w26492, w26493, w26494, w26495, w26496, w26497, w26498, w26499, w26500, w26501, w26502, w26503, w26504, w26505, w26506, w26507, w26508, w26509, w26510, w26511, w26512, w26513, w26514, w26515, w26516, w26517, w26518, w26519, w26520, w26521, w26522, w26523, w26524, w26525, w26526, w26527, w26528, w26529, w26530, w26531, w26532, w26533, w26534, w26535, w26536, w26537, w26538, w26539, w26540, w26541, w26542, w26543, w26544, w26545, w26546, w26547, w26548, w26549, w26550, w26551, w26552, w26553, w26554, w26555, w26556, w26557, w26558, w26559, w26560, w26561, w26562, w26563, w26564, w26565, w26566, w26567, w26568, w26569, w26570, w26571, w26572, w26573, w26574, w26575, w26576, w26577, w26578, w26579, w26580, w26581, w26582, w26583, w26584, w26585, w26586, w26587, w26588, w26589, w26590, w26591, w26592, w26593, w26594, w26595, w26596, w26597, w26598, w26599, w26600, w26601, w26602, w26603, w26604, w26605, w26606, w26607, w26608, w26609, w26610, w26611, w26612, w26613, w26614, w26615, w26616, w26617, w26618, w26619, w26620, w26621, w26622, w26623, w26624, w26625, w26626, w26627, w26628, w26629, w26630, w26631, w26632, w26633, w26634, w26635, w26636, w26637, w26638, w26639, w26640, w26641, w26642, w26643, w26644, w26645, w26646, w26647, w26648, w26649, w26650, w26651, w26652, w26653, w26654, w26655, w26656, w26657, w26658, w26659, w26660, w26661, w26662, w26663, w26664, w26665, w26666, w26667, w26668, w26669, w26670, w26671, w26672, w26673, w26674, w26675, w26676, w26677, w26678, w26679, w26680, w26681, w26682, w26683, w26684, w26685, w26686, w26687, w26688, w26689, w26690, w26691, w26692, w26693, w26694, w26695, w26696, w26697, w26698, w26699, w26700, w26701, w26702, w26703, w26704, w26705, w26706, w26707, w26708, w26709, w26710, w26711, w26712, w26713, w26714, w26715, w26716, w26717, w26718, w26719, w26720, w26721, w26722, w26723, w26724, w26725, w26726, w26727, w26728, w26729, w26730, w26731, w26732, w26733, w26734, w26735, w26736, w26737, w26738, w26739, w26740, w26741, w26742, w26743, w26744, w26745, w26746, w26747, w26748, w26749, w26750, w26751, w26752, w26753, w26754, w26755, w26756, w26757, w26758, w26759, w26760, w26761, w26762, w26763, w26764, w26765, w26766, w26767, w26768, w26769, w26770, w26771, w26772, w26773, w26774, w26775, w26776, w26777, w26778, w26779, w26780, w26781, w26782, w26783, w26784, w26785, w26786, w26787, w26788, w26789, w26790, w26791, w26792, w26793, w26794, w26795, w26796, w26797, w26798, w26799, w26800, w26801, w26802, w26803, w26804, w26805, w26806, w26807, w26808, w26809, w26810, w26811, w26812, w26813, w26814, w26815, w26816, w26817, w26818, w26819, w26820, w26821, w26822, w26823, w26824, w26825, w26826, w26827, w26828, w26829, w26830, w26831, w26832, w26833, w26834, w26835, w26836, w26837, w26838, w26839, w26840, w26841, w26842, w26843, w26844, w26845, w26846, w26847, w26848, w26849, w26850, w26851, w26852, w26853, w26854, w26855, w26856, w26857, w26858, w26859, w26860, w26861, w26862, w26863, w26864, w26865, w26866, w26867, w26868, w26869, w26870, w26871, w26872, w26873, w26874, w26875, w26876, w26877, w26878, w26879, w26880, w26881, w26882, w26883, w26884, w26885, w26886, w26887, w26888, w26889, w26890, w26891, w26892, w26893, w26894, w26895, w26896, w26897, w26898, w26899, w26900, w26901, w26902, w26903, w26904, w26905, w26906, w26907, w26908, w26909, w26910, w26911, w26912, w26913, w26914, w26915, w26916, w26917, w26918, w26919, w26920, w26921, w26922, w26923, w26924, w26925, w26926, w26927, w26928, w26929, w26930, w26931, w26932, w26933, w26934, w26935, w26936, w26937, w26938, w26939, w26940, w26941, w26942, w26943, w26944, w26945, w26946, w26947, w26948, w26949, w26950, w26951, w26952, w26953, w26954, w26955, w26956, w26957, w26958, w26959, w26960, w26961, w26962, w26963, w26964, w26965, w26966, w26967, w26968, w26969, w26970, w26971, w26972, w26973, w26974, w26975, w26976, w26977, w26978, w26979, w26980, w26981, w26982, w26983, w26984, w26985, w26986, w26987, w26988, w26989, w26990, w26991, w26992, w26993, w26994, w26995, w26996, w26997, w26998, w26999, w27000, w27001, w27002, w27003, w27004, w27005, w27006, w27007, w27008, w27009, w27010, w27011, w27012, w27013, w27014, w27015, w27016, w27017, w27018, w27019, w27020, w27021, w27022, w27023, w27024, w27025, w27026, w27027, w27028, w27029, w27030, w27031, w27032, w27033, w27034, w27035, w27036, w27037, w27038, w27039, w27040, w27041, w27042, w27043, w27044, w27045, w27046, w27047, w27048, w27049, w27050, w27051, w27052, w27053, w27054, w27055, w27056, w27057, w27058, w27059, w27060, w27061, w27062, w27063, w27064, w27065, w27066, w27067, w27068, w27069, w27070, w27071, w27072, w27073, w27074, w27075, w27076, w27077, w27078, w27079, w27080, w27081, w27082, w27083, w27084, w27085, w27086, w27087, w27088, w27089, w27090, w27091, w27092, w27093, w27094, w27095, w27096, w27097, w27098, w27099, w27100, w27101, w27102, w27103, w27104, w27105, w27106, w27107, w27108, w27109, w27110, w27111, w27112, w27113, w27114, w27115, w27116, w27117, w27118, w27119, w27120, w27121, w27122, w27123, w27124, w27125, w27126, w27127, w27128, w27129, w27130, w27131, w27132, w27133, w27134, w27135, w27136, w27137, w27138, w27139, w27140, w27141, w27142, w27143, w27144, w27145, w27146, w27147, w27148, w27149, w27150, w27151, w27152, w27153, w27154, w27155, w27156, w27157, w27158, w27159, w27160, w27161, w27162, w27163, w27164, w27165, w27166, w27167, w27168, w27169, w27170, w27171, w27172, w27173, w27174, w27175, w27176, w27177, w27178, w27179, w27180, w27181, w27182, w27183, w27184, w27185, w27186, w27187, w27188, w27189, w27190, w27191, w27192, w27193, w27194, w27195, w27196, w27197, w27198, w27199, w27200, w27201, w27202, w27203, w27204, w27205, w27206, w27207, w27208, w27209, w27210, w27211, w27212, w27213, w27214, w27215, w27216, w27217, w27218, w27219, w27220, w27221, w27222, w27223, w27224, w27225, w27226, w27227, w27228, w27229, w27230, w27231, w27232, w27233, w27234, w27235, w27236, w27237, w27238, w27239, w27240, w27241, w27242, w27243, w27244, w27245, w27246, w27247, w27248, w27249, w27250, w27251, w27252, w27253, w27254, w27255, w27256, w27257, w27258, w27259, w27260, w27261, w27262, w27263, w27264, w27265, w27266, w27267, w27268, w27269, w27270, w27271, w27272, w27273, w27274, w27275, w27276, w27277, w27278, w27279, w27280, w27281, w27282, w27283, w27284, w27285, w27286, w27287, w27288, w27289, w27290, w27291, w27292, w27293, w27294, w27295, w27296, w27297, w27298, w27299, w27300, w27301, w27302, w27303, w27304, w27305, w27306, w27307, w27308, w27309, w27310, w27311, w27312, w27313, w27314, w27315, w27316, w27317, w27318, w27319, w27320, w27321, w27322, w27323, w27324, w27325, w27326, w27327, w27328, w27329, w27330, w27331, w27332, w27333, w27334, w27335, w27336, w27337, w27338, w27339, w27340, w27341, w27342, w27343, w27344, w27345, w27346, w27347, w27348, w27349, w27350, w27351, w27352, w27353, w27354, w27355, w27356, w27357, w27358, w27359, w27360, w27361, w27362, w27363, w27364, w27365, w27366, w27367, w27368, w27369, w27370, w27371, w27372, w27373, w27374, w27375, w27376, w27377, w27378, w27379, w27380, w27381, w27382, w27383, w27384, w27385, w27386, w27387, w27388, w27389, w27390, w27391, w27392, w27393, w27394, w27395, w27396, w27397, w27398, w27399, w27400, w27401, w27402, w27403, w27404, w27405, w27406, w27407, w27408, w27409, w27410, w27411, w27412, w27413, w27414, w27415, w27416, w27417, w27418, w27419, w27420, w27421, w27422, w27423, w27424, w27425, w27426, w27427, w27428, w27429, w27430, w27431, w27432, w27433, w27434, w27435, w27436, w27437, w27438, w27439, w27440, w27441, w27442, w27443, w27444, w27445, w27446, w27447, w27448, w27449, w27450, w27451, w27452, w27453, w27454, w27455, w27456, w27457, w27458, w27459, w27460, w27461, w27462, w27463, w27464, w27465, w27466, w27467, w27468, w27469, w27470, w27471, w27472, w27473, w27474, w27475, w27476, w27477, w27478, w27479, w27480, w27481, w27482, w27483, w27484, w27485, w27486, w27487, w27488, w27489, w27490, w27491, w27492, w27493, w27494, w27495, w27496, w27497, w27498, w27499, w27500, w27501, w27502, w27503, w27504, w27505, w27506, w27507, w27508, w27509, w27510, w27511, w27512, w27513, w27514, w27515, w27516, w27517, w27518, w27519, w27520, w27521, w27522, w27523, w27524, w27525, w27526, w27527, w27528, w27529, w27530, w27531, w27532, w27533, w27534, w27535, w27536, w27537, w27538, w27539, w27540, w27541, w27542, w27543, w27544, w27545, w27546, w27547, w27548, w27549, w27550, w27551, w27552, w27553, w27554, w27555, w27556, w27557, w27558, w27559, w27560, w27561, w27562, w27563, w27564, w27565, w27566, w27567, w27568, w27569, w27570, w27571, w27572, w27573, w27574, w27575, w27576, w27577, w27578, w27579, w27580, w27581, w27582, w27583, w27584, w27585, w27586, w27587, w27588, w27589, w27590, w27591, w27592, w27593, w27594, w27595, w27596, w27597, w27598, w27599, w27600, w27601, w27602, w27603, w27604, w27605, w27606, w27607, w27608, w27609, w27610, w27611, w27612, w27613, w27614, w27615, w27616, w27617, w27618, w27619, w27620, w27621, w27622, w27623, w27624, w27625, w27626, w27627, w27628, w27629, w27630, w27631, w27632, w27633, w27634, w27635, w27636, w27637, w27638, w27639, w27640, w27641, w27642, w27643, w27644, w27645, w27646, w27647, w27648, w27649, w27650, w27651, w27652, w27653, w27654, w27655, w27656, w27657, w27658, w27659, w27660, w27661, w27662, w27663, w27664, w27665, w27666, w27667, w27668, w27669, w27670, w27671, w27672, w27673, w27674, w27675, w27676, w27677, w27678, w27679, w27680, w27681, w27682, w27683, w27684, w27685, w27686, w27687, w27688, w27689, w27690, w27691, w27692, w27693, w27694, w27695, w27696, w27697, w27698, w27699, w27700, w27701, w27702, w27703, w27704, w27705, w27706, w27707, w27708, w27709, w27710, w27711, w27712, w27713, w27714, w27715, w27716, w27717, w27718, w27719, w27720, w27721, w27722, w27723, w27724, w27725, w27726, w27727, w27728, w27729, w27730, w27731, w27732, w27733, w27734, w27735, w27736, w27737, w27738, w27739, w27740, w27741, w27742, w27743, w27744, w27745, w27746, w27747, w27748, w27749, w27750, w27751, w27752, w27753, w27754, w27755, w27756, w27757, w27758, w27759, w27760, w27761, w27762, w27763, w27764, w27765, w27766, w27767, w27768, w27769, w27770, w27771, w27772, w27773, w27774, w27775, w27776, w27777, w27778, w27779, w27780, w27781, w27782, w27783, w27784, w27785, w27786, w27787, w27788, w27789, w27790, w27791, w27792, w27793, w27794, w27795, w27796, w27797, w27798, w27799, w27800, w27801, w27802, w27803, w27804, w27805, w27806, w27807, w27808, w27809, w27810, w27811, w27812, w27813, w27814, w27815, w27816, w27817, w27818, w27819, w27820, w27821, w27822, w27823, w27824, w27825, w27826, w27827, w27828, w27829, w27830, w27831, w27832, w27833, w27834, w27835, w27836, w27837, w27838, w27839, w27840, w27841, w27842, w27843, w27844, w27845, w27846, w27847, w27848, w27849, w27850, w27851, w27852, w27853, w27854, w27855, w27856, w27857, w27858, w27859, w27860, w27861, w27862, w27863, w27864, w27865, w27866, w27867, w27868, w27869, w27870, w27871, w27872, w27873, w27874, w27875, w27876, w27877, w27878, w27879, w27880, w27881, w27882, w27883, w27884, w27885, w27886, w27887, w27888, w27889, w27890, w27891, w27892, w27893, w27894, w27895, w27896, w27897, w27898, w27899, w27900, w27901, w27902, w27903, w27904, w27905, w27906, w27907, w27908, w27909, w27910, w27911, w27912, w27913, w27914, w27915, w27916, w27917, w27918, w27919, w27920, w27921, w27922, w27923, w27924, w27925, w27926, w27927, w27928, w27929, w27930, w27931, w27932, w27933, w27934, w27935, w27936, w27937, w27938, w27939, w27940, w27941, w27942, w27943, w27944, w27945, w27946, w27947, w27948, w27949, w27950, w27951, w27952, w27953, w27954, w27955, w27956, w27957, w27958, w27959, w27960, w27961, w27962, w27963, w27964, w27965, w27966, w27967, w27968, w27969, w27970, w27971, w27972, w27973, w27974, w27975, w27976, w27977, w27978, w27979, w27980, w27981, w27982, w27983, w27984, w27985, w27986, w27987, w27988, w27989, w27990, w27991, w27992, w27993, w27994, w27995, w27996, w27997, w27998, w27999, w28000, w28001, w28002, w28003, w28004, w28005, w28006, w28007, w28008, w28009, w28010, w28011, w28012, w28013, w28014, w28015, w28016, w28017, w28018, w28019, w28020, w28021, w28022, w28023, w28024, w28025, w28026, w28027, w28028, w28029, w28030, w28031, w28032, w28033, w28034, w28035, w28036, w28037, w28038, w28039, w28040, w28041, w28042, w28043, w28044, w28045, w28046, w28047, w28048, w28049, w28050, w28051, w28052, w28053, w28054, w28055, w28056, w28057, w28058, w28059, w28060, w28061, w28062, w28063, w28064, w28065, w28066, w28067, w28068, w28069, w28070, w28071, w28072, w28073, w28074, w28075, w28076, w28077, w28078, w28079, w28080, w28081, w28082, w28083, w28084, w28085, w28086, w28087, w28088, w28089, w28090, w28091, w28092, w28093, w28094, w28095, w28096, w28097, w28098, w28099, w28100, w28101, w28102, w28103, w28104, w28105, w28106, w28107, w28108, w28109, w28110, w28111, w28112, w28113, w28114, w28115, w28116, w28117, w28118, w28119, w28120, w28121, w28122, w28123, w28124, w28125, w28126, w28127, w28128, w28129, w28130, w28131, w28132, w28133, w28134, w28135, w28136, w28137, w28138, w28139, w28140, w28141, w28142, w28143, w28144, w28145, w28146, w28147, w28148, w28149, w28150, w28151, w28152, w28153, w28154, w28155, w28156, w28157, w28158, w28159, w28160, w28161, w28162, w28163, w28164, w28165, w28166, w28167, w28168, w28169, w28170, w28171, w28172, w28173, w28174, w28175, w28176, w28177, w28178, w28179, w28180, w28181, w28182, w28183, w28184, w28185, w28186, w28187, w28188, w28189, w28190, w28191, w28192, w28193, w28194, w28195, w28196, w28197, w28198, w28199, w28200, w28201, w28202, w28203, w28204, w28205, w28206, w28207, w28208, w28209, w28210, w28211, w28212, w28213, w28214, w28215, w28216, w28217, w28218, w28219, w28220, w28221, w28222, w28223, w28224, w28225, w28226, w28227, w28228, w28229, w28230, w28231, w28232, w28233, w28234, w28235, w28236, w28237, w28238, w28239, w28240, w28241, w28242, w28243, w28244, w28245, w28246, w28247, w28248, w28249, w28250, w28251, w28252, w28253, w28254, w28255, w28256, w28257, w28258, w28259, w28260, w28261, w28262, w28263, w28264, w28265, w28266, w28267, w28268, w28269, w28270, w28271, w28272, w28273, w28274, w28275, w28276, w28277, w28278, w28279, w28280, w28281, w28282, w28283, w28284, w28285, w28286, w28287, w28288, w28289, w28290, w28291, w28292, w28293, w28294, w28295, w28296, w28297, w28298, w28299, w28300, w28301, w28302, w28303, w28304, w28305, w28306, w28307, w28308, w28309, w28310, w28311, w28312, w28313, w28314, w28315, w28316, w28317, w28318, w28319, w28320, w28321, w28322, w28323, w28324, w28325, w28326, w28327, w28328, w28329, w28330, w28331, w28332, w28333, w28334, w28335, w28336, w28337, w28338, w28339, w28340, w28341, w28342, w28343, w28344, w28345, w28346, w28347, w28348, w28349, w28350, w28351, w28352, w28353, w28354, w28355, w28356, w28357, w28358, w28359, w28360, w28361, w28362, w28363, w28364, w28365, w28366, w28367, w28368, w28369, w28370, w28371, w28372, w28373, w28374, w28375, w28376, w28377, w28378, w28379, w28380, w28381, w28382, w28383, w28384, w28385, w28386, w28387, w28388, w28389, w28390, w28391, w28392, w28393, w28394, w28395, w28396, w28397, w28398, w28399, w28400, w28401, w28402, w28403, w28404, w28405, w28406, w28407, w28408, w28409, w28410, w28411, w28412, w28413, w28414, w28415, w28416, w28417, w28418, w28419, w28420, w28421, w28422, w28423, w28424, w28425, w28426, w28427, w28428, w28429, w28430, w28431, w28432, w28433, w28434, w28435, w28436, w28437, w28438, w28439, w28440, w28441, w28442, w28443, w28444, w28445, w28446, w28447, w28448, w28449, w28450, w28451, w28452, w28453, w28454, w28455, w28456, w28457, w28458, w28459, w28460, w28461, w28462, w28463, w28464, w28465, w28466, w28467, w28468, w28469, w28470, w28471, w28472, w28473, w28474, w28475, w28476, w28477, w28478, w28479, w28480, w28481, w28482, w28483, w28484, w28485, w28486, w28487, w28488, w28489, w28490, w28491, w28492, w28493, w28494, w28495, w28496, w28497, w28498, w28499, w28500, w28501, w28502, w28503, w28504, w28505, w28506, w28507, w28508, w28509, w28510, w28511, w28512, w28513, w28514, w28515, w28516, w28517, w28518, w28519, w28520, w28521, w28522, w28523, w28524, w28525, w28526, w28527, w28528, w28529, w28530, w28531, w28532, w28533, w28534, w28535, w28536, w28537, w28538, w28539, w28540, w28541, w28542, w28543, w28544, w28545, w28546, w28547, w28548, w28549, w28550, w28551, w28552, w28553, w28554, w28555, w28556, w28557, w28558, w28559, w28560, w28561, w28562, w28563, w28564, w28565, w28566, w28567, w28568, w28569, w28570, w28571, w28572, w28573, w28574, w28575, w28576, w28577, w28578, w28579, w28580, w28581, w28582, w28583, w28584, w28585, w28586, w28587, w28588, w28589, w28590, w28591, w28592, w28593, w28594, w28595, w28596, w28597, w28598, w28599, w28600, w28601, w28602, w28603, w28604, w28605, w28606, w28607, w28608, w28609, w28610, w28611, w28612, w28613, w28614, w28615, w28616, w28617, w28618, w28619, w28620, w28621, w28622, w28623, w28624, w28625, w28626, w28627, w28628, w28629, w28630, w28631, w28632, w28633, w28634, w28635, w28636, w28637, w28638, w28639, w28640, w28641, w28642, w28643, w28644, w28645, w28646, w28647, w28648, w28649, w28650, w28651, w28652, w28653, w28654, w28655, w28656, w28657, w28658, w28659, w28660, w28661, w28662, w28663, w28664, w28665, w28666, w28667, w28668, w28669, w28670, w28671, w28672, w28673, w28674, w28675, w28676, w28677, w28678, w28679, w28680, w28681, w28682, w28683, w28684, w28685, w28686, w28687, w28688, w28689, w28690, w28691, w28692, w28693, w28694, w28695, w28696, w28697, w28698, w28699, w28700, w28701, w28702, w28703, w28704, w28705, w28706, w28707, w28708, w28709, w28710, w28711, w28712, w28713, w28714, w28715, w28716, w28717, w28718, w28719, w28720, w28721, w28722, w28723, w28724, w28725, w28726, w28727, w28728, w28729, w28730, w28731, w28732, w28733, w28734, w28735, w28736, w28737, w28738, w28739, w28740, w28741, w28742, w28743, w28744, w28745, w28746, w28747, w28748, w28749, w28750, w28751, w28752, w28753, w28754, w28755, w28756, w28757, w28758, w28759, w28760, w28761, w28762, w28763, w28764, w28765, w28766, w28767, w28768, w28769, w28770, w28771, w28772, w28773, w28774, w28775, w28776, w28777, w28778, w28779, w28780, w28781, w28782, w28783, w28784, w28785, w28786, w28787, w28788, w28789, w28790, w28791, w28792, w28793, w28794, w28795, w28796, w28797, w28798, w28799, w28800, w28801, w28802, w28803, w28804, w28805, w28806, w28807, w28808, w28809, w28810, w28811, w28812, w28813, w28814, w28815, w28816, w28817, w28818, w28819, w28820, w28821, w28822, w28823, w28824, w28825, w28826, w28827, w28828, w28829, w28830, w28831, w28832, w28833, w28834, w28835, w28836, w28837, w28838, w28839, w28840, w28841, w28842, w28843, w28844, w28845, w28846, w28847, w28848, w28849, w28850, w28851, w28852, w28853, w28854, w28855, w28856, w28857, w28858, w28859, w28860, w28861, w28862, w28863, w28864, w28865, w28866, w28867, w28868, w28869, w28870, w28871, w28872, w28873, w28874, w28875, w28876, w28877, w28878, w28879, w28880, w28881, w28882, w28883, w28884, w28885, w28886, w28887, w28888, w28889, w28890, w28891, w28892, w28893, w28894, w28895, w28896, w28897, w28898, w28899, w28900, w28901, w28902, w28903, w28904, w28905, w28906, w28907, w28908, w28909, w28910, w28911, w28912, w28913, w28914, w28915, w28916, w28917, w28918, w28919, w28920, w28921, w28922, w28923, w28924, w28925, w28926, w28927, w28928, w28929, w28930, w28931, w28932, w28933, w28934, w28935, w28936, w28937, w28938, w28939, w28940, w28941, w28942, w28943, w28944, w28945, w28946, w28947, w28948, w28949, w28950, w28951, w28952, w28953, w28954, w28955, w28956, w28957, w28958, w28959, w28960, w28961, w28962, w28963, w28964, w28965, w28966, w28967, w28968, w28969, w28970, w28971, w28972, w28973, w28974, w28975, w28976, w28977, w28978, w28979, w28980, w28981, w28982, w28983, w28984, w28985, w28986, w28987, w28988, w28989, w28990, w28991, w28992, w28993, w28994, w28995, w28996, w28997, w28998, w28999, w29000, w29001, w29002, w29003, w29004, w29005, w29006, w29007, w29008, w29009, w29010, w29011, w29012, w29013, w29014, w29015, w29016, w29017, w29018, w29019, w29020, w29021, w29022, w29023, w29024, w29025, w29026, w29027, w29028, w29029, w29030, w29031, w29032, w29033, w29034, w29035, w29036, w29037, w29038, w29039, w29040, w29041, w29042, w29043, w29044, w29045, w29046, w29047, w29048, w29049, w29050, w29051, w29052, w29053, w29054, w29055, w29056, w29057, w29058, w29059, w29060, w29061, w29062, w29063, w29064, w29065, w29066, w29067, w29068, w29069, w29070, w29071, w29072, w29073, w29074, w29075, w29076, w29077, w29078, w29079, w29080, w29081, w29082, w29083, w29084, w29085, w29086, w29087, w29088, w29089, w29090, w29091, w29092, w29093, w29094, w29095, w29096, w29097, w29098, w29099, w29100, w29101, w29102, w29103, w29104, w29105, w29106, w29107, w29108, w29109, w29110, w29111, w29112, w29113, w29114, w29115, w29116, w29117, w29118, w29119, w29120, w29121, w29122, w29123, w29124, w29125, w29126, w29127, w29128, w29129, w29130, w29131, w29132, w29133, w29134, w29135, w29136, w29137, w29138, w29139, w29140, w29141, w29142, w29143, w29144, w29145, w29146, w29147, w29148, w29149, w29150, w29151, w29152, w29153, w29154, w29155, w29156, w29157, w29158, w29159, w29160, w29161, w29162, w29163, w29164, w29165, w29166, w29167, w29168, w29169, w29170, w29171, w29172, w29173, w29174, w29175, w29176, w29177, w29178, w29179, w29180, w29181, w29182, w29183, w29184, w29185, w29186, w29187, w29188, w29189, w29190, w29191, w29192, w29193, w29194, w29195, w29196, w29197, w29198, w29199, w29200, w29201, w29202, w29203, w29204, w29205, w29206, w29207, w29208, w29209, w29210, w29211, w29212, w29213, w29214, w29215, w29216, w29217, w29218, w29219, w29220, w29221, w29222, w29223, w29224, w29225, w29226, w29227, w29228, w29229, w29230, w29231, w29232, w29233, w29234, w29235, w29236, w29237, w29238, w29239, w29240, w29241, w29242, w29243, w29244, w29245, w29246, w29247, w29248, w29249, w29250, w29251, w29252, w29253, w29254, w29255, w29256, w29257, w29258, w29259, w29260, w29261, w29262, w29263, w29264, w29265, w29266, w29267, w29268, w29269, w29270, w29271, w29272, w29273, w29274, w29275, w29276, w29277, w29278, w29279, w29280, w29281, w29282, w29283, w29284, w29285, w29286, w29287, w29288, w29289, w29290, w29291, w29292, w29293, w29294, w29295, w29296, w29297, w29298, w29299, w29300, w29301, w29302, w29303, w29304, w29305, w29306, w29307, w29308, w29309, w29310, w29311, w29312, w29313, w29314, w29315, w29316, w29317, w29318, w29319, w29320, w29321, w29322, w29323, w29324, w29325, w29326, w29327, w29328, w29329, w29330, w29331, w29332, w29333, w29334, w29335, w29336, w29337, w29338, w29339, w29340, w29341, w29342, w29343, w29344, w29345, w29346, w29347, w29348, w29349, w29350, w29351, w29352, w29353, w29354, w29355, w29356, w29357, w29358, w29359, w29360, w29361, w29362, w29363, w29364, w29365, w29366, w29367, w29368, w29369, w29370, w29371, w29372, w29373, w29374, w29375, w29376, w29377, w29378, w29379, w29380, w29381, w29382, w29383, w29384, w29385, w29386, w29387, w29388, w29389, w29390, w29391, w29392, w29393, w29394, w29395, w29396, w29397, w29398, w29399, w29400, w29401, w29402, w29403, w29404, w29405, w29406, w29407, w29408, w29409, w29410, w29411, w29412, w29413, w29414, w29415, w29416, w29417, w29418, w29419, w29420, w29421, w29422, w29423, w29424, w29425, w29426, w29427, w29428, w29429, w29430, w29431, w29432, w29433, w29434, w29435, w29436, w29437, w29438, w29439, w29440, w29441, w29442, w29443, w29444, w29445, w29446, w29447, w29448, w29449, w29450, w29451, w29452, w29453, w29454, w29455, w29456, w29457, w29458, w29459, w29460, w29461, w29462, w29463, w29464, w29465, w29466, w29467, w29468, w29469, w29470, w29471, w29472, w29473, w29474, w29475, w29476, w29477, w29478, w29479, w29480, w29481, w29482, w29483, w29484, w29485, w29486, w29487, w29488, w29489, w29490, w29491, w29492, w29493, w29494, w29495, w29496, w29497, w29498, w29499, w29500, w29501, w29502, w29503, w29504, w29505, w29506, w29507, w29508, w29509, w29510, w29511, w29512, w29513, w29514, w29515, w29516, w29517, w29518, w29519, w29520, w29521, w29522, w29523, w29524, w29525, w29526, w29527, w29528, w29529, w29530, w29531, w29532, w29533, w29534, w29535, w29536, w29537, w29538, w29539, w29540, w29541, w29542, w29543, w29544, w29545, w29546, w29547, w29548, w29549, w29550, w29551, w29552, w29553, w29554, w29555, w29556, w29557, w29558, w29559, w29560, w29561, w29562, w29563, w29564, w29565, w29566, w29567, w29568, w29569, w29570, w29571, w29572, w29573, w29574, w29575, w29576, w29577, w29578, w29579, w29580, w29581, w29582, w29583, w29584, w29585, w29586, w29587, w29588, w29589, w29590, w29591, w29592, w29593, w29594, w29595, w29596, w29597, w29598, w29599, w29600, w29601, w29602, w29603, w29604, w29605, w29606, w29607, w29608, w29609, w29610, w29611, w29612, w29613, w29614, w29615, w29616, w29617, w29618, w29619, w29620, w29621, w29622, w29623, w29624, w29625, w29626, w29627, w29628, w29629, w29630, w29631, w29632, w29633, w29634, w29635, w29636, w29637, w29638, w29639, w29640, w29641, w29642, w29643, w29644, w29645, w29646, w29647, w29648, w29649, w29650, w29651, w29652, w29653, w29654, w29655, w29656, w29657, w29658, w29659, w29660, w29661, w29662, w29663, w29664, w29665, w29666, w29667, w29668, w29669, w29670, w29671, w29672, w29673, w29674, w29675, w29676, w29677, w29678, w29679, w29680, w29681, w29682, w29683, w29684, w29685, w29686, w29687, w29688, w29689, w29690, w29691, w29692, w29693, w29694, w29695, w29696, w29697, w29698, w29699, w29700, w29701, w29702, w29703, w29704, w29705, w29706, w29707, w29708, w29709, w29710, w29711, w29712, w29713, w29714, w29715, w29716, w29717, w29718, w29719, w29720, w29721, w29722, w29723, w29724, w29725, w29726, w29727, w29728, w29729, w29730, w29731, w29732, w29733, w29734, w29735, w29736, w29737, w29738, w29739, w29740, w29741, w29742, w29743, w29744, w29745, w29746, w29747, w29748, w29749, w29750, w29751, w29752, w29753, w29754, w29755, w29756, w29757, w29758, w29759, w29760, w29761, w29762, w29763, w29764, w29765, w29766, w29767, w29768, w29769, w29770, w29771, w29772, w29773, w29774, w29775, w29776, w29777, w29778, w29779, w29780, w29781, w29782, w29783, w29784, w29785, w29786, w29787, w29788, w29789, w29790, w29791, w29792, w29793, w29794, w29795, w29796, w29797, w29798, w29799, w29800, w29801, w29802, w29803, w29804, w29805, w29806, w29807, w29808, w29809, w29810, w29811, w29812, w29813, w29814, w29815, w29816, w29817, w29818, w29819, w29820, w29821, w29822, w29823, w29824, w29825, w29826, w29827, w29828, w29829, w29830, w29831, w29832, w29833, w29834, w29835, w29836, w29837, w29838, w29839, w29840, w29841, w29842, w29843, w29844, w29845, w29846, w29847, w29848, w29849, w29850, w29851, w29852, w29853, w29854, w29855, w29856, w29857, w29858, w29859, w29860, w29861, w29862, w29863, w29864, w29865, w29866, w29867, w29868, w29869, w29870, w29871, w29872, w29873, w29874, w29875, w29876, w29877, w29878, w29879, w29880, w29881, w29882, w29883, w29884, w29885, w29886, w29887, w29888, w29889, w29890, w29891, w29892, w29893, w29894, w29895, w29896, w29897, w29898, w29899, w29900, w29901, w29902, w29903, w29904, w29905, w29906, w29907, w29908, w29909, w29910, w29911, w29912, w29913, w29914, w29915, w29916, w29917, w29918, w29919, w29920, w29921, w29922, w29923, w29924, w29925, w29926, w29927, w29928, w29929, w29930, w29931, w29932, w29933, w29934, w29935, w29936, w29937, w29938, w29939, w29940, w29941, w29942, w29943, w29944, w29945, w29946, w29947, w29948, w29949, w29950, w29951, w29952, w29953, w29954, w29955, w29956, w29957, w29958, w29959, w29960, w29961, w29962, w29963, w29964, w29965, w29966, w29967, w29968, w29969, w29970, w29971, w29972, w29973, w29974, w29975, w29976, w29977, w29978, w29979, w29980, w29981, w29982, w29983, w29984, w29985, w29986, w29987, w29988, w29989, w29990, w29991, w29992, w29993, w29994, w29995, w29996, w29997, w29998, w29999, w30000, w30001, w30002, w30003, w30004, w30005, w30006, w30007, w30008, w30009, w30010, w30011, w30012, w30013, w30014, w30015, w30016, w30017, w30018, w30019, w30020, w30021, w30022, w30023, w30024, w30025, w30026, w30027, w30028, w30029, w30030, w30031, w30032, w30033, w30034, w30035, w30036, w30037, w30038, w30039, w30040, w30041, w30042, w30043, w30044, w30045, w30046, w30047, w30048, w30049, w30050, w30051, w30052, w30053, w30054, w30055, w30056, w30057, w30058, w30059, w30060, w30061, w30062, w30063, w30064, w30065, w30066, w30067, w30068, w30069, w30070, w30071, w30072, w30073, w30074, w30075, w30076, w30077, w30078, w30079, w30080, w30081, w30082, w30083, w30084, w30085, w30086, w30087, w30088, w30089, w30090, w30091, w30092, w30093, w30094, w30095, w30096, w30097, w30098, w30099, w30100, w30101, w30102, w30103, w30104, w30105, w30106, w30107, w30108, w30109, w30110, w30111, w30112, w30113, w30114, w30115, w30116, w30117, w30118, w30119, w30120, w30121, w30122, w30123, w30124, w30125, w30126, w30127, w30128, w30129, w30130, w30131, w30132, w30133, w30134, w30135, w30136, w30137, w30138, w30139, w30140, w30141, w30142, w30143, w30144, w30145, w30146, w30147, w30148, w30149, w30150, w30151, w30152, w30153, w30154, w30155, w30156, w30157, w30158, w30159, w30160, w30161, w30162, w30163, w30164, w30165, w30166, w30167, w30168, w30169, w30170, w30171, w30172, w30173, w30174, w30175, w30176, w30177, w30178, w30179, w30180, w30181, w30182, w30183, w30184, w30185, w30186, w30187, w30188, w30189, w30190, w30191, w30192, w30193, w30194, w30195, w30196, w30197, w30198, w30199, w30200, w30201, w30202, w30203, w30204, w30205, w30206, w30207, w30208, w30209, w30210, w30211, w30212, w30213, w30214, w30215, w30216, w30217, w30218, w30219, w30220, w30221, w30222, w30223, w30224, w30225, w30226, w30227, w30228, w30229, w30230, w30231, w30232, w30233, w30234, w30235, w30236, w30237, w30238, w30239, w30240, w30241, w30242, w30243, w30244, w30245, w30246, w30247, w30248, w30249, w30250, w30251, w30252, w30253, w30254, w30255, w30256, w30257, w30258, w30259, w30260, w30261, w30262, w30263, w30264, w30265, w30266, w30267, w30268, w30269, w30270, w30271, w30272, w30273, w30274, w30275, w30276, w30277, w30278, w30279, w30280, w30281, w30282, w30283, w30284, w30285, w30286, w30287, w30288, w30289, w30290, w30291, w30292, w30293, w30294, w30295, w30296, w30297, w30298, w30299, w30300, w30301, w30302, w30303, w30304, w30305, w30306, w30307, w30308, w30309, w30310, w30311, w30312, w30313, w30314, w30315, w30316, w30317, w30318, w30319, w30320, w30321, w30322, w30323, w30324, w30325, w30326, w30327, w30328, w30329, w30330, w30331, w30332, w30333, w30334, w30335, w30336, w30337, w30338, w30339, w30340, w30341, w30342, w30343, w30344, w30345, w30346, w30347, w30348, w30349, w30350, w30351, w30352, w30353, w30354, w30355, w30356, w30357, w30358, w30359, w30360, w30361, w30362, w30363, w30364, w30365, w30366, w30367, w30368, w30369, w30370, w30371, w30372, w30373, w30374, w30375, w30376, w30377, w30378, w30379, w30380, w30381, w30382, w30383, w30384, w30385, w30386, w30387, w30388, w30389, w30390, w30391, w30392, w30393, w30394, w30395, w30396, w30397, w30398, w30399, w30400, w30401, w30402, w30403, w30404, w30405, w30406, w30407, w30408, w30409, w30410, w30411, w30412, w30413, w30414, w30415, w30416, w30417, w30418, w30419, w30420, w30421, w30422, w30423, w30424, w30425, w30426, w30427, w30428, w30429, w30430, w30431, w30432, w30433, w30434, w30435, w30436, w30437, w30438, w30439, w30440, w30441, w30442, w30443, w30444, w30445, w30446, w30447, w30448, w30449, w30450, w30451, w30452, w30453, w30454, w30455, w30456, w30457, w30458, w30459, w30460, w30461, w30462, w30463, w30464, w30465, w30466, w30467, w30468, w30469, w30470, w30471, w30472, w30473, w30474, w30475, w30476, w30477, w30478, w30479, w30480, w30481, w30482, w30483, w30484, w30485, w30486, w30487, w30488, w30489, w30490, w30491, w30492, w30493, w30494, w30495, w30496, w30497, w30498, w30499, w30500, w30501, w30502, w30503, w30504, w30505, w30506, w30507, w30508, w30509, w30510, w30511, w30512, w30513, w30514, w30515, w30516, w30517, w30518, w30519, w30520, w30521, w30522, w30523, w30524, w30525, w30526, w30527, w30528, w30529, w30530, w30531, w30532, w30533, w30534, w30535, w30536, w30537, w30538, w30539, w30540, w30541, w30542, w30543, w30544, w30545, w30546, w30547, w30548, w30549, w30550, w30551, w30552, w30553, w30554, w30555, w30556, w30557, w30558, w30559, w30560, w30561, w30562, w30563, w30564, w30565, w30566, w30567, w30568, w30569, w30570, w30571, w30572, w30573, w30574, w30575, w30576, w30577, w30578, w30579, w30580, w30581, w30582, w30583, w30584, w30585, w30586, w30587, w30588, w30589, w30590, w30591, w30592, w30593, w30594, w30595, w30596, w30597, w30598, w30599, w30600, w30601, w30602, w30603, w30604, w30605, w30606, w30607, w30608, w30609, w30610, w30611, w30612, w30613, w30614, w30615, w30616, w30617, w30618, w30619, w30620, w30621, w30622, w30623, w30624, w30625, w30626, w30627, w30628, w30629, w30630, w30631, w30632, w30633, w30634, w30635, w30636, w30637, w30638, w30639, w30640, w30641, w30642, w30643, w30644, w30645, w30646, w30647, w30648, w30649, w30650, w30651, w30652, w30653, w30654, w30655, w30656, w30657, w30658, w30659, w30660, w30661, w30662, w30663, w30664, w30665, w30666, w30667, w30668, w30669, w30670, w30671, w30672, w30673, w30674, w30675, w30676, w30677, w30678, w30679, w30680, w30681, w30682, w30683, w30684, w30685, w30686, w30687, w30688, w30689, w30690, w30691, w30692, w30693, w30694, w30695, w30696, w30697, w30698, w30699, w30700, w30701, w30702, w30703, w30704, w30705, w30706, w30707, w30708, w30709, w30710, w30711, w30712, w30713, w30714, w30715, w30716, w30717, w30718, w30719, w30720, w30721, w30722, w30723, w30724, w30725, w30726, w30727, w30728, w30729, w30730, w30731, w30732, w30733, w30734, w30735, w30736, w30737, w30738, w30739, w30740, w30741, w30742, w30743, w30744, w30745, w30746, w30747, w30748, w30749, w30750, w30751, w30752, w30753, w30754, w30755, w30756, w30757, w30758, w30759, w30760, w30761, w30762, w30763, w30764, w30765, w30766, w30767, w30768, w30769, w30770, w30771, w30772, w30773, w30774, w30775, w30776, w30777, w30778, w30779, w30780, w30781, w30782, w30783, w30784, w30785, w30786, w30787, w30788, w30789, w30790, w30791, w30792, w30793, w30794, w30795, w30796, w30797, w30798, w30799, w30800, w30801, w30802, w30803, w30804, w30805, w30806, w30807, w30808, w30809, w30810, w30811, w30812, w30813, w30814, w30815, w30816, w30817, w30818, w30819, w30820, w30821, w30822, w30823, w30824, w30825, w30826, w30827, w30828, w30829, w30830, w30831, w30832, w30833, w30834, w30835, w30836, w30837, w30838, w30839, w30840, w30841, w30842, w30843, w30844, w30845, w30846, w30847, w30848, w30849, w30850, w30851, w30852, w30853, w30854, w30855, w30856, w30857, w30858, w30859, w30860, w30861, w30862, w30863, w30864, w30865, w30866, w30867, w30868, w30869, w30870, w30871, w30872, w30873, w30874, w30875, w30876, w30877, w30878, w30879, w30880, w30881, w30882, w30883, w30884, w30885, w30886, w30887, w30888, w30889, w30890, w30891, w30892, w30893, w30894, w30895, w30896, w30897, w30898, w30899, w30900, w30901, w30902, w30903, w30904, w30905, w30906, w30907, w30908, w30909, w30910, w30911, w30912, w30913, w30914, w30915, w30916, w30917, w30918, w30919, w30920, w30921, w30922, w30923, w30924, w30925, w30926, w30927, w30928, w30929, w30930, w30931, w30932, w30933, w30934, w30935, w30936, w30937, w30938, w30939, w30940, w30941, w30942, w30943, w30944, w30945, w30946, w30947, w30948, w30949, w30950, w30951, w30952, w30953, w30954, w30955, w30956, w30957, w30958, w30959, w30960, w30961, w30962, w30963, w30964, w30965, w30966, w30967, w30968, w30969, w30970, w30971, w30972, w30973, w30974, w30975, w30976, w30977, w30978, w30979, w30980, w30981, w30982, w30983, w30984, w30985, w30986, w30987, w30988, w30989, w30990, w30991, w30992, w30993, w30994, w30995, w30996, w30997, w30998, w30999, w31000, w31001, w31002, w31003, w31004, w31005, w31006, w31007, w31008, w31009, w31010, w31011, w31012, w31013, w31014, w31015, w31016, w31017, w31018, w31019, w31020, w31021, w31022, w31023, w31024, w31025, w31026, w31027, w31028, w31029, w31030, w31031, w31032, w31033, w31034, w31035, w31036, w31037, w31038, w31039, w31040, w31041, w31042, w31043, w31044, w31045, w31046, w31047, w31048, w31049, w31050, w31051, w31052, w31053, w31054, w31055, w31056, w31057, w31058, w31059, w31060, w31061, w31062, w31063, w31064, w31065, w31066, w31067, w31068, w31069, w31070, w31071, w31072, w31073, w31074, w31075, w31076, w31077, w31078, w31079, w31080, w31081, w31082, w31083, w31084, w31085, w31086, w31087, w31088, w31089, w31090, w31091, w31092, w31093, w31094, w31095, w31096, w31097, w31098, w31099, w31100, w31101, w31102, w31103, w31104, w31105, w31106, w31107, w31108, w31109, w31110, w31111, w31112, w31113, w31114, w31115, w31116, w31117, w31118, w31119, w31120, w31121, w31122, w31123, w31124, w31125, w31126, w31127, w31128, w31129, w31130, w31131, w31132, w31133, w31134, w31135, w31136, w31137, w31138, w31139, w31140, w31141, w31142, w31143, w31144, w31145, w31146, w31147, w31148, w31149, w31150, w31151, w31152, w31153, w31154, w31155, w31156, w31157, w31158, w31159, w31160, w31161, w31162, w31163, w31164, w31165, w31166, w31167, w31168, w31169, w31170, w31171, w31172, w31173, w31174, w31175, w31176, w31177, w31178, w31179, w31180, w31181, w31182, w31183, w31184, w31185, w31186, w31187, w31188, w31189, w31190, w31191, w31192, w31193, w31194, w31195, w31196, w31197, w31198, w31199, w31200, w31201, w31202, w31203, w31204, w31205, w31206, w31207, w31208, w31209, w31210, w31211, w31212, w31213, w31214, w31215, w31216, w31217, w31218, w31219, w31220, w31221, w31222, w31223, w31224, w31225, w31226, w31227, w31228, w31229, w31230, w31231, w31232, w31233, w31234, w31235, w31236, w31237, w31238, w31239, w31240, w31241, w31242, w31243, w31244, w31245, w31246, w31247, w31248, w31249, w31250, w31251, w31252, w31253, w31254, w31255, w31256, w31257, w31258, w31259, w31260, w31261, w31262, w31263, w31264, w31265, w31266, w31267, w31268, w31269, w31270, w31271, w31272, w31273, w31274, w31275, w31276, w31277, w31278, w31279, w31280, w31281, w31282, w31283, w31284, w31285, w31286, w31287, w31288, w31289, w31290, w31291, w31292, w31293, w31294, w31295, w31296, w31297, w31298, w31299, w31300, w31301, w31302, w31303, w31304, w31305, w31306, w31307, w31308, w31309, w31310, w31311, w31312, w31313, w31314, w31315, w31316, w31317, w31318, w31319, w31320, w31321, w31322, w31323, w31324, w31325, w31326, w31327, w31328, w31329, w31330, w31331, w31332, w31333, w31334, w31335, w31336, w31337, w31338, w31339, w31340, w31341, w31342, w31343, w31344, w31345, w31346, w31347, w31348, w31349, w31350, w31351, w31352, w31353, w31354, w31355, w31356, w31357, w31358, w31359, w31360, w31361, w31362, w31363, w31364, w31365, w31366, w31367, w31368, w31369, w31370, w31371, w31372, w31373, w31374, w31375, w31376, w31377, w31378, w31379, w31380, w31381, w31382, w31383, w31384, w31385, w31386, w31387, w31388, w31389, w31390, w31391, w31392, w31393, w31394, w31395, w31396, w31397, w31398, w31399, w31400, w31401, w31402, w31403, w31404, w31405, w31406, w31407, w31408, w31409, w31410, w31411, w31412, w31413, w31414, w31415, w31416, w31417, w31418, w31419, w31420, w31421, w31422, w31423, w31424, w31425, w31426, w31427, w31428, w31429, w31430, w31431, w31432, w31433, w31434, w31435, w31436, w31437, w31438, w31439, w31440, w31441, w31442, w31443, w31444, w31445, w31446, w31447, w31448, w31449, w31450, w31451, w31452, w31453, w31454, w31455, w31456, w31457, w31458, w31459, w31460, w31461, w31462, w31463, w31464, w31465, w31466, w31467, w31468, w31469, w31470, w31471, w31472, w31473, w31474, w31475, w31476, w31477, w31478, w31479, w31480, w31481, w31482, w31483, w31484, w31485, w31486, w31487, w31488, w31489, w31490, w31491, w31492, w31493, w31494, w31495, w31496, w31497, w31498, w31499, w31500, w31501, w31502, w31503, w31504, w31505, w31506, w31507, w31508, w31509, w31510, w31511, w31512, w31513, w31514, w31515, w31516, w31517, w31518, w31519, w31520, w31521, w31522, w31523, w31524, w31525, w31526, w31527, w31528, w31529, w31530, w31531, w31532, w31533, w31534, w31535, w31536, w31537, w31538, w31539, w31540, w31541, w31542, w31543, w31544, w31545, w31546, w31547, w31548, w31549, w31550, w31551, w31552, w31553, w31554, w31555, w31556, w31557, w31558, w31559, w31560, w31561, w31562, w31563, w31564, w31565, w31566, w31567, w31568, w31569, w31570, w31571, w31572, w31573, w31574, w31575, w31576, w31577, w31578, w31579, w31580, w31581, w31582, w31583, w31584, w31585, w31586, w31587, w31588, w31589, w31590, w31591, w31592, w31593, w31594, w31595, w31596, w31597, w31598, w31599, w31600, w31601, w31602, w31603, w31604, w31605, w31606, w31607, w31608, w31609, w31610, w31611, w31612, w31613, w31614, w31615, w31616, w31617, w31618, w31619, w31620, w31621, w31622, w31623, w31624, w31625, w31626, w31627, w31628, w31629, w31630, w31631, w31632, w31633, w31634, w31635, w31636, w31637, w31638, w31639, w31640, w31641, w31642, w31643, w31644, w31645, w31646, w31647, w31648, w31649, w31650, w31651, w31652, w31653, w31654, w31655, w31656, w31657, w31658, w31659, w31660, w31661, w31662, w31663, w31664, w31665, w31666, w31667, w31668, w31669, w31670, w31671, w31672, w31673, w31674, w31675, w31676, w31677, w31678, w31679, w31680, w31681, w31682, w31683, w31684, w31685, w31686, w31687, w31688, w31689, w31690, w31691, w31692, w31693, w31694, w31695, w31696, w31697, w31698, w31699, w31700, w31701, w31702, w31703, w31704, w31705, w31706, w31707, w31708, w31709, w31710, w31711, w31712, w31713, w31714, w31715, w31716, w31717, w31718, w31719, w31720, w31721, w31722, w31723, w31724, w31725, w31726, w31727, w31728, w31729, w31730, w31731, w31732, w31733, w31734, w31735, w31736, w31737, w31738, w31739, w31740, w31741, w31742, w31743, w31744, w31745, w31746, w31747, w31748, w31749, w31750, w31751, w31752, w31753, w31754, w31755, w31756, w31757, w31758, w31759, w31760, w31761, w31762, w31763, w31764, w31765, w31766, w31767, w31768, w31769, w31770, w31771, w31772, w31773, w31774, w31775, w31776, w31777, w31778, w31779, w31780, w31781, w31782, w31783, w31784, w31785, w31786, w31787, w31788, w31789, w31790, w31791, w31792, w31793, w31794, w31795, w31796, w31797, w31798, w31799, w31800, w31801, w31802, w31803, w31804, w31805, w31806, w31807, w31808, w31809, w31810, w31811, w31812, w31813, w31814, w31815, w31816, w31817, w31818, w31819, w31820, w31821, w31822, w31823, w31824, w31825, w31826, w31827, w31828, w31829, w31830, w31831, w31832, w31833, w31834, w31835, w31836, w31837, w31838, w31839, w31840, w31841, w31842, w31843, w31844, w31845, w31846, w31847, w31848, w31849, w31850, w31851, w31852, w31853, w31854, w31855, w31856, w31857, w31858, w31859, w31860, w31861, w31862, w31863, w31864, w31865, w31866, w31867, w31868, w31869, w31870, w31871, w31872, w31873, w31874, w31875, w31876, w31877, w31878, w31879, w31880, w31881, w31882, w31883, w31884, w31885, w31886, w31887, w31888, w31889, w31890, w31891, w31892, w31893, w31894, w31895, w31896, w31897, w31898, w31899, w31900, w31901, w31902, w31903, w31904, w31905, w31906, w31907, w31908, w31909, w31910, w31911, w31912, w31913, w31914, w31915, w31916, w31917, w31918, w31919, w31920, w31921, w31922, w31923, w31924, w31925, w31926, w31927, w31928, w31929, w31930, w31931, w31932, w31933, w31934, w31935, w31936, w31937, w31938, w31939, w31940, w31941, w31942, w31943, w31944, w31945, w31946, w31947, w31948, w31949, w31950, w31951, w31952, w31953, w31954, w31955, w31956, w31957, w31958, w31959, w31960, w31961, w31962, w31963, w31964, w31965, w31966, w31967, w31968, w31969, w31970, w31971, w31972, w31973, w31974, w31975, w31976, w31977, w31978, w31979, w31980, w31981, w31982, w31983, w31984, w31985, w31986, w31987, w31988, w31989, w31990, w31991, w31992, w31993, w31994, w31995, w31996, w31997, w31998, w31999, w32000, w32001, w32002, w32003, w32004, w32005, w32006, w32007, w32008, w32009, w32010, w32011, w32012, w32013, w32014, w32015, w32016, w32017, w32018, w32019, w32020, w32021, w32022, w32023, w32024, w32025, w32026, w32027, w32028, w32029, w32030, w32031, w32032, w32033, w32034, w32035, w32036, w32037, w32038, w32039, w32040, w32041, w32042, w32043, w32044, w32045, w32046, w32047, w32048, w32049, w32050, w32051, w32052, w32053, w32054, w32055, w32056, w32057, w32058, w32059, w32060, w32061, w32062, w32063, w32064, w32065, w32066, w32067, w32068, w32069, w32070, w32071, w32072, w32073, w32074, w32075, w32076, w32077, w32078, w32079, w32080, w32081, w32082, w32083, w32084, w32085, w32086, w32087, w32088, w32089, w32090, w32091, w32092, w32093, w32094, w32095, w32096, w32097, w32098, w32099, w32100, w32101, w32102, w32103, w32104, w32105, w32106, w32107, w32108, w32109, w32110, w32111, w32112, w32113, w32114, w32115, w32116, w32117, w32118, w32119, w32120, w32121, w32122, w32123, w32124, w32125, w32126, w32127, w32128, w32129, w32130, w32131, w32132, w32133, w32134, w32135, w32136, w32137, w32138, w32139, w32140, w32141, w32142, w32143, w32144, w32145, w32146, w32147, w32148, w32149, w32150, w32151, w32152, w32153, w32154, w32155, w32156, w32157, w32158, w32159, w32160, w32161, w32162, w32163, w32164, w32165, w32166, w32167, w32168, w32169, w32170, w32171, w32172, w32173, w32174, w32175, w32176, w32177, w32178, w32179, w32180, w32181, w32182, w32183, w32184, w32185, w32186, w32187, w32188, w32189, w32190, w32191, w32192, w32193, w32194, w32195, w32196, w32197, w32198, w32199, w32200, w32201, w32202, w32203, w32204, w32205, w32206, w32207, w32208, w32209, w32210, w32211, w32212, w32213, w32214, w32215, w32216, w32217, w32218, w32219, w32220, w32221, w32222, w32223, w32224, w32225, w32226, w32227, w32228, w32229, w32230, w32231, w32232, w32233, w32234, w32235, w32236, w32237, w32238, w32239, w32240, w32241, w32242, w32243, w32244, w32245, w32246, w32247, w32248, w32249, w32250, w32251, w32252, w32253, w32254, w32255, w32256, w32257, w32258, w32259, w32260, w32261, w32262, w32263, w32264, w32265, w32266, w32267, w32268, w32269, w32270, w32271, w32272, w32273, w32274, w32275, w32276, w32277, w32278, w32279, w32280, w32281, w32282, w32283, w32284, w32285, w32286, w32287, w32288, w32289, w32290, w32291, w32292, w32293, w32294, w32295, w32296, w32297, w32298, w32299, w32300, w32301, w32302, w32303, w32304, w32305, w32306, w32307, w32308, w32309, w32310, w32311, w32312, w32313, w32314, w32315, w32316, w32317, w32318, w32319, w32320, w32321, w32322, w32323, w32324, w32325, w32326, w32327, w32328, w32329, w32330, w32331, w32332, w32333, w32334, w32335, w32336, w32337, w32338, w32339, w32340, w32341, w32342, w32343, w32344, w32345, w32346, w32347, w32348, w32349, w32350, w32351, w32352, w32353, w32354, w32355, w32356, w32357, w32358, w32359, w32360, w32361, w32362, w32363, w32364, w32365, w32366, w32367, w32368, w32369, w32370, w32371, w32372, w32373, w32374, w32375, w32376, w32377, w32378, w32379, w32380, w32381, w32382, w32383, w32384, w32385, w32386, w32387, w32388, w32389, w32390, w32391, w32392, w32393, w32394, w32395, w32396, w32397, w32398, w32399, w32400, w32401, w32402, w32403, w32404, w32405, w32406, w32407, w32408, w32409, w32410, w32411, w32412, w32413, w32414, w32415, w32416, w32417, w32418, w32419, w32420, w32421, w32422, w32423, w32424, w32425, w32426, w32427, w32428, w32429, w32430, w32431, w32432, w32433, w32434, w32435, w32436, w32437, w32438, w32439, w32440, w32441, w32442, w32443, w32444, w32445, w32446, w32447, w32448, w32449, w32450, w32451, w32452, w32453, w32454, w32455, w32456, w32457, w32458, w32459, w32460, w32461, w32462, w32463, w32464, w32465, w32466, w32467, w32468, w32469, w32470, w32471, w32472, w32473, w32474, w32475, w32476, w32477, w32478, w32479, w32480, w32481, w32482, w32483, w32484, w32485, w32486, w32487, w32488, w32489, w32490, w32491, w32492, w32493, w32494, w32495, w32496, w32497, w32498, w32499, w32500, w32501, w32502, w32503, w32504, w32505, w32506, w32507, w32508, w32509, w32510, w32511, w32512, w32513, w32514, w32515, w32516, w32517, w32518, w32519, w32520, w32521, w32522, w32523, w32524, w32525, w32526, w32527, w32528, w32529, w32530, w32531, w32532, w32533, w32534, w32535, w32536, w32537, w32538, w32539, w32540, w32541, w32542, w32543, w32544, w32545, w32546, w32547, w32548, w32549, w32550, w32551, w32552, w32553, w32554, w32555, w32556, w32557, w32558, w32559, w32560, w32561, w32562, w32563, w32564, w32565, w32566, w32567, w32568, w32569, w32570, w32571, w32572, w32573, w32574, w32575, w32576, w32577, w32578, w32579, w32580, w32581, w32582, w32583, w32584, w32585, w32586, w32587, w32588, w32589, w32590, w32591, w32592, w32593, w32594, w32595, w32596, w32597, w32598, w32599, w32600, w32601, w32602, w32603, w32604, w32605, w32606, w32607, w32608, w32609, w32610, w32611, w32612, w32613, w32614, w32615, w32616, w32617, w32618, w32619, w32620, w32621, w32622, w32623, w32624, w32625, w32626, w32627, w32628, w32629, w32630, w32631, w32632, w32633, w32634, w32635, w32636, w32637, w32638, w32639, w32640, w32641, w32642, w32643, w32644, w32645, w32646, w32647, w32648, w32649, w32650, w32651, w32652, w32653, w32654, w32655, w32656, w32657, w32658, w32659, w32660, w32661, w32662, w32663, w32664, w32665, w32666, w32667, w32668, w32669, w32670, w32671, w32672, w32673, w32674, w32675, w32676, w32677, w32678, w32679, w32680, w32681, w32682, w32683, w32684, w32685, w32686, w32687, w32688, w32689, w32690, w32691, w32692, w32693, w32694, w32695, w32696, w32697, w32698, w32699, w32700, w32701, w32702, w32703, w32704, w32705, w32706, w32707, w32708, w32709, w32710, w32711, w32712, w32713, w32714, w32715, w32716, w32717, w32718, w32719, w32720, w32721, w32722, w32723, w32724, w32725, w32726, w32727, w32728, w32729, w32730, w32731, w32732, w32733, w32734, w32735, w32736, w32737, w32738, w32739, w32740, w32741, w32742, w32743, w32744, w32745, w32746, w32747, w32748, w32749, w32750, w32751, w32752, w32753, w32754, w32755, w32756, w32757, w32758, w32759, w32760, w32761, w32762, w32763, w32764, w32765, w32766, w32767, w32768, w32769, w32770, w32771, w32772, w32773, w32774, w32775, w32776, w32777, w32778, w32779, w32780, w32781, w32782, w32783, w32784, w32785, w32786, w32787, w32788, w32789, w32790, w32791, w32792, w32793, w32794, w32795, w32796, w32797, w32798, w32799, w32800, w32801, w32802, w32803, w32804, w32805, w32806, w32807, w32808, w32809, w32810, w32811, w32812, w32813, w32814, w32815, w32816, w32817, w32818, w32819, w32820, w32821, w32822, w32823, w32824, w32825, w32826, w32827, w32828, w32829, w32830, w32831, w32832, w32833, w32834, w32835, w32836, w32837, w32838, w32839, w32840, w32841, w32842, w32843, w32844, w32845, w32846, w32847, w32848, w32849, w32850, w32851, w32852, w32853, w32854, w32855, w32856, w32857, w32858, w32859, w32860, w32861, w32862, w32863, w32864, w32865, w32866, w32867, w32868, w32869, w32870, w32871, w32872, w32873, w32874, w32875, w32876, w32877, w32878, w32879, w32880, w32881, w32882, w32883, w32884, w32885, w32886, w32887, w32888, w32889, w32890, w32891, w32892, w32893, w32894, w32895, w32896, w32897, w32898, w32899, w32900, w32901, w32902, w32903, w32904, w32905, w32906, w32907, w32908, w32909, w32910, w32911, w32912, w32913, w32914, w32915, w32916, w32917, w32918, w32919, w32920, w32921, w32922, w32923, w32924, w32925, w32926, w32927, w32928, w32929, w32930, w32931, w32932, w32933, w32934, w32935, w32936, w32937, w32938, w32939, w32940, w32941, w32942, w32943, w32944, w32945, w32946, w32947, w32948, w32949, w32950, w32951, w32952, w32953, w32954, w32955, w32956, w32957, w32958, w32959, w32960, w32961, w32962, w32963, w32964, w32965, w32966, w32967, w32968, w32969, w32970, w32971, w32972, w32973, w32974, w32975, w32976, w32977, w32978, w32979, w32980, w32981, w32982, w32983, w32984, w32985, w32986, w32987, w32988, w32989, w32990, w32991, w32992, w32993, w32994, w32995, w32996, w32997, w32998, w32999, w33000, w33001, w33002, w33003, w33004, w33005, w33006, w33007, w33008, w33009, w33010, w33011, w33012, w33013, w33014, w33015, w33016, w33017, w33018, w33019, w33020, w33021, w33022, w33023, w33024, w33025, w33026, w33027, w33028, w33029, w33030, w33031, w33032, w33033, w33034, w33035, w33036, w33037, w33038, w33039, w33040, w33041, w33042, w33043, w33044, w33045, w33046, w33047, w33048, w33049, w33050, w33051, w33052, w33053, w33054, w33055, w33056, w33057, w33058, w33059, w33060, w33061, w33062, w33063, w33064, w33065, w33066, w33067, w33068, w33069, w33070, w33071, w33072, w33073, w33074, w33075, w33076, w33077, w33078, w33079, w33080, w33081, w33082, w33083, w33084, w33085, w33086, w33087, w33088, w33089, w33090, w33091, w33092, w33093, w33094, w33095, w33096, w33097, w33098, w33099, w33100, w33101, w33102, w33103, w33104, w33105, w33106, w33107, w33108, w33109, w33110, w33111, w33112, w33113, w33114, w33115, w33116, w33117, w33118, w33119, w33120, w33121, w33122, w33123, w33124, w33125, w33126, w33127, w33128, w33129, w33130, w33131, w33132, w33133, w33134, w33135, w33136, w33137, w33138, w33139, w33140, w33141, w33142, w33143, w33144, w33145, w33146, w33147, w33148, w33149, w33150, w33151, w33152, w33153, w33154, w33155, w33156, w33157, w33158, w33159, w33160, w33161, w33162, w33163, w33164, w33165, w33166, w33167, w33168, w33169, w33170, w33171, w33172, w33173, w33174, w33175, w33176, w33177, w33178, w33179, w33180, w33181, w33182, w33183, w33184, w33185, w33186, w33187, w33188, w33189, w33190, w33191, w33192, w33193, w33194, w33195, w33196, w33197, w33198, w33199, w33200, w33201, w33202, w33203, w33204, w33205, w33206, w33207, w33208, w33209, w33210, w33211, w33212, w33213, w33214, w33215, w33216, w33217, w33218, w33219, w33220, w33221, w33222, w33223, w33224, w33225, w33226, w33227, w33228, w33229, w33230, w33231, w33232, w33233, w33234, w33235, w33236, w33237, w33238, w33239, w33240, w33241, w33242, w33243, w33244, w33245, w33246, w33247, w33248, w33249, w33250, w33251, w33252, w33253, w33254, w33255, w33256, w33257, w33258, w33259, w33260, w33261, w33262, w33263, w33264, w33265, w33266, w33267, w33268, w33269, w33270, w33271, w33272, w33273, w33274, w33275, w33276, w33277, w33278, w33279, w33280, w33281, w33282, w33283, w33284, w33285, w33286, w33287, w33288, w33289, w33290, w33291, w33292, w33293, w33294, w33295, w33296, w33297, w33298, w33299, w33300, w33301, w33302, w33303, w33304, w33305, w33306, w33307, w33308, w33309, w33310, w33311, w33312, w33313, w33314, w33315, w33316, w33317, w33318, w33319, w33320, w33321, w33322, w33323, w33324, w33325, w33326, w33327, w33328, w33329, w33330, w33331, w33332, w33333, w33334, w33335, w33336, w33337, w33338, w33339, w33340, w33341, w33342, w33343, w33344, w33345, w33346, w33347, w33348, w33349, w33350, w33351, w33352, w33353, w33354, w33355, w33356, w33357, w33358, w33359, w33360, w33361, w33362, w33363, w33364, w33365, w33366, w33367, w33368, w33369, w33370, w33371, w33372, w33373, w33374, w33375, w33376, w33377, w33378, w33379, w33380, w33381, w33382, w33383, w33384, w33385, w33386, w33387, w33388, w33389, w33390, w33391, w33392, w33393, w33394, w33395, w33396, w33397, w33398, w33399, w33400, w33401, w33402, w33403, w33404, w33405, w33406, w33407, w33408, w33409, w33410, w33411, w33412, w33413, w33414, w33415, w33416, w33417, w33418, w33419, w33420, w33421, w33422, w33423, w33424, w33425, w33426, w33427, w33428, w33429, w33430, w33431, w33432, w33433, w33434, w33435, w33436, w33437, w33438, w33439, w33440, w33441, w33442, w33443, w33444, w33445, w33446, w33447, w33448, w33449, w33450, w33451, w33452, w33453, w33454, w33455, w33456, w33457, w33458, w33459, w33460, w33461, w33462, w33463, w33464, w33465, w33466, w33467, w33468, w33469, w33470, w33471, w33472, w33473, w33474, w33475, w33476, w33477, w33478, w33479, w33480, w33481, w33482, w33483, w33484, w33485, w33486, w33487, w33488, w33489, w33490, w33491, w33492, w33493, w33494, w33495, w33496, w33497, w33498, w33499, w33500, w33501, w33502, w33503, w33504, w33505, w33506, w33507, w33508, w33509, w33510, w33511, w33512, w33513, w33514, w33515, w33516, w33517, w33518, w33519, w33520, w33521, w33522, w33523, w33524, w33525, w33526, w33527, w33528, w33529, w33530, w33531, w33532, w33533, w33534, w33535, w33536, w33537, w33538, w33539, w33540, w33541, w33542, w33543, w33544, w33545, w33546, w33547, w33548, w33549, w33550, w33551, w33552, w33553, w33554, w33555, w33556, w33557, w33558, w33559, w33560, w33561, w33562, w33563, w33564, w33565, w33566, w33567, w33568, w33569, w33570, w33571, w33572, w33573, w33574, w33575, w33576, w33577, w33578, w33579, w33580, w33581, w33582, w33583, w33584, w33585, w33586, w33587, w33588, w33589, w33590, w33591, w33592, w33593, w33594, w33595, w33596, w33597, w33598, w33599, w33600, w33601, w33602, w33603, w33604, w33605, w33606, w33607, w33608, w33609, w33610, w33611, w33612, w33613, w33614, w33615, w33616, w33617, w33618, w33619, w33620, w33621, w33622, w33623, w33624, w33625, w33626, w33627, w33628, w33629, w33630, w33631, w33632, w33633, w33634, w33635, w33636, w33637, w33638, w33639, w33640, w33641, w33642, w33643, w33644, w33645, w33646, w33647, w33648, w33649, w33650, w33651, w33652, w33653, w33654, w33655, w33656, w33657, w33658, w33659, w33660, w33661, w33662, w33663, w33664, w33665, w33666, w33667, w33668, w33669, w33670, w33671, w33672, w33673, w33674, w33675, w33676, w33677, w33678, w33679, w33680, w33681, w33682, w33683, w33684, w33685, w33686, w33687, w33688, w33689, w33690, w33691, w33692, w33693, w33694, w33695, w33696, w33697, w33698, w33699, w33700, w33701, w33702, w33703, w33704, w33705, w33706, w33707, w33708, w33709, w33710, w33711, w33712, w33713, w33714, w33715, w33716, w33717, w33718, w33719, w33720, w33721, w33722, w33723, w33724, w33725, w33726, w33727, w33728, w33729, w33730, w33731, w33732, w33733, w33734, w33735, w33736, w33737, w33738, w33739, w33740, w33741, w33742, w33743, w33744, w33745, w33746, w33747, w33748, w33749, w33750, w33751, w33752, w33753, w33754, w33755, w33756, w33757, w33758, w33759, w33760, w33761, w33762, w33763, w33764, w33765, w33766, w33767, w33768, w33769, w33770, w33771, w33772, w33773, w33774, w33775, w33776, w33777, w33778, w33779, w33780, w33781, w33782, w33783, w33784, w33785, w33786, w33787, w33788, w33789, w33790, w33791, w33792, w33793, w33794, w33795, w33796, w33797, w33798, w33799, w33800, w33801, w33802, w33803, w33804, w33805, w33806, w33807, w33808, w33809, w33810, w33811, w33812, w33813, w33814, w33815, w33816, w33817, w33818, w33819, w33820, w33821, w33822, w33823, w33824, w33825, w33826, w33827, w33828, w33829, w33830, w33831, w33832, w33833, w33834, w33835, w33836, w33837, w33838, w33839, w33840, w33841, w33842, w33843, w33844, w33845, w33846, w33847, w33848, w33849, w33850, w33851, w33852, w33853, w33854, w33855, w33856, w33857, w33858, w33859, w33860, w33861, w33862, w33863, w33864, w33865, w33866, w33867, w33868, w33869, w33870, w33871, w33872, w33873, w33874, w33875, w33876, w33877, w33878, w33879, w33880, w33881, w33882, w33883, w33884, w33885, w33886, w33887, w33888, w33889, w33890, w33891, w33892, w33893, w33894, w33895, w33896, w33897, w33898, w33899, w33900, w33901, w33902, w33903, w33904, w33905, w33906, w33907, w33908, w33909, w33910, w33911, w33912, w33913, w33914, w33915, w33916, w33917, w33918, w33919, w33920, w33921, w33922, w33923, w33924, w33925, w33926, w33927, w33928, w33929, w33930, w33931, w33932, w33933, w33934, w33935, w33936, w33937, w33938, w33939, w33940, w33941, w33942, w33943, w33944, w33945, w33946, w33947, w33948, w33949, w33950, w33951, w33952, w33953, w33954, w33955, w33956, w33957, w33958, w33959, w33960, w33961, w33962, w33963, w33964, w33965, w33966, w33967, w33968, w33969, w33970, w33971, w33972, w33973, w33974, w33975, w33976, w33977, w33978, w33979, w33980, w33981, w33982, w33983, w33984, w33985, w33986, w33987, w33988, w33989, w33990, w33991, w33992, w33993, w33994, w33995, w33996, w33997, w33998, w33999, w34000, w34001, w34002, w34003, w34004, w34005, w34006, w34007, w34008, w34009, w34010, w34011, w34012, w34013, w34014, w34015, w34016, w34017, w34018, w34019, w34020, w34021, w34022, w34023, w34024, w34025, w34026, w34027, w34028, w34029, w34030, w34031, w34032, w34033, w34034, w34035, w34036, w34037, w34038, w34039, w34040, w34041, w34042, w34043, w34044, w34045, w34046, w34047, w34048, w34049, w34050, w34051, w34052, w34053, w34054, w34055, w34056, w34057, w34058, w34059, w34060, w34061, w34062, w34063, w34064, w34065, w34066, w34067, w34068, w34069, w34070, w34071, w34072, w34073, w34074, w34075, w34076, w34077, w34078, w34079, w34080, w34081, w34082, w34083, w34084, w34085, w34086, w34087, w34088, w34089, w34090, w34091, w34092, w34093, w34094, w34095, w34096, w34097, w34098, w34099, w34100, w34101, w34102, w34103, w34104, w34105, w34106, w34107, w34108, w34109, w34110, w34111, w34112, w34113, w34114, w34115, w34116, w34117, w34118, w34119, w34120, w34121, w34122, w34123, w34124, w34125, w34126, w34127, w34128, w34129, w34130, w34131, w34132, w34133, w34134, w34135, w34136, w34137, w34138, w34139, w34140, w34141, w34142, w34143, w34144, w34145, w34146, w34147, w34148, w34149, w34150, w34151, w34152, w34153, w34154, w34155, w34156, w34157, w34158, w34159, w34160, w34161, w34162, w34163, w34164, w34165, w34166, w34167, w34168, w34169, w34170, w34171, w34172, w34173, w34174, w34175, w34176, w34177, w34178, w34179, w34180, w34181, w34182, w34183, w34184, w34185, w34186, w34187, w34188, w34189, w34190, w34191, w34192, w34193, w34194, w34195, w34196, w34197, w34198, w34199, w34200, w34201, w34202, w34203, w34204, w34205, w34206, w34207, w34208, w34209, w34210, w34211, w34212, w34213, w34214, w34215, w34216, w34217, w34218, w34219, w34220, w34221, w34222, w34223, w34224, w34225, w34226, w34227, w34228, w34229, w34230, w34231, w34232, w34233, w34234, w34235, w34236, w34237, w34238, w34239, w34240, w34241, w34242, w34243, w34244, w34245, w34246, w34247, w34248, w34249, w34250, w34251, w34252, w34253, w34254, w34255, w34256, w34257, w34258, w34259, w34260, w34261, w34262, w34263, w34264, w34265, w34266, w34267, w34268, w34269, w34270, w34271, w34272, w34273, w34274, w34275, w34276, w34277, w34278, w34279, w34280, w34281, w34282, w34283, w34284, w34285, w34286, w34287, w34288, w34289, w34290, w34291, w34292, w34293, w34294, w34295, w34296, w34297, w34298, w34299, w34300, w34301, w34302, w34303, w34304, w34305, w34306, w34307, w34308, w34309, w34310, w34311, w34312, w34313, w34314, w34315, w34316, w34317, w34318, w34319, w34320, w34321, w34322, w34323, w34324, w34325, w34326, w34327, w34328, w34329, w34330, w34331, w34332, w34333, w34334, w34335, w34336, w34337, w34338, w34339, w34340, w34341, w34342, w34343, w34344, w34345, w34346, w34347, w34348, w34349, w34350, w34351, w34352, w34353, w34354, w34355, w34356, w34357, w34358, w34359, w34360, w34361, w34362, w34363, w34364, w34365, w34366, w34367, w34368, w34369, w34370, w34371, w34372, w34373, w34374, w34375, w34376, w34377, w34378, w34379, w34380, w34381, w34382, w34383, w34384, w34385, w34386, w34387, w34388, w34389, w34390, w34391, w34392, w34393, w34394, w34395, w34396, w34397, w34398, w34399, w34400, w34401, w34402, w34403, w34404, w34405, w34406, w34407, w34408, w34409, w34410, w34411, w34412, w34413, w34414, w34415, w34416, w34417, w34418, w34419, w34420, w34421, w34422, w34423, w34424, w34425, w34426, w34427, w34428, w34429, w34430, w34431, w34432, w34433, w34434, w34435, w34436, w34437, w34438, w34439, w34440, w34441, w34442, w34443, w34444, w34445, w34446, w34447, w34448, w34449, w34450, w34451, w34452, w34453, w34454, w34455, w34456, w34457, w34458, w34459, w34460, w34461, w34462, w34463, w34464, w34465, w34466, w34467, w34468, w34469, w34470, w34471, w34472, w34473, w34474, w34475, w34476, w34477, w34478, w34479, w34480, w34481, w34482, w34483, w34484, w34485, w34486, w34487, w34488, w34489, w34490, w34491, w34492, w34493, w34494, w34495, w34496, w34497, w34498, w34499, w34500, w34501, w34502, w34503, w34504, w34505, w34506, w34507, w34508, w34509, w34510, w34511, w34512, w34513, w34514, w34515, w34516, w34517, w34518, w34519, w34520, w34521, w34522, w34523, w34524, w34525, w34526, w34527, w34528, w34529, w34530, w34531, w34532, w34533, w34534, w34535, w34536, w34537, w34538, w34539, w34540, w34541, w34542, w34543, w34544, w34545, w34546, w34547, w34548, w34549, w34550, w34551, w34552, w34553, w34554, w34555, w34556, w34557, w34558, w34559, w34560, w34561, w34562, w34563, w34564, w34565, w34566, w34567, w34568, w34569, w34570, w34571, w34572, w34573, w34574, w34575, w34576, w34577, w34578, w34579, w34580, w34581, w34582, w34583, w34584, w34585, w34586, w34587, w34588, w34589, w34590, w34591, w34592, w34593, w34594, w34595, w34596, w34597, w34598, w34599, w34600, w34601, w34602, w34603, w34604, w34605, w34606, w34607, w34608, w34609, w34610, w34611, w34612, w34613, w34614, w34615, w34616, w34617, w34618, w34619, w34620, w34621, w34622, w34623, w34624, w34625, w34626, w34627, w34628, w34629, w34630, w34631, w34632, w34633, w34634, w34635, w34636, w34637, w34638, w34639, w34640, w34641, w34642, w34643, w34644, w34645, w34646, w34647, w34648, w34649, w34650, w34651, w34652, w34653, w34654, w34655, w34656, w34657, w34658, w34659, w34660, w34661, w34662, w34663, w34664, w34665, w34666, w34667, w34668, w34669, w34670, w34671, w34672, w34673, w34674, w34675, w34676, w34677, w34678, w34679, w34680, w34681, w34682, w34683, w34684, w34685, w34686, w34687, w34688, w34689, w34690, w34691, w34692, w34693, w34694, w34695, w34696, w34697, w34698, w34699, w34700, w34701, w34702, w34703, w34704, w34705, w34706, w34707, w34708, w34709, w34710, w34711, w34712, w34713, w34714, w34715, w34716, w34717, w34718, w34719, w34720, w34721, w34722, w34723, w34724, w34725, w34726, w34727, w34728, w34729, w34730, w34731, w34732, w34733, w34734, w34735, w34736, w34737, w34738, w34739, w34740, w34741, w34742, w34743, w34744, w34745, w34746, w34747, w34748, w34749, w34750, w34751, w34752, w34753, w34754, w34755, w34756, w34757, w34758, w34759, w34760, w34761, w34762, w34763, w34764, w34765, w34766, w34767, w34768, w34769, w34770, w34771, w34772, w34773, w34774, w34775, w34776, w34777, w34778, w34779, w34780, w34781, w34782, w34783, w34784, w34785, w34786, w34787, w34788, w34789, w34790, w34791, w34792, w34793, w34794, w34795, w34796, w34797, w34798, w34799, w34800, w34801, w34802, w34803, w34804, w34805, w34806, w34807, w34808, w34809, w34810, w34811, w34812, w34813, w34814, w34815, w34816, w34817, w34818, w34819, w34820, w34821, w34822, w34823, w34824, w34825, w34826, w34827, w34828, w34829, w34830, w34831, w34832, w34833, w34834, w34835, w34836, w34837, w34838, w34839, w34840, w34841, w34842, w34843, w34844, w34845, w34846, w34847, w34848, w34849, w34850, w34851, w34852, w34853, w34854, w34855, w34856, w34857, w34858, w34859, w34860, w34861, w34862, w34863, w34864, w34865, w34866, w34867, w34868, w34869, w34870, w34871, w34872, w34873, w34874, w34875, w34876, w34877, w34878, w34879, w34880, w34881, w34882, w34883, w34884, w34885, w34886, w34887, w34888, w34889, w34890, w34891, w34892, w34893, w34894, w34895, w34896, w34897, w34898, w34899, w34900, w34901, w34902, w34903, w34904, w34905, w34906, w34907, w34908, w34909, w34910, w34911, w34912, w34913, w34914, w34915, w34916, w34917, w34918, w34919, w34920, w34921, w34922, w34923, w34924, w34925, w34926, w34927, w34928, w34929, w34930, w34931, w34932, w34933, w34934, w34935, w34936, w34937, w34938, w34939, w34940, w34941, w34942, w34943, w34944, w34945, w34946, w34947, w34948, w34949, w34950, w34951, w34952, w34953, w34954, w34955, w34956, w34957, w34958, w34959, w34960, w34961, w34962, w34963, w34964, w34965, w34966, w34967, w34968, w34969, w34970, w34971, w34972, w34973, w34974, w34975, w34976, w34977, w34978, w34979, w34980, w34981, w34982, w34983, w34984, w34985, w34986, w34987, w34988, w34989, w34990, w34991, w34992, w34993, w34994, w34995, w34996, w34997, w34998, w34999, w35000, w35001, w35002, w35003, w35004, w35005, w35006, w35007, w35008, w35009, w35010, w35011, w35012, w35013, w35014, w35015, w35016, w35017, w35018, w35019, w35020, w35021, w35022, w35023, w35024, w35025, w35026, w35027, w35028, w35029, w35030, w35031, w35032, w35033, w35034, w35035, w35036, w35037, w35038, w35039, w35040, w35041, w35042, w35043, w35044, w35045, w35046, w35047, w35048, w35049, w35050, w35051, w35052, w35053, w35054, w35055, w35056, w35057, w35058, w35059, w35060, w35061, w35062, w35063, w35064, w35065, w35066, w35067, w35068, w35069, w35070, w35071, w35072, w35073, w35074, w35075, w35076, w35077, w35078, w35079, w35080, w35081, w35082, w35083, w35084, w35085, w35086, w35087, w35088, w35089, w35090, w35091, w35092, w35093, w35094, w35095, w35096, w35097, w35098, w35099, w35100, w35101, w35102, w35103, w35104, w35105, w35106, w35107, w35108, w35109, w35110, w35111, w35112, w35113, w35114, w35115, w35116, w35117, w35118, w35119, w35120, w35121, w35122, w35123, w35124, w35125, w35126, w35127, w35128, w35129, w35130, w35131, w35132, w35133, w35134, w35135, w35136, w35137, w35138, w35139, w35140, w35141, w35142, w35143, w35144, w35145, w35146, w35147, w35148, w35149, w35150, w35151, w35152, w35153, w35154, w35155, w35156, w35157, w35158, w35159, w35160, w35161, w35162, w35163, w35164, w35165, w35166, w35167, w35168, w35169, w35170, w35171, w35172, w35173, w35174, w35175, w35176, w35177, w35178, w35179, w35180, w35181, w35182, w35183, w35184, w35185, w35186, w35187, w35188, w35189, w35190, w35191, w35192, w35193, w35194, w35195, w35196, w35197, w35198, w35199, w35200, w35201, w35202, w35203, w35204, w35205, w35206, w35207, w35208, w35209, w35210, w35211, w35212, w35213, w35214, w35215, w35216, w35217, w35218, w35219, w35220, w35221, w35222, w35223, w35224, w35225, w35226, w35227, w35228, w35229, w35230, w35231, w35232, w35233, w35234, w35235, w35236, w35237, w35238, w35239, w35240, w35241, w35242, w35243, w35244, w35245, w35246, w35247, w35248, w35249, w35250, w35251, w35252, w35253, w35254, w35255, w35256, w35257, w35258, w35259, w35260, w35261, w35262, w35263, w35264, w35265, w35266, w35267, w35268, w35269, w35270, w35271, w35272, w35273, w35274, w35275, w35276, w35277, w35278, w35279, w35280, w35281, w35282, w35283, w35284, w35285, w35286, w35287, w35288, w35289, w35290, w35291, w35292, w35293, w35294, w35295, w35296, w35297, w35298, w35299, w35300, w35301, w35302, w35303, w35304, w35305, w35306, w35307, w35308, w35309, w35310, w35311, w35312, w35313, w35314, w35315, w35316, w35317, w35318, w35319, w35320, w35321, w35322, w35323, w35324, w35325, w35326, w35327, w35328, w35329, w35330, w35331, w35332, w35333, w35334, w35335, w35336, w35337, w35338, w35339, w35340, w35341, w35342, w35343, w35344, w35345, w35346, w35347, w35348, w35349, w35350, w35351, w35352, w35353, w35354, w35355, w35356, w35357, w35358, w35359, w35360, w35361, w35362, w35363, w35364, w35365, w35366, w35367, w35368, w35369, w35370, w35371, w35372, w35373, w35374, w35375, w35376, w35377, w35378, w35379, w35380, w35381, w35382, w35383, w35384, w35385, w35386, w35387, w35388, w35389, w35390, w35391, w35392, w35393, w35394, w35395, w35396, w35397, w35398, w35399, w35400, w35401, w35402, w35403, w35404, w35405, w35406, w35407, w35408, w35409, w35410, w35411, w35412, w35413, w35414, w35415, w35416, w35417, w35418, w35419, w35420, w35421, w35422, w35423, w35424, w35425, w35426, w35427, w35428, w35429, w35430, w35431, w35432, w35433, w35434, w35435, w35436, w35437, w35438, w35439, w35440, w35441, w35442, w35443, w35444, w35445, w35446, w35447, w35448, w35449, w35450, w35451, w35452, w35453, w35454, w35455, w35456, w35457, w35458, w35459, w35460, w35461, w35462, w35463, w35464, w35465, w35466, w35467, w35468, w35469, w35470, w35471, w35472, w35473, w35474, w35475, w35476, w35477, w35478, w35479, w35480, w35481, w35482, w35483, w35484, w35485, w35486, w35487, w35488, w35489, w35490, w35491, w35492, w35493, w35494, w35495, w35496, w35497, w35498, w35499, w35500, w35501, w35502, w35503, w35504, w35505, w35506, w35507, w35508, w35509, w35510, w35511, w35512, w35513, w35514, w35515, w35516, w35517, w35518, w35519, w35520, w35521, w35522, w35523, w35524, w35525, w35526, w35527, w35528, w35529, w35530, w35531, w35532, w35533, w35534, w35535, w35536, w35537, w35538, w35539, w35540, w35541, w35542, w35543, w35544, w35545, w35546, w35547, w35548, w35549, w35550, w35551, w35552, w35553, w35554, w35555, w35556, w35557, w35558, w35559, w35560, w35561, w35562, w35563, w35564, w35565, w35566, w35567, w35568, w35569, w35570, w35571, w35572, w35573, w35574, w35575, w35576, w35577, w35578, w35579, w35580, w35581, w35582, w35583, w35584, w35585, w35586, w35587, w35588, w35589, w35590, w35591, w35592, w35593, w35594, w35595, w35596, w35597, w35598, w35599, w35600, w35601, w35602, w35603, w35604, w35605, w35606, w35607, w35608, w35609, w35610, w35611, w35612, w35613, w35614, w35615, w35616, w35617, w35618, w35619, w35620, w35621, w35622, w35623, w35624, w35625, w35626, w35627, w35628, w35629, w35630, w35631, w35632, w35633, w35634, w35635, w35636, w35637, w35638, w35639, w35640, w35641, w35642, w35643, w35644, w35645, w35646, w35647, w35648, w35649, w35650, w35651, w35652, w35653, w35654, w35655, w35656, w35657, w35658, w35659, w35660, w35661, w35662, w35663, w35664, w35665, w35666, w35667, w35668, w35669, w35670, w35671, w35672, w35673, w35674, w35675, w35676, w35677, w35678, w35679, w35680, w35681, w35682, w35683, w35684, w35685, w35686, w35687, w35688, w35689, w35690, w35691, w35692, w35693, w35694, w35695, w35696, w35697, w35698, w35699, w35700, w35701, w35702, w35703, w35704, w35705, w35706, w35707, w35708, w35709, w35710, w35711, w35712, w35713, w35714, w35715, w35716, w35717, w35718, w35719, w35720, w35721, w35722, w35723, w35724, w35725, w35726, w35727, w35728, w35729, w35730, w35731, w35732, w35733, w35734, w35735, w35736, w35737, w35738, w35739, w35740, w35741, w35742, w35743, w35744, w35745, w35746, w35747, w35748, w35749, w35750, w35751, w35752, w35753, w35754, w35755, w35756, w35757, w35758, w35759, w35760, w35761, w35762, w35763, w35764, w35765, w35766, w35767, w35768, w35769, w35770, w35771, w35772, w35773, w35774, w35775, w35776, w35777, w35778, w35779, w35780, w35781, w35782, w35783, w35784, w35785, w35786, w35787, w35788, w35789, w35790, w35791, w35792, w35793, w35794, w35795, w35796, w35797, w35798, w35799, w35800, w35801, w35802, w35803, w35804, w35805, w35806, w35807, w35808, w35809, w35810, w35811, w35812, w35813, w35814, w35815, w35816, w35817, w35818, w35819, w35820, w35821, w35822, w35823, w35824, w35825, w35826, w35827, w35828, w35829, w35830, w35831, w35832, w35833, w35834, w35835, w35836, w35837, w35838, w35839, w35840, w35841, w35842, w35843, w35844, w35845, w35846, w35847, w35848, w35849, w35850, w35851, w35852, w35853, w35854, w35855, w35856, w35857, w35858, w35859, w35860, w35861, w35862, w35863, w35864, w35865, w35866, w35867, w35868, w35869, w35870, w35871, w35872, w35873, w35874, w35875, w35876, w35877, w35878, w35879, w35880, w35881, w35882, w35883, w35884, w35885, w35886, w35887, w35888, w35889, w35890, w35891, w35892, w35893, w35894, w35895, w35896, w35897, w35898, w35899, w35900, w35901, w35902, w35903, w35904, w35905, w35906, w35907, w35908, w35909, w35910, w35911, w35912, w35913, w35914, w35915, w35916, w35917, w35918, w35919, w35920, w35921, w35922, w35923, w35924, w35925, w35926, w35927, w35928, w35929, w35930, w35931, w35932, w35933, w35934, w35935, w35936, w35937, w35938, w35939, w35940, w35941, w35942, w35943, w35944, w35945, w35946, w35947, w35948, w35949, w35950, w35951, w35952, w35953, w35954, w35955, w35956, w35957, w35958, w35959, w35960, w35961, w35962, w35963, w35964, w35965, w35966, w35967, w35968, w35969, w35970, w35971, w35972, w35973, w35974, w35975, w35976, w35977, w35978, w35979, w35980, w35981, w35982, w35983, w35984, w35985, w35986, w35987, w35988, w35989, w35990, w35991, w35992, w35993, w35994, w35995, w35996, w35997, w35998, w35999, w36000, w36001, w36002, w36003, w36004, w36005, w36006, w36007, w36008, w36009, w36010, w36011, w36012, w36013, w36014, w36015, w36016, w36017, w36018, w36019, w36020, w36021, w36022, w36023, w36024, w36025, w36026, w36027, w36028, w36029, w36030, w36031, w36032, w36033, w36034, w36035, w36036, w36037, w36038, w36039, w36040, w36041, w36042, w36043, w36044, w36045, w36046, w36047, w36048, w36049, w36050, w36051, w36052, w36053, w36054, w36055, w36056, w36057, w36058, w36059, w36060, w36061, w36062, w36063, w36064, w36065, w36066, w36067, w36068, w36069, w36070, w36071, w36072, w36073, w36074, w36075, w36076, w36077, w36078, w36079, w36080, w36081, w36082, w36083, w36084, w36085, w36086, w36087, w36088, w36089, w36090, w36091, w36092, w36093, w36094, w36095, w36096, w36097, w36098, w36099, w36100, w36101, w36102, w36103, w36104, w36105, w36106, w36107, w36108, w36109, w36110, w36111, w36112, w36113, w36114, w36115, w36116, w36117, w36118, w36119, w36120, w36121, w36122, w36123, w36124, w36125, w36126, w36127, w36128, w36129, w36130, w36131, w36132, w36133, w36134, w36135, w36136, w36137, w36138, w36139, w36140, w36141, w36142, w36143, w36144, w36145, w36146, w36147, w36148, w36149, w36150, w36151, w36152, w36153, w36154, w36155, w36156, w36157, w36158, w36159, w36160, w36161, w36162, w36163, w36164, w36165, w36166, w36167, w36168, w36169, w36170, w36171, w36172, w36173, w36174, w36175, w36176, w36177, w36178, w36179, w36180, w36181, w36182, w36183, w36184, w36185, w36186, w36187, w36188, w36189, w36190, w36191, w36192, w36193, w36194, w36195, w36196, w36197, w36198, w36199, w36200, w36201, w36202, w36203, w36204, w36205, w36206, w36207, w36208, w36209, w36210, w36211, w36212, w36213, w36214, w36215, w36216, w36217, w36218, w36219, w36220, w36221, w36222, w36223, w36224, w36225, w36226, w36227, w36228, w36229, w36230, w36231, w36232, w36233, w36234, w36235, w36236, w36237, w36238, w36239, w36240, w36241, w36242, w36243, w36244, w36245, w36246, w36247, w36248, w36249, w36250, w36251, w36252, w36253, w36254, w36255, w36256, w36257, w36258, w36259, w36260, w36261, w36262, w36263, w36264, w36265, w36266, w36267, w36268, w36269, w36270, w36271, w36272, w36273, w36274, w36275, w36276, w36277, w36278, w36279, w36280, w36281, w36282, w36283, w36284, w36285, w36286, w36287, w36288, w36289, w36290, w36291, w36292, w36293, w36294, w36295, w36296, w36297, w36298, w36299, w36300, w36301, w36302, w36303, w36304, w36305, w36306, w36307, w36308, w36309, w36310, w36311, w36312, w36313, w36314, w36315, w36316, w36317, w36318, w36319, w36320, w36321, w36322, w36323, w36324, w36325, w36326, w36327, w36328, w36329, w36330, w36331, w36332, w36333, w36334, w36335, w36336, w36337, w36338, w36339, w36340, w36341, w36342, w36343, w36344, w36345, w36346, w36347, w36348, w36349, w36350, w36351, w36352, w36353, w36354, w36355, w36356, w36357, w36358, w36359, w36360, w36361, w36362, w36363, w36364, w36365, w36366, w36367, w36368, w36369, w36370, w36371, w36372, w36373, w36374, w36375, w36376, w36377, w36378, w36379, w36380, w36381, w36382, w36383, w36384, w36385, w36386, w36387, w36388, w36389, w36390, w36391, w36392, w36393, w36394, w36395, w36396, w36397, w36398, w36399, w36400, w36401, w36402, w36403, w36404, w36405, w36406, w36407, w36408, w36409, w36410, w36411, w36412, w36413, w36414, w36415, w36416, w36417, w36418, w36419, w36420, w36421, w36422, w36423, w36424, w36425, w36426, w36427, w36428, w36429, w36430, w36431, w36432, w36433, w36434, w36435, w36436, w36437, w36438, w36439, w36440, w36441, w36442, w36443, w36444, w36445, w36446, w36447, w36448, w36449, w36450, w36451, w36452, w36453, w36454, w36455, w36456, w36457, w36458, w36459, w36460, w36461, w36462, w36463, w36464, w36465, w36466, w36467, w36468, w36469, w36470, w36471, w36472, w36473, w36474, w36475, w36476, w36477, w36478, w36479, w36480, w36481, w36482, w36483, w36484, w36485, w36486, w36487, w36488, w36489, w36490, w36491, w36492, w36493, w36494, w36495, w36496, w36497, w36498, w36499, w36500, w36501, w36502, w36503, w36504, w36505, w36506, w36507, w36508, w36509, w36510, w36511, w36512, w36513, w36514, w36515, w36516, w36517, w36518, w36519, w36520, w36521, w36522, w36523, w36524, w36525, w36526, w36527, w36528, w36529, w36530, w36531, w36532, w36533, w36534, w36535, w36536, w36537, w36538, w36539, w36540, w36541, w36542, w36543, w36544, w36545, w36546, w36547, w36548, w36549, w36550, w36551, w36552, w36553, w36554, w36555, w36556, w36557, w36558, w36559, w36560, w36561, w36562, w36563, w36564, w36565, w36566, w36567, w36568, w36569, w36570, w36571, w36572, w36573, w36574, w36575, w36576, w36577, w36578, w36579, w36580, w36581, w36582, w36583, w36584, w36585, w36586, w36587, w36588, w36589, w36590, w36591, w36592, w36593, w36594, w36595, w36596, w36597, w36598, w36599, w36600, w36601, w36602, w36603, w36604, w36605, w36606, w36607, w36608, w36609, w36610, w36611, w36612, w36613, w36614, w36615, w36616, w36617, w36618, w36619, w36620, w36621, w36622, w36623, w36624, w36625, w36626, w36627, w36628, w36629, w36630, w36631, w36632, w36633, w36634, w36635, w36636, w36637, w36638, w36639, w36640, w36641, w36642, w36643, w36644, w36645, w36646, w36647, w36648, w36649, w36650, w36651, w36652, w36653, w36654, w36655, w36656, w36657, w36658, w36659, w36660, w36661, w36662, w36663, w36664, w36665, w36666, w36667, w36668, w36669, w36670, w36671, w36672, w36673, w36674, w36675, w36676, w36677, w36678, w36679, w36680, w36681, w36682, w36683, w36684, w36685, w36686, w36687, w36688, w36689, w36690, w36691, w36692, w36693, w36694, w36695, w36696, w36697, w36698, w36699, w36700, w36701, w36702, w36703, w36704, w36705, w36706, w36707, w36708, w36709, w36710, w36711, w36712, w36713, w36714, w36715, w36716, w36717, w36718, w36719, w36720, w36721, w36722, w36723, w36724, w36725, w36726, w36727, w36728, w36729, w36730, w36731, w36732, w36733, w36734, w36735, w36736, w36737, w36738, w36739, w36740, w36741, w36742, w36743, w36744, w36745, w36746, w36747, w36748, w36749, w36750, w36751, w36752, w36753, w36754, w36755, w36756, w36757, w36758, w36759, w36760, w36761, w36762, w36763, w36764, w36765, w36766, w36767, w36768, w36769, w36770, w36771, w36772, w36773, w36774, w36775, w36776, w36777, w36778, w36779, w36780, w36781, w36782, w36783, w36784, w36785, w36786, w36787, w36788, w36789, w36790, w36791, w36792, w36793, w36794, w36795, w36796, w36797, w36798, w36799, w36800, w36801, w36802, w36803, w36804, w36805, w36806, w36807, w36808, w36809, w36810, w36811, w36812, w36813, w36814, w36815, w36816, w36817, w36818, w36819, w36820, w36821, w36822, w36823, w36824, w36825, w36826, w36827, w36828, w36829, w36830, w36831, w36832, w36833, w36834, w36835, w36836, w36837, w36838, w36839, w36840, w36841, w36842, w36843, w36844, w36845, w36846, w36847, w36848, w36849, w36850, w36851, w36852, w36853, w36854, w36855, w36856, w36857, w36858, w36859, w36860, w36861, w36862, w36863, w36864, w36865, w36866, w36867, w36868, w36869, w36870, w36871, w36872, w36873, w36874, w36875, w36876, w36877, w36878, w36879, w36880, w36881, w36882, w36883, w36884, w36885, w36886, w36887, w36888, w36889, w36890, w36891, w36892, w36893, w36894, w36895, w36896, w36897, w36898, w36899, w36900, w36901, w36902, w36903, w36904, w36905, w36906, w36907, w36908, w36909, w36910, w36911, w36912, w36913, w36914, w36915, w36916, w36917, w36918, w36919, w36920, w36921, w36922, w36923, w36924, w36925, w36926, w36927, w36928, w36929, w36930, w36931, w36932, w36933, w36934, w36935, w36936, w36937, w36938, w36939, w36940, w36941, w36942, w36943, w36944, w36945, w36946, w36947, w36948, w36949, w36950, w36951, w36952, w36953, w36954, w36955, w36956, w36957, w36958, w36959, w36960, w36961, w36962, w36963, w36964, w36965, w36966, w36967, w36968, w36969, w36970, w36971, w36972, w36973, w36974, w36975, w36976, w36977, w36978, w36979, w36980, w36981, w36982, w36983, w36984, w36985, w36986, w36987, w36988, w36989, w36990, w36991, w36992, w36993, w36994, w36995, w36996, w36997, w36998, w36999, w37000, w37001, w37002, w37003, w37004, w37005, w37006, w37007, w37008, w37009, w37010, w37011, w37012, w37013, w37014, w37015, w37016, w37017, w37018, w37019, w37020, w37021, w37022, w37023, w37024, w37025, w37026, w37027, w37028, w37029, w37030, w37031, w37032, w37033, w37034, w37035, w37036, w37037, w37038, w37039, w37040, w37041, w37042, w37043, w37044, w37045, w37046, w37047, w37048, w37049, w37050, w37051, w37052, w37053, w37054, w37055, w37056, w37057, w37058, w37059, w37060, w37061, w37062, w37063, w37064, w37065, w37066, w37067, w37068, w37069, w37070, w37071, w37072, w37073, w37074, w37075, w37076, w37077, w37078, w37079, w37080, w37081, w37082, w37083, w37084, w37085, w37086, w37087, w37088, w37089, w37090, w37091, w37092, w37093, w37094, w37095, w37096, w37097, w37098, w37099, w37100, w37101, w37102, w37103, w37104, w37105, w37106, w37107, w37108, w37109, w37110, w37111, w37112, w37113, w37114, w37115, w37116, w37117, w37118, w37119, w37120, w37121, w37122, w37123, w37124, w37125, w37126, w37127, w37128, w37129, w37130, w37131, w37132, w37133, w37134, w37135, w37136, w37137, w37138, w37139, w37140, w37141, w37142, w37143, w37144, w37145, w37146, w37147, w37148, w37149, w37150, w37151, w37152, w37153, w37154, w37155, w37156, w37157, w37158, w37159, w37160, w37161, w37162, w37163, w37164, w37165, w37166, w37167, w37168, w37169, w37170, w37171, w37172, w37173, w37174, w37175, w37176, w37177, w37178, w37179, w37180, w37181, w37182, w37183, w37184, w37185, w37186, w37187, w37188, w37189, w37190, w37191, w37192, w37193, w37194, w37195, w37196, w37197, w37198, w37199, w37200, w37201, w37202, w37203, w37204, w37205, w37206, w37207, w37208, w37209, w37210, w37211, w37212, w37213, w37214, w37215, w37216, w37217, w37218, w37219, w37220, w37221, w37222, w37223, w37224, w37225, w37226, w37227, w37228, w37229, w37230, w37231, w37232, w37233, w37234, w37235, w37236, w37237, w37238, w37239, w37240, w37241, w37242, w37243, w37244, w37245, w37246, w37247, w37248, w37249, w37250, w37251, w37252, w37253, w37254, w37255, w37256, w37257, w37258, w37259, w37260, w37261, w37262, w37263, w37264, w37265, w37266, w37267, w37268, w37269, w37270, w37271, w37272, w37273, w37274, w37275, w37276, w37277, w37278, w37279, w37280, w37281, w37282, w37283, w37284, w37285, w37286, w37287, w37288, w37289, w37290, w37291, w37292, w37293, w37294, w37295, w37296, w37297, w37298, w37299, w37300, w37301, w37302, w37303, w37304, w37305, w37306, w37307, w37308, w37309, w37310, w37311, w37312, w37313, w37314, w37315, w37316, w37317, w37318, w37319, w37320, w37321, w37322, w37323, w37324, w37325, w37326, w37327, w37328, w37329, w37330, w37331, w37332, w37333, w37334, w37335, w37336, w37337, w37338, w37339, w37340, w37341, w37342, w37343, w37344, w37345, w37346, w37347, w37348, w37349, w37350, w37351, w37352, w37353, w37354, w37355, w37356, w37357, w37358, w37359, w37360, w37361, w37362, w37363, w37364, w37365, w37366, w37367, w37368, w37369, w37370, w37371, w37372, w37373, w37374, w37375, w37376, w37377, w37378, w37379, w37380, w37381, w37382, w37383, w37384, w37385, w37386, w37387, w37388, w37389, w37390, w37391, w37392, w37393, w37394, w37395, w37396, w37397, w37398, w37399, w37400, w37401, w37402, w37403, w37404, w37405, w37406, w37407, w37408, w37409, w37410, w37411, w37412, w37413, w37414, w37415, w37416, w37417, w37418, w37419, w37420, w37421, w37422, w37423, w37424, w37425, w37426, w37427, w37428, w37429, w37430, w37431, w37432, w37433, w37434, w37435, w37436, w37437, w37438, w37439, w37440, w37441, w37442, w37443, w37444, w37445, w37446, w37447, w37448, w37449, w37450, w37451, w37452, w37453, w37454, w37455, w37456, w37457, w37458, w37459, w37460, w37461, w37462, w37463, w37464, w37465, w37466, w37467, w37468, w37469, w37470, w37471, w37472, w37473, w37474, w37475, w37476, w37477, w37478, w37479, w37480, w37481, w37482, w37483, w37484, w37485, w37486, w37487, w37488, w37489, w37490, w37491, w37492, w37493, w37494, w37495, w37496, w37497, w37498, w37499, w37500, w37501, w37502, w37503, w37504, w37505, w37506, w37507, w37508, w37509, w37510, w37511, w37512, w37513, w37514, w37515, w37516, w37517, w37518, w37519, w37520, w37521, w37522, w37523, w37524, w37525, w37526, w37527, w37528, w37529, w37530, w37531, w37532, w37533, w37534, w37535, w37536, w37537, w37538, w37539, w37540, w37541, w37542, w37543, w37544, w37545, w37546, w37547, w37548, w37549, w37550, w37551, w37552, w37553, w37554, w37555, w37556, w37557, w37558, w37559, w37560, w37561, w37562, w37563, w37564, w37565, w37566, w37567, w37568, w37569, w37570, w37571, w37572, w37573, w37574, w37575, w37576, w37577, w37578, w37579, w37580, w37581, w37582, w37583, w37584, w37585, w37586, w37587, w37588, w37589, w37590, w37591, w37592, w37593, w37594, w37595, w37596, w37597, w37598, w37599, w37600, w37601, w37602, w37603, w37604, w37605, w37606, w37607, w37608, w37609, w37610, w37611, w37612, w37613, w37614, w37615, w37616, w37617, w37618, w37619, w37620, w37621, w37622, w37623, w37624, w37625, w37626, w37627, w37628, w37629, w37630, w37631, w37632, w37633, w37634, w37635, w37636, w37637, w37638, w37639, w37640, w37641, w37642, w37643, w37644, w37645, w37646, w37647, w37648, w37649, w37650, w37651, w37652, w37653, w37654, w37655, w37656, w37657, w37658, w37659, w37660, w37661, w37662, w37663, w37664, w37665, w37666, w37667, w37668, w37669, w37670, w37671, w37672, w37673, w37674, w37675, w37676, w37677, w37678, w37679, w37680, w37681, w37682, w37683, w37684, w37685, w37686, w37687, w37688, w37689, w37690, w37691, w37692, w37693, w37694, w37695, w37696, w37697, w37698, w37699, w37700, w37701, w37702, w37703, w37704, w37705, w37706, w37707, w37708, w37709, w37710, w37711, w37712, w37713, w37714, w37715, w37716, w37717, w37718, w37719, w37720, w37721, w37722, w37723, w37724, w37725, w37726, w37727, w37728, w37729, w37730, w37731, w37732, w37733, w37734, w37735, w37736, w37737, w37738, w37739, w37740, w37741, w37742, w37743, w37744, w37745, w37746, w37747, w37748, w37749, w37750, w37751, w37752, w37753, w37754, w37755, w37756, w37757, w37758, w37759, w37760, w37761, w37762, w37763, w37764, w37765, w37766, w37767, w37768, w37769, w37770, w37771, w37772, w37773, w37774, w37775, w37776, w37777, w37778, w37779, w37780, w37781, w37782, w37783, w37784, w37785, w37786, w37787, w37788, w37789, w37790, w37791, w37792, w37793, w37794, w37795, w37796, w37797, w37798, w37799, w37800, w37801, w37802, w37803, w37804, w37805, w37806, w37807, w37808, w37809, w37810, w37811, w37812, w37813, w37814, w37815, w37816, w37817, w37818, w37819, w37820, w37821, w37822, w37823, w37824, w37825, w37826, w37827, w37828, w37829, w37830, w37831, w37832, w37833, w37834, w37835, w37836, w37837, w37838, w37839, w37840, w37841, w37842, w37843, w37844, w37845, w37846, w37847, w37848, w37849, w37850, w37851, w37852, w37853, w37854, w37855, w37856, w37857, w37858, w37859, w37860, w37861, w37862, w37863, w37864, w37865, w37866, w37867, w37868, w37869, w37870, w37871, w37872, w37873, w37874, w37875, w37876, w37877, w37878, w37879, w37880, w37881, w37882, w37883, w37884, w37885, w37886, w37887, w37888, w37889, w37890, w37891, w37892, w37893, w37894, w37895, w37896, w37897, w37898, w37899, w37900, w37901, w37902, w37903, w37904, w37905, w37906, w37907, w37908, w37909, w37910, w37911, w37912, w37913, w37914, w37915, w37916, w37917, w37918, w37919, w37920, w37921, w37922, w37923, w37924, w37925, w37926, w37927, w37928, w37929, w37930, w37931, w37932, w37933, w37934, w37935, w37936, w37937, w37938, w37939, w37940, w37941, w37942, w37943, w37944, w37945, w37946, w37947, w37948, w37949, w37950, w37951, w37952, w37953, w37954, w37955, w37956, w37957, w37958, w37959, w37960, w37961, w37962, w37963, w37964, w37965, w37966, w37967, w37968, w37969, w37970, w37971, w37972, w37973, w37974, w37975, w37976, w37977, w37978, w37979, w37980, w37981, w37982, w37983, w37984, w37985, w37986, w37987, w37988, w37989, w37990, w37991, w37992, w37993, w37994, w37995, w37996, w37997, w37998, w37999, w38000, w38001, w38002, w38003, w38004, w38005, w38006, w38007, w38008, w38009, w38010, w38011, w38012, w38013, w38014, w38015, w38016, w38017, w38018, w38019, w38020, w38021, w38022, w38023, w38024, w38025, w38026, w38027, w38028, w38029, w38030, w38031, w38032, w38033, w38034, w38035, w38036, w38037, w38038, w38039, w38040, w38041, w38042, w38043, w38044, w38045, w38046, w38047, w38048, w38049, w38050, w38051, w38052, w38053, w38054, w38055, w38056, w38057, w38058, w38059, w38060, w38061, w38062, w38063, w38064, w38065, w38066, w38067, w38068, w38069, w38070, w38071, w38072, w38073, w38074, w38075, w38076, w38077, w38078, w38079, w38080, w38081, w38082, w38083, w38084, w38085, w38086, w38087, w38088, w38089, w38090, w38091, w38092, w38093, w38094, w38095, w38096, w38097, w38098, w38099, w38100, w38101, w38102, w38103, w38104, w38105, w38106, w38107, w38108, w38109, w38110, w38111, w38112, w38113, w38114, w38115, w38116, w38117, w38118, w38119, w38120, w38121, w38122, w38123, w38124, w38125, w38126, w38127, w38128, w38129, w38130, w38131, w38132, w38133, w38134, w38135, w38136, w38137, w38138, w38139, w38140, w38141, w38142, w38143, w38144, w38145, w38146, w38147, w38148, w38149, w38150, w38151, w38152, w38153, w38154, w38155, w38156, w38157, w38158, w38159, w38160, w38161, w38162, w38163, w38164, w38165, w38166, w38167, w38168, w38169, w38170, w38171, w38172, w38173, w38174, w38175, w38176, w38177, w38178, w38179, w38180, w38181, w38182, w38183, w38184, w38185, w38186, w38187, w38188, w38189, w38190, w38191, w38192, w38193, w38194, w38195, w38196, w38197, w38198, w38199, w38200, w38201, w38202, w38203, w38204, w38205, w38206, w38207, w38208, w38209, w38210, w38211, w38212, w38213, w38214, w38215, w38216, w38217, w38218, w38219, w38220, w38221, w38222, w38223, w38224, w38225, w38226, w38227, w38228, w38229, w38230, w38231, w38232, w38233, w38234, w38235, w38236, w38237, w38238, w38239, w38240, w38241, w38242, w38243, w38244, w38245, w38246, w38247, w38248, w38249, w38250, w38251, w38252, w38253, w38254, w38255, w38256, w38257, w38258, w38259, w38260, w38261, w38262, w38263, w38264, w38265, w38266, w38267, w38268, w38269, w38270, w38271, w38272, w38273, w38274, w38275, w38276, w38277, w38278, w38279, w38280, w38281, w38282, w38283, w38284, w38285, w38286, w38287, w38288, w38289, w38290, w38291, w38292, w38293, w38294, w38295, w38296, w38297, w38298, w38299, w38300, w38301, w38302, w38303, w38304, w38305, w38306, w38307, w38308, w38309, w38310, w38311, w38312, w38313, w38314, w38315, w38316, w38317, w38318, w38319, w38320, w38321, w38322, w38323, w38324, w38325, w38326, w38327, w38328, w38329, w38330, w38331, w38332, w38333, w38334, w38335, w38336, w38337, w38338, w38339, w38340, w38341, w38342, w38343, w38344, w38345, w38346, w38347, w38348, w38349, w38350, w38351, w38352, w38353, w38354, w38355, w38356, w38357, w38358, w38359, w38360, w38361, w38362, w38363, w38364, w38365, w38366, w38367, w38368, w38369, w38370, w38371, w38372, w38373, w38374, w38375, w38376, w38377, w38378, w38379, w38380, w38381, w38382, w38383, w38384, w38385, w38386, w38387, w38388, w38389, w38390, w38391, w38392, w38393, w38394, w38395, w38396, w38397, w38398, w38399, w38400, w38401, w38402, w38403, w38404, w38405, w38406, w38407, w38408, w38409, w38410, w38411, w38412, w38413, w38414, w38415, w38416, w38417, w38418, w38419, w38420, w38421, w38422, w38423, w38424, w38425, w38426, w38427, w38428, w38429, w38430, w38431, w38432, w38433, w38434, w38435, w38436, w38437, w38438, w38439, w38440, w38441, w38442, w38443, w38444, w38445, w38446, w38447, w38448, w38449, w38450, w38451, w38452, w38453, w38454, w38455, w38456, w38457, w38458, w38459, w38460, w38461, w38462, w38463, w38464, w38465, w38466, w38467, w38468, w38469, w38470, w38471, w38472, w38473, w38474, w38475, w38476, w38477, w38478, w38479, w38480, w38481, w38482, w38483, w38484, w38485, w38486, w38487, w38488, w38489, w38490, w38491, w38492, w38493, w38494, w38495, w38496, w38497, w38498, w38499, w38500, w38501, w38502, w38503, w38504, w38505, w38506, w38507, w38508, w38509, w38510, w38511, w38512, w38513, w38514, w38515, w38516, w38517, w38518, w38519, w38520, w38521, w38522, w38523, w38524, w38525, w38526, w38527, w38528, w38529, w38530, w38531, w38532, w38533, w38534, w38535, w38536, w38537, w38538, w38539, w38540, w38541, w38542, w38543, w38544, w38545, w38546, w38547, w38548, w38549, w38550, w38551, w38552, w38553, w38554, w38555, w38556, w38557, w38558, w38559, w38560, w38561, w38562, w38563, w38564, w38565, w38566, w38567, w38568, w38569, w38570, w38571, w38572, w38573, w38574, w38575, w38576, w38577, w38578, w38579, w38580, w38581, w38582, w38583, w38584, w38585, w38586, w38587, w38588, w38589, w38590, w38591, w38592, w38593, w38594, w38595, w38596, w38597, w38598, w38599, w38600, w38601, w38602, w38603, w38604, w38605, w38606, w38607, w38608, w38609, w38610, w38611, w38612, w38613, w38614, w38615, w38616, w38617, w38618, w38619, w38620, w38621, w38622, w38623, w38624, w38625, w38626, w38627, w38628, w38629, w38630, w38631, w38632, w38633, w38634, w38635, w38636, w38637, w38638, w38639, w38640, w38641, w38642, w38643, w38644, w38645, w38646, w38647, w38648, w38649, w38650, w38651, w38652, w38653, w38654, w38655, w38656, w38657, w38658, w38659, w38660, w38661, w38662, w38663, w38664, w38665, w38666, w38667, w38668, w38669, w38670, w38671, w38672, w38673, w38674, w38675, w38676, w38677, w38678, w38679, w38680, w38681, w38682, w38683, w38684, w38685, w38686, w38687, w38688, w38689, w38690, w38691, w38692, w38693, w38694, w38695, w38696, w38697, w38698, w38699, w38700, w38701, w38702, w38703, w38704, w38705, w38706, w38707, w38708, w38709, w38710, w38711, w38712, w38713, w38714, w38715, w38716, w38717, w38718, w38719, w38720, w38721, w38722, w38723, w38724, w38725, w38726, w38727, w38728, w38729, w38730, w38731, w38732, w38733, w38734, w38735, w38736, w38737, w38738, w38739, w38740, w38741, w38742, w38743, w38744, w38745, w38746, w38747, w38748, w38749, w38750, w38751, w38752, w38753, w38754, w38755, w38756, w38757, w38758, w38759, w38760, w38761, w38762, w38763, w38764, w38765, w38766, w38767, w38768, w38769, w38770, w38771, w38772, w38773, w38774, w38775, w38776, w38777, w38778, w38779, w38780, w38781, w38782, w38783, w38784, w38785, w38786, w38787, w38788, w38789, w38790, w38791, w38792, w38793, w38794, w38795, w38796, w38797, w38798, w38799, w38800, w38801, w38802, w38803, w38804, w38805, w38806, w38807, w38808, w38809, w38810, w38811, w38812, w38813, w38814, w38815, w38816, w38817, w38818, w38819, w38820, w38821, w38822, w38823, w38824, w38825, w38826, w38827, w38828, w38829, w38830, w38831, w38832, w38833, w38834, w38835, w38836, w38837, w38838, w38839, w38840, w38841, w38842, w38843, w38844, w38845, w38846, w38847, w38848, w38849, w38850, w38851, w38852, w38853, w38854, w38855, w38856, w38857, w38858, w38859, w38860, w38861, w38862, w38863, w38864, w38865, w38866, w38867, w38868, w38869, w38870, w38871, w38872, w38873, w38874, w38875, w38876, w38877, w38878, w38879, w38880, w38881, w38882, w38883, w38884, w38885, w38886, w38887, w38888, w38889, w38890, w38891, w38892, w38893, w38894, w38895, w38896, w38897, w38898, w38899, w38900, w38901, w38902, w38903, w38904, w38905, w38906, w38907, w38908, w38909, w38910, w38911, w38912, w38913, w38914, w38915, w38916, w38917, w38918, w38919, w38920, w38921, w38922, w38923, w38924, w38925, w38926, w38927, w38928, w38929, w38930, w38931, w38932, w38933, w38934, w38935, w38936, w38937, w38938, w38939, w38940, w38941, w38942, w38943, w38944, w38945, w38946, w38947, w38948, w38949, w38950, w38951, w38952, w38953, w38954, w38955, w38956, w38957, w38958, w38959, w38960, w38961, w38962, w38963, w38964, w38965, w38966, w38967, w38968, w38969, w38970, w38971, w38972, w38973, w38974, w38975, w38976, w38977, w38978, w38979, w38980, w38981, w38982, w38983, w38984, w38985, w38986, w38987, w38988, w38989, w38990, w38991, w38992, w38993, w38994, w38995, w38996, w38997, w38998, w38999, w39000, w39001, w39002, w39003, w39004, w39005, w39006, w39007, w39008, w39009, w39010, w39011, w39012, w39013, w39014, w39015, w39016, w39017, w39018, w39019, w39020, w39021, w39022, w39023, w39024, w39025, w39026, w39027, w39028, w39029, w39030, w39031, w39032, w39033, w39034, w39035, w39036, w39037, w39038, w39039, w39040, w39041, w39042, w39043, w39044, w39045, w39046, w39047, w39048, w39049, w39050, w39051, w39052, w39053, w39054, w39055, w39056, w39057, w39058, w39059, w39060, w39061, w39062, w39063, w39064, w39065, w39066, w39067, w39068, w39069, w39070, w39071, w39072, w39073, w39074, w39075, w39076, w39077, w39078, w39079, w39080, w39081, w39082, w39083, w39084, w39085, w39086, w39087, w39088, w39089, w39090, w39091, w39092, w39093, w39094, w39095, w39096, w39097, w39098, w39099, w39100, w39101, w39102, w39103, w39104, w39105, w39106, w39107, w39108, w39109, w39110, w39111, w39112, w39113, w39114, w39115, w39116, w39117, w39118, w39119, w39120, w39121, w39122, w39123, w39124, w39125, w39126, w39127, w39128, w39129, w39130, w39131, w39132, w39133, w39134, w39135, w39136, w39137, w39138, w39139, w39140, w39141, w39142, w39143, w39144, w39145, w39146, w39147, w39148, w39149, w39150, w39151, w39152, w39153, w39154, w39155, w39156, w39157, w39158, w39159, w39160, w39161, w39162, w39163, w39164, w39165, w39166, w39167, w39168, w39169, w39170, w39171, w39172, w39173, w39174, w39175, w39176, w39177, w39178, w39179, w39180, w39181, w39182, w39183, w39184, w39185, w39186, w39187, w39188, w39189, w39190, w39191, w39192, w39193, w39194, w39195, w39196, w39197, w39198, w39199, w39200, w39201, w39202, w39203, w39204, w39205, w39206, w39207, w39208, w39209, w39210, w39211, w39212, w39213, w39214, w39215, w39216, w39217, w39218, w39219, w39220, w39221, w39222, w39223, w39224, w39225, w39226, w39227, w39228, w39229, w39230, w39231, w39232, w39233, w39234, w39235, w39236, w39237, w39238, w39239, w39240, w39241, w39242, w39243, w39244, w39245, w39246, w39247, w39248, w39249, w39250, w39251, w39252, w39253, w39254, w39255, w39256, w39257, w39258, w39259, w39260, w39261, w39262, w39263, w39264, w39265, w39266, w39267, w39268, w39269, w39270, w39271, w39272, w39273, w39274, w39275, w39276, w39277, w39278, w39279, w39280, w39281, w39282, w39283, w39284, w39285, w39286, w39287, w39288, w39289, w39290, w39291, w39292, w39293, w39294, w39295, w39296, w39297, w39298, w39299, w39300, w39301, w39302, w39303, w39304, w39305, w39306, w39307, w39308, w39309, w39310, w39311, w39312, w39313, w39314, w39315, w39316, w39317, w39318, w39319, w39320, w39321, w39322, w39323, w39324, w39325, w39326, w39327, w39328, w39329, w39330, w39331, w39332, w39333, w39334, w39335, w39336, w39337, w39338, w39339, w39340, w39341, w39342, w39343, w39344, w39345, w39346, w39347, w39348, w39349, w39350, w39351, w39352, w39353, w39354, w39355, w39356, w39357, w39358, w39359, w39360, w39361, w39362, w39363, w39364, w39365, w39366, w39367, w39368, w39369, w39370, w39371, w39372, w39373, w39374, w39375, w39376, w39377, w39378, w39379, w39380, w39381, w39382, w39383, w39384, w39385, w39386, w39387, w39388, w39389, w39390, w39391, w39392, w39393, w39394, w39395, w39396, w39397, w39398, w39399, w39400, w39401, w39402, w39403, w39404, w39405, w39406, w39407, w39408, w39409, w39410, w39411, w39412, w39413, w39414, w39415, w39416, w39417, w39418, w39419, w39420, w39421, w39422, w39423, w39424, w39425, w39426, w39427, w39428, w39429, w39430, w39431, w39432, w39433, w39434, w39435, w39436, w39437, w39438, w39439, w39440, w39441, w39442, w39443, w39444, w39445, w39446, w39447, w39448, w39449, w39450, w39451, w39452, w39453, w39454, w39455, w39456, w39457, w39458, w39459, w39460, w39461, w39462, w39463, w39464, w39465, w39466, w39467, w39468, w39469, w39470, w39471, w39472, w39473, w39474, w39475, w39476, w39477, w39478, w39479, w39480, w39481, w39482, w39483, w39484, w39485, w39486, w39487, w39488, w39489, w39490, w39491, w39492, w39493, w39494, w39495, w39496, w39497, w39498, w39499, w39500, w39501, w39502, w39503, w39504, w39505, w39506, w39507, w39508, w39509, w39510, w39511, w39512, w39513, w39514, w39515, w39516, w39517, w39518, w39519, w39520, w39521, w39522, w39523, w39524, w39525, w39526, w39527, w39528, w39529, w39530, w39531, w39532, w39533, w39534, w39535, w39536, w39537, w39538, w39539, w39540, w39541, w39542, w39543, w39544, w39545, w39546, w39547, w39548, w39549, w39550, w39551, w39552, w39553, w39554, w39555, w39556, w39557, w39558, w39559, w39560, w39561, w39562, w39563, w39564, w39565, w39566, w39567, w39568, w39569, w39570, w39571, w39572, w39573, w39574, w39575, w39576, w39577, w39578, w39579, w39580, w39581, w39582, w39583, w39584, w39585, w39586, w39587, w39588, w39589, w39590, w39591, w39592, w39593, w39594, w39595, w39596, w39597, w39598, w39599, w39600, w39601, w39602, w39603, w39604, w39605, w39606, w39607, w39608, w39609, w39610, w39611, w39612, w39613, w39614, w39615, w39616, w39617, w39618, w39619, w39620, w39621, w39622, w39623, w39624, w39625, w39626, w39627, w39628, w39629, w39630, w39631, w39632, w39633, w39634, w39635, w39636, w39637, w39638, w39639, w39640, w39641, w39642, w39643, w39644, w39645, w39646, w39647, w39648, w39649, w39650, w39651, w39652, w39653, w39654, w39655, w39656, w39657, w39658, w39659, w39660, w39661, w39662, w39663, w39664, w39665, w39666, w39667, w39668, w39669, w39670, w39671, w39672, w39673, w39674, w39675, w39676, w39677, w39678, w39679, w39680, w39681, w39682, w39683, w39684, w39685, w39686, w39687, w39688, w39689, w39690, w39691, w39692, w39693, w39694, w39695, w39696, w39697, w39698, w39699, w39700, w39701, w39702, w39703, w39704, w39705, w39706, w39707, w39708, w39709, w39710, w39711, w39712, w39713, w39714, w39715, w39716, w39717, w39718, w39719, w39720, w39721, w39722, w39723, w39724, w39725, w39726, w39727, w39728, w39729, w39730, w39731, w39732, w39733, w39734, w39735, w39736, w39737, w39738, w39739, w39740, w39741, w39742, w39743, w39744, w39745, w39746, w39747, w39748, w39749, w39750, w39751, w39752, w39753, w39754, w39755, w39756, w39757, w39758, w39759, w39760, w39761, w39762, w39763, w39764, w39765, w39766, w39767, w39768, w39769, w39770, w39771, w39772, w39773, w39774, w39775, w39776, w39777, w39778, w39779, w39780, w39781, w39782, w39783, w39784, w39785, w39786, w39787, w39788, w39789, w39790, w39791, w39792, w39793, w39794, w39795, w39796, w39797, w39798, w39799, w39800, w39801, w39802, w39803, w39804, w39805, w39806, w39807, w39808, w39809, w39810, w39811, w39812, w39813, w39814, w39815, w39816, w39817, w39818, w39819, w39820, w39821, w39822, w39823, w39824, w39825, w39826, w39827, w39828, w39829, w39830, w39831, w39832, w39833, w39834, w39835, w39836, w39837, w39838, w39839, w39840, w39841, w39842, w39843, w39844, w39845, w39846, w39847, w39848, w39849, w39850, w39851, w39852, w39853, w39854, w39855, w39856, w39857, w39858, w39859, w39860, w39861, w39862, w39863, w39864, w39865, w39866, w39867, w39868, w39869, w39870, w39871, w39872, w39873, w39874, w39875, w39876, w39877, w39878, w39879, w39880, w39881, w39882, w39883, w39884, w39885, w39886, w39887, w39888, w39889, w39890, w39891, w39892, w39893, w39894, w39895, w39896, w39897, w39898, w39899, w39900, w39901, w39902, w39903, w39904, w39905, w39906, w39907, w39908, w39909, w39910, w39911, w39912, w39913, w39914, w39915, w39916, w39917, w39918, w39919, w39920, w39921, w39922, w39923, w39924, w39925, w39926, w39927, w39928, w39929, w39930, w39931, w39932, w39933, w39934, w39935, w39936, w39937, w39938, w39939, w39940, w39941, w39942, w39943, w39944, w39945, w39946, w39947, w39948, w39949, w39950, w39951, w39952, w39953, w39954, w39955, w39956, w39957, w39958, w39959, w39960, w39961, w39962, w39963, w39964, w39965, w39966, w39967, w39968, w39969, w39970, w39971, w39972, w39973, w39974, w39975, w39976, w39977, w39978, w39979, w39980, w39981, w39982, w39983, w39984, w39985, w39986, w39987, w39988, w39989, w39990, w39991, w39992, w39993, w39994, w39995, w39996, w39997, w39998, w39999, w40000, w40001, w40002, w40003, w40004, w40005, w40006, w40007, w40008, w40009, w40010, w40011, w40012, w40013, w40014, w40015, w40016, w40017, w40018, w40019, w40020, w40021, w40022, w40023, w40024, w40025, w40026, w40027, w40028, w40029, w40030, w40031, w40032, w40033, w40034, w40035, w40036, w40037, w40038, w40039, w40040, w40041, w40042, w40043, w40044, w40045, w40046, w40047, w40048, w40049, w40050, w40051, w40052, w40053, w40054, w40055, w40056, w40057, w40058, w40059, w40060, w40061, w40062, w40063, w40064, w40065, w40066, w40067, w40068, w40069, w40070, w40071, w40072, w40073, w40074, w40075, w40076, w40077, w40078, w40079, w40080, w40081, w40082, w40083, w40084, w40085, w40086, w40087, w40088, w40089, w40090, w40091, w40092, w40093, w40094, w40095, w40096, w40097, w40098, w40099, w40100, w40101, w40102, w40103, w40104, w40105, w40106, w40107, w40108, w40109, w40110, w40111, w40112, w40113, w40114, w40115, w40116, w40117, w40118, w40119, w40120, w40121, w40122, w40123, w40124, w40125, w40126, w40127, w40128, w40129, w40130, w40131, w40132, w40133, w40134, w40135, w40136, w40137, w40138, w40139, w40140, w40141, w40142, w40143, w40144, w40145, w40146, w40147, w40148, w40149, w40150, w40151, w40152, w40153, w40154, w40155, w40156, w40157, w40158, w40159, w40160, w40161, w40162, w40163, w40164, w40165, w40166, w40167, w40168, w40169, w40170, w40171, w40172, w40173, w40174, w40175, w40176, w40177, w40178, w40179, w40180, w40181, w40182, w40183, w40184, w40185, w40186, w40187, w40188, w40189, w40190, w40191, w40192, w40193, w40194, w40195, w40196, w40197, w40198, w40199, w40200, w40201, w40202, w40203, w40204, w40205, w40206, w40207, w40208, w40209, w40210, w40211, w40212, w40213, w40214, w40215, w40216, w40217, w40218, w40219, w40220, w40221, w40222, w40223, w40224, w40225, w40226, w40227, w40228, w40229, w40230, w40231, w40232, w40233, w40234, w40235, w40236, w40237, w40238, w40239, w40240, w40241, w40242, w40243, w40244, w40245, w40246, w40247, w40248, w40249, w40250, w40251, w40252, w40253, w40254, w40255, w40256, w40257, w40258, w40259, w40260, w40261, w40262, w40263, w40264, w40265, w40266, w40267, w40268, w40269, w40270, w40271, w40272, w40273, w40274, w40275, w40276, w40277, w40278, w40279, w40280, w40281, w40282, w40283, w40284, w40285, w40286, w40287, w40288, w40289, w40290, w40291, w40292, w40293, w40294, w40295, w40296, w40297, w40298, w40299, w40300, w40301, w40302, w40303, w40304, w40305, w40306, w40307, w40308, w40309, w40310, w40311, w40312, w40313, w40314, w40315, w40316, w40317, w40318, w40319, w40320, w40321, w40322, w40323, w40324, w40325, w40326, w40327, w40328, w40329, w40330, w40331, w40332, w40333, w40334, w40335, w40336, w40337, w40338, w40339, w40340, w40341, w40342, w40343, w40344, w40345, w40346, w40347, w40348, w40349, w40350, w40351, w40352, w40353, w40354, w40355, w40356, w40357, w40358, w40359, w40360, w40361, w40362, w40363, w40364, w40365, w40366, w40367, w40368, w40369, w40370, w40371, w40372, w40373, w40374, w40375, w40376, w40377, w40378, w40379, w40380, w40381, w40382, w40383, w40384, w40385, w40386, w40387, w40388, w40389, w40390, w40391, w40392, w40393, w40394, w40395, w40396, w40397, w40398, w40399, w40400, w40401, w40402, w40403, w40404, w40405, w40406, w40407, w40408, w40409, w40410, w40411, w40412, w40413, w40414, w40415, w40416, w40417, w40418, w40419, w40420, w40421, w40422, w40423, w40424, w40425, w40426, w40427, w40428, w40429, w40430, w40431, w40432, w40433, w40434, w40435, w40436, w40437, w40438, w40439, w40440, w40441, w40442, w40443, w40444, w40445, w40446, w40447, w40448, w40449, w40450, w40451, w40452, w40453, w40454, w40455, w40456, w40457, w40458, w40459, w40460, w40461, w40462, w40463, w40464, w40465, w40466, w40467, w40468, w40469, w40470, w40471, w40472, w40473, w40474, w40475, w40476, w40477, w40478, w40479, w40480, w40481, w40482, w40483, w40484, w40485, w40486, w40487, w40488, w40489, w40490, w40491, w40492, w40493, w40494, w40495, w40496, w40497, w40498, w40499, w40500, w40501, w40502, w40503, w40504, w40505, w40506, w40507, w40508, w40509, w40510, w40511, w40512, w40513, w40514, w40515, w40516, w40517, w40518, w40519, w40520, w40521, w40522, w40523, w40524, w40525, w40526, w40527, w40528, w40529, w40530, w40531, w40532, w40533, w40534, w40535, w40536, w40537, w40538, w40539, w40540, w40541, w40542, w40543, w40544, w40545, w40546, w40547, w40548, w40549, w40550, w40551, w40552, w40553, w40554, w40555, w40556, w40557, w40558, w40559, w40560, w40561, w40562, w40563, w40564, w40565, w40566, w40567, w40568, w40569, w40570, w40571, w40572, w40573, w40574, w40575, w40576, w40577, w40578, w40579, w40580, w40581, w40582, w40583, w40584, w40585, w40586, w40587, w40588, w40589, w40590, w40591, w40592, w40593, w40594, w40595, w40596, w40597, w40598, w40599, w40600, w40601, w40602, w40603, w40604, w40605, w40606, w40607, w40608, w40609, w40610, w40611, w40612, w40613, w40614, w40615, w40616, w40617, w40618, w40619, w40620, w40621, w40622, w40623, w40624, w40625, w40626, w40627, w40628, w40629, w40630, w40631, w40632, w40633, w40634, w40635, w40636, w40637, w40638, w40639, w40640, w40641, w40642, w40643, w40644, w40645, w40646, w40647, w40648, w40649, w40650, w40651, w40652, w40653, w40654, w40655, w40656, w40657, w40658, w40659, w40660, w40661, w40662, w40663, w40664, w40665, w40666, w40667, w40668, w40669, w40670, w40671, w40672, w40673, w40674, w40675, w40676, w40677, w40678, w40679, w40680, w40681, w40682, w40683, w40684, w40685, w40686, w40687, w40688, w40689, w40690, w40691, w40692, w40693, w40694, w40695, w40696, w40697, w40698, w40699, w40700, w40701, w40702, w40703, w40704, w40705, w40706, w40707, w40708, w40709, w40710, w40711, w40712, w40713, w40714, w40715, w40716, w40717, w40718, w40719, w40720, w40721, w40722, w40723, w40724, w40725, w40726, w40727, w40728, w40729, w40730, w40731, w40732, w40733, w40734, w40735, w40736, w40737, w40738, w40739, w40740, w40741, w40742, w40743, w40744, w40745, w40746, w40747, w40748, w40749, w40750, w40751, w40752, w40753, w40754, w40755, w40756, w40757, w40758, w40759, w40760, w40761, w40762, w40763, w40764, w40765, w40766, w40767, w40768, w40769, w40770, w40771, w40772, w40773, w40774, w40775, w40776, w40777, w40778, w40779, w40780, w40781, w40782, w40783, w40784, w40785, w40786, w40787, w40788, w40789, w40790, w40791, w40792, w40793, w40794, w40795, w40796, w40797, w40798, w40799, w40800, w40801, w40802, w40803, w40804, w40805, w40806, w40807, w40808, w40809, w40810, w40811, w40812, w40813, w40814, w40815, w40816, w40817, w40818, w40819, w40820, w40821, w40822, w40823, w40824, w40825, w40826, w40827, w40828, w40829, w40830, w40831, w40832, w40833, w40834, w40835, w40836, w40837, w40838, w40839, w40840, w40841, w40842, w40843, w40844, w40845, w40846, w40847, w40848, w40849, w40850, w40851, w40852, w40853, w40854, w40855, w40856, w40857, w40858, w40859, w40860, w40861, w40862, w40863, w40864, w40865, w40866, w40867, w40868, w40869, w40870, w40871, w40872, w40873, w40874, w40875, w40876, w40877, w40878, w40879, w40880, w40881, w40882, w40883, w40884, w40885, w40886, w40887, w40888, w40889, w40890, w40891, w40892, w40893, w40894, w40895, w40896, w40897, w40898, w40899, w40900, w40901, w40902, w40903, w40904, w40905, w40906, w40907, w40908, w40909, w40910, w40911, w40912, w40913, w40914, w40915, w40916, w40917, w40918, w40919, w40920, w40921, w40922, w40923, w40924, w40925, w40926, w40927, w40928, w40929, w40930, w40931, w40932, w40933, w40934, w40935, w40936, w40937, w40938, w40939, w40940, w40941, w40942, w40943, w40944, w40945, w40946, w40947, w40948, w40949, w40950, w40951, w40952, w40953, w40954, w40955, w40956, w40957, w40958, w40959, w40960, w40961, w40962, w40963, w40964, w40965, w40966, w40967, w40968, w40969, w40970, w40971, w40972, w40973, w40974, w40975, w40976, w40977, w40978, w40979, w40980, w40981, w40982, w40983, w40984, w40985, w40986, w40987, w40988, w40989, w40990, w40991, w40992, w40993, w40994, w40995, w40996, w40997, w40998, w40999, w41000, w41001, w41002, w41003, w41004, w41005, w41006, w41007, w41008, w41009, w41010, w41011, w41012, w41013, w41014, w41015, w41016, w41017, w41018, w41019, w41020, w41021, w41022, w41023, w41024, w41025, w41026, w41027, w41028, w41029, w41030, w41031, w41032, w41033, w41034, w41035, w41036, w41037, w41038, w41039, w41040, w41041, w41042, w41043, w41044, w41045, w41046, w41047, w41048, w41049, w41050, w41051, w41052, w41053, w41054, w41055, w41056, w41057, w41058, w41059, w41060, w41061, w41062, w41063, w41064, w41065, w41066, w41067, w41068, w41069, w41070, w41071, w41072, w41073, w41074, w41075, w41076, w41077, w41078, w41079, w41080, w41081, w41082, w41083, w41084, w41085, w41086, w41087, w41088, w41089, w41090, w41091, w41092, w41093, w41094, w41095, w41096, w41097, w41098, w41099, w41100, w41101, w41102, w41103, w41104, w41105, w41106, w41107, w41108, w41109, w41110, w41111, w41112, w41113, w41114, w41115, w41116, w41117, w41118, w41119, w41120, w41121, w41122, w41123, w41124, w41125, w41126, w41127, w41128, w41129, w41130, w41131, w41132, w41133, w41134, w41135, w41136, w41137, w41138, w41139, w41140, w41141, w41142, w41143, w41144, w41145, w41146, w41147, w41148, w41149, w41150, w41151, w41152, w41153, w41154, w41155, w41156, w41157, w41158, w41159, w41160, w41161, w41162, w41163, w41164, w41165, w41166, w41167, w41168, w41169, w41170, w41171, w41172, w41173, w41174, w41175, w41176, w41177, w41178, w41179, w41180, w41181, w41182, w41183, w41184, w41185, w41186, w41187, w41188, w41189, w41190, w41191, w41192, w41193, w41194, w41195, w41196, w41197, w41198, w41199, w41200, w41201, w41202, w41203, w41204, w41205, w41206, w41207, w41208, w41209, w41210, w41211, w41212, w41213, w41214, w41215, w41216, w41217, w41218, w41219, w41220, w41221, w41222, w41223, w41224, w41225, w41226, w41227, w41228, w41229, w41230, w41231, w41232, w41233, w41234, w41235, w41236, w41237, w41238, w41239, w41240, w41241, w41242, w41243, w41244, w41245, w41246, w41247, w41248, w41249, w41250, w41251, w41252, w41253, w41254, w41255, w41256, w41257, w41258, w41259, w41260, w41261, w41262, w41263, w41264, w41265, w41266, w41267, w41268, w41269, w41270, w41271, w41272, w41273, w41274, w41275, w41276, w41277, w41278, w41279, w41280, w41281, w41282, w41283, w41284, w41285, w41286, w41287, w41288, w41289, w41290, w41291, w41292, w41293, w41294, w41295, w41296, w41297, w41298, w41299, w41300, w41301, w41302, w41303, w41304, w41305, w41306, w41307, w41308, w41309, w41310, w41311, w41312, w41313, w41314, w41315, w41316, w41317, w41318, w41319, w41320, w41321, w41322, w41323, w41324, w41325, w41326, w41327, w41328, w41329, w41330, w41331, w41332, w41333, w41334, w41335, w41336, w41337, w41338, w41339, w41340, w41341, w41342, w41343, w41344, w41345, w41346, w41347, w41348, w41349, w41350, w41351, w41352, w41353, w41354, w41355, w41356, w41357, w41358, w41359, w41360, w41361, w41362, w41363, w41364, w41365, w41366, w41367, w41368, w41369, w41370, w41371, w41372, w41373, w41374, w41375, w41376, w41377, w41378, w41379, w41380, w41381, w41382, w41383, w41384, w41385, w41386, w41387, w41388, w41389, w41390, w41391, w41392, w41393, w41394, w41395, w41396, w41397, w41398, w41399, w41400, w41401, w41402, w41403, w41404, w41405, w41406, w41407, w41408, w41409, w41410, w41411, w41412, w41413, w41414, w41415, w41416, w41417, w41418, w41419, w41420, w41421, w41422, w41423, w41424, w41425, w41426, w41427, w41428, w41429, w41430, w41431, w41432, w41433, w41434, w41435, w41436, w41437, w41438, w41439, w41440, w41441, w41442, w41443, w41444, w41445, w41446, w41447, w41448, w41449, w41450, w41451, w41452, w41453, w41454, w41455, w41456, w41457, w41458, w41459, w41460, w41461, w41462, w41463, w41464, w41465, w41466, w41467, w41468, w41469, w41470, w41471, w41472, w41473, w41474, w41475, w41476, w41477, w41478, w41479, w41480, w41481, w41482, w41483, w41484, w41485, w41486, w41487, w41488, w41489, w41490, w41491, w41492, w41493, w41494, w41495, w41496, w41497, w41498, w41499, w41500, w41501, w41502, w41503, w41504, w41505, w41506, w41507, w41508, w41509, w41510, w41511, w41512, w41513, w41514, w41515, w41516, w41517, w41518, w41519, w41520, w41521, w41522, w41523, w41524, w41525, w41526, w41527, w41528, w41529, w41530, w41531, w41532, w41533, w41534, w41535, w41536, w41537, w41538, w41539, w41540, w41541, w41542, w41543, w41544, w41545, w41546, w41547, w41548, w41549, w41550, w41551, w41552, w41553, w41554, w41555, w41556, w41557, w41558, w41559, w41560, w41561, w41562, w41563, w41564, w41565, w41566, w41567, w41568, w41569, w41570, w41571, w41572, w41573, w41574, w41575, w41576, w41577, w41578, w41579, w41580, w41581, w41582, w41583, w41584, w41585, w41586, w41587, w41588, w41589, w41590, w41591, w41592, w41593, w41594, w41595, w41596, w41597, w41598, w41599, w41600, w41601, w41602, w41603, w41604, w41605, w41606, w41607, w41608, w41609, w41610, w41611, w41612, w41613, w41614, w41615, w41616, w41617, w41618, w41619, w41620, w41621, w41622, w41623, w41624, w41625, w41626, w41627, w41628, w41629, w41630, w41631, w41632, w41633, w41634, w41635, w41636, w41637, w41638, w41639, w41640, w41641, w41642, w41643, w41644, w41645, w41646, w41647, w41648, w41649, w41650, w41651, w41652, w41653, w41654, w41655, w41656, w41657, w41658, w41659, w41660, w41661, w41662, w41663, w41664, w41665, w41666, w41667, w41668, w41669, w41670, w41671, w41672, w41673, w41674, w41675, w41676, w41677, w41678, w41679, w41680, w41681, w41682, w41683, w41684, w41685, w41686, w41687, w41688, w41689, w41690, w41691, w41692, w41693, w41694, w41695, w41696, w41697, w41698, w41699, w41700, w41701, w41702, w41703, w41704, w41705, w41706, w41707, w41708, w41709, w41710, w41711, w41712, w41713, w41714, w41715, w41716, w41717, w41718, w41719, w41720, w41721, w41722, w41723, w41724, w41725, w41726, w41727, w41728, w41729, w41730, w41731, w41732, w41733, w41734, w41735, w41736, w41737, w41738, w41739, w41740, w41741, w41742, w41743, w41744, w41745, w41746, w41747, w41748, w41749, w41750, w41751, w41752, w41753, w41754, w41755, w41756, w41757, w41758, w41759, w41760, w41761, w41762, w41763, w41764, w41765, w41766, w41767, w41768, w41769, w41770, w41771, w41772, w41773, w41774, w41775, w41776, w41777, w41778, w41779, w41780, w41781, w41782, w41783, w41784, w41785, w41786, w41787, w41788, w41789, w41790, w41791, w41792, w41793, w41794, w41795, w41796, w41797, w41798, w41799, w41800, w41801, w41802, w41803, w41804, w41805, w41806, w41807, w41808, w41809, w41810, w41811, w41812, w41813, w41814, w41815, w41816, w41817, w41818, w41819, w41820, w41821, w41822, w41823, w41824, w41825, w41826, w41827, w41828, w41829, w41830, w41831, w41832, w41833, w41834, w41835, w41836, w41837, w41838, w41839, w41840, w41841, w41842, w41843, w41844, w41845, w41846, w41847, w41848, w41849, w41850, w41851, w41852, w41853, w41854, w41855, w41856, w41857, w41858, w41859, w41860, w41861, w41862, w41863, w41864, w41865, w41866, w41867, w41868, w41869, w41870, w41871, w41872, w41873, w41874, w41875, w41876, w41877, w41878, w41879, w41880, w41881, w41882, w41883, w41884, w41885, w41886, w41887, w41888, w41889, w41890, w41891, w41892, w41893, w41894, w41895, w41896, w41897, w41898, w41899, w41900, w41901, w41902, w41903, w41904, w41905, w41906, w41907, w41908, w41909, w41910, w41911, w41912, w41913, w41914, w41915, w41916, w41917, w41918, w41919, w41920, w41921, w41922, w41923, w41924, w41925, w41926, w41927, w41928, w41929, w41930, w41931, w41932, w41933, w41934, w41935, w41936, w41937, w41938, w41939, w41940, w41941, w41942, w41943, w41944, w41945, w41946, w41947, w41948, w41949, w41950, w41951, w41952, w41953, w41954, w41955, w41956, w41957, w41958, w41959, w41960, w41961, w41962, w41963, w41964, w41965, w41966, w41967, w41968, w41969, w41970, w41971, w41972, w41973, w41974, w41975, w41976, w41977, w41978, w41979, w41980, w41981, w41982, w41983, w41984, w41985, w41986, w41987, w41988, w41989, w41990, w41991, w41992, w41993, w41994, w41995, w41996, w41997, w41998, w41999, w42000, w42001, w42002, w42003, w42004, w42005, w42006, w42007, w42008, w42009, w42010, w42011, w42012, w42013, w42014, w42015, w42016, w42017, w42018, w42019, w42020, w42021, w42022, w42023, w42024, w42025, w42026, w42027, w42028, w42029, w42030, w42031, w42032, w42033, w42034, w42035, w42036, w42037, w42038, w42039, w42040, w42041, w42042, w42043, w42044, w42045, w42046, w42047, w42048, w42049, w42050, w42051, w42052, w42053, w42054, w42055, w42056, w42057, w42058, w42059, w42060, w42061, w42062, w42063, w42064, w42065, w42066, w42067, w42068, w42069, w42070, w42071, w42072, w42073, w42074, w42075, w42076, w42077, w42078, w42079, w42080, w42081, w42082, w42083, w42084, w42085, w42086, w42087, w42088, w42089, w42090, w42091, w42092, w42093, w42094, w42095, w42096, w42097, w42098, w42099, w42100, w42101, w42102, w42103, w42104, w42105, w42106, w42107, w42108, w42109, w42110, w42111, w42112, w42113, w42114, w42115, w42116, w42117, w42118, w42119, w42120, w42121, w42122, w42123, w42124, w42125, w42126, w42127, w42128, w42129, w42130, w42131, w42132, w42133, w42134, w42135, w42136, w42137, w42138, w42139, w42140, w42141, w42142, w42143, w42144, w42145, w42146, w42147, w42148, w42149, w42150, w42151, w42152, w42153, w42154, w42155, w42156, w42157, w42158, w42159, w42160, w42161, w42162, w42163, w42164, w42165, w42166, w42167, w42168, w42169, w42170, w42171, w42172, w42173, w42174, w42175, w42176, w42177, w42178, w42179, w42180, w42181, w42182, w42183, w42184, w42185, w42186, w42187, w42188, w42189, w42190, w42191, w42192, w42193, w42194, w42195, w42196, w42197, w42198, w42199, w42200, w42201, w42202, w42203, w42204, w42205, w42206, w42207, w42208, w42209, w42210, w42211, w42212, w42213, w42214, w42215, w42216, w42217, w42218, w42219, w42220, w42221, w42222, w42223, w42224, w42225, w42226, w42227, w42228, w42229, w42230, w42231, w42232, w42233, w42234, w42235, w42236, w42237, w42238, w42239, w42240, w42241, w42242, w42243, w42244, w42245, w42246, w42247, w42248, w42249, w42250, w42251, w42252, w42253, w42254, w42255, w42256, w42257, w42258, w42259, w42260, w42261, w42262, w42263, w42264, w42265, w42266, w42267, w42268, w42269, w42270, w42271, w42272, w42273, w42274, w42275, w42276, w42277, w42278, w42279, w42280, w42281, w42282, w42283, w42284, w42285, w42286, w42287, w42288, w42289, w42290, w42291, w42292, w42293, w42294, w42295, w42296, w42297, w42298, w42299, w42300, w42301, w42302, w42303, w42304, w42305, w42306, w42307, w42308, w42309, w42310, w42311, w42312, w42313, w42314, w42315, w42316, w42317, w42318, w42319, w42320, w42321, w42322, w42323, w42324, w42325, w42326, w42327, w42328, w42329, w42330, w42331, w42332, w42333, w42334, w42335, w42336, w42337, w42338, w42339, w42340, w42341, w42342, w42343, w42344, w42345, w42346, w42347, w42348, w42349, w42350, w42351, w42352, w42353, w42354, w42355, w42356, w42357, w42358, w42359, w42360, w42361, w42362, w42363, w42364, w42365, w42366, w42367, w42368, w42369, w42370, w42371, w42372, w42373, w42374, w42375, w42376, w42377, w42378, w42379, w42380, w42381, w42382, w42383, w42384, w42385, w42386, w42387, w42388, w42389, w42390, w42391, w42392, w42393, w42394, w42395, w42396, w42397, w42398, w42399, w42400, w42401, w42402, w42403, w42404, w42405, w42406, w42407, w42408, w42409, w42410, w42411, w42412, w42413, w42414, w42415, w42416, w42417, w42418, w42419, w42420, w42421, w42422, w42423, w42424, w42425, w42426, w42427, w42428, w42429, w42430, w42431, w42432, w42433, w42434, w42435, w42436, w42437, w42438, w42439, w42440, w42441, w42442, w42443, w42444, w42445, w42446, w42447, w42448, w42449, w42450, w42451, w42452, w42453, w42454, w42455, w42456, w42457, w42458, w42459, w42460, w42461, w42462, w42463, w42464, w42465, w42466, w42467, w42468, w42469, w42470, w42471, w42472, w42473, w42474, w42475, w42476, w42477, w42478, w42479, w42480, w42481, w42482, w42483, w42484, w42485, w42486, w42487, w42488, w42489, w42490, w42491, w42492, w42493, w42494, w42495, w42496, w42497, w42498, w42499, w42500, w42501, w42502, w42503, w42504, w42505, w42506, w42507, w42508, w42509, w42510, w42511, w42512, w42513, w42514, w42515, w42516, w42517, w42518, w42519, w42520, w42521, w42522, w42523, w42524, w42525, w42526, w42527, w42528, w42529, w42530, w42531, w42532, w42533, w42534, w42535, w42536, w42537, w42538, w42539, w42540, w42541, w42542, w42543, w42544, w42545, w42546, w42547, w42548, w42549, w42550, w42551, w42552, w42553, w42554, w42555, w42556, w42557, w42558, w42559, w42560, w42561, w42562, w42563, w42564, w42565, w42566, w42567, w42568, w42569, w42570, w42571, w42572, w42573, w42574, w42575, w42576, w42577, w42578, w42579, w42580, w42581, w42582, w42583, w42584, w42585, w42586, w42587, w42588, w42589, w42590, w42591, w42592, w42593, w42594, w42595, w42596, w42597, w42598, w42599, w42600, w42601, w42602, w42603, w42604, w42605, w42606, w42607, w42608, w42609, w42610, w42611, w42612, w42613, w42614, w42615, w42616, w42617, w42618, w42619, w42620, w42621, w42622, w42623, w42624, w42625, w42626, w42627, w42628, w42629, w42630, w42631, w42632, w42633, w42634, w42635, w42636, w42637, w42638, w42639, w42640, w42641, w42642, w42643, w42644, w42645, w42646, w42647, w42648, w42649, w42650, w42651, w42652, w42653, w42654, w42655, w42656, w42657, w42658, w42659, w42660, w42661, w42662, w42663, w42664, w42665, w42666, w42667, w42668, w42669, w42670, w42671, w42672, w42673, w42674, w42675, w42676, w42677, w42678, w42679, w42680, w42681, w42682, w42683, w42684, w42685, w42686, w42687, w42688, w42689, w42690, w42691, w42692, w42693, w42694, w42695, w42696, w42697, w42698, w42699, w42700, w42701, w42702, w42703, w42704, w42705, w42706, w42707, w42708, w42709, w42710, w42711, w42712, w42713, w42714, w42715, w42716, w42717, w42718, w42719, w42720, w42721, w42722, w42723, w42724, w42725, w42726, w42727, w42728, w42729, w42730, w42731, w42732, w42733, w42734, w42735, w42736, w42737, w42738, w42739, w42740, w42741, w42742, w42743, w42744, w42745, w42746, w42747, w42748, w42749, w42750, w42751, w42752, w42753, w42754, w42755, w42756, w42757, w42758, w42759, w42760, w42761, w42762, w42763, w42764, w42765, w42766, w42767, w42768, w42769, w42770, w42771, w42772, w42773, w42774, w42775, w42776, w42777, w42778, w42779, w42780, w42781, w42782, w42783, w42784, w42785, w42786, w42787, w42788, w42789, w42790, w42791, w42792, w42793, w42794, w42795, w42796, w42797, w42798, w42799, w42800, w42801, w42802, w42803, w42804, w42805, w42806, w42807, w42808, w42809, w42810, w42811, w42812, w42813, w42814, w42815, w42816, w42817, w42818, w42819, w42820, w42821, w42822, w42823, w42824, w42825, w42826, w42827, w42828, w42829, w42830, w42831, w42832, w42833, w42834, w42835, w42836, w42837, w42838, w42839, w42840, w42841, w42842, w42843, w42844, w42845, w42846, w42847, w42848, w42849, w42850, w42851, w42852, w42853, w42854, w42855, w42856, w42857, w42858, w42859, w42860, w42861, w42862, w42863, w42864, w42865, w42866, w42867, w42868, w42869, w42870, w42871, w42872, w42873, w42874, w42875, w42876, w42877, w42878, w42879, w42880, w42881, w42882, w42883, w42884, w42885, w42886, w42887, w42888, w42889, w42890, w42891, w42892, w42893, w42894, w42895, w42896, w42897, w42898, w42899, w42900, w42901, w42902, w42903, w42904, w42905, w42906, w42907, w42908, w42909, w42910, w42911, w42912, w42913, w42914, w42915, w42916, w42917, w42918, w42919, w42920, w42921, w42922, w42923, w42924, w42925, w42926, w42927, w42928, w42929, w42930, w42931, w42932, w42933, w42934, w42935, w42936, w42937, w42938, w42939, w42940, w42941, w42942, w42943, w42944, w42945, w42946, w42947, w42948, w42949, w42950, w42951, w42952, w42953, w42954, w42955, w42956, w42957, w42958, w42959, w42960, w42961, w42962, w42963, w42964, w42965, w42966, w42967, w42968, w42969, w42970, w42971, w42972, w42973, w42974, w42975, w42976, w42977, w42978, w42979, w42980, w42981, w42982, w42983, w42984, w42985, w42986, w42987, w42988, w42989, w42990, w42991, w42992, w42993, w42994, w42995, w42996, w42997, w42998, w42999, w43000, w43001, w43002, w43003, w43004, w43005, w43006, w43007, w43008, w43009, w43010, w43011, w43012, w43013, w43014, w43015, w43016, w43017, w43018, w43019, w43020, w43021, w43022, w43023, w43024, w43025, w43026, w43027, w43028, w43029, w43030, w43031, w43032, w43033, w43034, w43035, w43036, w43037, w43038, w43039, w43040, w43041, w43042, w43043, w43044, w43045, w43046, w43047, w43048, w43049, w43050, w43051, w43052, w43053, w43054, w43055, w43056, w43057, w43058, w43059, w43060, w43061, w43062, w43063, w43064, w43065, w43066, w43067, w43068, w43069, w43070, w43071, w43072, w43073, w43074, w43075, w43076, w43077, w43078, w43079, w43080, w43081, w43082, w43083, w43084, w43085, w43086, w43087, w43088, w43089, w43090, w43091, w43092, w43093, w43094, w43095, w43096, w43097, w43098, w43099, w43100, w43101, w43102, w43103, w43104, w43105, w43106, w43107, w43108, w43109, w43110, w43111, w43112, w43113, w43114, w43115, w43116, w43117, w43118, w43119, w43120, w43121, w43122, w43123, w43124, w43125, w43126, w43127, w43128, w43129, w43130, w43131, w43132, w43133, w43134, w43135, w43136, w43137, w43138, w43139, w43140, w43141, w43142, w43143, w43144, w43145, w43146, w43147, w43148, w43149, w43150, w43151, w43152, w43153, w43154, w43155, w43156, w43157, w43158, w43159, w43160, w43161, w43162, w43163, w43164, w43165, w43166, w43167, w43168, w43169, w43170, w43171, w43172, w43173, w43174, w43175, w43176, w43177, w43178, w43179, w43180, w43181, w43182, w43183, w43184, w43185, w43186, w43187, w43188, w43189, w43190, w43191, w43192, w43193, w43194, w43195, w43196, w43197, w43198, w43199, w43200, w43201, w43202, w43203, w43204, w43205, w43206, w43207, w43208, w43209, w43210, w43211, w43212, w43213, w43214, w43215, w43216, w43217, w43218, w43219, w43220, w43221, w43222, w43223, w43224, w43225, w43226, w43227, w43228, w43229, w43230, w43231, w43232, w43233, w43234, w43235, w43236, w43237, w43238, w43239, w43240, w43241, w43242, w43243, w43244, w43245, w43246, w43247, w43248, w43249, w43250, w43251, w43252, w43253, w43254, w43255, w43256, w43257, w43258, w43259, w43260, w43261, w43262, w43263, w43264, w43265, w43266, w43267, w43268, w43269, w43270, w43271, w43272, w43273, w43274, w43275, w43276, w43277, w43278, w43279, w43280, w43281, w43282, w43283, w43284, w43285, w43286, w43287, w43288, w43289, w43290, w43291, w43292, w43293, w43294, w43295, w43296, w43297, w43298, w43299, w43300, w43301, w43302, w43303, w43304, w43305, w43306, w43307, w43308, w43309, w43310, w43311, w43312, w43313, w43314, w43315, w43316, w43317, w43318, w43319, w43320, w43321, w43322, w43323, w43324, w43325, w43326, w43327, w43328, w43329, w43330, w43331, w43332, w43333, w43334, w43335, w43336, w43337, w43338, w43339, w43340, w43341, w43342, w43343, w43344, w43345, w43346, w43347, w43348, w43349, w43350, w43351, w43352, w43353, w43354, w43355, w43356, w43357, w43358, w43359, w43360, w43361, w43362, w43363, w43364, w43365, w43366, w43367, w43368, w43369, w43370, w43371, w43372, w43373, w43374, w43375, w43376, w43377, w43378, w43379, w43380, w43381, w43382, w43383, w43384, w43385, w43386, w43387, w43388, w43389, w43390, w43391, w43392, w43393, w43394, w43395, w43396, w43397, w43398, w43399, w43400, w43401, w43402, w43403, w43404, w43405, w43406, w43407, w43408, w43409, w43410, w43411, w43412, w43413, w43414, w43415, w43416, w43417, w43418, w43419, w43420, w43421, w43422, w43423, w43424, w43425, w43426, w43427, w43428, w43429, w43430, w43431, w43432, w43433, w43434, w43435, w43436, w43437, w43438, w43439, w43440, w43441, w43442, w43443, w43444, w43445, w43446, w43447, w43448, w43449, w43450, w43451, w43452, w43453, w43454, w43455, w43456, w43457, w43458, w43459, w43460, w43461, w43462, w43463, w43464, w43465, w43466, w43467, w43468, w43469, w43470, w43471, w43472, w43473, w43474, w43475, w43476, w43477, w43478, w43479, w43480, w43481, w43482, w43483, w43484, w43485, w43486, w43487, w43488, w43489, w43490, w43491, w43492, w43493, w43494, w43495, w43496, w43497, w43498, w43499, w43500, w43501, w43502, w43503, w43504, w43505, w43506, w43507, w43508, w43509, w43510, w43511, w43512, w43513, w43514, w43515, w43516, w43517, w43518, w43519, w43520, w43521, w43522, w43523, w43524, w43525, w43526, w43527, w43528, w43529, w43530, w43531, w43532, w43533, w43534, w43535, w43536, w43537, w43538, w43539, w43540, w43541, w43542, w43543, w43544, w43545, w43546, w43547, w43548, w43549, w43550, w43551, w43552, w43553, w43554, w43555, w43556, w43557, w43558, w43559, w43560, w43561, w43562, w43563, w43564, w43565, w43566, w43567, w43568, w43569, w43570, w43571, w43572, w43573, w43574, w43575, w43576, w43577, w43578, w43579, w43580, w43581, w43582, w43583, w43584, w43585, w43586, w43587, w43588, w43589, w43590, w43591, w43592, w43593, w43594, w43595, w43596, w43597, w43598, w43599, w43600, w43601, w43602, w43603, w43604, w43605, w43606, w43607, w43608, w43609, w43610, w43611, w43612, w43613, w43614, w43615, w43616, w43617, w43618, w43619, w43620, w43621, w43622, w43623, w43624, w43625, w43626, w43627, w43628, w43629, w43630, w43631, w43632, w43633, w43634, w43635, w43636, w43637, w43638, w43639, w43640, w43641, w43642, w43643, w43644, w43645, w43646, w43647, w43648, w43649, w43650, w43651, w43652, w43653, w43654, w43655, w43656, w43657, w43658, w43659, w43660, w43661, w43662, w43663, w43664, w43665, w43666, w43667, w43668, w43669, w43670, w43671, w43672, w43673, w43674, w43675, w43676, w43677, w43678, w43679, w43680, w43681, w43682, w43683, w43684, w43685, w43686, w43687, w43688, w43689, w43690, w43691, w43692, w43693, w43694, w43695, w43696, w43697, w43698, w43699, w43700, w43701, w43702, w43703, w43704, w43705, w43706, w43707, w43708, w43709, w43710, w43711, w43712, w43713, w43714, w43715, w43716, w43717, w43718, w43719, w43720, w43721, w43722, w43723, w43724, w43725, w43726, w43727, w43728, w43729, w43730, w43731, w43732, w43733, w43734, w43735, w43736, w43737, w43738, w43739, w43740, w43741, w43742, w43743, w43744, w43745, w43746, w43747, w43748, w43749, w43750, w43751, w43752, w43753, w43754, w43755, w43756, w43757, w43758, w43759, w43760, w43761, w43762, w43763, w43764, w43765, w43766, w43767, w43768, w43769, w43770, w43771, w43772, w43773, w43774, w43775, w43776, w43777, w43778, w43779, w43780, w43781, w43782, w43783, w43784, w43785, w43786, w43787, w43788, w43789, w43790, w43791, w43792, w43793, w43794, w43795, w43796, w43797, w43798, w43799, w43800, w43801, w43802, w43803, w43804, w43805, w43806, w43807, w43808, w43809, w43810, w43811, w43812, w43813, w43814, w43815, w43816, w43817, w43818, w43819, w43820, w43821, w43822, w43823, w43824, w43825, w43826, w43827, w43828, w43829, w43830, w43831, w43832, w43833, w43834, w43835, w43836, w43837, w43838, w43839, w43840, w43841, w43842, w43843, w43844, w43845, w43846, w43847, w43848, w43849, w43850, w43851, w43852, w43853, w43854, w43855, w43856, w43857, w43858, w43859, w43860, w43861, w43862, w43863, w43864, w43865, w43866, w43867, w43868, w43869, w43870, w43871, w43872, w43873, w43874, w43875, w43876, w43877, w43878, w43879, w43880, w43881, w43882, w43883, w43884, w43885, w43886, w43887, w43888, w43889, w43890, w43891, w43892, w43893, w43894, w43895, w43896, w43897, w43898, w43899, w43900, w43901, w43902, w43903, w43904, w43905, w43906, w43907, w43908, w43909, w43910, w43911, w43912, w43913, w43914, w43915, w43916, w43917, w43918, w43919, w43920, w43921, w43922, w43923, w43924, w43925, w43926, w43927, w43928, w43929, w43930, w43931, w43932, w43933, w43934, w43935, w43936, w43937, w43938, w43939, w43940, w43941, w43942, w43943, w43944, w43945, w43946, w43947, w43948, w43949, w43950, w43951, w43952, w43953, w43954, w43955, w43956, w43957, w43958, w43959, w43960, w43961, w43962, w43963, w43964, w43965, w43966, w43967, w43968, w43969, w43970, w43971, w43972, w43973, w43974, w43975, w43976, w43977, w43978, w43979, w43980, w43981, w43982, w43983, w43984, w43985, w43986, w43987, w43988, w43989, w43990, w43991, w43992, w43993, w43994, w43995, w43996, w43997, w43998, w43999, w44000, w44001, w44002, w44003, w44004, w44005, w44006, w44007, w44008, w44009, w44010, w44011, w44012, w44013, w44014, w44015, w44016, w44017, w44018, w44019, w44020, w44021, w44022, w44023, w44024, w44025, w44026, w44027, w44028, w44029, w44030, w44031, w44032, w44033, w44034, w44035, w44036, w44037, w44038, w44039, w44040, w44041, w44042, w44043, w44044, w44045, w44046, w44047, w44048, w44049, w44050, w44051, w44052, w44053, w44054, w44055, w44056, w44057, w44058, w44059, w44060, w44061, w44062, w44063, w44064, w44065, w44066, w44067, w44068, w44069, w44070, w44071, w44072, w44073, w44074, w44075, w44076, w44077, w44078, w44079, w44080, w44081, w44082, w44083, w44084, w44085, w44086, w44087, w44088, w44089, w44090, w44091, w44092, w44093, w44094, w44095, w44096, w44097, w44098, w44099, w44100, w44101, w44102, w44103, w44104, w44105, w44106, w44107, w44108, w44109, w44110, w44111, w44112, w44113, w44114, w44115, w44116, w44117, w44118, w44119, w44120, w44121, w44122, w44123, w44124, w44125, w44126, w44127, w44128, w44129, w44130, w44131, w44132, w44133, w44134, w44135, w44136, w44137, w44138, w44139, w44140, w44141, w44142, w44143, w44144, w44145, w44146, w44147, w44148, w44149, w44150, w44151, w44152, w44153, w44154, w44155, w44156, w44157, w44158, w44159, w44160, w44161, w44162, w44163, w44164, w44165, w44166, w44167, w44168, w44169, w44170, w44171, w44172, w44173, w44174, w44175, w44176, w44177, w44178, w44179, w44180, w44181, w44182, w44183, w44184, w44185, w44186, w44187, w44188, w44189, w44190, w44191, w44192, w44193, w44194, w44195, w44196, w44197, w44198, w44199, w44200, w44201, w44202, w44203, w44204, w44205, w44206, w44207, w44208, w44209, w44210, w44211, w44212, w44213, w44214, w44215, w44216, w44217, w44218, w44219, w44220, w44221, w44222, w44223, w44224, w44225, w44226, w44227, w44228, w44229, w44230, w44231, w44232, w44233, w44234, w44235, w44236, w44237, w44238, w44239, w44240, w44241, w44242, w44243, w44244, w44245, w44246, w44247, w44248, w44249, w44250, w44251, w44252, w44253, w44254, w44255, w44256, w44257, w44258, w44259, w44260, w44261, w44262, w44263, w44264, w44265, w44266, w44267, w44268, w44269, w44270, w44271, w44272, w44273, w44274, w44275, w44276, w44277, w44278, w44279, w44280, w44281, w44282, w44283, w44284, w44285, w44286, w44287, w44288, w44289, w44290, w44291, w44292, w44293, w44294, w44295, w44296, w44297, w44298, w44299, w44300, w44301, w44302, w44303, w44304, w44305, w44306, w44307, w44308, w44309, w44310, w44311, w44312, w44313, w44314, w44315, w44316, w44317, w44318, w44319, w44320, w44321, w44322, w44323, w44324, w44325, w44326, w44327, w44328, w44329, w44330, w44331, w44332, w44333, w44334, w44335, w44336, w44337, w44338, w44339, w44340, w44341, w44342, w44343, w44344, w44345, w44346, w44347, w44348, w44349, w44350, w44351, w44352, w44353, w44354, w44355, w44356, w44357, w44358, w44359, w44360, w44361, w44362, w44363, w44364, w44365, w44366, w44367, w44368, w44369, w44370, w44371, w44372, w44373, w44374, w44375, w44376, w44377, w44378, w44379, w44380, w44381, w44382, w44383, w44384, w44385, w44386, w44387, w44388, w44389, w44390, w44391, w44392, w44393, w44394, w44395, w44396, w44397, w44398, w44399, w44400, w44401, w44402, w44403, w44404, w44405, w44406, w44407, w44408, w44409, w44410, w44411, w44412, w44413, w44414, w44415, w44416, w44417, w44418, w44419, w44420, w44421, w44422, w44423, w44424, w44425, w44426, w44427, w44428, w44429, w44430, w44431, w44432, w44433, w44434, w44435, w44436, w44437, w44438, w44439, w44440, w44441, w44442, w44443, w44444, w44445, w44446, w44447, w44448, w44449, w44450, w44451, w44452, w44453, w44454, w44455, w44456, w44457, w44458, w44459, w44460, w44461, w44462, w44463, w44464, w44465, w44466, w44467, w44468, w44469, w44470, w44471, w44472, w44473, w44474, w44475, w44476, w44477, w44478, w44479, w44480, w44481, w44482, w44483, w44484, w44485, w44486, w44487, w44488, w44489, w44490, w44491, w44492, w44493, w44494, w44495, w44496, w44497, w44498, w44499, w44500, w44501, w44502, w44503, w44504, w44505, w44506, w44507, w44508, w44509, w44510, w44511, w44512, w44513, w44514, w44515, w44516, w44517, w44518, w44519, w44520, w44521, w44522, w44523, w44524, w44525, w44526, w44527, w44528, w44529, w44530, w44531, w44532, w44533, w44534, w44535, w44536, w44537, w44538, w44539, w44540, w44541, w44542, w44543, w44544, w44545, w44546, w44547, w44548, w44549, w44550, w44551, w44552, w44553, w44554, w44555, w44556, w44557, w44558, w44559, w44560, w44561, w44562, w44563, w44564, w44565, w44566, w44567, w44568, w44569, w44570, w44571, w44572, w44573, w44574, w44575, w44576, w44577, w44578, w44579, w44580, w44581, w44582, w44583, w44584, w44585, w44586, w44587, w44588, w44589, w44590, w44591, w44592, w44593, w44594, w44595, w44596, w44597, w44598, w44599, w44600, w44601, w44602, w44603, w44604, w44605, w44606, w44607, w44608, w44609, w44610, w44611, w44612, w44613, w44614, w44615, w44616, w44617, w44618, w44619, w44620, w44621, w44622, w44623, w44624, w44625, w44626, w44627, w44628, w44629, w44630, w44631, w44632, w44633, w44634, w44635, w44636, w44637, w44638, w44639, w44640, w44641, w44642, w44643, w44644, w44645, w44646, w44647, w44648, w44649, w44650, w44651, w44652, w44653, w44654, w44655, w44656, w44657, w44658, w44659, w44660, w44661, w44662, w44663, w44664, w44665, w44666, w44667, w44668, w44669, w44670, w44671, w44672, w44673, w44674, w44675, w44676, w44677, w44678, w44679, w44680, w44681, w44682, w44683, w44684, w44685, w44686, w44687, w44688, w44689, w44690, w44691, w44692, w44693, w44694, w44695, w44696, w44697, w44698, w44699, w44700, w44701, w44702, w44703, w44704, w44705, w44706, w44707, w44708, w44709, w44710, w44711, w44712, w44713, w44714, w44715, w44716, w44717, w44718, w44719, w44720, w44721, w44722, w44723, w44724, w44725, w44726, w44727, w44728, w44729, w44730, w44731, w44732, w44733, w44734, w44735, w44736, w44737, w44738, w44739, w44740, w44741, w44742, w44743, w44744, w44745, w44746, w44747, w44748, w44749, w44750, w44751, w44752, w44753, w44754, w44755, w44756, w44757, w44758, w44759, w44760, w44761, w44762, w44763, w44764, w44765, w44766, w44767, w44768, w44769, w44770, w44771, w44772, w44773, w44774, w44775, w44776, w44777, w44778, w44779, w44780, w44781, w44782, w44783, w44784, w44785, w44786, w44787, w44788, w44789, w44790, w44791, w44792, w44793, w44794, w44795, w44796, w44797, w44798, w44799, w44800, w44801, w44802, w44803, w44804, w44805, w44806, w44807, w44808, w44809, w44810, w44811, w44812, w44813, w44814, w44815, w44816, w44817, w44818, w44819, w44820, w44821, w44822, w44823, w44824, w44825, w44826, w44827, w44828, w44829, w44830, w44831, w44832, w44833, w44834, w44835, w44836, w44837, w44838, w44839, w44840, w44841, w44842, w44843, w44844, w44845, w44846, w44847, w44848, w44849, w44850, w44851, w44852, w44853, w44854, w44855, w44856, w44857, w44858, w44859, w44860, w44861, w44862, w44863, w44864, w44865, w44866, w44867, w44868, w44869, w44870, w44871, w44872, w44873, w44874, w44875, w44876, w44877, w44878, w44879, w44880, w44881, w44882, w44883, w44884, w44885, w44886, w44887, w44888, w44889, w44890, w44891, w44892, w44893, w44894, w44895, w44896, w44897, w44898, w44899, w44900, w44901, w44902, w44903, w44904, w44905, w44906, w44907, w44908, w44909, w44910, w44911, w44912, w44913, w44914, w44915, w44916, w44917, w44918, w44919, w44920, w44921, w44922, w44923, w44924, w44925, w44926, w44927, w44928, w44929, w44930, w44931, w44932, w44933, w44934, w44935, w44936, w44937, w44938, w44939, w44940, w44941, w44942, w44943, w44944, w44945, w44946, w44947, w44948, w44949, w44950, w44951, w44952, w44953, w44954, w44955, w44956, w44957, w44958, w44959, w44960, w44961, w44962, w44963, w44964, w44965, w44966, w44967, w44968, w44969, w44970, w44971, w44972, w44973, w44974, w44975, w44976, w44977, w44978, w44979, w44980, w44981, w44982, w44983, w44984, w44985, w44986, w44987, w44988, w44989, w44990, w44991, w44992, w44993, w44994, w44995, w44996, w44997, w44998, w44999, w45000, w45001, w45002, w45003, w45004, w45005, w45006, w45007, w45008, w45009, w45010, w45011, w45012, w45013, w45014, w45015, w45016, w45017, w45018, w45019, w45020, w45021, w45022, w45023, w45024, w45025, w45026, w45027, w45028, w45029, w45030, w45031, w45032, w45033, w45034, w45035, w45036, w45037, w45038, w45039, w45040, w45041, w45042, w45043, w45044, w45045, w45046, w45047, w45048, w45049, w45050, w45051, w45052, w45053, w45054, w45055, w45056, w45057, w45058, w45059, w45060, w45061, w45062, w45063, w45064, w45065, w45066, w45067, w45068, w45069, w45070, w45071, w45072, w45073, w45074, w45075, w45076, w45077, w45078, w45079, w45080, w45081, w45082, w45083, w45084, w45085, w45086, w45087, w45088, w45089, w45090, w45091, w45092, w45093, w45094, w45095, w45096, w45097, w45098, w45099, w45100, w45101, w45102, w45103, w45104, w45105, w45106, w45107, w45108, w45109, w45110, w45111, w45112, w45113, w45114, w45115, w45116, w45117, w45118, w45119, w45120, w45121, w45122, w45123, w45124, w45125, w45126, w45127, w45128, w45129, w45130, w45131, w45132, w45133, w45134, w45135, w45136, w45137, w45138, w45139, w45140, w45141, w45142, w45143, w45144, w45145, w45146, w45147, w45148, w45149, w45150, w45151, w45152, w45153, w45154, w45155, w45156, w45157, w45158, w45159, w45160, w45161, w45162, w45163, w45164, w45165, w45166, w45167, w45168, w45169, w45170, w45171, w45172, w45173, w45174, w45175, w45176, w45177, w45178, w45179, w45180, w45181, w45182, w45183, w45184, w45185, w45186, w45187, w45188, w45189, w45190, w45191, w45192, w45193, w45194, w45195, w45196, w45197, w45198, w45199, w45200, w45201, w45202, w45203, w45204, w45205, w45206, w45207, w45208, w45209, w45210, w45211, w45212, w45213, w45214, w45215, w45216, w45217, w45218, w45219, w45220, w45221, w45222, w45223, w45224, w45225, w45226, w45227, w45228, w45229, w45230, w45231, w45232, w45233, w45234, w45235, w45236, w45237, w45238, w45239, w45240, w45241, w45242, w45243, w45244, w45245, w45246, w45247, w45248, w45249, w45250, w45251, w45252, w45253, w45254, w45255, w45256, w45257, w45258, w45259, w45260, w45261, w45262, w45263, w45264, w45265, w45266, w45267, w45268, w45269, w45270, w45271, w45272, w45273, w45274, w45275, w45276, w45277, w45278, w45279, w45280, w45281, w45282, w45283, w45284, w45285, w45286, w45287, w45288, w45289, w45290, w45291, w45292, w45293, w45294, w45295, w45296, w45297, w45298, w45299, w45300, w45301, w45302, w45303, w45304, w45305, w45306, w45307, w45308, w45309, w45310, w45311, w45312, w45313, w45314, w45315, w45316, w45317, w45318, w45319, w45320, w45321, w45322, w45323, w45324, w45325, w45326, w45327, w45328, w45329, w45330, w45331, w45332, w45333, w45334, w45335, w45336, w45337, w45338, w45339, w45340, w45341, w45342, w45343, w45344, w45345, w45346, w45347, w45348, w45349, w45350, w45351, w45352, w45353, w45354, w45355, w45356, w45357, w45358, w45359, w45360, w45361, w45362, w45363, w45364, w45365, w45366, w45367, w45368, w45369, w45370, w45371, w45372, w45373, w45374, w45375, w45376, w45377, w45378, w45379, w45380, w45381, w45382, w45383, w45384, w45385, w45386, w45387, w45388, w45389, w45390, w45391, w45392, w45393, w45394, w45395, w45396, w45397, w45398, w45399, w45400, w45401, w45402, w45403, w45404, w45405, w45406, w45407, w45408, w45409, w45410, w45411, w45412, w45413, w45414, w45415, w45416, w45417, w45418, w45419, w45420, w45421, w45422, w45423, w45424, w45425, w45426, w45427, w45428, w45429, w45430, w45431, w45432, w45433, w45434, w45435, w45436, w45437, w45438, w45439, w45440, w45441, w45442, w45443, w45444, w45445, w45446, w45447, w45448, w45449, w45450, w45451, w45452, w45453, w45454, w45455, w45456, w45457, w45458, w45459, w45460, w45461, w45462, w45463, w45464, w45465, w45466, w45467, w45468, w45469, w45470, w45471, w45472, w45473, w45474, w45475, w45476, w45477, w45478, w45479, w45480, w45481, w45482, w45483, w45484, w45485, w45486, w45487, w45488, w45489, w45490, w45491, w45492, w45493, w45494, w45495, w45496, w45497, w45498, w45499, w45500, w45501, w45502, w45503, w45504, w45505, w45506, w45507, w45508, w45509, w45510, w45511, w45512, w45513, w45514, w45515, w45516, w45517, w45518, w45519, w45520, w45521, w45522, w45523, w45524, w45525, w45526, w45527, w45528, w45529, w45530, w45531, w45532, w45533, w45534, w45535, w45536, w45537, w45538, w45539, w45540, w45541, w45542, w45543, w45544, w45545, w45546, w45547, w45548, w45549, w45550, w45551, w45552, w45553, w45554, w45555, w45556, w45557, w45558, w45559, w45560, w45561, w45562, w45563, w45564, w45565, w45566, w45567, w45568, w45569, w45570, w45571, w45572, w45573, w45574, w45575, w45576, w45577, w45578, w45579, w45580, w45581, w45582, w45583, w45584, w45585, w45586, w45587, w45588, w45589, w45590, w45591, w45592, w45593, w45594, w45595, w45596, w45597, w45598, w45599, w45600, w45601, w45602, w45603, w45604, w45605, w45606, w45607, w45608, w45609, w45610, w45611, w45612, w45613, w45614, w45615, w45616, w45617, w45618, w45619, w45620, w45621, w45622, w45623, w45624, w45625, w45626, w45627, w45628, w45629, w45630, w45631, w45632, w45633, w45634, w45635, w45636, w45637, w45638, w45639, w45640, w45641, w45642, w45643, w45644, w45645, w45646, w45647, w45648, w45649, w45650, w45651, w45652, w45653, w45654, w45655, w45656, w45657, w45658, w45659, w45660, w45661, w45662, w45663, w45664, w45665, w45666, w45667, w45668, w45669, w45670, w45671, w45672, w45673, w45674, w45675, w45676, w45677, w45678, w45679, w45680, w45681, w45682, w45683, w45684, w45685, w45686, w45687, w45688, w45689, w45690, w45691, w45692, w45693, w45694, w45695, w45696, w45697, w45698, w45699, w45700, w45701, w45702, w45703, w45704, w45705, w45706, w45707, w45708, w45709, w45710, w45711, w45712, w45713, w45714, w45715, w45716, w45717, w45718, w45719, w45720, w45721, w45722, w45723, w45724, w45725, w45726, w45727, w45728, w45729, w45730, w45731, w45732, w45733, w45734, w45735, w45736, w45737, w45738, w45739, w45740, w45741, w45742, w45743, w45744, w45745, w45746, w45747, w45748, w45749, w45750, w45751, w45752, w45753, w45754, w45755, w45756, w45757, w45758, w45759, w45760, w45761, w45762, w45763, w45764, w45765, w45766, w45767, w45768, w45769, w45770, w45771, w45772, w45773, w45774, w45775, w45776, w45777, w45778, w45779, w45780, w45781, w45782, w45783, w45784, w45785, w45786, w45787, w45788, w45789, w45790, w45791, w45792, w45793, w45794, w45795, w45796, w45797, w45798, w45799, w45800, w45801, w45802, w45803, w45804, w45805, w45806, w45807, w45808, w45809, w45810, w45811, w45812, w45813, w45814, w45815, w45816, w45817, w45818, w45819, w45820, w45821, w45822, w45823, w45824, w45825, w45826, w45827, w45828, w45829, w45830, w45831, w45832, w45833, w45834, w45835, w45836, w45837, w45838, w45839, w45840, w45841, w45842, w45843, w45844, w45845, w45846, w45847, w45848, w45849, w45850, w45851, w45852, w45853, w45854, w45855, w45856, w45857, w45858, w45859, w45860, w45861, w45862, w45863, w45864, w45865, w45866, w45867, w45868, w45869, w45870, w45871, w45872, w45873, w45874, w45875, w45876, w45877, w45878, w45879, w45880, w45881, w45882, w45883, w45884, w45885, w45886, w45887, w45888, w45889, w45890, w45891, w45892, w45893, w45894, w45895, w45896, w45897, w45898, w45899, w45900, w45901, w45902, w45903, w45904, w45905, w45906, w45907, w45908, w45909, w45910, w45911, w45912, w45913, w45914, w45915, w45916, w45917, w45918, w45919, w45920, w45921, w45922, w45923, w45924, w45925, w45926, w45927, w45928, w45929, w45930, w45931, w45932, w45933, w45934, w45935, w45936, w45937, w45938, w45939, w45940, w45941, w45942, w45943, w45944, w45945, w45946, w45947, w45948, w45949, w45950, w45951, w45952, w45953, w45954, w45955, w45956, w45957, w45958, w45959, w45960, w45961, w45962, w45963, w45964, w45965, w45966, w45967, w45968, w45969, w45970, w45971, w45972, w45973, w45974, w45975, w45976, w45977, w45978, w45979, w45980, w45981, w45982, w45983, w45984, w45985, w45986, w45987, w45988, w45989, w45990, w45991, w45992, w45993, w45994, w45995, w45996, w45997, w45998, w45999, w46000, w46001, w46002, w46003, w46004, w46005, w46006, w46007, w46008, w46009, w46010, w46011, w46012, w46013, w46014, w46015, w46016, w46017, w46018, w46019, w46020, w46021, w46022, w46023, w46024, w46025, w46026, w46027, w46028, w46029, w46030, w46031, w46032, w46033, w46034, w46035, w46036, w46037, w46038, w46039, w46040, w46041, w46042, w46043, w46044, w46045, w46046, w46047, w46048, w46049, w46050, w46051, w46052, w46053, w46054, w46055, w46056, w46057, w46058, w46059, w46060, w46061, w46062, w46063, w46064, w46065, w46066, w46067, w46068, w46069, w46070, w46071, w46072, w46073, w46074, w46075, w46076, w46077, w46078, w46079, w46080, w46081, w46082, w46083, w46084, w46085, w46086, w46087, w46088, w46089, w46090, w46091, w46092, w46093, w46094, w46095, w46096, w46097, w46098, w46099, w46100, w46101, w46102, w46103, w46104, w46105, w46106, w46107, w46108, w46109, w46110, w46111, w46112, w46113, w46114, w46115, w46116, w46117, w46118, w46119, w46120, w46121, w46122, w46123, w46124, w46125, w46126, w46127, w46128, w46129, w46130, w46131, w46132, w46133, w46134, w46135, w46136, w46137, w46138, w46139, w46140, w46141, w46142, w46143, w46144, w46145, w46146, w46147, w46148, w46149, w46150, w46151, w46152, w46153, w46154, w46155, w46156, w46157, w46158, w46159, w46160, w46161, w46162, w46163, w46164, w46165, w46166, w46167, w46168, w46169, w46170, w46171, w46172, w46173, w46174, w46175, w46176, w46177, w46178, w46179, w46180, w46181, w46182, w46183, w46184, w46185, w46186, w46187, w46188, w46189, w46190, w46191, w46192, w46193, w46194, w46195, w46196, w46197, w46198, w46199, w46200, w46201, w46202, w46203, w46204, w46205, w46206, w46207, w46208, w46209, w46210, w46211, w46212, w46213, w46214, w46215, w46216, w46217, w46218, w46219, w46220, w46221, w46222, w46223, w46224, w46225, w46226, w46227, w46228, w46229, w46230, w46231, w46232, w46233, w46234, w46235, w46236, w46237, w46238, w46239, w46240, w46241, w46242, w46243, w46244, w46245, w46246, w46247, w46248, w46249, w46250, w46251, w46252, w46253, w46254, w46255, w46256, w46257, w46258, w46259, w46260, w46261, w46262, w46263, w46264, w46265, w46266, w46267, w46268, w46269, w46270, w46271, w46272, w46273, w46274, w46275, w46276, w46277, w46278, w46279, w46280, w46281, w46282, w46283, w46284, w46285, w46286, w46287, w46288, w46289, w46290, w46291, w46292, w46293, w46294, w46295, w46296, w46297, w46298, w46299, w46300, w46301, w46302, w46303, w46304, w46305, w46306, w46307, w46308, w46309, w46310, w46311, w46312, w46313, w46314, w46315, w46316, w46317, w46318, w46319, w46320, w46321, w46322, w46323, w46324, w46325, w46326, w46327, w46328, w46329, w46330, w46331, w46332, w46333, w46334, w46335, w46336, w46337, w46338, w46339, w46340, w46341, w46342, w46343, w46344, w46345, w46346, w46347, w46348, w46349, w46350, w46351, w46352, w46353, w46354, w46355, w46356, w46357, w46358, w46359, w46360, w46361, w46362, w46363, w46364, w46365, w46366, w46367, w46368, w46369, w46370, w46371, w46372, w46373, w46374, w46375, w46376, w46377, w46378, w46379, w46380, w46381, w46382, w46383, w46384, w46385, w46386, w46387, w46388, w46389, w46390, w46391, w46392, w46393, w46394, w46395, w46396, w46397, w46398, w46399, w46400, w46401, w46402, w46403, w46404, w46405, w46406, w46407, w46408, w46409, w46410, w46411, w46412, w46413, w46414, w46415, w46416, w46417, w46418, w46419, w46420, w46421, w46422, w46423, w46424, w46425, w46426, w46427, w46428, w46429, w46430, w46431, w46432, w46433, w46434, w46435, w46436, w46437, w46438, w46439, w46440, w46441, w46442, w46443, w46444, w46445, w46446, w46447, w46448, w46449, w46450, w46451, w46452, w46453, w46454, w46455, w46456, w46457, w46458, w46459, w46460, w46461, w46462, w46463, w46464, w46465, w46466, w46467, w46468, w46469, w46470, w46471, w46472, w46473, w46474, w46475, w46476, w46477, w46478, w46479, w46480, w46481, w46482, w46483, w46484, w46485, w46486, w46487, w46488, w46489, w46490, w46491, w46492, w46493, w46494, w46495, w46496, w46497, w46498, w46499, w46500, w46501, w46502, w46503, w46504, w46505, w46506, w46507, w46508, w46509, w46510, w46511, w46512, w46513, w46514, w46515, w46516, w46517, w46518, w46519, w46520, w46521, w46522, w46523, w46524, w46525, w46526, w46527, w46528, w46529, w46530, w46531, w46532, w46533, w46534, w46535, w46536, w46537, w46538, w46539, w46540, w46541, w46542, w46543, w46544, w46545, w46546, w46547, w46548, w46549, w46550, w46551, w46552, w46553, w46554, w46555, w46556, w46557, w46558, w46559, w46560, w46561, w46562, w46563, w46564, w46565, w46566, w46567, w46568, w46569, w46570, w46571, w46572, w46573, w46574, w46575, w46576, w46577, w46578, w46579, w46580, w46581, w46582, w46583, w46584, w46585, w46586, w46587, w46588, w46589, w46590, w46591, w46592, w46593, w46594, w46595, w46596, w46597, w46598, w46599, w46600, w46601, w46602, w46603, w46604, w46605, w46606, w46607, w46608, w46609, w46610, w46611, w46612, w46613, w46614, w46615, w46616, w46617, w46618, w46619, w46620, w46621, w46622, w46623, w46624, w46625, w46626, w46627, w46628, w46629, w46630, w46631, w46632, w46633, w46634, w46635, w46636, w46637, w46638, w46639, w46640, w46641, w46642, w46643, w46644, w46645, w46646, w46647, w46648, w46649, w46650, w46651, w46652, w46653, w46654, w46655, w46656, w46657, w46658, w46659, w46660, w46661, w46662, w46663, w46664, w46665, w46666, w46667, w46668, w46669, w46670, w46671, w46672, w46673, w46674, w46675, w46676, w46677, w46678, w46679, w46680, w46681, w46682, w46683, w46684, w46685, w46686, w46687, w46688, w46689, w46690, w46691, w46692, w46693, w46694, w46695, w46696, w46697, w46698, w46699, w46700, w46701, w46702, w46703, w46704, w46705, w46706, w46707, w46708, w46709, w46710, w46711, w46712, w46713, w46714, w46715, w46716, w46717, w46718, w46719, w46720, w46721, w46722, w46723, w46724, w46725, w46726, w46727, w46728, w46729, w46730, w46731, w46732, w46733, w46734, w46735, w46736, w46737, w46738, w46739, w46740, w46741, w46742, w46743, w46744, w46745, w46746, w46747, w46748, w46749, w46750, w46751, w46752, w46753, w46754, w46755, w46756, w46757, w46758, w46759, w46760, w46761, w46762, w46763, w46764, w46765, w46766, w46767, w46768, w46769, w46770, w46771, w46772, w46773, w46774, w46775, w46776, w46777, w46778, w46779, w46780, w46781, w46782, w46783, w46784, w46785, w46786, w46787, w46788, w46789, w46790, w46791, w46792, w46793, w46794, w46795, w46796, w46797, w46798, w46799, w46800, w46801, w46802, w46803, w46804, w46805, w46806, w46807, w46808, w46809, w46810, w46811, w46812, w46813, w46814, w46815, w46816, w46817, w46818, w46819, w46820, w46821, w46822, w46823, w46824, w46825, w46826, w46827, w46828, w46829, w46830, w46831, w46832, w46833, w46834, w46835, w46836, w46837, w46838, w46839, w46840, w46841, w46842, w46843, w46844, w46845, w46846, w46847, w46848, w46849, w46850, w46851, w46852, w46853, w46854, w46855, w46856, w46857, w46858, w46859, w46860, w46861, w46862, w46863, w46864, w46865, w46866, w46867, w46868, w46869, w46870, w46871, w46872, w46873, w46874, w46875, w46876, w46877, w46878, w46879, w46880, w46881, w46882, w46883, w46884, w46885, w46886, w46887, w46888, w46889, w46890, w46891, w46892, w46893, w46894, w46895, w46896, w46897, w46898, w46899, w46900, w46901, w46902, w46903, w46904, w46905, w46906, w46907, w46908, w46909, w46910, w46911, w46912, w46913, w46914, w46915, w46916, w46917, w46918, w46919, w46920, w46921, w46922, w46923, w46924, w46925, w46926, w46927, w46928, w46929, w46930, w46931, w46932, w46933, w46934, w46935, w46936, w46937, w46938, w46939, w46940, w46941, w46942, w46943, w46944, w46945, w46946, w46947, w46948, w46949, w46950, w46951, w46952, w46953, w46954, w46955, w46956, w46957, w46958, w46959, w46960, w46961, w46962, w46963, w46964, w46965, w46966, w46967, w46968, w46969, w46970, w46971, w46972, w46973, w46974, w46975, w46976, w46977, w46978, w46979, w46980, w46981, w46982, w46983, w46984, w46985, w46986, w46987, w46988, w46989, w46990, w46991, w46992, w46993, w46994, w46995, w46996, w46997, w46998, w46999, w47000, w47001, w47002, w47003, w47004, w47005, w47006, w47007, w47008, w47009, w47010, w47011, w47012, w47013, w47014, w47015, w47016, w47017, w47018, w47019, w47020, w47021, w47022, w47023, w47024, w47025, w47026, w47027, w47028, w47029, w47030, w47031, w47032, w47033, w47034, w47035, w47036, w47037, w47038, w47039, w47040, w47041, w47042, w47043, w47044, w47045, w47046, w47047, w47048, w47049, w47050, w47051, w47052, w47053, w47054, w47055, w47056, w47057, w47058, w47059, w47060, w47061, w47062, w47063, w47064, w47065, w47066, w47067, w47068, w47069, w47070, w47071, w47072, w47073, w47074, w47075, w47076, w47077, w47078, w47079, w47080, w47081, w47082, w47083, w47084, w47085, w47086, w47087, w47088, w47089, w47090, w47091, w47092, w47093, w47094, w47095, w47096, w47097, w47098, w47099, w47100, w47101, w47102, w47103, w47104, w47105, w47106, w47107, w47108, w47109, w47110, w47111, w47112, w47113, w47114, w47115, w47116, w47117, w47118, w47119, w47120, w47121, w47122, w47123, w47124, w47125, w47126, w47127, w47128, w47129, w47130, w47131, w47132, w47133, w47134, w47135, w47136, w47137, w47138, w47139, w47140, w47141, w47142, w47143, w47144, w47145, w47146, w47147, w47148, w47149, w47150, w47151, w47152, w47153, w47154, w47155, w47156, w47157, w47158, w47159, w47160, w47161, w47162, w47163, w47164, w47165, w47166, w47167, w47168, w47169, w47170, w47171, w47172, w47173, w47174, w47175, w47176, w47177, w47178, w47179, w47180, w47181, w47182, w47183, w47184, w47185, w47186, w47187, w47188, w47189, w47190, w47191, w47192, w47193, w47194, w47195, w47196, w47197, w47198, w47199, w47200, w47201, w47202, w47203, w47204, w47205, w47206, w47207, w47208, w47209, w47210, w47211, w47212, w47213, w47214, w47215, w47216, w47217, w47218, w47219, w47220, w47221, w47222, w47223, w47224, w47225, w47226, w47227, w47228, w47229, w47230, w47231, w47232, w47233, w47234, w47235, w47236, w47237, w47238, w47239, w47240, w47241, w47242, w47243, w47244, w47245, w47246, w47247, w47248, w47249, w47250, w47251, w47252, w47253, w47254, w47255, w47256, w47257, w47258, w47259, w47260, w47261, w47262, w47263, w47264, w47265, w47266, w47267, w47268, w47269, w47270, w47271, w47272, w47273, w47274, w47275, w47276, w47277, w47278, w47279, w47280, w47281, w47282, w47283, w47284, w47285, w47286, w47287, w47288, w47289, w47290, w47291, w47292, w47293, w47294, w47295, w47296, w47297, w47298, w47299, w47300, w47301, w47302, w47303, w47304, w47305, w47306, w47307, w47308, w47309, w47310, w47311, w47312, w47313, w47314, w47315, w47316, w47317, w47318, w47319, w47320, w47321, w47322, w47323, w47324, w47325, w47326, w47327, w47328, w47329, w47330, w47331, w47332, w47333, w47334, w47335, w47336, w47337, w47338, w47339, w47340, w47341, w47342, w47343, w47344, w47345, w47346, w47347, w47348, w47349, w47350, w47351, w47352, w47353, w47354, w47355, w47356, w47357, w47358, w47359, w47360, w47361, w47362, w47363, w47364, w47365, w47366, w47367, w47368, w47369, w47370, w47371, w47372, w47373, w47374, w47375, w47376, w47377, w47378, w47379, w47380, w47381, w47382, w47383, w47384, w47385, w47386, w47387, w47388, w47389, w47390, w47391, w47392, w47393, w47394, w47395, w47396, w47397, w47398, w47399, w47400, w47401, w47402, w47403, w47404, w47405, w47406, w47407, w47408, w47409, w47410, w47411, w47412, w47413, w47414, w47415, w47416, w47417, w47418, w47419, w47420, w47421, w47422, w47423, w47424, w47425, w47426, w47427, w47428, w47429, w47430, w47431, w47432, w47433, w47434, w47435, w47436, w47437, w47438, w47439, w47440, w47441, w47442, w47443, w47444, w47445, w47446, w47447, w47448, w47449, w47450, w47451, w47452, w47453, w47454, w47455, w47456, w47457, w47458, w47459, w47460, w47461, w47462, w47463, w47464, w47465, w47466, w47467, w47468, w47469, w47470, w47471, w47472, w47473, w47474, w47475, w47476, w47477, w47478, w47479, w47480, w47481, w47482, w47483, w47484, w47485, w47486, w47487, w47488, w47489, w47490, w47491, w47492, w47493, w47494, w47495, w47496, w47497, w47498, w47499, w47500, w47501, w47502, w47503, w47504, w47505, w47506, w47507, w47508, w47509, w47510, w47511, w47512, w47513, w47514, w47515, w47516, w47517, w47518, w47519, w47520, w47521, w47522, w47523, w47524, w47525, w47526, w47527, w47528, w47529, w47530, w47531, w47532, w47533, w47534, w47535, w47536, w47537, w47538, w47539, w47540, w47541, w47542, w47543, w47544, w47545, w47546, w47547, w47548, w47549, w47550, w47551, w47552, w47553, w47554, w47555, w47556, w47557, w47558, w47559, w47560, w47561, w47562, w47563, w47564, w47565, w47566, w47567, w47568, w47569, w47570, w47571, w47572, w47573, w47574, w47575, w47576, w47577, w47578, w47579, w47580, w47581, w47582, w47583, w47584, w47585, w47586, w47587, w47588, w47589, w47590, w47591, w47592, w47593, w47594, w47595, w47596, w47597, w47598, w47599, w47600, w47601, w47602, w47603, w47604, w47605, w47606, w47607, w47608, w47609, w47610, w47611, w47612, w47613, w47614, w47615, w47616, w47617, w47618, w47619, w47620, w47621, w47622, w47623, w47624, w47625, w47626, w47627, w47628, w47629, w47630, w47631, w47632, w47633, w47634, w47635, w47636, w47637, w47638, w47639, w47640, w47641, w47642, w47643, w47644, w47645, w47646, w47647, w47648, w47649, w47650, w47651, w47652, w47653, w47654, w47655, w47656, w47657, w47658, w47659, w47660, w47661, w47662, w47663, w47664, w47665, w47666, w47667, w47668, w47669, w47670, w47671, w47672, w47673, w47674, w47675, w47676, w47677, w47678, w47679, w47680, w47681, w47682, w47683, w47684, w47685, w47686, w47687, w47688, w47689, w47690, w47691, w47692, w47693, w47694, w47695, w47696, w47697, w47698, w47699, w47700, w47701, w47702, w47703, w47704, w47705, w47706, w47707, w47708, w47709, w47710, w47711, w47712, w47713, w47714, w47715, w47716, w47717, w47718, w47719, w47720, w47721, w47722, w47723, w47724, w47725, w47726, w47727, w47728, w47729, w47730, w47731, w47732, w47733, w47734, w47735, w47736, w47737, w47738, w47739, w47740, w47741, w47742, w47743, w47744, w47745, w47746, w47747, w47748, w47749, w47750, w47751, w47752, w47753, w47754, w47755, w47756, w47757, w47758, w47759, w47760, w47761, w47762, w47763, w47764, w47765, w47766, w47767, w47768, w47769, w47770, w47771, w47772, w47773, w47774, w47775, w47776, w47777, w47778, w47779, w47780, w47781, w47782, w47783, w47784, w47785, w47786, w47787, w47788, w47789, w47790, w47791, w47792, w47793, w47794, w47795, w47796, w47797, w47798, w47799, w47800, w47801, w47802, w47803, w47804, w47805, w47806, w47807, w47808, w47809, w47810, w47811, w47812, w47813, w47814, w47815, w47816, w47817, w47818, w47819, w47820, w47821, w47822, w47823, w47824, w47825, w47826, w47827, w47828, w47829, w47830, w47831, w47832, w47833, w47834, w47835, w47836, w47837, w47838, w47839, w47840, w47841, w47842, w47843, w47844, w47845, w47846, w47847, w47848, w47849, w47850, w47851, w47852, w47853, w47854, w47855, w47856, w47857, w47858, w47859, w47860, w47861, w47862, w47863, w47864, w47865, w47866, w47867, w47868, w47869, w47870, w47871, w47872, w47873, w47874, w47875, w47876, w47877, w47878, w47879, w47880, w47881, w47882, w47883, w47884, w47885, w47886, w47887, w47888, w47889, w47890, w47891, w47892, w47893, w47894, w47895, w47896, w47897, w47898, w47899, w47900, w47901, w47902, w47903, w47904, w47905, w47906, w47907, w47908, w47909, w47910, w47911, w47912, w47913, w47914, w47915, w47916, w47917, w47918, w47919, w47920, w47921, w47922, w47923, w47924, w47925, w47926, w47927, w47928, w47929, w47930, w47931, w47932, w47933, w47934, w47935, w47936, w47937, w47938, w47939, w47940, w47941, w47942, w47943, w47944, w47945, w47946, w47947, w47948, w47949, w47950, w47951, w47952, w47953, w47954, w47955, w47956, w47957, w47958, w47959, w47960, w47961, w47962, w47963, w47964, w47965, w47966, w47967, w47968, w47969, w47970, w47971, w47972, w47973, w47974, w47975, w47976, w47977, w47978, w47979, w47980, w47981, w47982, w47983, w47984, w47985, w47986, w47987, w47988, w47989, w47990, w47991, w47992, w47993, w47994, w47995, w47996, w47997, w47998, w47999, w48000, w48001, w48002, w48003, w48004, w48005, w48006, w48007, w48008, w48009, w48010, w48011, w48012, w48013, w48014, w48015, w48016, w48017, w48018, w48019, w48020, w48021, w48022, w48023, w48024, w48025, w48026, w48027, w48028, w48029, w48030, w48031, w48032, w48033, w48034, w48035, w48036, w48037, w48038, w48039, w48040, w48041, w48042, w48043, w48044, w48045, w48046, w48047, w48048, w48049, w48050, w48051, w48052, w48053, w48054, w48055, w48056, w48057, w48058, w48059, w48060, w48061, w48062, w48063, w48064, w48065, w48066, w48067, w48068, w48069, w48070, w48071, w48072, w48073, w48074, w48075, w48076, w48077, w48078, w48079, w48080, w48081, w48082, w48083, w48084, w48085, w48086, w48087, w48088, w48089, w48090, w48091, w48092, w48093, w48094, w48095, w48096, w48097, w48098, w48099, w48100, w48101, w48102, w48103, w48104, w48105, w48106, w48107, w48108, w48109, w48110, w48111, w48112, w48113, w48114, w48115, w48116, w48117, w48118, w48119, w48120, w48121, w48122, w48123, w48124, w48125, w48126, w48127, w48128, w48129, w48130, w48131, w48132, w48133, w48134, w48135, w48136, w48137, w48138, w48139, w48140, w48141, w48142, w48143, w48144, w48145, w48146, w48147, w48148, w48149, w48150, w48151, w48152, w48153, w48154, w48155, w48156, w48157, w48158, w48159, w48160, w48161, w48162, w48163, w48164, w48165, w48166, w48167, w48168, w48169, w48170, w48171, w48172, w48173, w48174, w48175, w48176, w48177, w48178, w48179, w48180, w48181, w48182, w48183, w48184, w48185, w48186, w48187, w48188, w48189, w48190, w48191, w48192, w48193, w48194, w48195, w48196, w48197, w48198, w48199, w48200, w48201, w48202, w48203, w48204, w48205, w48206, w48207, w48208, w48209, w48210, w48211, w48212, w48213, w48214, w48215, w48216, w48217, w48218, w48219, w48220, w48221, w48222, w48223, w48224, w48225, w48226, w48227, w48228, w48229, w48230, w48231, w48232, w48233, w48234, w48235, w48236, w48237, w48238, w48239, w48240, w48241, w48242, w48243, w48244, w48245, w48246, w48247, w48248, w48249, w48250, w48251, w48252, w48253, w48254, w48255, w48256, w48257, w48258, w48259, w48260, w48261, w48262, w48263, w48264, w48265, w48266, w48267, w48268, w48269, w48270, w48271, w48272, w48273, w48274, w48275, w48276, w48277, w48278, w48279, w48280, w48281, w48282, w48283, w48284, w48285, w48286, w48287, w48288, w48289, w48290, w48291, w48292, w48293, w48294, w48295, w48296, w48297, w48298, w48299, w48300, w48301, w48302, w48303, w48304, w48305, w48306, w48307, w48308, w48309, w48310, w48311, w48312, w48313, w48314, w48315, w48316, w48317, w48318, w48319, w48320, w48321, w48322, w48323, w48324, w48325, w48326, w48327, w48328, w48329, w48330, w48331, w48332, w48333, w48334, w48335, w48336, w48337, w48338, w48339, w48340, w48341, w48342, w48343, w48344, w48345, w48346, w48347, w48348, w48349, w48350, w48351, w48352, w48353, w48354, w48355, w48356, w48357, w48358, w48359, w48360, w48361, w48362, w48363, w48364, w48365, w48366, w48367, w48368, w48369, w48370, w48371, w48372, w48373, w48374, w48375, w48376, w48377, w48378, w48379, w48380, w48381, w48382, w48383, w48384, w48385, w48386, w48387, w48388, w48389, w48390, w48391, w48392, w48393, w48394, w48395, w48396, w48397, w48398, w48399, w48400, w48401, w48402, w48403, w48404, w48405, w48406, w48407, w48408, w48409, w48410, w48411, w48412, w48413, w48414, w48415, w48416, w48417, w48418, w48419, w48420, w48421, w48422, w48423, w48424, w48425, w48426, w48427, w48428, w48429, w48430, w48431, w48432, w48433, w48434, w48435, w48436, w48437, w48438, w48439, w48440, w48441, w48442, w48443, w48444, w48445, w48446, w48447, w48448, w48449, w48450, w48451, w48452, w48453, w48454, w48455, w48456, w48457, w48458, w48459, w48460, w48461, w48462, w48463, w48464, w48465, w48466, w48467, w48468, w48469, w48470, w48471, w48472, w48473, w48474, w48475, w48476, w48477, w48478, w48479, w48480, w48481, w48482, w48483, w48484, w48485, w48486, w48487, w48488, w48489, w48490, w48491, w48492, w48493, w48494, w48495, w48496, w48497, w48498, w48499, w48500, w48501, w48502, w48503, w48504, w48505, w48506, w48507, w48508, w48509, w48510, w48511, w48512, w48513, w48514, w48515, w48516, w48517, w48518, w48519, w48520, w48521, w48522, w48523, w48524, w48525, w48526, w48527, w48528, w48529, w48530, w48531, w48532, w48533, w48534, w48535, w48536, w48537, w48538, w48539, w48540, w48541, w48542, w48543, w48544, w48545, w48546, w48547, w48548, w48549, w48550, w48551, w48552, w48553, w48554, w48555, w48556, w48557, w48558, w48559, w48560, w48561, w48562, w48563, w48564, w48565, w48566, w48567, w48568, w48569, w48570, w48571, w48572, w48573, w48574, w48575, w48576, w48577, w48578, w48579, w48580, w48581, w48582, w48583, w48584, w48585, w48586, w48587, w48588, w48589, w48590, w48591, w48592, w48593, w48594, w48595, w48596, w48597, w48598, w48599, w48600, w48601, w48602, w48603, w48604, w48605, w48606, w48607, w48608, w48609, w48610, w48611, w48612, w48613, w48614, w48615, w48616, w48617, w48618, w48619, w48620, w48621, w48622, w48623, w48624, w48625, w48626, w48627, w48628, w48629, w48630, w48631, w48632, w48633, w48634, w48635, w48636, w48637, w48638, w48639, w48640, w48641, w48642, w48643, w48644, w48645, w48646, w48647, w48648, w48649, w48650, w48651, w48652, w48653, w48654, w48655, w48656, w48657, w48658, w48659, w48660, w48661, w48662, w48663, w48664, w48665, w48666, w48667, w48668, w48669, w48670, w48671, w48672, w48673, w48674, w48675, w48676, w48677, w48678, w48679, w48680, w48681, w48682, w48683, w48684, w48685, w48686, w48687, w48688, w48689, w48690, w48691, w48692, w48693, w48694, w48695, w48696, w48697, w48698, w48699, w48700, w48701, w48702, w48703, w48704, w48705, w48706, w48707, w48708, w48709, w48710, w48711, w48712, w48713, w48714, w48715, w48716, w48717, w48718, w48719, w48720, w48721, w48722, w48723, w48724, w48725, w48726, w48727, w48728, w48729, w48730, w48731, w48732, w48733, w48734, w48735, w48736, w48737, w48738, w48739, w48740, w48741, w48742, w48743, w48744, w48745, w48746, w48747, w48748, w48749, w48750, w48751, w48752, w48753, w48754, w48755, w48756, w48757, w48758, w48759, w48760, w48761, w48762, w48763, w48764, w48765, w48766, w48767, w48768, w48769, w48770, w48771, w48772, w48773, w48774, w48775, w48776, w48777, w48778, w48779, w48780, w48781, w48782, w48783, w48784, w48785, w48786, w48787, w48788, w48789, w48790, w48791, w48792, w48793, w48794, w48795, w48796, w48797, w48798, w48799, w48800, w48801, w48802, w48803, w48804, w48805, w48806, w48807, w48808, w48809, w48810, w48811, w48812, w48813, w48814, w48815, w48816, w48817, w48818, w48819, w48820, w48821, w48822, w48823, w48824, w48825, w48826, w48827, w48828, w48829, w48830, w48831, w48832, w48833, w48834, w48835, w48836, w48837, w48838, w48839, w48840, w48841, w48842, w48843, w48844, w48845, w48846, w48847, w48848, w48849, w48850, w48851, w48852, w48853, w48854, w48855, w48856, w48857, w48858, w48859, w48860, w48861, w48862, w48863, w48864, w48865, w48866, w48867, w48868, w48869, w48870, w48871, w48872, w48873, w48874, w48875, w48876, w48877, w48878, w48879, w48880, w48881, w48882, w48883, w48884, w48885, w48886, w48887, w48888, w48889, w48890, w48891, w48892, w48893, w48894, w48895, w48896, w48897, w48898, w48899, w48900, w48901, w48902, w48903, w48904, w48905, w48906, w48907, w48908, w48909, w48910, w48911, w48912, w48913, w48914, w48915, w48916, w48917, w48918, w48919, w48920, w48921, w48922, w48923, w48924, w48925, w48926, w48927, w48928, w48929, w48930, w48931, w48932, w48933, w48934, w48935, w48936, w48937, w48938, w48939, w48940, w48941, w48942, w48943, w48944, w48945, w48946, w48947, w48948, w48949, w48950, w48951, w48952, w48953, w48954, w48955, w48956, w48957, w48958, w48959, w48960, w48961, w48962, w48963, w48964, w48965, w48966, w48967, w48968, w48969, w48970, w48971, w48972, w48973, w48974, w48975, w48976, w48977, w48978, w48979, w48980, w48981, w48982, w48983, w48984, w48985, w48986, w48987, w48988, w48989, w48990, w48991, w48992, w48993, w48994, w48995, w48996, w48997, w48998, w48999, w49000, w49001, w49002, w49003, w49004, w49005, w49006, w49007, w49008, w49009, w49010, w49011, w49012, w49013, w49014, w49015, w49016, w49017, w49018, w49019, w49020, w49021, w49022, w49023, w49024, w49025, w49026, w49027, w49028, w49029, w49030, w49031, w49032, w49033, w49034, w49035, w49036, w49037, w49038, w49039, w49040, w49041, w49042, w49043, w49044, w49045, w49046, w49047, w49048, w49049, w49050, w49051, w49052, w49053, w49054, w49055, w49056, w49057, w49058, w49059, w49060, w49061, w49062, w49063, w49064, w49065, w49066, w49067, w49068, w49069, w49070, w49071, w49072, w49073, w49074, w49075, w49076, w49077, w49078, w49079, w49080, w49081, w49082, w49083, w49084, w49085, w49086, w49087, w49088, w49089, w49090, w49091, w49092, w49093, w49094, w49095, w49096, w49097, w49098, w49099, w49100, w49101, w49102, w49103, w49104, w49105, w49106, w49107, w49108, w49109, w49110, w49111, w49112, w49113, w49114, w49115, w49116, w49117, w49118, w49119, w49120, w49121, w49122, w49123, w49124, w49125, w49126, w49127, w49128, w49129, w49130, w49131, w49132, w49133, w49134, w49135, w49136, w49137, w49138, w49139, w49140, w49141, w49142, w49143, w49144, w49145, w49146, w49147, w49148, w49149, w49150, w49151, w49152, w49153, w49154, w49155, w49156, w49157, w49158, w49159, w49160, w49161, w49162, w49163, w49164, w49165, w49166, w49167, w49168, w49169, w49170, w49171, w49172, w49173, w49174, w49175, w49176, w49177, w49178, w49179, w49180, w49181, w49182, w49183, w49184, w49185, w49186, w49187, w49188, w49189, w49190, w49191, w49192, w49193, w49194, w49195, w49196, w49197, w49198, w49199, w49200, w49201, w49202, w49203, w49204, w49205, w49206, w49207, w49208, w49209, w49210, w49211, w49212, w49213, w49214, w49215, w49216, w49217, w49218, w49219, w49220, w49221, w49222, w49223, w49224, w49225, w49226, w49227, w49228, w49229, w49230, w49231, w49232, w49233, w49234, w49235, w49236, w49237, w49238, w49239, w49240, w49241, w49242, w49243, w49244, w49245, w49246, w49247, w49248, w49249, w49250, w49251, w49252, w49253, w49254, w49255, w49256, w49257, w49258, w49259, w49260, w49261, w49262, w49263, w49264, w49265, w49266, w49267, w49268, w49269, w49270, w49271, w49272, w49273, w49274, w49275, w49276, w49277, w49278, w49279, w49280, w49281, w49282, w49283, w49284, w49285, w49286, w49287, w49288, w49289, w49290, w49291, w49292, w49293, w49294, w49295, w49296, w49297, w49298, w49299, w49300, w49301, w49302, w49303, w49304, w49305, w49306, w49307, w49308, w49309, w49310, w49311, w49312, w49313, w49314, w49315, w49316, w49317, w49318, w49319, w49320, w49321, w49322, w49323, w49324, w49325, w49326, w49327, w49328, w49329, w49330, w49331, w49332, w49333, w49334, w49335, w49336, w49337, w49338, w49339, w49340, w49341, w49342, w49343, w49344, w49345, w49346, w49347, w49348, w49349, w49350, w49351, w49352, w49353, w49354, w49355, w49356, w49357, w49358, w49359, w49360, w49361, w49362, w49363, w49364, w49365, w49366, w49367, w49368, w49369, w49370, w49371, w49372, w49373, w49374, w49375, w49376, w49377, w49378, w49379, w49380, w49381, w49382, w49383, w49384, w49385, w49386, w49387, w49388, w49389, w49390, w49391, w49392, w49393, w49394, w49395, w49396, w49397, w49398, w49399, w49400, w49401, w49402, w49403, w49404, w49405, w49406, w49407, w49408, w49409, w49410, w49411, w49412, w49413, w49414, w49415, w49416, w49417, w49418, w49419, w49420, w49421, w49422, w49423, w49424, w49425, w49426, w49427, w49428, w49429, w49430, w49431, w49432, w49433, w49434, w49435, w49436, w49437, w49438, w49439, w49440, w49441, w49442, w49443, w49444, w49445, w49446, w49447, w49448, w49449, w49450, w49451, w49452, w49453, w49454, w49455, w49456, w49457, w49458, w49459, w49460, w49461, w49462, w49463, w49464, w49465, w49466, w49467, w49468, w49469, w49470, w49471, w49472, w49473, w49474, w49475, w49476, w49477, w49478, w49479, w49480, w49481, w49482, w49483, w49484, w49485, w49486, w49487, w49488, w49489, w49490, w49491, w49492, w49493, w49494, w49495, w49496, w49497, w49498, w49499, w49500, w49501, w49502, w49503, w49504, w49505, w49506, w49507, w49508, w49509, w49510, w49511, w49512, w49513, w49514, w49515, w49516, w49517, w49518, w49519, w49520, w49521, w49522, w49523, w49524, w49525, w49526, w49527, w49528, w49529, w49530, w49531, w49532, w49533, w49534, w49535, w49536, w49537, w49538, w49539, w49540, w49541, w49542, w49543, w49544, w49545, w49546, w49547, w49548, w49549, w49550, w49551, w49552, w49553, w49554, w49555, w49556, w49557, w49558, w49559, w49560, w49561, w49562, w49563, w49564, w49565, w49566, w49567, w49568, w49569, w49570, w49571, w49572, w49573, w49574, w49575, w49576, w49577, w49578, w49579, w49580, w49581, w49582, w49583, w49584, w49585, w49586, w49587, w49588, w49589, w49590, w49591, w49592, w49593, w49594, w49595, w49596, w49597, w49598, w49599, w49600, w49601, w49602, w49603, w49604, w49605, w49606, w49607, w49608, w49609, w49610, w49611, w49612, w49613, w49614, w49615, w49616, w49617, w49618, w49619, w49620, w49621, w49622, w49623, w49624, w49625, w49626, w49627, w49628, w49629, w49630, w49631, w49632, w49633, w49634, w49635, w49636, w49637, w49638, w49639, w49640, w49641, w49642, w49643, w49644, w49645, w49646, w49647, w49648, w49649, w49650, w49651, w49652, w49653, w49654, w49655, w49656, w49657, w49658, w49659, w49660, w49661, w49662, w49663, w49664, w49665, w49666, w49667, w49668, w49669, w49670, w49671, w49672, w49673, w49674, w49675, w49676, w49677, w49678, w49679, w49680, w49681, w49682, w49683, w49684, w49685, w49686, w49687, w49688, w49689, w49690, w49691, w49692, w49693, w49694, w49695, w49696, w49697, w49698, w49699, w49700, w49701, w49702, w49703, w49704, w49705, w49706, w49707, w49708, w49709, w49710, w49711, w49712, w49713, w49714, w49715, w49716, w49717, w49718, w49719, w49720, w49721, w49722, w49723, w49724, w49725, w49726, w49727, w49728, w49729, w49730, w49731, w49732, w49733, w49734, w49735, w49736, w49737, w49738, w49739, w49740, w49741, w49742, w49743, w49744, w49745, w49746, w49747, w49748, w49749, w49750, w49751, w49752, w49753, w49754, w49755, w49756, w49757, w49758, w49759, w49760, w49761, w49762, w49763, w49764, w49765, w49766, w49767, w49768, w49769, w49770, w49771, w49772, w49773, w49774, w49775, w49776, w49777, w49778, w49779, w49780, w49781, w49782, w49783, w49784, w49785, w49786, w49787, w49788, w49789, w49790, w49791, w49792, w49793, w49794, w49795, w49796, w49797, w49798, w49799, w49800, w49801, w49802, w49803, w49804, w49805, w49806, w49807, w49808, w49809, w49810, w49811, w49812, w49813, w49814, w49815, w49816, w49817, w49818, w49819, w49820, w49821, w49822, w49823, w49824, w49825, w49826, w49827, w49828, w49829, w49830, w49831, w49832, w49833, w49834, w49835, w49836, w49837, w49838, w49839, w49840, w49841, w49842, w49843, w49844, w49845, w49846, w49847, w49848, w49849, w49850, w49851, w49852, w49853, w49854, w49855, w49856, w49857, w49858, w49859, w49860, w49861, w49862, w49863, w49864, w49865, w49866, w49867, w49868, w49869, w49870, w49871, w49872, w49873, w49874, w49875, w49876, w49877, w49878, w49879, w49880, w49881, w49882, w49883, w49884, w49885, w49886, w49887, w49888, w49889, w49890, w49891, w49892, w49893, w49894, w49895, w49896, w49897, w49898, w49899, w49900, w49901, w49902, w49903, w49904, w49905, w49906, w49907, w49908, w49909, w49910, w49911, w49912, w49913, w49914, w49915, w49916, w49917, w49918, w49919, w49920, w49921, w49922, w49923, w49924, w49925, w49926, w49927, w49928, w49929, w49930, w49931, w49932, w49933, w49934, w49935, w49936, w49937, w49938, w49939, w49940, w49941, w49942, w49943, w49944, w49945, w49946, w49947, w49948, w49949, w49950, w49951, w49952, w49953, w49954, w49955, w49956, w49957, w49958, w49959, w49960, w49961, w49962, w49963, w49964, w49965, w49966, w49967, w49968, w49969, w49970, w49971, w49972, w49973, w49974, w49975, w49976, w49977, w49978, w49979, w49980, w49981, w49982, w49983, w49984, w49985, w49986, w49987, w49988, w49989, w49990, w49991, w49992, w49993, w49994, w49995, w49996, w49997, w49998, w49999, w50000, w50001, w50002, w50003, w50004, w50005, w50006, w50007, w50008, w50009, w50010, w50011, w50012, w50013, w50014, w50015, w50016, w50017, w50018, w50019, w50020, w50021, w50022, w50023, w50024, w50025, w50026, w50027, w50028, w50029, w50030, w50031, w50032, w50033, w50034, w50035, w50036, w50037, w50038, w50039, w50040, w50041, w50042, w50043, w50044, w50045, w50046, w50047, w50048, w50049, w50050, w50051, w50052, w50053, w50054, w50055, w50056, w50057, w50058, w50059, w50060, w50061, w50062, w50063, w50064, w50065, w50066, w50067, w50068, w50069, w50070, w50071, w50072, w50073, w50074, w50075, w50076, w50077, w50078, w50079, w50080, w50081, w50082, w50083, w50084, w50085, w50086, w50087, w50088, w50089, w50090, w50091, w50092, w50093, w50094, w50095, w50096, w50097, w50098, w50099, w50100, w50101, w50102, w50103, w50104, w50105, w50106, w50107, w50108, w50109, w50110, w50111, w50112, w50113, w50114, w50115, w50116, w50117, w50118, w50119, w50120, w50121, w50122, w50123, w50124, w50125, w50126, w50127, w50128, w50129, w50130, w50131, w50132, w50133, w50134, w50135, w50136, w50137, w50138, w50139, w50140, w50141, w50142, w50143, w50144, w50145, w50146, w50147, w50148, w50149, w50150, w50151, w50152, w50153, w50154, w50155, w50156, w50157, w50158, w50159, w50160, w50161, w50162, w50163, w50164, w50165, w50166, w50167, w50168, w50169, w50170, w50171, w50172, w50173, w50174, w50175, w50176, w50177, w50178, w50179, w50180, w50181, w50182, w50183, w50184, w50185, w50186, w50187, w50188, w50189, w50190, w50191, w50192, w50193, w50194, w50195, w50196, w50197, w50198, w50199, w50200, w50201, w50202, w50203, w50204, w50205, w50206, w50207, w50208, w50209, w50210, w50211, w50212, w50213, w50214, w50215, w50216, w50217, w50218, w50219, w50220, w50221, w50222, w50223, w50224, w50225, w50226, w50227, w50228, w50229, w50230, w50231, w50232, w50233, w50234, w50235, w50236, w50237, w50238, w50239, w50240, w50241, w50242, w50243, w50244, w50245, w50246, w50247, w50248, w50249, w50250, w50251, w50252, w50253, w50254, w50255, w50256, w50257, w50258, w50259, w50260, w50261, w50262, w50263, w50264, w50265, w50266, w50267, w50268, w50269, w50270, w50271, w50272, w50273, w50274, w50275, w50276, w50277, w50278, w50279, w50280, w50281, w50282, w50283, w50284, w50285, w50286, w50287, w50288, w50289, w50290, w50291, w50292, w50293, w50294, w50295, w50296, w50297, w50298, w50299, w50300, w50301, w50302, w50303, w50304, w50305, w50306, w50307, w50308, w50309, w50310, w50311, w50312, w50313, w50314, w50315, w50316, w50317, w50318, w50319, w50320, w50321, w50322, w50323, w50324, w50325, w50326, w50327, w50328, w50329, w50330, w50331, w50332, w50333, w50334, w50335, w50336, w50337, w50338, w50339, w50340, w50341, w50342, w50343, w50344, w50345, w50346, w50347, w50348, w50349, w50350, w50351, w50352, w50353, w50354, w50355, w50356, w50357, w50358, w50359, w50360, w50361, w50362, w50363, w50364, w50365, w50366, w50367, w50368, w50369, w50370, w50371, w50372, w50373, w50374, w50375, w50376, w50377, w50378, w50379, w50380, w50381, w50382, w50383, w50384, w50385, w50386, w50387, w50388, w50389, w50390, w50391, w50392, w50393, w50394, w50395, w50396, w50397, w50398, w50399, w50400, w50401, w50402, w50403, w50404, w50405, w50406, w50407, w50408, w50409, w50410, w50411, w50412, w50413, w50414, w50415, w50416, w50417, w50418, w50419, w50420, w50421, w50422, w50423, w50424, w50425, w50426, w50427, w50428, w50429, w50430, w50431, w50432, w50433, w50434, w50435, w50436, w50437, w50438, w50439, w50440, w50441, w50442, w50443, w50444, w50445, w50446, w50447, w50448, w50449, w50450, w50451, w50452, w50453, w50454, w50455, w50456, w50457, w50458, w50459, w50460, w50461, w50462, w50463, w50464, w50465, w50466, w50467, w50468, w50469, w50470, w50471, w50472, w50473, w50474, w50475, w50476, w50477, w50478, w50479, w50480, w50481, w50482, w50483, w50484, w50485, w50486, w50487, w50488, w50489, w50490, w50491, w50492, w50493, w50494, w50495, w50496, w50497, w50498, w50499, w50500, w50501, w50502, w50503, w50504, w50505, w50506, w50507, w50508, w50509, w50510, w50511, w50512, w50513, w50514, w50515, w50516, w50517, w50518, w50519, w50520, w50521, w50522, w50523, w50524, w50525, w50526, w50527, w50528, w50529, w50530, w50531, w50532, w50533, w50534, w50535, w50536, w50537, w50538, w50539, w50540, w50541, w50542, w50543, w50544, w50545, w50546, w50547, w50548, w50549, w50550, w50551, w50552, w50553, w50554, w50555, w50556, w50557, w50558, w50559, w50560, w50561, w50562, w50563, w50564, w50565, w50566, w50567, w50568, w50569, w50570, w50571, w50572, w50573, w50574, w50575, w50576, w50577, w50578, w50579, w50580, w50581, w50582, w50583, w50584, w50585, w50586, w50587, w50588, w50589, w50590, w50591, w50592, w50593, w50594, w50595, w50596, w50597, w50598, w50599, w50600, w50601, w50602, w50603, w50604, w50605, w50606, w50607, w50608, w50609, w50610, w50611, w50612, w50613, w50614, w50615, w50616, w50617, w50618, w50619, w50620, w50621, w50622, w50623, w50624, w50625, w50626, w50627, w50628, w50629, w50630, w50631, w50632, w50633, w50634, w50635, w50636, w50637, w50638, w50639, w50640, w50641, w50642, w50643, w50644, w50645, w50646, w50647, w50648, w50649, w50650, w50651, w50652, w50653, w50654, w50655, w50656, w50657, w50658, w50659, w50660, w50661, w50662, w50663, w50664, w50665, w50666, w50667, w50668, w50669, w50670, w50671, w50672, w50673, w50674, w50675, w50676, w50677, w50678, w50679, w50680, w50681, w50682, w50683, w50684, w50685, w50686, w50687, w50688, w50689, w50690, w50691, w50692, w50693, w50694, w50695, w50696, w50697, w50698, w50699, w50700, w50701, w50702, w50703, w50704, w50705, w50706, w50707, w50708, w50709, w50710, w50711, w50712, w50713, w50714, w50715, w50716, w50717, w50718, w50719, w50720, w50721, w50722, w50723, w50724, w50725, w50726, w50727, w50728, w50729, w50730, w50731, w50732, w50733, w50734, w50735, w50736, w50737, w50738, w50739, w50740, w50741, w50742, w50743, w50744, w50745, w50746, w50747, w50748, w50749, w50750, w50751, w50752, w50753, w50754, w50755, w50756, w50757, w50758, w50759, w50760, w50761, w50762, w50763, w50764, w50765, w50766, w50767, w50768, w50769, w50770, w50771, w50772, w50773, w50774, w50775, w50776, w50777, w50778, w50779, w50780, w50781, w50782, w50783, w50784, w50785, w50786, w50787, w50788, w50789, w50790, w50791, w50792, w50793, w50794, w50795, w50796, w50797, w50798, w50799, w50800, w50801, w50802, w50803, w50804, w50805, w50806, w50807, w50808, w50809, w50810, w50811, w50812, w50813, w50814, w50815, w50816, w50817, w50818, w50819, w50820, w50821, w50822, w50823, w50824, w50825, w50826, w50827, w50828, w50829, w50830, w50831, w50832, w50833, w50834, w50835, w50836, w50837, w50838, w50839, w50840, w50841, w50842, w50843, w50844, w50845, w50846, w50847, w50848, w50849, w50850, w50851, w50852, w50853, w50854, w50855, w50856, w50857, w50858, w50859, w50860, w50861, w50862, w50863, w50864, w50865, w50866, w50867, w50868, w50869, w50870, w50871, w50872, w50873, w50874, w50875, w50876, w50877, w50878, w50879, w50880, w50881, w50882, w50883, w50884, w50885, w50886, w50887, w50888, w50889, w50890, w50891, w50892, w50893, w50894, w50895, w50896, w50897, w50898, w50899, w50900, w50901, w50902, w50903, w50904, w50905, w50906, w50907, w50908, w50909, w50910, w50911, w50912, w50913, w50914, w50915, w50916, w50917, w50918, w50919, w50920, w50921, w50922, w50923, w50924, w50925, w50926, w50927, w50928, w50929, w50930, w50931, w50932, w50933, w50934, w50935, w50936, w50937, w50938, w50939, w50940, w50941, w50942, w50943, w50944, w50945, w50946, w50947, w50948, w50949, w50950, w50951, w50952, w50953, w50954, w50955, w50956, w50957, w50958, w50959, w50960, w50961, w50962, w50963, w50964, w50965, w50966, w50967, w50968, w50969, w50970, w50971, w50972, w50973, w50974, w50975, w50976, w50977, w50978, w50979, w50980, w50981, w50982, w50983, w50984, w50985, w50986, w50987, w50988, w50989, w50990, w50991, w50992, w50993, w50994, w50995, w50996, w50997, w50998, w50999, w51000, w51001, w51002, w51003, w51004, w51005, w51006, w51007, w51008, w51009, w51010, w51011, w51012, w51013, w51014, w51015, w51016, w51017, w51018, w51019, w51020, w51021, w51022, w51023, w51024, w51025, w51026, w51027, w51028, w51029, w51030, w51031, w51032, w51033, w51034, w51035, w51036, w51037, w51038, w51039, w51040, w51041, w51042, w51043, w51044, w51045, w51046, w51047, w51048, w51049, w51050, w51051, w51052, w51053, w51054, w51055, w51056, w51057, w51058, w51059, w51060, w51061, w51062, w51063, w51064, w51065, w51066, w51067, w51068, w51069, w51070, w51071, w51072, w51073, w51074, w51075, w51076, w51077, w51078, w51079, w51080, w51081, w51082, w51083, w51084, w51085, w51086, w51087, w51088, w51089, w51090, w51091, w51092, w51093, w51094, w51095, w51096, w51097, w51098, w51099, w51100, w51101, w51102, w51103, w51104, w51105, w51106, w51107, w51108, w51109, w51110, w51111, w51112, w51113, w51114, w51115, w51116, w51117, w51118, w51119, w51120, w51121, w51122, w51123, w51124, w51125, w51126, w51127, w51128, w51129, w51130, w51131, w51132, w51133, w51134, w51135, w51136, w51137, w51138, w51139, w51140, w51141, w51142, w51143, w51144, w51145, w51146, w51147, w51148, w51149, w51150, w51151, w51152, w51153, w51154, w51155, w51156, w51157, w51158, w51159, w51160, w51161, w51162, w51163, w51164, w51165, w51166, w51167, w51168, w51169, w51170, w51171, w51172, w51173, w51174, w51175, w51176, w51177, w51178, w51179, w51180, w51181, w51182, w51183, w51184, w51185, w51186, w51187, w51188, w51189, w51190, w51191, w51192, w51193, w51194, w51195, w51196, w51197, w51198, w51199, w51200, w51201, w51202, w51203, w51204, w51205, w51206, w51207, w51208, w51209, w51210, w51211, w51212, w51213, w51214, w51215, w51216, w51217, w51218, w51219, w51220, w51221, w51222, w51223, w51224, w51225, w51226, w51227, w51228, w51229, w51230, w51231, w51232, w51233, w51234, w51235, w51236, w51237, w51238, w51239, w51240, w51241, w51242, w51243, w51244, w51245, w51246, w51247, w51248, w51249, w51250, w51251, w51252, w51253, w51254, w51255, w51256, w51257, w51258, w51259, w51260, w51261, w51262, w51263, w51264, w51265, w51266, w51267, w51268, w51269, w51270, w51271, w51272, w51273, w51274, w51275, w51276, w51277, w51278, w51279, w51280, w51281, w51282, w51283, w51284, w51285, w51286, w51287, w51288, w51289, w51290, w51291, w51292, w51293, w51294, w51295, w51296, w51297, w51298, w51299, w51300, w51301, w51302, w51303, w51304, w51305, w51306, w51307, w51308, w51309, w51310, w51311, w51312, w51313, w51314, w51315, w51316, w51317, w51318, w51319, w51320, w51321, w51322, w51323, w51324, w51325, w51326, w51327, w51328, w51329, w51330, w51331, w51332, w51333, w51334, w51335, w51336, w51337, w51338, w51339, w51340, w51341, w51342, w51343, w51344, w51345, w51346, w51347, w51348, w51349, w51350, w51351, w51352, w51353, w51354, w51355, w51356, w51357, w51358, w51359, w51360, w51361, w51362, w51363, w51364, w51365, w51366, w51367, w51368, w51369, w51370, w51371, w51372, w51373, w51374, w51375, w51376, w51377, w51378, w51379, w51380, w51381, w51382, w51383, w51384, w51385, w51386, w51387, w51388, w51389, w51390, w51391, w51392, w51393, w51394, w51395, w51396, w51397, w51398, w51399, w51400, w51401, w51402, w51403, w51404, w51405, w51406, w51407, w51408, w51409, w51410, w51411, w51412, w51413, w51414, w51415, w51416, w51417, w51418, w51419, w51420, w51421, w51422, w51423, w51424, w51425, w51426, w51427, w51428, w51429, w51430, w51431, w51432, w51433, w51434, w51435, w51436, w51437, w51438, w51439, w51440, w51441, w51442, w51443, w51444, w51445, w51446, w51447, w51448, w51449, w51450, w51451, w51452, w51453, w51454, w51455, w51456, w51457, w51458, w51459, w51460, w51461, w51462, w51463, w51464, w51465, w51466, w51467, w51468, w51469, w51470, w51471, w51472, w51473, w51474, w51475, w51476, w51477, w51478, w51479, w51480, w51481, w51482, w51483, w51484, w51485, w51486, w51487, w51488, w51489, w51490, w51491, w51492, w51493, w51494, w51495, w51496, w51497, w51498, w51499, w51500, w51501, w51502, w51503, w51504, w51505, w51506, w51507, w51508, w51509, w51510, w51511, w51512, w51513, w51514, w51515, w51516, w51517, w51518, w51519, w51520, w51521, w51522, w51523, w51524, w51525, w51526, w51527, w51528, w51529, w51530, w51531, w51532, w51533, w51534, w51535, w51536, w51537, w51538, w51539, w51540, w51541, w51542, w51543, w51544, w51545, w51546, w51547, w51548, w51549, w51550, w51551, w51552, w51553, w51554, w51555, w51556, w51557, w51558, w51559, w51560, w51561, w51562, w51563, w51564, w51565, w51566, w51567, w51568, w51569, w51570, w51571, w51572, w51573, w51574, w51575, w51576, w51577, w51578, w51579, w51580, w51581, w51582, w51583, w51584, w51585, w51586, w51587, w51588, w51589, w51590, w51591, w51592, w51593, w51594, w51595, w51596, w51597, w51598, w51599, w51600, w51601, w51602, w51603, w51604, w51605, w51606, w51607, w51608, w51609, w51610, w51611, w51612, w51613, w51614, w51615, w51616, w51617, w51618, w51619, w51620, w51621, w51622, w51623, w51624, w51625, w51626, w51627, w51628, w51629, w51630, w51631, w51632, w51633, w51634, w51635, w51636, w51637, w51638, w51639, w51640, w51641, w51642, w51643, w51644, w51645, w51646, w51647, w51648, w51649, w51650, w51651, w51652, w51653, w51654, w51655, w51656, w51657, w51658, w51659, w51660, w51661, w51662, w51663, w51664, w51665, w51666, w51667, w51668, w51669, w51670, w51671, w51672, w51673, w51674, w51675, w51676, w51677, w51678, w51679, w51680, w51681, w51682, w51683, w51684, w51685, w51686, w51687, w51688, w51689, w51690, w51691, w51692, w51693, w51694, w51695, w51696, w51697, w51698, w51699, w51700, w51701, w51702, w51703, w51704, w51705, w51706, w51707, w51708, w51709, w51710, w51711, w51712, w51713, w51714, w51715, w51716, w51717, w51718, w51719, w51720, w51721, w51722, w51723, w51724, w51725, w51726, w51727, w51728, w51729, w51730, w51731, w51732, w51733, w51734, w51735, w51736, w51737, w51738, w51739, w51740, w51741, w51742, w51743, w51744, w51745, w51746, w51747, w51748, w51749, w51750, w51751, w51752, w51753, w51754, w51755, w51756, w51757, w51758, w51759, w51760, w51761, w51762, w51763, w51764, w51765, w51766, w51767, w51768, w51769, w51770, w51771, w51772, w51773, w51774, w51775, w51776, w51777, w51778, w51779, w51780, w51781, w51782, w51783, w51784, w51785, w51786, w51787, w51788, w51789, w51790, w51791, w51792, w51793, w51794, w51795, w51796, w51797, w51798, w51799, w51800, w51801, w51802, w51803, w51804, w51805, w51806, w51807, w51808, w51809, w51810, w51811, w51812, w51813, w51814, w51815, w51816, w51817, w51818, w51819, w51820, w51821, w51822, w51823, w51824, w51825, w51826, w51827, w51828, w51829, w51830, w51831, w51832, w51833, w51834, w51835, w51836, w51837, w51838, w51839, w51840, w51841, w51842, w51843, w51844, w51845, w51846, w51847, w51848, w51849, w51850, w51851, w51852, w51853, w51854, w51855, w51856, w51857, w51858, w51859, w51860, w51861, w51862, w51863, w51864, w51865, w51866, w51867, w51868, w51869, w51870, w51871, w51872, w51873, w51874, w51875, w51876, w51877, w51878, w51879, w51880, w51881, w51882, w51883, w51884, w51885, w51886, w51887, w51888, w51889, w51890, w51891, w51892, w51893, w51894, w51895, w51896, w51897, w51898, w51899, w51900, w51901, w51902, w51903, w51904, w51905, w51906, w51907, w51908, w51909, w51910, w51911, w51912, w51913, w51914, w51915, w51916, w51917, w51918, w51919, w51920, w51921, w51922, w51923, w51924, w51925, w51926, w51927, w51928, w51929, w51930, w51931, w51932, w51933, w51934, w51935, w51936, w51937, w51938, w51939, w51940, w51941, w51942, w51943, w51944, w51945, w51946, w51947, w51948, w51949, w51950, w51951, w51952, w51953, w51954, w51955, w51956, w51957, w51958, w51959, w51960, w51961, w51962, w51963, w51964, w51965, w51966, w51967, w51968, w51969, w51970, w51971, w51972, w51973, w51974, w51975, w51976, w51977, w51978, w51979, w51980, w51981, w51982, w51983, w51984, w51985, w51986, w51987, w51988, w51989, w51990, w51991, w51992, w51993, w51994, w51995, w51996, w51997, w51998, w51999, w52000, w52001, w52002, w52003, w52004, w52005, w52006, w52007, w52008, w52009, w52010, w52011, w52012, w52013, w52014, w52015, w52016, w52017, w52018, w52019, w52020, w52021, w52022, w52023, w52024, w52025, w52026, w52027, w52028, w52029, w52030, w52031, w52032, w52033, w52034, w52035, w52036, w52037, w52038, w52039, w52040, w52041, w52042, w52043, w52044, w52045, w52046, w52047, w52048, w52049, w52050, w52051, w52052, w52053, w52054, w52055, w52056, w52057, w52058, w52059, w52060, w52061, w52062, w52063, w52064, w52065, w52066, w52067, w52068, w52069, w52070, w52071, w52072, w52073, w52074, w52075, w52076, w52077, w52078, w52079, w52080, w52081, w52082, w52083, w52084, w52085, w52086, w52087, w52088, w52089, w52090, w52091, w52092, w52093, w52094, w52095, w52096, w52097, w52098, w52099, w52100, w52101, w52102, w52103, w52104, w52105, w52106, w52107, w52108, w52109, w52110, w52111, w52112, w52113, w52114, w52115, w52116, w52117, w52118, w52119, w52120, w52121, w52122, w52123, w52124, w52125, w52126, w52127, w52128, w52129, w52130, w52131, w52132, w52133, w52134, w52135, w52136, w52137, w52138, w52139, w52140, w52141, w52142, w52143, w52144, w52145, w52146, w52147, w52148, w52149, w52150, w52151, w52152, w52153, w52154, w52155, w52156, w52157, w52158, w52159, w52160, w52161, w52162, w52163, w52164, w52165, w52166, w52167, w52168, w52169, w52170, w52171, w52172, w52173, w52174, w52175, w52176, w52177, w52178, w52179, w52180, w52181, w52182, w52183, w52184, w52185, w52186, w52187, w52188, w52189, w52190, w52191, w52192, w52193, w52194, w52195, w52196, w52197, w52198, w52199, w52200, w52201, w52202, w52203, w52204, w52205, w52206, w52207, w52208, w52209, w52210, w52211, w52212, w52213, w52214, w52215, w52216, w52217, w52218, w52219, w52220, w52221, w52222, w52223, w52224, w52225, w52226, w52227, w52228, w52229, w52230, w52231, w52232, w52233, w52234, w52235, w52236, w52237, w52238, w52239, w52240, w52241, w52242, w52243, w52244, w52245, w52246, w52247, w52248, w52249, w52250, w52251, w52252, w52253, w52254, w52255, w52256, w52257, w52258, w52259, w52260, w52261, w52262, w52263, w52264, w52265, w52266, w52267, w52268, w52269, w52270, w52271, w52272, w52273, w52274, w52275, w52276, w52277, w52278, w52279, w52280, w52281, w52282, w52283, w52284, w52285, w52286, w52287, w52288, w52289, w52290, w52291, w52292, w52293, w52294, w52295, w52296, w52297, w52298, w52299, w52300, w52301, w52302, w52303, w52304, w52305, w52306, w52307, w52308, w52309, w52310, w52311, w52312, w52313, w52314, w52315, w52316, w52317, w52318, w52319, w52320, w52321, w52322, w52323, w52324, w52325, w52326, w52327, w52328, w52329, w52330, w52331, w52332, w52333, w52334, w52335, w52336, w52337, w52338, w52339, w52340, w52341, w52342, w52343, w52344, w52345, w52346, w52347, w52348, w52349, w52350, w52351, w52352, w52353, w52354, w52355, w52356, w52357, w52358, w52359, w52360, w52361, w52362, w52363, w52364, w52365, w52366, w52367, w52368, w52369, w52370, w52371, w52372, w52373, w52374, w52375, w52376, w52377, w52378, w52379, w52380, w52381, w52382, w52383, w52384, w52385, w52386, w52387, w52388, w52389, w52390, w52391, w52392, w52393, w52394, w52395, w52396, w52397, w52398, w52399, w52400, w52401, w52402, w52403, w52404, w52405, w52406, w52407, w52408, w52409, w52410, w52411, w52412, w52413, w52414, w52415, w52416, w52417, w52418, w52419, w52420, w52421, w52422, w52423, w52424, w52425, w52426, w52427, w52428, w52429, w52430, w52431, w52432, w52433, w52434, w52435, w52436, w52437, w52438, w52439, w52440, w52441, w52442, w52443, w52444, w52445, w52446, w52447, w52448, w52449, w52450, w52451, w52452, w52453, w52454, w52455, w52456, w52457, w52458, w52459, w52460, w52461, w52462, w52463, w52464, w52465, w52466, w52467, w52468, w52469, w52470, w52471, w52472, w52473, w52474, w52475, w52476, w52477, w52478, w52479, w52480, w52481, w52482, w52483, w52484, w52485, w52486, w52487, w52488, w52489, w52490, w52491, w52492, w52493, w52494, w52495, w52496, w52497, w52498, w52499, w52500, w52501, w52502, w52503, w52504, w52505, w52506, w52507, w52508, w52509, w52510, w52511, w52512, w52513, w52514, w52515, w52516, w52517, w52518, w52519, w52520, w52521, w52522, w52523, w52524, w52525, w52526, w52527, w52528, w52529, w52530, w52531, w52532, w52533, w52534, w52535, w52536, w52537, w52538, w52539, w52540, w52541, w52542, w52543, w52544, w52545, w52546, w52547, w52548, w52549, w52550, w52551, w52552, w52553, w52554, w52555, w52556, w52557, w52558, w52559, w52560, w52561, w52562, w52563, w52564, w52565, w52566, w52567, w52568, w52569, w52570, w52571, w52572, w52573, w52574, w52575, w52576, w52577, w52578, w52579, w52580, w52581, w52582, w52583, w52584, w52585, w52586, w52587, w52588, w52589, w52590, w52591, w52592, w52593, w52594, w52595, w52596, w52597, w52598, w52599, w52600, w52601, w52602, w52603, w52604, w52605, w52606, w52607, w52608, w52609, w52610, w52611, w52612, w52613, w52614, w52615, w52616, w52617, w52618, w52619, w52620, w52621, w52622, w52623, w52624, w52625, w52626, w52627, w52628, w52629, w52630, w52631, w52632, w52633, w52634, w52635, w52636, w52637, w52638, w52639, w52640, w52641, w52642, w52643, w52644, w52645, w52646, w52647, w52648, w52649, w52650, w52651, w52652, w52653, w52654, w52655, w52656, w52657, w52658, w52659, w52660, w52661, w52662, w52663, w52664, w52665, w52666, w52667, w52668, w52669, w52670, w52671, w52672, w52673, w52674, w52675, w52676, w52677, w52678, w52679, w52680, w52681, w52682, w52683, w52684, w52685, w52686, w52687, w52688, w52689, w52690, w52691, w52692, w52693, w52694, w52695, w52696, w52697, w52698, w52699, w52700, w52701, w52702, w52703, w52704, w52705, w52706, w52707, w52708, w52709, w52710, w52711, w52712, w52713, w52714, w52715, w52716, w52717, w52718, w52719, w52720, w52721, w52722, w52723, w52724, w52725, w52726, w52727, w52728, w52729, w52730, w52731, w52732, w52733, w52734, w52735, w52736, w52737, w52738, w52739, w52740, w52741, w52742, w52743, w52744, w52745, w52746, w52747, w52748, w52749, w52750, w52751, w52752, w52753, w52754, w52755, w52756, w52757, w52758, w52759, w52760, w52761, w52762, w52763, w52764, w52765, w52766, w52767, w52768, w52769, w52770, w52771, w52772, w52773, w52774, w52775, w52776, w52777, w52778, w52779, w52780, w52781, w52782, w52783, w52784, w52785, w52786, w52787, w52788, w52789, w52790, w52791, w52792, w52793, w52794, w52795, w52796, w52797, w52798, w52799, w52800, w52801, w52802, w52803, w52804, w52805, w52806, w52807, w52808, w52809, w52810, w52811, w52812, w52813, w52814, w52815, w52816, w52817, w52818, w52819, w52820, w52821, w52822, w52823, w52824, w52825, w52826, w52827, w52828, w52829, w52830, w52831, w52832, w52833, w52834, w52835, w52836, w52837, w52838, w52839, w52840, w52841, w52842, w52843, w52844, w52845, w52846, w52847, w52848, w52849, w52850, w52851, w52852, w52853, w52854, w52855, w52856, w52857, w52858, w52859, w52860, w52861, w52862, w52863, w52864, w52865, w52866, w52867, w52868, w52869, w52870, w52871, w52872, w52873, w52874, w52875, w52876, w52877, w52878, w52879, w52880, w52881, w52882, w52883, w52884, w52885, w52886, w52887, w52888, w52889, w52890, w52891, w52892, w52893, w52894, w52895, w52896, w52897, w52898, w52899, w52900, w52901, w52902, w52903, w52904, w52905, w52906, w52907, w52908, w52909, w52910, w52911, w52912, w52913, w52914, w52915, w52916, w52917, w52918, w52919, w52920, w52921, w52922, w52923, w52924, w52925, w52926, w52927, w52928, w52929, w52930, w52931, w52932, w52933, w52934, w52935, w52936, w52937, w52938, w52939, w52940, w52941, w52942, w52943, w52944, w52945, w52946, w52947, w52948, w52949, w52950, w52951, w52952, w52953, w52954, w52955, w52956, w52957, w52958, w52959, w52960, w52961, w52962, w52963, w52964, w52965, w52966, w52967, w52968, w52969, w52970, w52971, w52972, w52973, w52974, w52975, w52976, w52977, w52978, w52979, w52980, w52981, w52982, w52983, w52984, w52985, w52986, w52987, w52988, w52989, w52990, w52991, w52992, w52993, w52994, w52995, w52996, w52997, w52998, w52999, w53000, w53001, w53002, w53003, w53004, w53005, w53006, w53007, w53008, w53009, w53010, w53011, w53012, w53013, w53014, w53015, w53016, w53017, w53018, w53019, w53020, w53021, w53022, w53023, w53024, w53025, w53026, w53027, w53028, w53029, w53030, w53031, w53032, w53033, w53034, w53035, w53036, w53037, w53038, w53039, w53040, w53041, w53042, w53043, w53044, w53045, w53046, w53047, w53048, w53049, w53050, w53051, w53052, w53053, w53054, w53055, w53056, w53057, w53058, w53059, w53060, w53061, w53062, w53063, w53064, w53065, w53066, w53067, w53068, w53069, w53070, w53071, w53072, w53073, w53074, w53075, w53076, w53077, w53078, w53079, w53080, w53081, w53082, w53083, w53084, w53085, w53086, w53087, w53088, w53089, w53090, w53091, w53092, w53093, w53094, w53095, w53096, w53097, w53098, w53099, w53100, w53101, w53102, w53103, w53104, w53105, w53106, w53107, w53108, w53109, w53110, w53111, w53112, w53113, w53114, w53115, w53116, w53117, w53118, w53119, w53120, w53121, w53122, w53123, w53124, w53125, w53126, w53127, w53128, w53129, w53130, w53131, w53132, w53133, w53134, w53135, w53136, w53137, w53138, w53139, w53140, w53141, w53142, w53143, w53144, w53145, w53146, w53147, w53148, w53149, w53150, w53151, w53152, w53153, w53154, w53155, w53156, w53157, w53158, w53159, w53160, w53161, w53162, w53163, w53164, w53165, w53166, w53167, w53168, w53169, w53170, w53171, w53172, w53173, w53174, w53175, w53176, w53177, w53178, w53179, w53180, w53181, w53182, w53183, w53184, w53185, w53186, w53187, w53188, w53189, w53190, w53191, w53192, w53193, w53194, w53195, w53196, w53197, w53198, w53199, w53200, w53201, w53202, w53203, w53204, w53205, w53206, w53207, w53208, w53209, w53210, w53211, w53212, w53213, w53214, w53215, w53216, w53217, w53218, w53219, w53220, w53221, w53222, w53223, w53224, w53225, w53226, w53227, w53228, w53229, w53230, w53231, w53232, w53233, w53234, w53235, w53236, w53237, w53238, w53239, w53240, w53241, w53242, w53243, w53244, w53245, w53246, w53247, w53248, w53249, w53250, w53251, w53252, w53253, w53254, w53255, w53256, w53257, w53258, w53259, w53260, w53261, w53262, w53263, w53264, w53265, w53266, w53267, w53268, w53269, w53270, w53271, w53272, w53273, w53274, w53275, w53276, w53277, w53278, w53279, w53280, w53281, w53282, w53283, w53284, w53285, w53286, w53287, w53288, w53289, w53290, w53291, w53292, w53293, w53294, w53295, w53296, w53297, w53298, w53299, w53300, w53301, w53302, w53303, w53304, w53305, w53306, w53307, w53308, w53309, w53310, w53311, w53312, w53313, w53314, w53315, w53316, w53317, w53318, w53319, w53320, w53321, w53322, w53323, w53324, w53325, w53326, w53327, w53328, w53329, w53330, w53331, w53332, w53333, w53334, w53335, w53336, w53337, w53338, w53339, w53340, w53341, w53342, w53343, w53344, w53345, w53346, w53347, w53348, w53349, w53350, w53351, w53352, w53353, w53354, w53355, w53356, w53357, w53358, w53359, w53360, w53361, w53362, w53363, w53364, w53365, w53366, w53367, w53368, w53369, w53370, w53371, w53372, w53373, w53374, w53375, w53376, w53377, w53378, w53379, w53380, w53381, w53382, w53383, w53384, w53385, w53386, w53387, w53388, w53389, w53390, w53391, w53392, w53393, w53394, w53395, w53396, w53397, w53398, w53399, w53400, w53401, w53402, w53403, w53404, w53405, w53406, w53407, w53408, w53409, w53410, w53411, w53412, w53413, w53414, w53415, w53416, w53417, w53418, w53419, w53420, w53421, w53422, w53423, w53424, w53425, w53426, w53427, w53428, w53429, w53430, w53431, w53432, w53433, w53434, w53435, w53436, w53437, w53438, w53439, w53440, w53441, w53442, w53443, w53444, w53445, w53446, w53447, w53448, w53449, w53450, w53451, w53452, w53453, w53454, w53455, w53456, w53457, w53458, w53459, w53460, w53461, w53462, w53463, w53464, w53465, w53466, w53467, w53468, w53469, w53470, w53471, w53472, w53473, w53474, w53475, w53476, w53477, w53478, w53479, w53480, w53481, w53482, w53483, w53484, w53485, w53486, w53487, w53488, w53489, w53490, w53491, w53492, w53493, w53494, w53495, w53496, w53497, w53498, w53499, w53500, w53501, w53502, w53503, w53504, w53505, w53506, w53507, w53508, w53509, w53510, w53511, w53512, w53513, w53514, w53515, w53516, w53517, w53518, w53519, w53520, w53521, w53522, w53523, w53524, w53525, w53526, w53527, w53528, w53529, w53530, w53531, w53532, w53533, w53534, w53535, w53536, w53537, w53538, w53539, w53540, w53541, w53542, w53543, w53544, w53545, w53546, w53547, w53548, w53549, w53550, w53551, w53552, w53553, w53554, w53555, w53556, w53557, w53558, w53559, w53560, w53561, w53562, w53563, w53564, w53565, w53566, w53567, w53568, w53569, w53570, w53571, w53572, w53573, w53574, w53575, w53576, w53577, w53578, w53579, w53580, w53581, w53582, w53583, w53584, w53585, w53586, w53587, w53588, w53589, w53590, w53591, w53592, w53593, w53594, w53595, w53596, w53597, w53598, w53599, w53600, w53601, w53602, w53603, w53604, w53605, w53606, w53607, w53608, w53609, w53610, w53611, w53612, w53613, w53614, w53615, w53616, w53617, w53618, w53619, w53620, w53621, w53622, w53623, w53624, w53625, w53626, w53627, w53628, w53629, w53630, w53631, w53632, w53633, w53634, w53635, w53636, w53637, w53638, w53639, w53640, w53641, w53642, w53643, w53644, w53645, w53646, w53647, w53648, w53649, w53650, w53651, w53652, w53653, w53654, w53655, w53656, w53657, w53658, w53659, w53660, w53661, w53662, w53663, w53664, w53665, w53666, w53667, w53668, w53669, w53670, w53671, w53672, w53673, w53674, w53675, w53676, w53677, w53678, w53679, w53680, w53681, w53682, w53683, w53684, w53685, w53686, w53687, w53688, w53689, w53690, w53691, w53692, w53693, w53694, w53695, w53696, w53697, w53698, w53699, w53700, w53701, w53702, w53703, w53704, w53705, w53706, w53707, w53708, w53709, w53710, w53711, w53712, w53713, w53714, w53715, w53716, w53717, w53718, w53719, w53720, w53721, w53722, w53723, w53724, w53725, w53726, w53727, w53728, w53729, w53730, w53731, w53732, w53733, w53734, w53735, w53736, w53737, w53738, w53739, w53740, w53741, w53742, w53743, w53744, w53745, w53746, w53747, w53748, w53749, w53750, w53751, w53752, w53753, w53754, w53755, w53756, w53757, w53758, w53759, w53760, w53761, w53762, w53763, w53764, w53765, w53766, w53767, w53768, w53769, w53770, w53771, w53772, w53773, w53774, w53775, w53776, w53777, w53778, w53779, w53780, w53781, w53782, w53783, w53784, w53785, w53786, w53787, w53788, w53789, w53790, w53791, w53792, w53793, w53794, w53795, w53796, w53797, w53798, w53799, w53800, w53801, w53802, w53803, w53804, w53805, w53806, w53807, w53808, w53809, w53810, w53811, w53812, w53813, w53814, w53815, w53816, w53817, w53818, w53819, w53820, w53821, w53822, w53823, w53824, w53825, w53826, w53827, w53828, w53829, w53830, w53831, w53832, w53833, w53834, w53835, w53836, w53837, w53838, w53839, w53840, w53841, w53842, w53843, w53844, w53845, w53846, w53847, w53848, w53849, w53850, w53851, w53852, w53853, w53854, w53855, w53856, w53857, w53858, w53859, w53860, w53861, w53862, w53863, w53864, w53865, w53866, w53867, w53868, w53869, w53870, w53871, w53872, w53873, w53874, w53875, w53876, w53877, w53878, w53879, w53880, w53881, w53882, w53883, w53884, w53885, w53886, w53887, w53888, w53889, w53890, w53891, w53892, w53893, w53894, w53895, w53896, w53897, w53898, w53899, w53900, w53901, w53902, w53903, w53904, w53905, w53906, w53907, w53908, w53909, w53910, w53911, w53912, w53913, w53914, w53915, w53916, w53917, w53918, w53919, w53920, w53921, w53922, w53923, w53924, w53925, w53926, w53927, w53928, w53929, w53930, w53931, w53932, w53933, w53934, w53935, w53936, w53937, w53938, w53939, w53940, w53941, w53942, w53943, w53944, w53945, w53946, w53947, w53948, w53949, w53950, w53951, w53952, w53953, w53954, w53955, w53956, w53957, w53958, w53959, w53960, w53961, w53962, w53963, w53964, w53965, w53966, w53967, w53968, w53969, w53970, w53971, w53972, w53973, w53974, w53975, w53976, w53977, w53978, w53979, w53980, w53981, w53982, w53983, w53984, w53985, w53986, w53987, w53988, w53989, w53990, w53991, w53992, w53993, w53994, w53995, w53996, w53997, w53998, w53999, w54000, w54001, w54002, w54003, w54004, w54005, w54006, w54007, w54008, w54009, w54010, w54011, w54012, w54013, w54014, w54015, w54016, w54017, w54018, w54019, w54020, w54021, w54022, w54023, w54024, w54025, w54026, w54027, w54028, w54029, w54030, w54031, w54032, w54033, w54034, w54035, w54036, w54037, w54038, w54039, w54040, w54041, w54042, w54043, w54044, w54045, w54046, w54047, w54048, w54049, w54050, w54051, w54052, w54053, w54054, w54055, w54056, w54057, w54058, w54059, w54060, w54061, w54062, w54063, w54064, w54065, w54066, w54067, w54068, w54069, w54070, w54071, w54072, w54073, w54074, w54075, w54076, w54077, w54078, w54079, w54080, w54081, w54082, w54083, w54084, w54085, w54086, w54087, w54088, w54089, w54090, w54091, w54092, w54093, w54094, w54095, w54096, w54097, w54098, w54099, w54100, w54101, w54102, w54103, w54104, w54105, w54106, w54107, w54108, w54109, w54110, w54111, w54112, w54113, w54114, w54115, w54116, w54117, w54118, w54119, w54120, w54121, w54122, w54123, w54124, w54125, w54126, w54127, w54128, w54129, w54130, w54131, w54132, w54133, w54134, w54135, w54136, w54137, w54138, w54139, w54140, w54141, w54142, w54143, w54144, w54145, w54146, w54147, w54148, w54149, w54150, w54151, w54152, w54153, w54154, w54155, w54156, w54157, w54158, w54159, w54160, w54161, w54162, w54163, w54164, w54165, w54166, w54167, w54168, w54169, w54170, w54171, w54172, w54173, w54174, w54175, w54176, w54177, w54178, w54179, w54180, w54181, w54182, w54183, w54184, w54185, w54186, w54187, w54188, w54189, w54190, w54191, w54192, w54193, w54194, w54195, w54196, w54197, w54198, w54199, w54200, w54201, w54202, w54203, w54204, w54205, w54206, w54207, w54208, w54209, w54210, w54211, w54212, w54213, w54214, w54215, w54216, w54217, w54218, w54219, w54220, w54221, w54222, w54223, w54224, w54225, w54226, w54227, w54228, w54229, w54230, w54231, w54232, w54233, w54234, w54235, w54236, w54237, w54238, w54239, w54240, w54241, w54242, w54243, w54244, w54245, w54246, w54247, w54248, w54249, w54250, w54251, w54252, w54253, w54254, w54255, w54256, w54257, w54258, w54259, w54260, w54261, w54262, w54263, w54264, w54265, w54266, w54267, w54268, w54269, w54270, w54271, w54272, w54273, w54274, w54275, w54276, w54277, w54278, w54279, w54280, w54281, w54282, w54283, w54284, w54285, w54286, w54287, w54288, w54289, w54290, w54291, w54292, w54293, w54294, w54295, w54296, w54297, w54298, w54299, w54300, w54301, w54302, w54303, w54304, w54305, w54306, w54307, w54308, w54309, w54310, w54311, w54312, w54313, w54314, w54315, w54316, w54317, w54318, w54319, w54320, w54321, w54322, w54323, w54324, w54325, w54326, w54327, w54328, w54329, w54330, w54331, w54332, w54333, w54334, w54335, w54336, w54337, w54338, w54339, w54340, w54341, w54342, w54343, w54344, w54345, w54346, w54347, w54348, w54349, w54350, w54351, w54352, w54353, w54354, w54355, w54356, w54357, w54358, w54359, w54360, w54361, w54362, w54363, w54364, w54365, w54366, w54367, w54368, w54369, w54370, w54371, w54372, w54373, w54374, w54375, w54376, w54377, w54378, w54379, w54380, w54381, w54382, w54383, w54384, w54385, w54386, w54387, w54388, w54389, w54390, w54391, w54392, w54393, w54394, w54395, w54396, w54397, w54398, w54399, w54400, w54401, w54402, w54403, w54404, w54405, w54406, w54407, w54408, w54409, w54410, w54411, w54412, w54413, w54414, w54415, w54416, w54417, w54418, w54419, w54420, w54421, w54422, w54423, w54424, w54425, w54426, w54427, w54428, w54429, w54430, w54431, w54432, w54433, w54434, w54435, w54436, w54437, w54438, w54439, w54440, w54441, w54442, w54443, w54444, w54445, w54446, w54447, w54448, w54449, w54450, w54451, w54452, w54453, w54454, w54455, w54456, w54457, w54458, w54459, w54460, w54461, w54462, w54463, w54464, w54465, w54466, w54467, w54468, w54469, w54470, w54471, w54472, w54473, w54474, w54475, w54476, w54477, w54478, w54479, w54480, w54481, w54482, w54483, w54484, w54485, w54486, w54487, w54488, w54489, w54490, w54491, w54492, w54493, w54494, w54495, w54496, w54497, w54498, w54499, w54500, w54501, w54502, w54503, w54504, w54505, w54506, w54507, w54508, w54509, w54510, w54511, w54512, w54513, w54514, w54515, w54516, w54517, w54518, w54519, w54520, w54521, w54522, w54523, w54524, w54525, w54526, w54527, w54528, w54529, w54530, w54531, w54532, w54533, w54534, w54535, w54536, w54537, w54538, w54539, w54540, w54541, w54542, w54543, w54544, w54545, w54546, w54547, w54548, w54549, w54550, w54551, w54552, w54553, w54554, w54555, w54556, w54557, w54558, w54559, w54560, w54561, w54562, w54563, w54564, w54565, w54566, w54567, w54568, w54569, w54570, w54571, w54572, w54573, w54574, w54575, w54576, w54577, w54578, w54579, w54580, w54581, w54582, w54583, w54584, w54585, w54586, w54587, w54588, w54589, w54590, w54591, w54592, w54593, w54594, w54595, w54596, w54597, w54598, w54599, w54600, w54601, w54602, w54603, w54604, w54605, w54606, w54607, w54608, w54609, w54610, w54611, w54612, w54613, w54614, w54615, w54616, w54617, w54618, w54619, w54620, w54621, w54622, w54623, w54624, w54625, w54626, w54627, w54628, w54629, w54630, w54631, w54632, w54633, w54634, w54635, w54636, w54637, w54638, w54639, w54640, w54641, w54642, w54643, w54644, w54645, w54646, w54647, w54648, w54649, w54650, w54651, w54652, w54653, w54654, w54655, w54656, w54657, w54658, w54659, w54660, w54661, w54662, w54663, w54664, w54665, w54666, w54667, w54668, w54669, w54670, w54671, w54672, w54673, w54674, w54675, w54676, w54677, w54678, w54679, w54680, w54681, w54682, w54683, w54684, w54685, w54686, w54687, w54688, w54689, w54690, w54691, w54692, w54693, w54694, w54695, w54696, w54697, w54698, w54699, w54700, w54701, w54702, w54703, w54704, w54705, w54706, w54707, w54708, w54709, w54710, w54711, w54712, w54713, w54714, w54715, w54716, w54717, w54718, w54719, w54720, w54721, w54722, w54723, w54724, w54725, w54726, w54727, w54728, w54729, w54730, w54731, w54732, w54733, w54734, w54735, w54736, w54737, w54738, w54739, w54740, w54741, w54742, w54743, w54744, w54745, w54746, w54747, w54748, w54749, w54750, w54751, w54752, w54753, w54754, w54755, w54756, w54757, w54758, w54759, w54760, w54761, w54762, w54763, w54764, w54765, w54766, w54767, w54768, w54769, w54770, w54771, w54772, w54773, w54774, w54775, w54776, w54777, w54778, w54779, w54780, w54781, w54782, w54783, w54784, w54785, w54786, w54787, w54788, w54789, w54790, w54791, w54792, w54793, w54794, w54795, w54796, w54797, w54798, w54799, w54800, w54801, w54802, w54803, w54804, w54805, w54806, w54807, w54808, w54809, w54810, w54811, w54812, w54813, w54814, w54815, w54816, w54817, w54818, w54819, w54820, w54821, w54822, w54823, w54824, w54825, w54826, w54827, w54828, w54829, w54830, w54831, w54832, w54833, w54834, w54835, w54836, w54837, w54838, w54839, w54840, w54841, w54842, w54843, w54844, w54845, w54846, w54847, w54848, w54849, w54850, w54851, w54852, w54853, w54854, w54855, w54856, w54857, w54858, w54859, w54860, w54861, w54862, w54863, w54864, w54865, w54866, w54867, w54868, w54869, w54870, w54871, w54872, w54873, w54874, w54875, w54876, w54877, w54878, w54879, w54880, w54881, w54882, w54883, w54884, w54885, w54886, w54887, w54888, w54889, w54890, w54891, w54892, w54893, w54894, w54895, w54896, w54897, w54898, w54899, w54900, w54901, w54902, w54903, w54904, w54905, w54906, w54907, w54908, w54909, w54910, w54911, w54912, w54913, w54914, w54915, w54916, w54917, w54918, w54919, w54920, w54921, w54922, w54923, w54924, w54925, w54926, w54927, w54928, w54929, w54930, w54931, w54932, w54933, w54934, w54935, w54936, w54937, w54938, w54939, w54940, w54941, w54942, w54943, w54944, w54945, w54946, w54947, w54948, w54949, w54950, w54951, w54952, w54953, w54954, w54955, w54956, w54957, w54958, w54959, w54960, w54961, w54962, w54963, w54964, w54965, w54966, w54967, w54968, w54969, w54970, w54971, w54972, w54973, w54974, w54975, w54976, w54977, w54978, w54979, w54980, w54981, w54982, w54983, w54984, w54985, w54986, w54987, w54988, w54989, w54990, w54991, w54992, w54993, w54994, w54995, w54996, w54997, w54998, w54999, w55000, w55001, w55002, w55003, w55004, w55005, w55006, w55007, w55008, w55009, w55010, w55011, w55012, w55013, w55014, w55015, w55016, w55017, w55018, w55019, w55020, w55021, w55022, w55023, w55024, w55025, w55026, w55027, w55028, w55029, w55030, w55031, w55032, w55033, w55034, w55035, w55036, w55037, w55038, w55039, w55040, w55041, w55042, w55043, w55044, w55045, w55046, w55047, w55048, w55049, w55050, w55051, w55052, w55053, w55054, w55055, w55056, w55057, w55058, w55059, w55060, w55061, w55062, w55063, w55064, w55065, w55066, w55067, w55068, w55069, w55070, w55071, w55072, w55073, w55074, w55075, w55076, w55077, w55078, w55079, w55080, w55081, w55082, w55083, w55084, w55085, w55086, w55087, w55088, w55089, w55090, w55091, w55092, w55093, w55094, w55095, w55096, w55097, w55098, w55099, w55100, w55101, w55102, w55103, w55104, w55105, w55106, w55107, w55108, w55109, w55110, w55111, w55112, w55113, w55114, w55115, w55116, w55117, w55118, w55119, w55120, w55121, w55122, w55123, w55124, w55125, w55126, w55127, w55128, w55129, w55130, w55131, w55132, w55133, w55134, w55135, w55136, w55137, w55138, w55139, w55140, w55141, w55142, w55143, w55144, w55145, w55146, w55147, w55148, w55149, w55150, w55151, w55152, w55153, w55154, w55155, w55156, w55157, w55158, w55159, w55160, w55161, w55162, w55163, w55164, w55165, w55166, w55167, w55168, w55169, w55170, w55171, w55172, w55173, w55174, w55175, w55176, w55177, w55178, w55179, w55180, w55181, w55182, w55183, w55184, w55185, w55186, w55187, w55188, w55189, w55190, w55191, w55192, w55193, w55194, w55195, w55196, w55197, w55198, w55199, w55200, w55201, w55202, w55203, w55204, w55205, w55206, w55207, w55208, w55209, w55210, w55211, w55212, w55213, w55214, w55215, w55216, w55217, w55218, w55219, w55220, w55221, w55222, w55223, w55224, w55225, w55226, w55227, w55228, w55229, w55230, w55231, w55232, w55233, w55234, w55235, w55236, w55237, w55238, w55239, w55240, w55241, w55242, w55243, w55244, w55245, w55246, w55247, w55248, w55249, w55250, w55251, w55252, w55253, w55254, w55255, w55256, w55257, w55258, w55259, w55260, w55261, w55262, w55263, w55264, w55265, w55266, w55267, w55268, w55269, w55270, w55271, w55272, w55273, w55274, w55275, w55276, w55277, w55278, w55279, w55280, w55281, w55282, w55283, w55284, w55285, w55286, w55287, w55288, w55289, w55290, w55291, w55292, w55293, w55294, w55295, w55296, w55297, w55298, w55299, w55300, w55301, w55302, w55303, w55304, w55305, w55306, w55307, w55308, w55309, w55310, w55311, w55312, w55313, w55314, w55315, w55316, w55317, w55318, w55319, w55320, w55321, w55322, w55323, w55324, w55325, w55326, w55327, w55328, w55329, w55330, w55331, w55332, w55333, w55334, w55335, w55336, w55337, w55338, w55339, w55340, w55341, w55342, w55343, w55344, w55345, w55346, w55347, w55348, w55349, w55350, w55351, w55352, w55353, w55354, w55355, w55356, w55357, w55358, w55359, w55360, w55361, w55362, w55363, w55364, w55365, w55366, w55367, w55368, w55369, w55370, w55371, w55372, w55373, w55374, w55375, w55376, w55377, w55378, w55379, w55380, w55381, w55382, w55383, w55384, w55385, w55386, w55387, w55388, w55389, w55390, w55391, w55392, w55393, w55394, w55395, w55396, w55397, w55398, w55399, w55400, w55401, w55402, w55403, w55404, w55405, w55406, w55407, w55408, w55409, w55410, w55411, w55412, w55413, w55414, w55415, w55416, w55417, w55418, w55419, w55420, w55421, w55422, w55423, w55424, w55425, w55426, w55427, w55428, w55429, w55430, w55431, w55432, w55433, w55434, w55435, w55436, w55437, w55438, w55439, w55440, w55441, w55442, w55443, w55444, w55445, w55446, w55447, w55448, w55449, w55450, w55451, w55452, w55453, w55454, w55455, w55456, w55457, w55458, w55459, w55460, w55461, w55462, w55463, w55464, w55465, w55466, w55467, w55468, w55469, w55470, w55471, w55472, w55473, w55474, w55475, w55476, w55477, w55478, w55479, w55480, w55481, w55482, w55483, w55484, w55485, w55486, w55487, w55488, w55489, w55490, w55491, w55492, w55493, w55494, w55495, w55496, w55497, w55498, w55499, w55500, w55501, w55502, w55503, w55504, w55505, w55506, w55507, w55508, w55509, w55510, w55511, w55512, w55513, w55514, w55515, w55516, w55517, w55518, w55519, w55520, w55521, w55522, w55523, w55524, w55525, w55526, w55527, w55528, w55529, w55530, w55531, w55532, w55533, w55534, w55535, w55536, w55537, w55538, w55539, w55540, w55541, w55542, w55543, w55544, w55545, w55546, w55547, w55548, w55549, w55550, w55551, w55552, w55553, w55554, w55555, w55556, w55557, w55558, w55559, w55560, w55561, w55562, w55563, w55564, w55565, w55566, w55567, w55568, w55569, w55570, w55571, w55572, w55573, w55574, w55575, w55576, w55577, w55578, w55579, w55580, w55581, w55582, w55583, w55584, w55585, w55586, w55587, w55588, w55589, w55590, w55591, w55592, w55593, w55594, w55595, w55596, w55597, w55598, w55599, w55600, w55601, w55602, w55603, w55604, w55605, w55606, w55607, w55608, w55609, w55610, w55611, w55612, w55613, w55614, w55615, w55616, w55617, w55618, w55619, w55620, w55621, w55622, w55623, w55624, w55625, w55626, w55627, w55628, w55629, w55630, w55631, w55632, w55633, w55634, w55635, w55636, w55637, w55638, w55639, w55640, w55641, w55642, w55643, w55644, w55645, w55646, w55647, w55648, w55649, w55650, w55651, w55652, w55653, w55654, w55655, w55656, w55657, w55658, w55659, w55660, w55661, w55662, w55663, w55664, w55665, w55666, w55667, w55668, w55669, w55670, w55671, w55672, w55673, w55674, w55675, w55676, w55677, w55678, w55679, w55680, w55681, w55682, w55683, w55684, w55685, w55686, w55687, w55688, w55689, w55690, w55691, w55692, w55693, w55694, w55695, w55696, w55697, w55698, w55699, w55700, w55701, w55702, w55703, w55704, w55705, w55706, w55707, w55708, w55709, w55710, w55711, w55712, w55713, w55714, w55715, w55716, w55717, w55718, w55719, w55720, w55721, w55722, w55723, w55724, w55725, w55726, w55727, w55728, w55729, w55730, w55731, w55732, w55733, w55734, w55735, w55736, w55737, w55738, w55739, w55740, w55741, w55742, w55743, w55744, w55745, w55746, w55747, w55748, w55749, w55750, w55751, w55752, w55753, w55754, w55755, w55756, w55757, w55758, w55759, w55760, w55761, w55762, w55763, w55764, w55765, w55766, w55767, w55768, w55769, w55770, w55771, w55772, w55773, w55774, w55775, w55776, w55777, w55778, w55779, w55780, w55781, w55782, w55783, w55784, w55785, w55786, w55787, w55788, w55789, w55790, w55791, w55792, w55793, w55794, w55795, w55796, w55797, w55798, w55799, w55800, w55801, w55802, w55803, w55804, w55805, w55806, w55807, w55808, w55809, w55810, w55811, w55812, w55813, w55814, w55815, w55816, w55817, w55818, w55819, w55820, w55821, w55822, w55823, w55824, w55825, w55826, w55827, w55828, w55829, w55830, w55831, w55832, w55833, w55834, w55835, w55836, w55837, w55838, w55839, w55840, w55841, w55842, w55843, w55844, w55845, w55846, w55847, w55848, w55849, w55850, w55851, w55852, w55853, w55854, w55855, w55856, w55857, w55858, w55859, w55860, w55861, w55862, w55863, w55864, w55865, w55866, w55867, w55868, w55869, w55870, w55871, w55872, w55873, w55874, w55875, w55876, w55877, w55878, w55879, w55880, w55881, w55882, w55883, w55884, w55885, w55886, w55887, w55888, w55889, w55890, w55891, w55892, w55893, w55894, w55895, w55896, w55897, w55898, w55899, w55900, w55901, w55902, w55903, w55904, w55905, w55906, w55907, w55908, w55909, w55910, w55911, w55912, w55913, w55914, w55915, w55916, w55917, w55918, w55919, w55920, w55921, w55922, w55923, w55924, w55925, w55926, w55927, w55928, w55929, w55930, w55931, w55932, w55933, w55934, w55935, w55936, w55937, w55938, w55939, w55940, w55941, w55942, w55943, w55944, w55945, w55946, w55947, w55948, w55949, w55950, w55951, w55952, w55953, w55954, w55955, w55956, w55957, w55958, w55959, w55960, w55961, w55962, w55963, w55964, w55965, w55966, w55967, w55968, w55969, w55970, w55971, w55972, w55973, w55974, w55975, w55976, w55977, w55978, w55979, w55980, w55981, w55982, w55983, w55984, w55985, w55986, w55987, w55988, w55989, w55990, w55991, w55992, w55993, w55994, w55995, w55996, w55997, w55998, w55999, w56000, w56001, w56002, w56003, w56004, w56005, w56006, w56007, w56008, w56009, w56010, w56011, w56012, w56013, w56014, w56015, w56016, w56017, w56018, w56019, w56020, w56021, w56022, w56023, w56024, w56025, w56026, w56027, w56028, w56029, w56030, w56031, w56032, w56033, w56034, w56035, w56036, w56037, w56038, w56039, w56040, w56041, w56042, w56043, w56044, w56045, w56046, w56047, w56048, w56049, w56050, w56051, w56052, w56053, w56054, w56055, w56056, w56057, w56058, w56059, w56060, w56061, w56062, w56063, w56064, w56065, w56066, w56067, w56068, w56069, w56070, w56071, w56072, w56073, w56074, w56075, w56076, w56077, w56078, w56079, w56080, w56081, w56082, w56083, w56084, w56085, w56086, w56087, w56088, w56089, w56090, w56091, w56092, w56093, w56094, w56095, w56096, w56097, w56098, w56099, w56100, w56101, w56102, w56103, w56104, w56105, w56106, w56107, w56108, w56109, w56110, w56111, w56112, w56113, w56114, w56115, w56116, w56117, w56118, w56119, w56120, w56121, w56122, w56123, w56124, w56125, w56126, w56127, w56128, w56129, w56130, w56131, w56132, w56133, w56134, w56135, w56136, w56137, w56138, w56139, w56140, w56141, w56142, w56143, w56144, w56145, w56146, w56147, w56148, w56149, w56150, w56151, w56152, w56153, w56154, w56155, w56156, w56157, w56158, w56159, w56160, w56161, w56162, w56163, w56164, w56165, w56166, w56167, w56168, w56169, w56170, w56171, w56172, w56173, w56174, w56175, w56176, w56177, w56178, w56179, w56180, w56181, w56182, w56183, w56184, w56185, w56186, w56187, w56188, w56189, w56190, w56191, w56192, w56193, w56194, w56195, w56196, w56197, w56198, w56199, w56200, w56201, w56202, w56203, w56204, w56205, w56206, w56207, w56208, w56209, w56210, w56211, w56212, w56213, w56214, w56215, w56216, w56217, w56218, w56219, w56220, w56221, w56222, w56223, w56224, w56225, w56226, w56227, w56228, w56229, w56230, w56231, w56232, w56233, w56234, w56235, w56236, w56237, w56238, w56239, w56240, w56241, w56242, w56243, w56244, w56245, w56246, w56247, w56248, w56249, w56250, w56251, w56252, w56253, w56254, w56255, w56256, w56257, w56258, w56259, w56260, w56261, w56262, w56263, w56264, w56265, w56266, w56267, w56268, w56269, w56270, w56271, w56272, w56273, w56274, w56275, w56276, w56277, w56278, w56279, w56280, w56281, w56282, w56283, w56284, w56285, w56286, w56287, w56288, w56289, w56290, w56291, w56292, w56293, w56294, w56295, w56296, w56297, w56298, w56299, w56300, w56301, w56302, w56303, w56304, w56305, w56306, w56307, w56308, w56309, w56310, w56311, w56312, w56313, w56314, w56315, w56316, w56317, w56318, w56319, w56320, w56321, w56322, w56323, w56324, w56325, w56326, w56327, w56328, w56329, w56330, w56331, w56332, w56333, w56334, w56335, w56336, w56337, w56338, w56339, w56340, w56341, w56342, w56343, w56344, w56345, w56346, w56347, w56348, w56349, w56350, w56351, w56352, w56353, w56354, w56355, w56356, w56357, w56358, w56359, w56360, w56361, w56362, w56363, w56364, w56365, w56366, w56367, w56368, w56369, w56370, w56371, w56372, w56373, w56374, w56375, w56376, w56377, w56378, w56379, w56380, w56381, w56382, w56383, w56384, w56385, w56386, w56387, w56388, w56389, w56390, w56391, w56392, w56393, w56394, w56395, w56396, w56397, w56398, w56399, w56400, w56401, w56402, w56403, w56404, w56405, w56406, w56407, w56408, w56409, w56410, w56411, w56412, w56413, w56414, w56415, w56416, w56417, w56418, w56419, w56420, w56421, w56422, w56423, w56424, w56425, w56426, w56427, w56428, w56429, w56430, w56431, w56432, w56433, w56434, w56435, w56436, w56437, w56438, w56439, w56440, w56441, w56442, w56443, w56444, w56445, w56446, w56447, w56448, w56449, w56450, w56451, w56452, w56453, w56454, w56455, w56456, w56457, w56458, w56459, w56460, w56461, w56462, w56463, w56464, w56465, w56466, w56467, w56468, w56469, w56470, w56471, w56472, w56473, w56474, w56475, w56476, w56477, w56478, w56479, w56480, w56481, w56482, w56483, w56484, w56485, w56486, w56487, w56488, w56489, w56490, w56491, w56492, w56493, w56494, w56495, w56496, w56497, w56498, w56499, w56500, w56501, w56502, w56503, w56504, w56505, w56506, w56507, w56508, w56509, w56510, w56511, w56512, w56513, w56514, w56515, w56516, w56517, w56518, w56519, w56520, w56521, w56522, w56523, w56524, w56525, w56526, w56527, w56528, w56529, w56530, w56531, w56532, w56533, w56534, w56535, w56536, w56537, w56538, w56539, w56540, w56541, w56542, w56543, w56544, w56545, w56546, w56547, w56548, w56549, w56550, w56551, w56552, w56553, w56554, w56555, w56556, w56557, w56558, w56559, w56560, w56561, w56562, w56563, w56564, w56565, w56566, w56567, w56568, w56569, w56570, w56571, w56572, w56573, w56574, w56575, w56576, w56577, w56578, w56579, w56580, w56581, w56582, w56583, w56584, w56585, w56586, w56587, w56588, w56589, w56590, w56591, w56592, w56593, w56594, w56595, w56596, w56597, w56598, w56599, w56600, w56601, w56602, w56603, w56604, w56605, w56606, w56607, w56608, w56609, w56610, w56611, w56612, w56613, w56614, w56615, w56616, w56617, w56618, w56619, w56620, w56621, w56622, w56623, w56624, w56625, w56626, w56627, w56628, w56629, w56630, w56631, w56632, w56633, w56634, w56635, w56636, w56637, w56638, w56639, w56640, w56641, w56642, w56643, w56644, w56645, w56646, w56647, w56648, w56649, w56650, w56651, w56652, w56653, w56654, w56655, w56656, w56657, w56658, w56659, w56660, w56661, w56662, w56663, w56664, w56665, w56666, w56667, w56668, w56669, w56670, w56671, w56672, w56673, w56674, w56675, w56676, w56677, w56678, w56679, w56680, w56681, w56682, w56683, w56684, w56685, w56686, w56687, w56688, w56689, w56690, w56691, w56692, w56693, w56694, w56695, w56696, w56697, w56698, w56699, w56700, w56701, w56702, w56703, w56704, w56705, w56706, w56707, w56708, w56709, w56710, w56711, w56712, w56713, w56714, w56715, w56716, w56717, w56718, w56719, w56720, w56721, w56722, w56723, w56724, w56725, w56726, w56727, w56728, w56729, w56730, w56731, w56732, w56733, w56734, w56735, w56736, w56737, w56738, w56739, w56740, w56741, w56742, w56743, w56744, w56745, w56746, w56747, w56748, w56749, w56750, w56751, w56752, w56753, w56754, w56755, w56756, w56757, w56758, w56759, w56760, w56761, w56762, w56763, w56764, w56765, w56766, w56767, w56768, w56769, w56770, w56771, w56772, w56773, w56774, w56775, w56776, w56777, w56778, w56779, w56780, w56781, w56782, w56783, w56784, w56785, w56786, w56787, w56788, w56789, w56790, w56791, w56792, w56793, w56794, w56795, w56796, w56797, w56798, w56799, w56800, w56801, w56802, w56803, w56804, w56805, w56806, w56807, w56808, w56809, w56810, w56811, w56812, w56813, w56814, w56815, w56816, w56817, w56818, w56819, w56820, w56821, w56822, w56823, w56824, w56825, w56826, w56827, w56828, w56829, w56830, w56831, w56832, w56833, w56834, w56835, w56836, w56837, w56838, w56839, w56840, w56841, w56842, w56843, w56844, w56845, w56846, w56847, w56848, w56849, w56850, w56851, w56852, w56853, w56854, w56855, w56856, w56857, w56858, w56859, w56860, w56861, w56862, w56863, w56864, w56865, w56866, w56867, w56868, w56869, w56870, w56871, w56872, w56873, w56874, w56875, w56876, w56877, w56878, w56879, w56880, w56881, w56882, w56883, w56884, w56885, w56886, w56887, w56888, w56889, w56890, w56891, w56892, w56893, w56894, w56895, w56896, w56897, w56898, w56899, w56900, w56901, w56902, w56903, w56904, w56905, w56906, w56907, w56908, w56909, w56910, w56911, w56912, w56913, w56914, w56915, w56916, w56917, w56918, w56919, w56920, w56921, w56922, w56923, w56924, w56925, w56926, w56927, w56928, w56929, w56930, w56931, w56932, w56933, w56934, w56935, w56936, w56937, w56938, w56939, w56940, w56941, w56942, w56943, w56944, w56945, w56946, w56947, w56948, w56949, w56950, w56951, w56952, w56953, w56954, w56955, w56956, w56957, w56958, w56959, w56960, w56961, w56962, w56963, w56964, w56965, w56966, w56967, w56968, w56969, w56970, w56971, w56972, w56973, w56974, w56975, w56976, w56977, w56978, w56979, w56980, w56981, w56982, w56983, w56984, w56985, w56986, w56987, w56988, w56989, w56990, w56991, w56992, w56993, w56994, w56995, w56996, w56997, w56998, w56999, w57000, w57001, w57002, w57003, w57004, w57005, w57006, w57007, w57008, w57009, w57010, w57011, w57012, w57013, w57014, w57015, w57016, w57017, w57018, w57019, w57020, w57021, w57022, w57023, w57024, w57025, w57026, w57027, w57028, w57029, w57030, w57031, w57032, w57033, w57034, w57035, w57036, w57037, w57038, w57039, w57040, w57041, w57042, w57043, w57044, w57045, w57046, w57047, w57048, w57049, w57050, w57051, w57052, w57053, w57054, w57055, w57056, w57057, w57058, w57059, w57060, w57061, w57062, w57063, w57064, w57065, w57066, w57067, w57068, w57069, w57070, w57071, w57072, w57073, w57074, w57075, w57076, w57077, w57078, w57079, w57080, w57081, w57082, w57083, w57084, w57085, w57086, w57087, w57088, w57089, w57090, w57091, w57092, w57093, w57094, w57095, w57096, w57097, w57098, w57099, w57100, w57101, w57102, w57103, w57104, w57105, w57106, w57107, w57108, w57109, w57110, w57111, w57112, w57113, w57114, w57115, w57116, w57117, w57118, w57119, w57120, w57121, w57122, w57123, w57124, w57125, w57126, w57127, w57128, w57129, w57130, w57131, w57132, w57133, w57134, w57135, w57136, w57137, w57138, w57139, w57140, w57141, w57142, w57143, w57144, w57145, w57146, w57147, w57148, w57149, w57150, w57151, w57152, w57153, w57154, w57155, w57156, w57157, w57158, w57159, w57160, w57161, w57162, w57163, w57164, w57165, w57166, w57167, w57168, w57169, w57170, w57171, w57172, w57173, w57174, w57175, w57176, w57177, w57178, w57179, w57180, w57181, w57182, w57183, w57184, w57185, w57186, w57187, w57188, w57189, w57190, w57191, w57192, w57193, w57194, w57195, w57196, w57197, w57198, w57199, w57200, w57201, w57202, w57203, w57204, w57205, w57206, w57207, w57208, w57209, w57210, w57211, w57212, w57213, w57214, w57215, w57216, w57217, w57218, w57219, w57220, w57221, w57222, w57223, w57224, w57225, w57226, w57227, w57228, w57229, w57230, w57231, w57232, w57233, w57234, w57235, w57236, w57237, w57238, w57239, w57240, w57241, w57242, w57243, w57244, w57245, w57246: std_logic;

begin

w0 <= not a(63) and b(0);
w1 <= b(0) and not b(1);
w2 <= not b(2) and not b(3);
w3 <= w1 and w2;
w4 <= not w0 and w3;
w5 <= not b(8) and not b(9);
w6 <= not b(10) and not b(11);
w7 <= w5 and w6;
w8 <= not b(4) and not b(5);
w9 <= not b(6) and not b(7);
w10 <= w8 and w9;
w11 <= w7 and w10;
w12 <= not b(16) and not b(17);
w13 <= not b(18) and not b(19);
w14 <= w12 and w13;
w15 <= not b(12) and not b(13);
w16 <= not b(14) and not b(15);
w17 <= w15 and w16;
w18 <= w14 and w17;
w19 <= w11 and w18;
w20 <= w4 and w19;
w21 <= not b(60) and not b(61);
w22 <= not b(62) and not b(63);
w23 <= w21 and w22;
w24 <= not b(56) and not b(57);
w25 <= not b(58) and not b(59);
w26 <= w24 and w25;
w27 <= not b(52) and not b(53);
w28 <= not b(54) and not b(55);
w29 <= w27 and w28;
w30 <= w26 and w29;
w31 <= w23 and w30;
w32 <= not b(40) and not b(41);
w33 <= not b(42) and not b(43);
w34 <= w32 and w33;
w35 <= not b(36) and not b(37);
w36 <= not b(38) and not b(39);
w37 <= w35 and w36;
w38 <= w34 and w37;
w39 <= not b(48) and not b(49);
w40 <= not b(50) and not b(51);
w41 <= w39 and w40;
w42 <= not b(44) and not b(45);
w43 <= not b(46) and not b(47);
w44 <= w42 and w43;
w45 <= w41 and w44;
w46 <= w38 and w45;
w47 <= not b(24) and not b(25);
w48 <= not b(26) and not b(27);
w49 <= w47 and w48;
w50 <= not b(20) and not b(21);
w51 <= not b(22) and not b(23);
w52 <= w50 and w51;
w53 <= w49 and w52;
w54 <= not b(32) and not b(33);
w55 <= not b(34) and not b(35);
w56 <= w54 and w55;
w57 <= not b(28) and not b(29);
w58 <= not b(30) and not b(31);
w59 <= w57 and w58;
w60 <= w56 and w59;
w61 <= w53 and w60;
w62 <= w46 and w61;
w63 <= w31 and w62;
w64 <= w20 and w63;
w65 <= not a(62) and b(0);
w66 <= b(1) and w65;
w67 <= a(63) and not w66;
w68 <= not w64 and w67;
w69 <= not b(1) and not w65;
w70 <= not w68 and not w69;
w71 <= a(63) and not w64;
w72 <= b(1) and not w65;
w73 <= not b(1) and w65;
w74 <= not w72 and not w73;
w75 <= w2 and w10;
w76 <= w7 and w17;
w77 <= w75 and w76;
w78 <= not w74 and w77;
w79 <= w29 and w41;
w80 <= w23 and w26;
w81 <= w79 and w80;
w82 <= w37 and w56;
w83 <= w34 and w44;
w84 <= w82 and w83;
w85 <= w14 and w52;
w86 <= w49 and w59;
w87 <= w85 and w86;
w88 <= w84 and w87;
w89 <= w81 and w88;
w90 <= w78 and w89;
w91 <= not w71 and w90;
w92 <= not w70 and w91;
w93 <= w76 and w85;
w94 <= w75 and w93;
w95 <= not w66 and not w69;
w96 <= w80 and w95;
w97 <= w79 and w83;
w98 <= w82 and w86;
w99 <= w97 and w98;
w100 <= w96 and w99;
w101 <= w94 and w100;
w102 <= not w70 and w101;
w103 <= w71 and not w102;
w104 <= not w92 and not w103;
w105 <= not a(61) and b(0);
w106 <= b(1) and w105;
w107 <= not b(21) and not b(22);
w108 <= not b(23) and not b(24);
w109 <= w107 and w108;
w110 <= not b(17) and not b(18);
w111 <= not b(19) and not b(20);
w112 <= w110 and w111;
w113 <= w109 and w112;
w114 <= not b(29) and not b(30);
w115 <= not b(31) and not b(32);
w116 <= w114 and w115;
w117 <= not b(25) and not b(26);
w118 <= not b(27) and not b(28);
w119 <= w117 and w118;
w120 <= w116 and w119;
w121 <= w113 and w120;
w122 <= not b(5) and not b(6);
w123 <= not b(7) and not b(8);
w124 <= w122 and w123;
w125 <= b(0) and not b(2);
w126 <= not b(3) and not b(4);
w127 <= w125 and w126;
w128 <= w124 and w127;
w129 <= not b(13) and not b(14);
w130 <= not b(15) and not b(16);
w131 <= w129 and w130;
w132 <= not b(9) and not b(10);
w133 <= not b(11) and not b(12);
w134 <= w132 and w133;
w135 <= w131 and w134;
w136 <= w128 and w135;
w137 <= w121 and w136;
w138 <= not b(53) and not b(54);
w139 <= not b(55) and not b(56);
w140 <= w138 and w139;
w141 <= not b(49) and not b(50);
w142 <= not b(51) and not b(52);
w143 <= w141 and w142;
w144 <= w140 and w143;
w145 <= not b(61) and not b(62);
w146 <= not b(63) and w145;
w147 <= not b(57) and not b(58);
w148 <= not b(59) and not b(60);
w149 <= w147 and w148;
w150 <= w146 and w149;
w151 <= w144 and w150;
w152 <= not b(37) and not b(38);
w153 <= not b(39) and not b(40);
w154 <= w152 and w153;
w155 <= not b(33) and not b(34);
w156 <= not b(35) and not b(36);
w157 <= w155 and w156;
w158 <= w154 and w157;
w159 <= not b(45) and not b(46);
w160 <= not b(47) and not b(48);
w161 <= w159 and w160;
w162 <= not b(41) and not b(42);
w163 <= not b(43) and not b(44);
w164 <= w162 and w163;
w165 <= w161 and w164;
w166 <= w158 and w165;
w167 <= w151 and w166;
w168 <= w137 and w167;
w169 <= not w70 and w168;
w170 <= a(62) and not w169;
w171 <= w2 and w65;
w172 <= w10 and w171;
w173 <= w76 and w172;
w174 <= w87 and w173;
w175 <= w81 and w84;
w176 <= w174 and w175;
w177 <= not w70 and w176;
w178 <= not w170 and not w177;
w179 <= not w106 and not w178;
w180 <= not b(1) and not w105;
w181 <= not w179 and not w180;
w182 <= b(2) and not w92;
w183 <= not w103 and w182;
w184 <= not b(2) and not w104;
w185 <= not w183 and not w184;
w186 <= w181 and not w185;
w187 <= not b(2) and not w186;
w188 <= not w181 and not w183;
w189 <= not w184 and not w188;
w190 <= w124 and w126;
w191 <= w135 and w190;
w192 <= w121 and w191;
w193 <= w167 and w192;
w194 <= not w189 and w193;
w195 <= not w187 and w194;
w196 <= not w104 and not w195;
w197 <= not w188 and w193;
w198 <= not w186 and w197;
w199 <= not w189 and w198;
w200 <= b(3) and not w199;
w201 <= not w196 and w200;
w202 <= w113 and w135;
w203 <= w190 and w202;
w204 <= not w106 and not w180;
w205 <= w150 and w204;
w206 <= w144 and w165;
w207 <= w120 and w158;
w208 <= w206 and w207;
w209 <= w205 and w208;
w210 <= w203 and w209;
w211 <= not w189 and w210;
w212 <= not w178 and not w211;
w213 <= b(1) and not w105;
w214 <= not b(1) and w105;
w215 <= not w213 and not w214;
w216 <= w191 and not w215;
w217 <= w121 and w166;
w218 <= w151 and w217;
w219 <= w216 and w218;
w220 <= not w177 and w219;
w221 <= not w170 and w220;
w222 <= not w189 and w221;
w223 <= not w212 and not w222;
w224 <= not b(2) and not w223;
w225 <= b(2) and not w222;
w226 <= not w212 and w225;
w227 <= b(0) and not b(3);
w228 <= w10 and w227;
w229 <= w76 and w228;
w230 <= w87 and w229;
w231 <= w175 and w230;
w232 <= not w189 and w231;
w233 <= a(61) and not w232;
w234 <= w105 and w126;
w235 <= w124 and w234;
w236 <= w135 and w235;
w237 <= w121 and w236;
w238 <= w167 and w237;
w239 <= not w189 and w238;
w240 <= not w233 and not w239;
w241 <= not a(60) and b(0);
w242 <= b(1) and w241;
w243 <= not w240 and not w242;
w244 <= not b(1) and not w241;
w245 <= not w243 and not w244;
w246 <= not w226 and not w245;
w247 <= not w224 and not w246;
w248 <= not w201 and not w247;
w249 <= not w196 and not w199;
w250 <= not b(3) and not w249;
w251 <= not w248 and not w250;
w252 <= not w201 and not w250;
w253 <= not w247 and w252;
w254 <= w19 and w61;
w255 <= w31 and w46;
w256 <= w254 and w255;
w257 <= w247 and not w252;
w258 <= w256 and not w257;
w259 <= not w253 and w258;
w260 <= not w251 and w259;
w261 <= not w251 and w256;
w262 <= not w249 and not w261;
w263 <= b(4) and not w262;
w264 <= not w260 and w263;
w265 <= not w224 and not w226;
w266 <= w245 and not w265;
w267 <= not w246 and w256;
w268 <= not w266 and w267;
w269 <= not w251 and w268;
w270 <= not b(2) and not w266;
w271 <= w256 and not w270;
w272 <= not w251 and w271;
w273 <= not w223 and not w272;
w274 <= not w269 and not w273;
w275 <= not b(3) and not w274;
w276 <= b(3) and not w269;
w277 <= not w273 and w276;
w278 <= w18 and w53;
w279 <= w11 and w278;
w280 <= w23 and not w242;
w281 <= not w244 and w280;
w282 <= w30 and w45;
w283 <= w38 and w60;
w284 <= w282 and w283;
w285 <= w281 and w284;
w286 <= w279 and w285;
w287 <= not w251 and w286;
w288 <= not w240 and not w287;
w289 <= b(1) and not w241;
w290 <= not b(1) and w241;
w291 <= not w289 and not w290;
w292 <= w19 and not w291;
w293 <= w63 and w292;
w294 <= not w239 and w293;
w295 <= not w233 and w294;
w296 <= not w251 and w295;
w297 <= not w288 and not w296;
w298 <= not b(2) and not w297;
w299 <= b(2) and not w296;
w300 <= not w288 and w299;
w301 <= not a(59) and b(0);
w302 <= b(1) and w301;
w303 <= b(0) and not b(4);
w304 <= w124 and w303;
w305 <= w135 and w304;
w306 <= w121 and w305;
w307 <= w167 and w306;
w308 <= not w251 and w307;
w309 <= a(60) and not w308;
w310 <= w10 and w241;
w311 <= w76 and w310;
w312 <= w87 and w311;
w313 <= w175 and w312;
w314 <= not w251 and w313;
w315 <= not w309 and not w314;
w316 <= not w302 and not w315;
w317 <= not b(1) and not w301;
w318 <= not w316 and not w317;
w319 <= not w300 and not w318;
w320 <= not w298 and not w319;
w321 <= not w277 and not w320;
w322 <= not w275 and not w321;
w323 <= not w264 and not w322;
w324 <= not w260 and not w262;
w325 <= not b(4) and not w324;
w326 <= not w323 and not w325;
w327 <= not w275 and not w277;
w328 <= not w298 and not w327;
w329 <= not w319 and w328;
w330 <= w109 and w119;
w331 <= w116 and w157;
w332 <= w330 and w331;
w333 <= w124 and w134;
w334 <= w112 and w131;
w335 <= w333 and w334;
w336 <= w332 and w335;
w337 <= w140 and w149;
w338 <= w146 and w337;
w339 <= w154 and w164;
w340 <= w143 and w161;
w341 <= w339 and w340;
w342 <= w338 and w341;
w343 <= w336 and w342;
w344 <= not w329 and w343;
w345 <= not w321 and w344;
w346 <= not w326 and w345;
w347 <= not b(3) and not w329;
w348 <= w343 and not w347;
w349 <= not w326 and w348;
w350 <= not w274 and not w349;
w351 <= not w346 and not w350;
w352 <= b(4) and not w351;
w353 <= not b(4) and not w346;
w354 <= not w350 and w353;
w355 <= not w352 and not w354;
w356 <= not w298 and not w300;
w357 <= w318 and not w356;
w358 <= not w319 and w343;
w359 <= not w357 and w358;
w360 <= not w326 and w359;
w361 <= not b(2) and not w357;
w362 <= w343 and not w361;
w363 <= not w326 and w362;
w364 <= not w297 and not w363;
w365 <= not w360 and not w364;
w366 <= b(3) and not w365;
w367 <= not b(3) and not w360;
w368 <= not w364 and w367;
w369 <= not w366 and not w368;
w370 <= w330 and w334;
w371 <= w333 and w370;
w372 <= w146 and not w302;
w373 <= not w317 and w372;
w374 <= w337 and w340;
w375 <= w331 and w339;
w376 <= w374 and w375;
w377 <= w373 and w376;
w378 <= w371 and w377;
w379 <= not w326 and w378;
w380 <= not w315 and not w379;
w381 <= b(1) and not w301;
w382 <= not b(1) and w301;
w383 <= not w381 and not w382;
w384 <= w335 and not w383;
w385 <= w332 and w341;
w386 <= w338 and w385;
w387 <= w384 and w386;
w388 <= not w314 and w387;
w389 <= not w309 and w388;
w390 <= not w326 and w389;
w391 <= not w380 and not w390;
w392 <= not b(2) and not w391;
w393 <= b(0) and not b(5);
w394 <= w9 and w393;
w395 <= w7 and w394;
w396 <= w18 and w395;
w397 <= w61 and w396;
w398 <= w255 and w397;
w399 <= not w326 and w398;
w400 <= a(59) and not w399;
w401 <= w124 and w301;
w402 <= w135 and w401;
w403 <= w121 and w402;
w404 <= w167 and w403;
w405 <= not w326 and w404;
w406 <= not w400 and not w405;
w407 <= b(1) and not w406;
w408 <= not b(1) and not w405;
w409 <= not w400 and w408;
w410 <= not w407 and not w409;
w411 <= not a(58) and b(0);
w412 <= not w410 and not w411;
w413 <= not b(1) and not w406;
w414 <= not w412 and not w413;
w415 <= b(2) and not w390;
w416 <= not w380 and w415;
w417 <= not w392 and not w416;
w418 <= not w414 and w417;
w419 <= not w392 and not w418;
w420 <= not w369 and not w419;
w421 <= not b(3) and not w365;
w422 <= not w420 and not w421;
w423 <= not w355 and not w422;
w424 <= not b(4) and not w351;
w425 <= not w423 and not w424;
w426 <= not w264 and not w325;
w427 <= not w275 and not w426;
w428 <= not w321 and w427;
w429 <= w343 and not w428;
w430 <= not w323 and w429;
w431 <= not w326 and w430;
w432 <= not b(4) and not w428;
w433 <= w343 and not w432;
w434 <= not w326 and w433;
w435 <= not w324 and not w434;
w436 <= not w431 and not w435;
w437 <= b(5) and not w436;
w438 <= not b(5) and not w431;
w439 <= not w435 and w438;
w440 <= not w437 and not w439;
w441 <= w7 and w9;
w442 <= w18 and w441;
w443 <= w61 and w442;
w444 <= w255 and w443;
w445 <= not w440 and w444;
w446 <= not w425 and w445;
w447 <= w343 and not w436;
w448 <= not w446 and not w447;
w449 <= w355 and not w421;
w450 <= not w420 and w449;
w451 <= not w423 and not w450;
w452 <= not w448 and w451;
w453 <= not w351 and not w447;
w454 <= not w446 and w453;
w455 <= not w452 and not w454;
w456 <= not w425 and not w440;
w457 <= not w424 and w440;
w458 <= not w423 and w457;
w459 <= not w456 and not w458;
w460 <= not w448 and w459;
w461 <= not w436 and not w447;
w462 <= not w446 and w461;
w463 <= not w460 and not w462;
w464 <= not b(6) and not w463;
w465 <= not b(5) and not w455;
w466 <= w369 and not w392;
w467 <= not w418 and w466;
w468 <= not w420 and not w467;
w469 <= not w448 and w468;
w470 <= not w365 and not w447;
w471 <= not w446 and w470;
w472 <= not w469 and not w471;
w473 <= not b(4) and not w472;
w474 <= not w413 and w417;
w475 <= not w412 and w474;
w476 <= not w414 and not w417;
w477 <= not w475 and not w476;
w478 <= not w448 and not w477;
w479 <= not w391 and not w447;
w480 <= not w446 and w479;
w481 <= not w478 and not w480;
w482 <= not b(3) and not w481;
w483 <= not w409 and w411;
w484 <= not w407 and w483;
w485 <= not w412 and not w484;
w486 <= not w448 and w485;
w487 <= not w406 and not w447;
w488 <= not w446 and w487;
w489 <= not w486 and not w488;
w490 <= not b(2) and not w489;
w491 <= b(0) and not w448;
w492 <= a(58) and not w491;
w493 <= w411 and not w448;
w494 <= not w492 and not w493;
w495 <= b(1) and not w494;
w496 <= not b(1) and not w493;
w497 <= not w492 and w496;
w498 <= not w495 and not w497;
w499 <= not a(57) and b(0);
w500 <= not w498 and not w499;
w501 <= not b(1) and not w494;
w502 <= not w500 and not w501;
w503 <= b(2) and not w488;
w504 <= not w486 and w503;
w505 <= not w490 and not w504;
w506 <= not w502 and w505;
w507 <= not w490 and not w506;
w508 <= b(3) and not w480;
w509 <= not w478 and w508;
w510 <= not w482 and not w509;
w511 <= not w507 and w510;
w512 <= not w482 and not w511;
w513 <= b(4) and not w471;
w514 <= not w469 and w513;
w515 <= not w473 and not w514;
w516 <= not w512 and w515;
w517 <= not w473 and not w516;
w518 <= b(5) and not w454;
w519 <= not w452 and w518;
w520 <= not w465 and not w519;
w521 <= not w517 and w520;
w522 <= not w465 and not w521;
w523 <= b(6) and not w462;
w524 <= not w460 and w523;
w525 <= not w464 and not w524;
w526 <= not w522 and w525;
w527 <= not w464 and not w526;
w528 <= w123 and w134;
w529 <= w334 and w528;
w530 <= w332 and w529;
w531 <= w342 and w530;
w532 <= not w527 and w531;
w533 <= not w455 and not w532;
w534 <= not w473 and w520;
w535 <= not w516 and w534;
w536 <= not w517 and not w520;
w537 <= not w535 and not w536;
w538 <= w531 and not w537;
w539 <= not w527 and w538;
w540 <= not w533 and not w539;
w541 <= not w463 and not w532;
w542 <= not w465 and w525;
w543 <= not w521 and w542;
w544 <= not w522 and not w525;
w545 <= not w543 and not w544;
w546 <= w532 and not w545;
w547 <= not w541 and not w546;
w548 <= not b(7) and not w547;
w549 <= not b(6) and not w540;
w550 <= not w472 and not w532;
w551 <= not w482 and w515;
w552 <= not w511 and w551;
w553 <= not w512 and not w515;
w554 <= not w552 and not w553;
w555 <= w531 and not w554;
w556 <= not w527 and w555;
w557 <= not w550 and not w556;
w558 <= not b(5) and not w557;
w559 <= not w481 and not w532;
w560 <= not w490 and w510;
w561 <= not w506 and w560;
w562 <= not w507 and not w510;
w563 <= not w561 and not w562;
w564 <= w531 and not w563;
w565 <= not w527 and w564;
w566 <= not w559 and not w565;
w567 <= not b(4) and not w566;
w568 <= not w489 and not w532;
w569 <= not w501 and w505;
w570 <= not w500 and w569;
w571 <= not w502 and not w505;
w572 <= not w570 and not w571;
w573 <= w531 and not w572;
w574 <= not w527 and w573;
w575 <= not w568 and not w574;
w576 <= not b(3) and not w575;
w577 <= not w494 and not w532;
w578 <= not w497 and w499;
w579 <= not w495 and w578;
w580 <= w531 and not w579;
w581 <= not w500 and w580;
w582 <= not w527 and w581;
w583 <= not w577 and not w582;
w584 <= not b(2) and not w583;
w585 <= b(0) and not b(7);
w586 <= w7 and w585;
w587 <= w18 and w586;
w588 <= w61 and w587;
w589 <= w255 and w588;
w590 <= not w527 and w589;
w591 <= a(57) and not w590;
w592 <= w123 and w499;
w593 <= w134 and w592;
w594 <= w334 and w593;
w595 <= w332 and w594;
w596 <= w342 and w595;
w597 <= not w527 and w596;
w598 <= not w591 and not w597;
w599 <= b(1) and not w598;
w600 <= not b(1) and not w597;
w601 <= not w591 and w600;
w602 <= not w599 and not w601;
w603 <= not a(56) and b(0);
w604 <= not w602 and not w603;
w605 <= not b(1) and not w598;
w606 <= not w604 and not w605;
w607 <= b(2) and not w582;
w608 <= not w577 and w607;
w609 <= not w584 and not w608;
w610 <= not w606 and w609;
w611 <= not w584 and not w610;
w612 <= b(3) and not w574;
w613 <= not w568 and w612;
w614 <= not w576 and not w613;
w615 <= not w611 and w614;
w616 <= not w576 and not w615;
w617 <= b(4) and not w565;
w618 <= not w559 and w617;
w619 <= not w567 and not w618;
w620 <= not w616 and w619;
w621 <= not w567 and not w620;
w622 <= b(5) and not w556;
w623 <= not w550 and w622;
w624 <= not w558 and not w623;
w625 <= not w621 and w624;
w626 <= not w558 and not w625;
w627 <= b(6) and not w539;
w628 <= not w533 and w627;
w629 <= not w549 and not w628;
w630 <= not w626 and w629;
w631 <= not w549 and not w630;
w632 <= b(7) and not w541;
w633 <= not w546 and w632;
w634 <= not w548 and not w633;
w635 <= not w631 and w634;
w636 <= not w548 and not w635;
w637 <= w76 and w87;
w638 <= w175 and w637;
w639 <= not w636 and w638;
w640 <= not w540 and not w639;
w641 <= not w558 and w629;
w642 <= not w625 and w641;
w643 <= not w626 and not w629;
w644 <= not w642 and not w643;
w645 <= w638 and not w644;
w646 <= not w636 and w645;
w647 <= not w640 and not w646;
w648 <= not b(7) and not w647;
w649 <= not w557 and not w639;
w650 <= not w567 and w624;
w651 <= not w620 and w650;
w652 <= not w621 and not w624;
w653 <= not w651 and not w652;
w654 <= w638 and not w653;
w655 <= not w636 and w654;
w656 <= not w649 and not w655;
w657 <= not b(6) and not w656;
w658 <= not w566 and not w639;
w659 <= not w576 and w619;
w660 <= not w615 and w659;
w661 <= not w616 and not w619;
w662 <= not w660 and not w661;
w663 <= w638 and not w662;
w664 <= not w636 and w663;
w665 <= not w658 and not w664;
w666 <= not b(5) and not w665;
w667 <= not w575 and not w639;
w668 <= not w584 and w614;
w669 <= not w610 and w668;
w670 <= not w611 and not w614;
w671 <= not w669 and not w670;
w672 <= w638 and not w671;
w673 <= not w636 and w672;
w674 <= not w667 and not w673;
w675 <= not b(4) and not w674;
w676 <= not w583 and not w639;
w677 <= not w605 and w609;
w678 <= not w604 and w677;
w679 <= not w606 and not w609;
w680 <= not w678 and not w679;
w681 <= w638 and not w680;
w682 <= not w636 and w681;
w683 <= not w676 and not w682;
w684 <= not b(3) and not w683;
w685 <= not w598 and not w639;
w686 <= not w601 and w603;
w687 <= not w599 and w686;
w688 <= w638 and not w687;
w689 <= not w604 and w688;
w690 <= not w636 and w689;
w691 <= not w685 and not w690;
w692 <= not b(2) and not w691;
w693 <= b(0) and not b(8);
w694 <= w134 and w693;
w695 <= w334 and w694;
w696 <= w332 and w695;
w697 <= w342 and w696;
w698 <= not w636 and w697;
w699 <= a(56) and not w698;
w700 <= w7 and w603;
w701 <= w18 and w700;
w702 <= w61 and w701;
w703 <= w255 and w702;
w704 <= not w636 and w703;
w705 <= not w699 and not w704;
w706 <= b(1) and not w705;
w707 <= not b(1) and not w704;
w708 <= not w699 and w707;
w709 <= not w706 and not w708;
w710 <= not a(55) and b(0);
w711 <= not w709 and not w710;
w712 <= not b(1) and not w705;
w713 <= not w711 and not w712;
w714 <= b(2) and not w690;
w715 <= not w685 and w714;
w716 <= not w692 and not w715;
w717 <= not w713 and w716;
w718 <= not w692 and not w717;
w719 <= b(3) and not w682;
w720 <= not w676 and w719;
w721 <= not w684 and not w720;
w722 <= not w718 and w721;
w723 <= not w684 and not w722;
w724 <= b(4) and not w673;
w725 <= not w667 and w724;
w726 <= not w675 and not w725;
w727 <= not w723 and w726;
w728 <= not w675 and not w727;
w729 <= b(5) and not w664;
w730 <= not w658 and w729;
w731 <= not w666 and not w730;
w732 <= not w728 and w731;
w733 <= not w666 and not w732;
w734 <= b(6) and not w655;
w735 <= not w649 and w734;
w736 <= not w657 and not w735;
w737 <= not w733 and w736;
w738 <= not w657 and not w737;
w739 <= b(7) and not w646;
w740 <= not w640 and w739;
w741 <= not w648 and not w740;
w742 <= not w738 and w741;
w743 <= not w648 and not w742;
w744 <= not w547 and not w639;
w745 <= not w549 and w634;
w746 <= not w630 and w745;
w747 <= not w631 and not w634;
w748 <= not w746 and not w747;
w749 <= w639 and not w748;
w750 <= not w744 and not w749;
w751 <= not b(8) and not w750;
w752 <= b(8) and not w744;
w753 <= not w749 and w752;
w754 <= w121 and w135;
w755 <= w167 and w754;
w756 <= not w753 and w755;
w757 <= not w751 and w756;
w758 <= not w743 and w757;
w759 <= w638 and not w750;
w760 <= not w758 and not w759;
w761 <= not w657 and w741;
w762 <= not w737 and w761;
w763 <= not w738 and not w741;
w764 <= not w762 and not w763;
w765 <= not w760 and not w764;
w766 <= not w647 and not w759;
w767 <= not w758 and w766;
w768 <= not w765 and not w767;
w769 <= not w648 and not w753;
w770 <= not w751 and w769;
w771 <= not w742 and w770;
w772 <= not w751 and not w753;
w773 <= not w743 and not w772;
w774 <= not w771 and not w773;
w775 <= not w760 and not w774;
w776 <= not w750 and not w759;
w777 <= not w758 and w776;
w778 <= not w775 and not w777;
w779 <= not b(9) and not w778;
w780 <= not b(8) and not w768;
w781 <= not w666 and w736;
w782 <= not w732 and w781;
w783 <= not w733 and not w736;
w784 <= not w782 and not w783;
w785 <= not w760 and not w784;
w786 <= not w656 and not w759;
w787 <= not w758 and w786;
w788 <= not w785 and not w787;
w789 <= not b(7) and not w788;
w790 <= not w675 and w731;
w791 <= not w727 and w790;
w792 <= not w728 and not w731;
w793 <= not w791 and not w792;
w794 <= not w760 and not w793;
w795 <= not w665 and not w759;
w796 <= not w758 and w795;
w797 <= not w794 and not w796;
w798 <= not b(6) and not w797;
w799 <= not w684 and w726;
w800 <= not w722 and w799;
w801 <= not w723 and not w726;
w802 <= not w800 and not w801;
w803 <= not w760 and not w802;
w804 <= not w674 and not w759;
w805 <= not w758 and w804;
w806 <= not w803 and not w805;
w807 <= not b(5) and not w806;
w808 <= not w692 and w721;
w809 <= not w717 and w808;
w810 <= not w718 and not w721;
w811 <= not w809 and not w810;
w812 <= not w760 and not w811;
w813 <= not w683 and not w759;
w814 <= not w758 and w813;
w815 <= not w812 and not w814;
w816 <= not b(4) and not w815;
w817 <= not w712 and w716;
w818 <= not w711 and w817;
w819 <= not w713 and not w716;
w820 <= not w818 and not w819;
w821 <= not w760 and not w820;
w822 <= not w691 and not w759;
w823 <= not w758 and w822;
w824 <= not w821 and not w823;
w825 <= not b(3) and not w824;
w826 <= not w708 and w710;
w827 <= not w706 and w826;
w828 <= not w711 and not w827;
w829 <= not w760 and w828;
w830 <= not w705 and not w759;
w831 <= not w758 and w830;
w832 <= not w829 and not w831;
w833 <= not b(2) and not w832;
w834 <= b(0) and not w760;
w835 <= a(55) and not w834;
w836 <= w710 and not w760;
w837 <= not w835 and not w836;
w838 <= b(1) and not w837;
w839 <= not b(1) and not w836;
w840 <= not w835 and w839;
w841 <= not w838 and not w840;
w842 <= not a(54) and b(0);
w843 <= not w841 and not w842;
w844 <= not b(1) and not w837;
w845 <= not w843 and not w844;
w846 <= b(2) and not w831;
w847 <= not w829 and w846;
w848 <= not w833 and not w847;
w849 <= not w845 and w848;
w850 <= not w833 and not w849;
w851 <= b(3) and not w823;
w852 <= not w821 and w851;
w853 <= not w825 and not w852;
w854 <= not w850 and w853;
w855 <= not w825 and not w854;
w856 <= b(4) and not w814;
w857 <= not w812 and w856;
w858 <= not w816 and not w857;
w859 <= not w855 and w858;
w860 <= not w816 and not w859;
w861 <= b(5) and not w805;
w862 <= not w803 and w861;
w863 <= not w807 and not w862;
w864 <= not w860 and w863;
w865 <= not w807 and not w864;
w866 <= b(6) and not w796;
w867 <= not w794 and w866;
w868 <= not w798 and not w867;
w869 <= not w865 and w868;
w870 <= not w798 and not w869;
w871 <= b(7) and not w787;
w872 <= not w785 and w871;
w873 <= not w789 and not w872;
w874 <= not w870 and w873;
w875 <= not w789 and not w874;
w876 <= b(8) and not w767;
w877 <= not w765 and w876;
w878 <= not w780 and not w877;
w879 <= not w875 and w878;
w880 <= not w780 and not w879;
w881 <= b(9) and not w777;
w882 <= not w775 and w881;
w883 <= not w779 and not w882;
w884 <= not w880 and w883;
w885 <= not w779 and not w884;
w886 <= w6 and w17;
w887 <= w87 and w886;
w888 <= w175 and w887;
w889 <= not w885 and w888;
w890 <= not w768 and not w889;
w891 <= not w789 and w878;
w892 <= not w874 and w891;
w893 <= not w875 and not w878;
w894 <= not w892 and not w893;
w895 <= w888 and not w894;
w896 <= not w885 and w895;
w897 <= not w890 and not w896;
w898 <= not w778 and not w889;
w899 <= not w780 and w883;
w900 <= not w879 and w899;
w901 <= not w880 and not w883;
w902 <= not w900 and not w901;
w903 <= w889 and not w902;
w904 <= not w898 and not w903;
w905 <= not b(10) and not w904;
w906 <= not b(9) and not w897;
w907 <= not w788 and not w889;
w908 <= not w798 and w873;
w909 <= not w869 and w908;
w910 <= not w870 and not w873;
w911 <= not w909 and not w910;
w912 <= w888 and not w911;
w913 <= not w885 and w912;
w914 <= not w907 and not w913;
w915 <= not b(8) and not w914;
w916 <= not w797 and not w889;
w917 <= not w807 and w868;
w918 <= not w864 and w917;
w919 <= not w865 and not w868;
w920 <= not w918 and not w919;
w921 <= w888 and not w920;
w922 <= not w885 and w921;
w923 <= not w916 and not w922;
w924 <= not b(7) and not w923;
w925 <= not w806 and not w889;
w926 <= not w816 and w863;
w927 <= not w859 and w926;
w928 <= not w860 and not w863;
w929 <= not w927 and not w928;
w930 <= w888 and not w929;
w931 <= not w885 and w930;
w932 <= not w925 and not w931;
w933 <= not b(6) and not w932;
w934 <= not w815 and not w889;
w935 <= not w825 and w858;
w936 <= not w854 and w935;
w937 <= not w855 and not w858;
w938 <= not w936 and not w937;
w939 <= w888 and not w938;
w940 <= not w885 and w939;
w941 <= not w934 and not w940;
w942 <= not b(5) and not w941;
w943 <= not w824 and not w889;
w944 <= not w833 and w853;
w945 <= not w849 and w944;
w946 <= not w850 and not w853;
w947 <= not w945 and not w946;
w948 <= w888 and not w947;
w949 <= not w885 and w948;
w950 <= not w943 and not w949;
w951 <= not b(4) and not w950;
w952 <= not w832 and not w889;
w953 <= not w844 and w848;
w954 <= not w843 and w953;
w955 <= not w845 and not w848;
w956 <= not w954 and not w955;
w957 <= w888 and not w956;
w958 <= not w885 and w957;
w959 <= not w952 and not w958;
w960 <= not b(3) and not w959;
w961 <= not w837 and not w889;
w962 <= not w840 and w842;
w963 <= not w838 and w962;
w964 <= w888 and not w963;
w965 <= not w843 and w964;
w966 <= not w885 and w965;
w967 <= not w961 and not w966;
w968 <= not b(2) and not w967;
w969 <= b(0) and not b(10);
w970 <= w133 and w969;
w971 <= w131 and w970;
w972 <= w121 and w971;
w973 <= w167 and w972;
w974 <= not w885 and w973;
w975 <= a(54) and not w974;
w976 <= w6 and w842;
w977 <= w17 and w976;
w978 <= w87 and w977;
w979 <= w175 and w978;
w980 <= not w885 and w979;
w981 <= not w975 and not w980;
w982 <= b(1) and not w981;
w983 <= not b(1) and not w980;
w984 <= not w975 and w983;
w985 <= not w982 and not w984;
w986 <= not a(53) and b(0);
w987 <= not w985 and not w986;
w988 <= not b(1) and not w981;
w989 <= not w987 and not w988;
w990 <= b(2) and not w966;
w991 <= not w961 and w990;
w992 <= not w968 and not w991;
w993 <= not w989 and w992;
w994 <= not w968 and not w993;
w995 <= b(3) and not w958;
w996 <= not w952 and w995;
w997 <= not w960 and not w996;
w998 <= not w994 and w997;
w999 <= not w960 and not w998;
w1000 <= b(4) and not w949;
w1001 <= not w943 and w1000;
w1002 <= not w951 and not w1001;
w1003 <= not w999 and w1002;
w1004 <= not w951 and not w1003;
w1005 <= b(5) and not w940;
w1006 <= not w934 and w1005;
w1007 <= not w942 and not w1006;
w1008 <= not w1004 and w1007;
w1009 <= not w942 and not w1008;
w1010 <= b(6) and not w931;
w1011 <= not w925 and w1010;
w1012 <= not w933 and not w1011;
w1013 <= not w1009 and w1012;
w1014 <= not w933 and not w1013;
w1015 <= b(7) and not w922;
w1016 <= not w916 and w1015;
w1017 <= not w924 and not w1016;
w1018 <= not w1014 and w1017;
w1019 <= not w924 and not w1018;
w1020 <= b(8) and not w913;
w1021 <= not w907 and w1020;
w1022 <= not w915 and not w1021;
w1023 <= not w1019 and w1022;
w1024 <= not w915 and not w1023;
w1025 <= b(9) and not w896;
w1026 <= not w890 and w1025;
w1027 <= not w906 and not w1026;
w1028 <= not w1024 and w1027;
w1029 <= not w906 and not w1028;
w1030 <= b(10) and not w898;
w1031 <= not w903 and w1030;
w1032 <= not w905 and not w1031;
w1033 <= not w1029 and w1032;
w1034 <= not w905 and not w1033;
w1035 <= w131 and w133;
w1036 <= w121 and w1035;
w1037 <= w167 and w1036;
w1038 <= not w1034 and w1037;
w1039 <= not w897 and not w1038;
w1040 <= not w915 and w1027;
w1041 <= not w1023 and w1040;
w1042 <= not w1024 and not w1027;
w1043 <= not w1041 and not w1042;
w1044 <= w1037 and not w1043;
w1045 <= not w1034 and w1044;
w1046 <= not w1039 and not w1045;
w1047 <= not b(10) and not w1046;
w1048 <= not w914 and not w1038;
w1049 <= not w924 and w1022;
w1050 <= not w1018 and w1049;
w1051 <= not w1019 and not w1022;
w1052 <= not w1050 and not w1051;
w1053 <= w1037 and not w1052;
w1054 <= not w1034 and w1053;
w1055 <= not w1048 and not w1054;
w1056 <= not b(9) and not w1055;
w1057 <= not w923 and not w1038;
w1058 <= not w933 and w1017;
w1059 <= not w1013 and w1058;
w1060 <= not w1014 and not w1017;
w1061 <= not w1059 and not w1060;
w1062 <= w1037 and not w1061;
w1063 <= not w1034 and w1062;
w1064 <= not w1057 and not w1063;
w1065 <= not b(8) and not w1064;
w1066 <= not w932 and not w1038;
w1067 <= not w942 and w1012;
w1068 <= not w1008 and w1067;
w1069 <= not w1009 and not w1012;
w1070 <= not w1068 and not w1069;
w1071 <= w1037 and not w1070;
w1072 <= not w1034 and w1071;
w1073 <= not w1066 and not w1072;
w1074 <= not b(7) and not w1073;
w1075 <= not w941 and not w1038;
w1076 <= not w951 and w1007;
w1077 <= not w1003 and w1076;
w1078 <= not w1004 and not w1007;
w1079 <= not w1077 and not w1078;
w1080 <= w1037 and not w1079;
w1081 <= not w1034 and w1080;
w1082 <= not w1075 and not w1081;
w1083 <= not b(6) and not w1082;
w1084 <= not w950 and not w1038;
w1085 <= not w960 and w1002;
w1086 <= not w998 and w1085;
w1087 <= not w999 and not w1002;
w1088 <= not w1086 and not w1087;
w1089 <= w1037 and not w1088;
w1090 <= not w1034 and w1089;
w1091 <= not w1084 and not w1090;
w1092 <= not b(5) and not w1091;
w1093 <= not w959 and not w1038;
w1094 <= not w968 and w997;
w1095 <= not w993 and w1094;
w1096 <= not w994 and not w997;
w1097 <= not w1095 and not w1096;
w1098 <= w1037 and not w1097;
w1099 <= not w1034 and w1098;
w1100 <= not w1093 and not w1099;
w1101 <= not b(4) and not w1100;
w1102 <= not w967 and not w1038;
w1103 <= not w988 and w992;
w1104 <= not w987 and w1103;
w1105 <= not w989 and not w992;
w1106 <= not w1104 and not w1105;
w1107 <= w1037 and not w1106;
w1108 <= not w1034 and w1107;
w1109 <= not w1102 and not w1108;
w1110 <= not b(3) and not w1109;
w1111 <= not w981 and not w1038;
w1112 <= not w984 and w986;
w1113 <= not w982 and w1112;
w1114 <= w1037 and not w1113;
w1115 <= not w987 and w1114;
w1116 <= not w1034 and w1115;
w1117 <= not w1111 and not w1116;
w1118 <= not b(2) and not w1117;
w1119 <= b(0) and not b(11);
w1120 <= w17 and w1119;
w1121 <= w87 and w1120;
w1122 <= w175 and w1121;
w1123 <= not w1034 and w1122;
w1124 <= a(53) and not w1123;
w1125 <= w133 and w986;
w1126 <= w131 and w1125;
w1127 <= w121 and w1126;
w1128 <= w167 and w1127;
w1129 <= not w1034 and w1128;
w1130 <= not w1124 and not w1129;
w1131 <= b(1) and not w1130;
w1132 <= not b(1) and not w1129;
w1133 <= not w1124 and w1132;
w1134 <= not w1131 and not w1133;
w1135 <= not a(52) and b(0);
w1136 <= not w1134 and not w1135;
w1137 <= not b(1) and not w1130;
w1138 <= not w1136 and not w1137;
w1139 <= b(2) and not w1116;
w1140 <= not w1111 and w1139;
w1141 <= not w1118 and not w1140;
w1142 <= not w1138 and w1141;
w1143 <= not w1118 and not w1142;
w1144 <= b(3) and not w1108;
w1145 <= not w1102 and w1144;
w1146 <= not w1110 and not w1145;
w1147 <= not w1143 and w1146;
w1148 <= not w1110 and not w1147;
w1149 <= b(4) and not w1099;
w1150 <= not w1093 and w1149;
w1151 <= not w1101 and not w1150;
w1152 <= not w1148 and w1151;
w1153 <= not w1101 and not w1152;
w1154 <= b(5) and not w1090;
w1155 <= not w1084 and w1154;
w1156 <= not w1092 and not w1155;
w1157 <= not w1153 and w1156;
w1158 <= not w1092 and not w1157;
w1159 <= b(6) and not w1081;
w1160 <= not w1075 and w1159;
w1161 <= not w1083 and not w1160;
w1162 <= not w1158 and w1161;
w1163 <= not w1083 and not w1162;
w1164 <= b(7) and not w1072;
w1165 <= not w1066 and w1164;
w1166 <= not w1074 and not w1165;
w1167 <= not w1163 and w1166;
w1168 <= not w1074 and not w1167;
w1169 <= b(8) and not w1063;
w1170 <= not w1057 and w1169;
w1171 <= not w1065 and not w1170;
w1172 <= not w1168 and w1171;
w1173 <= not w1065 and not w1172;
w1174 <= b(9) and not w1054;
w1175 <= not w1048 and w1174;
w1176 <= not w1056 and not w1175;
w1177 <= not w1173 and w1176;
w1178 <= not w1056 and not w1177;
w1179 <= b(10) and not w1045;
w1180 <= not w1039 and w1179;
w1181 <= not w1047 and not w1180;
w1182 <= not w1178 and w1181;
w1183 <= not w1047 and not w1182;
w1184 <= not w904 and not w1038;
w1185 <= not w906 and w1032;
w1186 <= not w1028 and w1185;
w1187 <= not w1029 and not w1032;
w1188 <= not w1186 and not w1187;
w1189 <= w1038 and not w1188;
w1190 <= not w1184 and not w1189;
w1191 <= not b(11) and not w1190;
w1192 <= b(11) and not w1184;
w1193 <= not w1189 and w1192;
w1194 <= w18 and w61;
w1195 <= w255 and w1194;
w1196 <= not w1193 and w1195;
w1197 <= not w1191 and w1196;
w1198 <= not w1183 and w1197;
w1199 <= w1037 and not w1190;
w1200 <= not w1198 and not w1199;
w1201 <= not w1056 and w1181;
w1202 <= not w1177 and w1201;
w1203 <= not w1178 and not w1181;
w1204 <= not w1202 and not w1203;
w1205 <= not w1200 and not w1204;
w1206 <= not w1046 and not w1199;
w1207 <= not w1198 and w1206;
w1208 <= not w1205 and not w1207;
w1209 <= not w1047 and not w1193;
w1210 <= not w1191 and w1209;
w1211 <= not w1182 and w1210;
w1212 <= not w1191 and not w1193;
w1213 <= not w1183 and not w1212;
w1214 <= not w1211 and not w1213;
w1215 <= not w1200 and not w1214;
w1216 <= not w1190 and not w1199;
w1217 <= not w1198 and w1216;
w1218 <= not w1215 and not w1217;
w1219 <= not b(12) and not w1218;
w1220 <= not b(11) and not w1208;
w1221 <= not w1065 and w1176;
w1222 <= not w1172 and w1221;
w1223 <= not w1173 and not w1176;
w1224 <= not w1222 and not w1223;
w1225 <= not w1200 and not w1224;
w1226 <= not w1055 and not w1199;
w1227 <= not w1198 and w1226;
w1228 <= not w1225 and not w1227;
w1229 <= not b(10) and not w1228;
w1230 <= not w1074 and w1171;
w1231 <= not w1167 and w1230;
w1232 <= not w1168 and not w1171;
w1233 <= not w1231 and not w1232;
w1234 <= not w1200 and not w1233;
w1235 <= not w1064 and not w1199;
w1236 <= not w1198 and w1235;
w1237 <= not w1234 and not w1236;
w1238 <= not b(9) and not w1237;
w1239 <= not w1083 and w1166;
w1240 <= not w1162 and w1239;
w1241 <= not w1163 and not w1166;
w1242 <= not w1240 and not w1241;
w1243 <= not w1200 and not w1242;
w1244 <= not w1073 and not w1199;
w1245 <= not w1198 and w1244;
w1246 <= not w1243 and not w1245;
w1247 <= not b(8) and not w1246;
w1248 <= not w1092 and w1161;
w1249 <= not w1157 and w1248;
w1250 <= not w1158 and not w1161;
w1251 <= not w1249 and not w1250;
w1252 <= not w1200 and not w1251;
w1253 <= not w1082 and not w1199;
w1254 <= not w1198 and w1253;
w1255 <= not w1252 and not w1254;
w1256 <= not b(7) and not w1255;
w1257 <= not w1101 and w1156;
w1258 <= not w1152 and w1257;
w1259 <= not w1153 and not w1156;
w1260 <= not w1258 and not w1259;
w1261 <= not w1200 and not w1260;
w1262 <= not w1091 and not w1199;
w1263 <= not w1198 and w1262;
w1264 <= not w1261 and not w1263;
w1265 <= not b(6) and not w1264;
w1266 <= not w1110 and w1151;
w1267 <= not w1147 and w1266;
w1268 <= not w1148 and not w1151;
w1269 <= not w1267 and not w1268;
w1270 <= not w1200 and not w1269;
w1271 <= not w1100 and not w1199;
w1272 <= not w1198 and w1271;
w1273 <= not w1270 and not w1272;
w1274 <= not b(5) and not w1273;
w1275 <= not w1118 and w1146;
w1276 <= not w1142 and w1275;
w1277 <= not w1143 and not w1146;
w1278 <= not w1276 and not w1277;
w1279 <= not w1200 and not w1278;
w1280 <= not w1109 and not w1199;
w1281 <= not w1198 and w1280;
w1282 <= not w1279 and not w1281;
w1283 <= not b(4) and not w1282;
w1284 <= not w1137 and w1141;
w1285 <= not w1136 and w1284;
w1286 <= not w1138 and not w1141;
w1287 <= not w1285 and not w1286;
w1288 <= not w1200 and not w1287;
w1289 <= not w1117 and not w1199;
w1290 <= not w1198 and w1289;
w1291 <= not w1288 and not w1290;
w1292 <= not b(3) and not w1291;
w1293 <= not w1133 and w1135;
w1294 <= not w1131 and w1293;
w1295 <= not w1136 and not w1294;
w1296 <= not w1200 and w1295;
w1297 <= not w1130 and not w1199;
w1298 <= not w1198 and w1297;
w1299 <= not w1296 and not w1298;
w1300 <= not b(2) and not w1299;
w1301 <= b(0) and not w1200;
w1302 <= a(52) and not w1301;
w1303 <= w1135 and not w1200;
w1304 <= not w1302 and not w1303;
w1305 <= b(1) and not w1304;
w1306 <= not b(1) and not w1303;
w1307 <= not w1302 and w1306;
w1308 <= not w1305 and not w1307;
w1309 <= not a(51) and b(0);
w1310 <= not w1308 and not w1309;
w1311 <= not b(1) and not w1304;
w1312 <= not w1310 and not w1311;
w1313 <= b(2) and not w1298;
w1314 <= not w1296 and w1313;
w1315 <= not w1300 and not w1314;
w1316 <= not w1312 and w1315;
w1317 <= not w1300 and not w1316;
w1318 <= b(3) and not w1290;
w1319 <= not w1288 and w1318;
w1320 <= not w1292 and not w1319;
w1321 <= not w1317 and w1320;
w1322 <= not w1292 and not w1321;
w1323 <= b(4) and not w1281;
w1324 <= not w1279 and w1323;
w1325 <= not w1283 and not w1324;
w1326 <= not w1322 and w1325;
w1327 <= not w1283 and not w1326;
w1328 <= b(5) and not w1272;
w1329 <= not w1270 and w1328;
w1330 <= not w1274 and not w1329;
w1331 <= not w1327 and w1330;
w1332 <= not w1274 and not w1331;
w1333 <= b(6) and not w1263;
w1334 <= not w1261 and w1333;
w1335 <= not w1265 and not w1334;
w1336 <= not w1332 and w1335;
w1337 <= not w1265 and not w1336;
w1338 <= b(7) and not w1254;
w1339 <= not w1252 and w1338;
w1340 <= not w1256 and not w1339;
w1341 <= not w1337 and w1340;
w1342 <= not w1256 and not w1341;
w1343 <= b(8) and not w1245;
w1344 <= not w1243 and w1343;
w1345 <= not w1247 and not w1344;
w1346 <= not w1342 and w1345;
w1347 <= not w1247 and not w1346;
w1348 <= b(9) and not w1236;
w1349 <= not w1234 and w1348;
w1350 <= not w1238 and not w1349;
w1351 <= not w1347 and w1350;
w1352 <= not w1238 and not w1351;
w1353 <= b(10) and not w1227;
w1354 <= not w1225 and w1353;
w1355 <= not w1229 and not w1354;
w1356 <= not w1352 and w1355;
w1357 <= not w1229 and not w1356;
w1358 <= b(11) and not w1207;
w1359 <= not w1205 and w1358;
w1360 <= not w1220 and not w1359;
w1361 <= not w1357 and w1360;
w1362 <= not w1220 and not w1361;
w1363 <= b(12) and not w1217;
w1364 <= not w1215 and w1363;
w1365 <= not w1219 and not w1364;
w1366 <= not w1362 and w1365;
w1367 <= not w1219 and not w1366;
w1368 <= w332 and w334;
w1369 <= w342 and w1368;
w1370 <= not w1367 and w1369;
w1371 <= not w1208 and not w1370;
w1372 <= not w1229 and w1360;
w1373 <= not w1356 and w1372;
w1374 <= not w1357 and not w1360;
w1375 <= not w1373 and not w1374;
w1376 <= w1369 and not w1375;
w1377 <= not w1367 and w1376;
w1378 <= not w1371 and not w1377;
w1379 <= not w1218 and not w1370;
w1380 <= not w1220 and w1365;
w1381 <= not w1361 and w1380;
w1382 <= not w1362 and not w1365;
w1383 <= not w1381 and not w1382;
w1384 <= w1370 and not w1383;
w1385 <= not w1379 and not w1384;
w1386 <= not b(13) and not w1385;
w1387 <= not b(12) and not w1378;
w1388 <= not w1228 and not w1370;
w1389 <= not w1238 and w1355;
w1390 <= not w1351 and w1389;
w1391 <= not w1352 and not w1355;
w1392 <= not w1390 and not w1391;
w1393 <= w1369 and not w1392;
w1394 <= not w1367 and w1393;
w1395 <= not w1388 and not w1394;
w1396 <= not b(11) and not w1395;
w1397 <= not w1237 and not w1370;
w1398 <= not w1247 and w1350;
w1399 <= not w1346 and w1398;
w1400 <= not w1347 and not w1350;
w1401 <= not w1399 and not w1400;
w1402 <= w1369 and not w1401;
w1403 <= not w1367 and w1402;
w1404 <= not w1397 and not w1403;
w1405 <= not b(10) and not w1404;
w1406 <= not w1246 and not w1370;
w1407 <= not w1256 and w1345;
w1408 <= not w1341 and w1407;
w1409 <= not w1342 and not w1345;
w1410 <= not w1408 and not w1409;
w1411 <= w1369 and not w1410;
w1412 <= not w1367 and w1411;
w1413 <= not w1406 and not w1412;
w1414 <= not b(9) and not w1413;
w1415 <= not w1255 and not w1370;
w1416 <= not w1265 and w1340;
w1417 <= not w1336 and w1416;
w1418 <= not w1337 and not w1340;
w1419 <= not w1417 and not w1418;
w1420 <= w1369 and not w1419;
w1421 <= not w1367 and w1420;
w1422 <= not w1415 and not w1421;
w1423 <= not b(8) and not w1422;
w1424 <= not w1264 and not w1370;
w1425 <= not w1274 and w1335;
w1426 <= not w1331 and w1425;
w1427 <= not w1332 and not w1335;
w1428 <= not w1426 and not w1427;
w1429 <= w1369 and not w1428;
w1430 <= not w1367 and w1429;
w1431 <= not w1424 and not w1430;
w1432 <= not b(7) and not w1431;
w1433 <= not w1273 and not w1370;
w1434 <= not w1283 and w1330;
w1435 <= not w1326 and w1434;
w1436 <= not w1327 and not w1330;
w1437 <= not w1435 and not w1436;
w1438 <= w1369 and not w1437;
w1439 <= not w1367 and w1438;
w1440 <= not w1433 and not w1439;
w1441 <= not b(6) and not w1440;
w1442 <= not w1282 and not w1370;
w1443 <= not w1292 and w1325;
w1444 <= not w1321 and w1443;
w1445 <= not w1322 and not w1325;
w1446 <= not w1444 and not w1445;
w1447 <= w1369 and not w1446;
w1448 <= not w1367 and w1447;
w1449 <= not w1442 and not w1448;
w1450 <= not b(5) and not w1449;
w1451 <= not w1291 and not w1370;
w1452 <= not w1300 and w1320;
w1453 <= not w1316 and w1452;
w1454 <= not w1317 and not w1320;
w1455 <= not w1453 and not w1454;
w1456 <= w1369 and not w1455;
w1457 <= not w1367 and w1456;
w1458 <= not w1451 and not w1457;
w1459 <= not b(4) and not w1458;
w1460 <= not w1299 and not w1370;
w1461 <= not w1311 and w1315;
w1462 <= not w1310 and w1461;
w1463 <= not w1312 and not w1315;
w1464 <= not w1462 and not w1463;
w1465 <= w1369 and not w1464;
w1466 <= not w1367 and w1465;
w1467 <= not w1460 and not w1466;
w1468 <= not b(3) and not w1467;
w1469 <= not w1304 and not w1370;
w1470 <= not w1307 and w1309;
w1471 <= not w1305 and w1470;
w1472 <= w1369 and not w1471;
w1473 <= not w1310 and w1472;
w1474 <= not w1367 and w1473;
w1475 <= not w1469 and not w1474;
w1476 <= not b(2) and not w1475;
w1477 <= b(0) and not b(13);
w1478 <= w16 and w1477;
w1479 <= w14 and w1478;
w1480 <= w61 and w1479;
w1481 <= w255 and w1480;
w1482 <= not w1367 and w1481;
w1483 <= a(51) and not w1482;
w1484 <= w131 and w1309;
w1485 <= w121 and w1484;
w1486 <= w167 and w1485;
w1487 <= not w1367 and w1486;
w1488 <= not w1483 and not w1487;
w1489 <= b(1) and not w1488;
w1490 <= not b(1) and not w1487;
w1491 <= not w1483 and w1490;
w1492 <= not w1489 and not w1491;
w1493 <= not a(50) and b(0);
w1494 <= not w1492 and not w1493;
w1495 <= not b(1) and not w1488;
w1496 <= not w1494 and not w1495;
w1497 <= b(2) and not w1474;
w1498 <= not w1469 and w1497;
w1499 <= not w1476 and not w1498;
w1500 <= not w1496 and w1499;
w1501 <= not w1476 and not w1500;
w1502 <= b(3) and not w1466;
w1503 <= not w1460 and w1502;
w1504 <= not w1468 and not w1503;
w1505 <= not w1501 and w1504;
w1506 <= not w1468 and not w1505;
w1507 <= b(4) and not w1457;
w1508 <= not w1451 and w1507;
w1509 <= not w1459 and not w1508;
w1510 <= not w1506 and w1509;
w1511 <= not w1459 and not w1510;
w1512 <= b(5) and not w1448;
w1513 <= not w1442 and w1512;
w1514 <= not w1450 and not w1513;
w1515 <= not w1511 and w1514;
w1516 <= not w1450 and not w1515;
w1517 <= b(6) and not w1439;
w1518 <= not w1433 and w1517;
w1519 <= not w1441 and not w1518;
w1520 <= not w1516 and w1519;
w1521 <= not w1441 and not w1520;
w1522 <= b(7) and not w1430;
w1523 <= not w1424 and w1522;
w1524 <= not w1432 and not w1523;
w1525 <= not w1521 and w1524;
w1526 <= not w1432 and not w1525;
w1527 <= b(8) and not w1421;
w1528 <= not w1415 and w1527;
w1529 <= not w1423 and not w1528;
w1530 <= not w1526 and w1529;
w1531 <= not w1423 and not w1530;
w1532 <= b(9) and not w1412;
w1533 <= not w1406 and w1532;
w1534 <= not w1414 and not w1533;
w1535 <= not w1531 and w1534;
w1536 <= not w1414 and not w1535;
w1537 <= b(10) and not w1403;
w1538 <= not w1397 and w1537;
w1539 <= not w1405 and not w1538;
w1540 <= not w1536 and w1539;
w1541 <= not w1405 and not w1540;
w1542 <= b(11) and not w1394;
w1543 <= not w1388 and w1542;
w1544 <= not w1396 and not w1543;
w1545 <= not w1541 and w1544;
w1546 <= not w1396 and not w1545;
w1547 <= b(12) and not w1377;
w1548 <= not w1371 and w1547;
w1549 <= not w1387 and not w1548;
w1550 <= not w1546 and w1549;
w1551 <= not w1387 and not w1550;
w1552 <= b(13) and not w1379;
w1553 <= not w1384 and w1552;
w1554 <= not w1386 and not w1553;
w1555 <= not w1551 and w1554;
w1556 <= not w1386 and not w1555;
w1557 <= w14 and w16;
w1558 <= w61 and w1557;
w1559 <= w255 and w1558;
w1560 <= not w1556 and w1559;
w1561 <= not w1378 and not w1560;
w1562 <= not w1396 and w1549;
w1563 <= not w1545 and w1562;
w1564 <= not w1546 and not w1549;
w1565 <= not w1563 and not w1564;
w1566 <= w1559 and not w1565;
w1567 <= not w1556 and w1566;
w1568 <= not w1561 and not w1567;
w1569 <= not b(13) and not w1568;
w1570 <= not w1395 and not w1560;
w1571 <= not w1405 and w1544;
w1572 <= not w1540 and w1571;
w1573 <= not w1541 and not w1544;
w1574 <= not w1572 and not w1573;
w1575 <= w1559 and not w1574;
w1576 <= not w1556 and w1575;
w1577 <= not w1570 and not w1576;
w1578 <= not b(12) and not w1577;
w1579 <= not w1404 and not w1560;
w1580 <= not w1414 and w1539;
w1581 <= not w1535 and w1580;
w1582 <= not w1536 and not w1539;
w1583 <= not w1581 and not w1582;
w1584 <= w1559 and not w1583;
w1585 <= not w1556 and w1584;
w1586 <= not w1579 and not w1585;
w1587 <= not b(11) and not w1586;
w1588 <= not w1413 and not w1560;
w1589 <= not w1423 and w1534;
w1590 <= not w1530 and w1589;
w1591 <= not w1531 and not w1534;
w1592 <= not w1590 and not w1591;
w1593 <= w1559 and not w1592;
w1594 <= not w1556 and w1593;
w1595 <= not w1588 and not w1594;
w1596 <= not b(10) and not w1595;
w1597 <= not w1422 and not w1560;
w1598 <= not w1432 and w1529;
w1599 <= not w1525 and w1598;
w1600 <= not w1526 and not w1529;
w1601 <= not w1599 and not w1600;
w1602 <= w1559 and not w1601;
w1603 <= not w1556 and w1602;
w1604 <= not w1597 and not w1603;
w1605 <= not b(9) and not w1604;
w1606 <= not w1431 and not w1560;
w1607 <= not w1441 and w1524;
w1608 <= not w1520 and w1607;
w1609 <= not w1521 and not w1524;
w1610 <= not w1608 and not w1609;
w1611 <= w1559 and not w1610;
w1612 <= not w1556 and w1611;
w1613 <= not w1606 and not w1612;
w1614 <= not b(8) and not w1613;
w1615 <= not w1440 and not w1560;
w1616 <= not w1450 and w1519;
w1617 <= not w1515 and w1616;
w1618 <= not w1516 and not w1519;
w1619 <= not w1617 and not w1618;
w1620 <= w1559 and not w1619;
w1621 <= not w1556 and w1620;
w1622 <= not w1615 and not w1621;
w1623 <= not b(7) and not w1622;
w1624 <= not w1449 and not w1560;
w1625 <= not w1459 and w1514;
w1626 <= not w1510 and w1625;
w1627 <= not w1511 and not w1514;
w1628 <= not w1626 and not w1627;
w1629 <= w1559 and not w1628;
w1630 <= not w1556 and w1629;
w1631 <= not w1624 and not w1630;
w1632 <= not b(6) and not w1631;
w1633 <= not w1458 and not w1560;
w1634 <= not w1468 and w1509;
w1635 <= not w1505 and w1634;
w1636 <= not w1506 and not w1509;
w1637 <= not w1635 and not w1636;
w1638 <= w1559 and not w1637;
w1639 <= not w1556 and w1638;
w1640 <= not w1633 and not w1639;
w1641 <= not b(5) and not w1640;
w1642 <= not w1467 and not w1560;
w1643 <= not w1476 and w1504;
w1644 <= not w1500 and w1643;
w1645 <= not w1501 and not w1504;
w1646 <= not w1644 and not w1645;
w1647 <= w1559 and not w1646;
w1648 <= not w1556 and w1647;
w1649 <= not w1642 and not w1648;
w1650 <= not b(4) and not w1649;
w1651 <= not w1475 and not w1560;
w1652 <= not w1495 and w1499;
w1653 <= not w1494 and w1652;
w1654 <= not w1496 and not w1499;
w1655 <= not w1653 and not w1654;
w1656 <= w1559 and not w1655;
w1657 <= not w1556 and w1656;
w1658 <= not w1651 and not w1657;
w1659 <= not b(3) and not w1658;
w1660 <= not w1488 and not w1560;
w1661 <= not w1491 and w1493;
w1662 <= not w1489 and w1661;
w1663 <= w1559 and not w1662;
w1664 <= not w1494 and w1663;
w1665 <= not w1556 and w1664;
w1666 <= not w1660 and not w1665;
w1667 <= not b(2) and not w1666;
w1668 <= b(0) and not b(14);
w1669 <= w130 and w1668;
w1670 <= w112 and w1669;
w1671 <= w332 and w1670;
w1672 <= w342 and w1671;
w1673 <= not w1556 and w1672;
w1674 <= a(50) and not w1673;
w1675 <= w16 and w1493;
w1676 <= w14 and w1675;
w1677 <= w61 and w1676;
w1678 <= w255 and w1677;
w1679 <= not w1556 and w1678;
w1680 <= not w1674 and not w1679;
w1681 <= b(1) and not w1680;
w1682 <= not b(1) and not w1679;
w1683 <= not w1674 and w1682;
w1684 <= not w1681 and not w1683;
w1685 <= not a(49) and b(0);
w1686 <= not w1684 and not w1685;
w1687 <= not b(1) and not w1680;
w1688 <= not w1686 and not w1687;
w1689 <= b(2) and not w1665;
w1690 <= not w1660 and w1689;
w1691 <= not w1667 and not w1690;
w1692 <= not w1688 and w1691;
w1693 <= not w1667 and not w1692;
w1694 <= b(3) and not w1657;
w1695 <= not w1651 and w1694;
w1696 <= not w1659 and not w1695;
w1697 <= not w1693 and w1696;
w1698 <= not w1659 and not w1697;
w1699 <= b(4) and not w1648;
w1700 <= not w1642 and w1699;
w1701 <= not w1650 and not w1700;
w1702 <= not w1698 and w1701;
w1703 <= not w1650 and not w1702;
w1704 <= b(5) and not w1639;
w1705 <= not w1633 and w1704;
w1706 <= not w1641 and not w1705;
w1707 <= not w1703 and w1706;
w1708 <= not w1641 and not w1707;
w1709 <= b(6) and not w1630;
w1710 <= not w1624 and w1709;
w1711 <= not w1632 and not w1710;
w1712 <= not w1708 and w1711;
w1713 <= not w1632 and not w1712;
w1714 <= b(7) and not w1621;
w1715 <= not w1615 and w1714;
w1716 <= not w1623 and not w1715;
w1717 <= not w1713 and w1716;
w1718 <= not w1623 and not w1717;
w1719 <= b(8) and not w1612;
w1720 <= not w1606 and w1719;
w1721 <= not w1614 and not w1720;
w1722 <= not w1718 and w1721;
w1723 <= not w1614 and not w1722;
w1724 <= b(9) and not w1603;
w1725 <= not w1597 and w1724;
w1726 <= not w1605 and not w1725;
w1727 <= not w1723 and w1726;
w1728 <= not w1605 and not w1727;
w1729 <= b(10) and not w1594;
w1730 <= not w1588 and w1729;
w1731 <= not w1596 and not w1730;
w1732 <= not w1728 and w1731;
w1733 <= not w1596 and not w1732;
w1734 <= b(11) and not w1585;
w1735 <= not w1579 and w1734;
w1736 <= not w1587 and not w1735;
w1737 <= not w1733 and w1736;
w1738 <= not w1587 and not w1737;
w1739 <= b(12) and not w1576;
w1740 <= not w1570 and w1739;
w1741 <= not w1578 and not w1740;
w1742 <= not w1738 and w1741;
w1743 <= not w1578 and not w1742;
w1744 <= b(13) and not w1567;
w1745 <= not w1561 and w1744;
w1746 <= not w1569 and not w1745;
w1747 <= not w1743 and w1746;
w1748 <= not w1569 and not w1747;
w1749 <= not w1385 and not w1560;
w1750 <= not w1387 and w1554;
w1751 <= not w1550 and w1750;
w1752 <= not w1551 and not w1554;
w1753 <= not w1751 and not w1752;
w1754 <= w1560 and not w1753;
w1755 <= not w1749 and not w1754;
w1756 <= not b(14) and not w1755;
w1757 <= b(14) and not w1749;
w1758 <= not w1754 and w1757;
w1759 <= w112 and w130;
w1760 <= w332 and w1759;
w1761 <= w342 and w1760;
w1762 <= not w1758 and w1761;
w1763 <= not w1756 and w1762;
w1764 <= not w1748 and w1763;
w1765 <= w1559 and not w1755;
w1766 <= not w1764 and not w1765;
w1767 <= not w1578 and w1746;
w1768 <= not w1742 and w1767;
w1769 <= not w1743 and not w1746;
w1770 <= not w1768 and not w1769;
w1771 <= not w1766 and not w1770;
w1772 <= not w1568 and not w1765;
w1773 <= not w1764 and w1772;
w1774 <= not w1771 and not w1773;
w1775 <= not w1569 and not w1758;
w1776 <= not w1756 and w1775;
w1777 <= not w1747 and w1776;
w1778 <= not w1756 and not w1758;
w1779 <= not w1748 and not w1778;
w1780 <= not w1777 and not w1779;
w1781 <= not w1766 and not w1780;
w1782 <= not w1755 and not w1765;
w1783 <= not w1764 and w1782;
w1784 <= not w1781 and not w1783;
w1785 <= not b(15) and not w1784;
w1786 <= not b(14) and not w1774;
w1787 <= not w1587 and w1741;
w1788 <= not w1737 and w1787;
w1789 <= not w1738 and not w1741;
w1790 <= not w1788 and not w1789;
w1791 <= not w1766 and not w1790;
w1792 <= not w1577 and not w1765;
w1793 <= not w1764 and w1792;
w1794 <= not w1791 and not w1793;
w1795 <= not b(13) and not w1794;
w1796 <= not w1596 and w1736;
w1797 <= not w1732 and w1796;
w1798 <= not w1733 and not w1736;
w1799 <= not w1797 and not w1798;
w1800 <= not w1766 and not w1799;
w1801 <= not w1586 and not w1765;
w1802 <= not w1764 and w1801;
w1803 <= not w1800 and not w1802;
w1804 <= not b(12) and not w1803;
w1805 <= not w1605 and w1731;
w1806 <= not w1727 and w1805;
w1807 <= not w1728 and not w1731;
w1808 <= not w1806 and not w1807;
w1809 <= not w1766 and not w1808;
w1810 <= not w1595 and not w1765;
w1811 <= not w1764 and w1810;
w1812 <= not w1809 and not w1811;
w1813 <= not b(11) and not w1812;
w1814 <= not w1614 and w1726;
w1815 <= not w1722 and w1814;
w1816 <= not w1723 and not w1726;
w1817 <= not w1815 and not w1816;
w1818 <= not w1766 and not w1817;
w1819 <= not w1604 and not w1765;
w1820 <= not w1764 and w1819;
w1821 <= not w1818 and not w1820;
w1822 <= not b(10) and not w1821;
w1823 <= not w1623 and w1721;
w1824 <= not w1717 and w1823;
w1825 <= not w1718 and not w1721;
w1826 <= not w1824 and not w1825;
w1827 <= not w1766 and not w1826;
w1828 <= not w1613 and not w1765;
w1829 <= not w1764 and w1828;
w1830 <= not w1827 and not w1829;
w1831 <= not b(9) and not w1830;
w1832 <= not w1632 and w1716;
w1833 <= not w1712 and w1832;
w1834 <= not w1713 and not w1716;
w1835 <= not w1833 and not w1834;
w1836 <= not w1766 and not w1835;
w1837 <= not w1622 and not w1765;
w1838 <= not w1764 and w1837;
w1839 <= not w1836 and not w1838;
w1840 <= not b(8) and not w1839;
w1841 <= not w1641 and w1711;
w1842 <= not w1707 and w1841;
w1843 <= not w1708 and not w1711;
w1844 <= not w1842 and not w1843;
w1845 <= not w1766 and not w1844;
w1846 <= not w1631 and not w1765;
w1847 <= not w1764 and w1846;
w1848 <= not w1845 and not w1847;
w1849 <= not b(7) and not w1848;
w1850 <= not w1650 and w1706;
w1851 <= not w1702 and w1850;
w1852 <= not w1703 and not w1706;
w1853 <= not w1851 and not w1852;
w1854 <= not w1766 and not w1853;
w1855 <= not w1640 and not w1765;
w1856 <= not w1764 and w1855;
w1857 <= not w1854 and not w1856;
w1858 <= not b(6) and not w1857;
w1859 <= not w1659 and w1701;
w1860 <= not w1697 and w1859;
w1861 <= not w1698 and not w1701;
w1862 <= not w1860 and not w1861;
w1863 <= not w1766 and not w1862;
w1864 <= not w1649 and not w1765;
w1865 <= not w1764 and w1864;
w1866 <= not w1863 and not w1865;
w1867 <= not b(5) and not w1866;
w1868 <= not w1667 and w1696;
w1869 <= not w1692 and w1868;
w1870 <= not w1693 and not w1696;
w1871 <= not w1869 and not w1870;
w1872 <= not w1766 and not w1871;
w1873 <= not w1658 and not w1765;
w1874 <= not w1764 and w1873;
w1875 <= not w1872 and not w1874;
w1876 <= not b(4) and not w1875;
w1877 <= not w1687 and w1691;
w1878 <= not w1686 and w1877;
w1879 <= not w1688 and not w1691;
w1880 <= not w1878 and not w1879;
w1881 <= not w1766 and not w1880;
w1882 <= not w1666 and not w1765;
w1883 <= not w1764 and w1882;
w1884 <= not w1881 and not w1883;
w1885 <= not b(3) and not w1884;
w1886 <= not w1683 and w1685;
w1887 <= not w1681 and w1886;
w1888 <= not w1686 and not w1887;
w1889 <= not w1766 and w1888;
w1890 <= not w1680 and not w1765;
w1891 <= not w1764 and w1890;
w1892 <= not w1889 and not w1891;
w1893 <= not b(2) and not w1892;
w1894 <= b(0) and not w1766;
w1895 <= a(49) and not w1894;
w1896 <= w1685 and not w1766;
w1897 <= not w1895 and not w1896;
w1898 <= b(1) and not w1897;
w1899 <= not b(1) and not w1896;
w1900 <= not w1895 and w1899;
w1901 <= not w1898 and not w1900;
w1902 <= not a(48) and b(0);
w1903 <= not w1901 and not w1902;
w1904 <= not b(1) and not w1897;
w1905 <= not w1903 and not w1904;
w1906 <= b(2) and not w1891;
w1907 <= not w1889 and w1906;
w1908 <= not w1893 and not w1907;
w1909 <= not w1905 and w1908;
w1910 <= not w1893 and not w1909;
w1911 <= b(3) and not w1883;
w1912 <= not w1881 and w1911;
w1913 <= not w1885 and not w1912;
w1914 <= not w1910 and w1913;
w1915 <= not w1885 and not w1914;
w1916 <= b(4) and not w1874;
w1917 <= not w1872 and w1916;
w1918 <= not w1876 and not w1917;
w1919 <= not w1915 and w1918;
w1920 <= not w1876 and not w1919;
w1921 <= b(5) and not w1865;
w1922 <= not w1863 and w1921;
w1923 <= not w1867 and not w1922;
w1924 <= not w1920 and w1923;
w1925 <= not w1867 and not w1924;
w1926 <= b(6) and not w1856;
w1927 <= not w1854 and w1926;
w1928 <= not w1858 and not w1927;
w1929 <= not w1925 and w1928;
w1930 <= not w1858 and not w1929;
w1931 <= b(7) and not w1847;
w1932 <= not w1845 and w1931;
w1933 <= not w1849 and not w1932;
w1934 <= not w1930 and w1933;
w1935 <= not w1849 and not w1934;
w1936 <= b(8) and not w1838;
w1937 <= not w1836 and w1936;
w1938 <= not w1840 and not w1937;
w1939 <= not w1935 and w1938;
w1940 <= not w1840 and not w1939;
w1941 <= b(9) and not w1829;
w1942 <= not w1827 and w1941;
w1943 <= not w1831 and not w1942;
w1944 <= not w1940 and w1943;
w1945 <= not w1831 and not w1944;
w1946 <= b(10) and not w1820;
w1947 <= not w1818 and w1946;
w1948 <= not w1822 and not w1947;
w1949 <= not w1945 and w1948;
w1950 <= not w1822 and not w1949;
w1951 <= b(11) and not w1811;
w1952 <= not w1809 and w1951;
w1953 <= not w1813 and not w1952;
w1954 <= not w1950 and w1953;
w1955 <= not w1813 and not w1954;
w1956 <= b(12) and not w1802;
w1957 <= not w1800 and w1956;
w1958 <= not w1804 and not w1957;
w1959 <= not w1955 and w1958;
w1960 <= not w1804 and not w1959;
w1961 <= b(13) and not w1793;
w1962 <= not w1791 and w1961;
w1963 <= not w1795 and not w1962;
w1964 <= not w1960 and w1963;
w1965 <= not w1795 and not w1964;
w1966 <= b(14) and not w1773;
w1967 <= not w1771 and w1966;
w1968 <= not w1786 and not w1967;
w1969 <= not w1965 and w1968;
w1970 <= not w1786 and not w1969;
w1971 <= b(15) and not w1783;
w1972 <= not w1781 and w1971;
w1973 <= not w1785 and not w1972;
w1974 <= not w1970 and w1973;
w1975 <= not w1785 and not w1974;
w1976 <= w89 and not w1975;
w1977 <= not w1774 and not w1976;
w1978 <= not w1795 and w1968;
w1979 <= not w1964 and w1978;
w1980 <= not w1965 and not w1968;
w1981 <= not w1979 and not w1980;
w1982 <= w89 and not w1981;
w1983 <= not w1975 and w1982;
w1984 <= not w1977 and not w1983;
w1985 <= not w1784 and not w1976;
w1986 <= not w1786 and w1973;
w1987 <= not w1969 and w1986;
w1988 <= not w1970 and not w1973;
w1989 <= not w1987 and not w1988;
w1990 <= w1976 and not w1989;
w1991 <= not w1985 and not w1990;
w1992 <= not b(16) and not w1991;
w1993 <= not b(15) and not w1984;
w1994 <= not w1794 and not w1976;
w1995 <= not w1804 and w1963;
w1996 <= not w1959 and w1995;
w1997 <= not w1960 and not w1963;
w1998 <= not w1996 and not w1997;
w1999 <= w89 and not w1998;
w2000 <= not w1975 and w1999;
w2001 <= not w1994 and not w2000;
w2002 <= not b(14) and not w2001;
w2003 <= not w1803 and not w1976;
w2004 <= not w1813 and w1958;
w2005 <= not w1954 and w2004;
w2006 <= not w1955 and not w1958;
w2007 <= not w2005 and not w2006;
w2008 <= w89 and not w2007;
w2009 <= not w1975 and w2008;
w2010 <= not w2003 and not w2009;
w2011 <= not b(13) and not w2010;
w2012 <= not w1812 and not w1976;
w2013 <= not w1822 and w1953;
w2014 <= not w1949 and w2013;
w2015 <= not w1950 and not w1953;
w2016 <= not w2014 and not w2015;
w2017 <= w89 and not w2016;
w2018 <= not w1975 and w2017;
w2019 <= not w2012 and not w2018;
w2020 <= not b(12) and not w2019;
w2021 <= not w1821 and not w1976;
w2022 <= not w1831 and w1948;
w2023 <= not w1944 and w2022;
w2024 <= not w1945 and not w1948;
w2025 <= not w2023 and not w2024;
w2026 <= w89 and not w2025;
w2027 <= not w1975 and w2026;
w2028 <= not w2021 and not w2027;
w2029 <= not b(11) and not w2028;
w2030 <= not w1830 and not w1976;
w2031 <= not w1840 and w1943;
w2032 <= not w1939 and w2031;
w2033 <= not w1940 and not w1943;
w2034 <= not w2032 and not w2033;
w2035 <= w89 and not w2034;
w2036 <= not w1975 and w2035;
w2037 <= not w2030 and not w2036;
w2038 <= not b(10) and not w2037;
w2039 <= not w1839 and not w1976;
w2040 <= not w1849 and w1938;
w2041 <= not w1934 and w2040;
w2042 <= not w1935 and not w1938;
w2043 <= not w2041 and not w2042;
w2044 <= w89 and not w2043;
w2045 <= not w1975 and w2044;
w2046 <= not w2039 and not w2045;
w2047 <= not b(9) and not w2046;
w2048 <= not w1848 and not w1976;
w2049 <= not w1858 and w1933;
w2050 <= not w1929 and w2049;
w2051 <= not w1930 and not w1933;
w2052 <= not w2050 and not w2051;
w2053 <= w89 and not w2052;
w2054 <= not w1975 and w2053;
w2055 <= not w2048 and not w2054;
w2056 <= not b(8) and not w2055;
w2057 <= not w1857 and not w1976;
w2058 <= not w1867 and w1928;
w2059 <= not w1924 and w2058;
w2060 <= not w1925 and not w1928;
w2061 <= not w2059 and not w2060;
w2062 <= w89 and not w2061;
w2063 <= not w1975 and w2062;
w2064 <= not w2057 and not w2063;
w2065 <= not b(7) and not w2064;
w2066 <= not w1866 and not w1976;
w2067 <= not w1876 and w1923;
w2068 <= not w1919 and w2067;
w2069 <= not w1920 and not w1923;
w2070 <= not w2068 and not w2069;
w2071 <= w89 and not w2070;
w2072 <= not w1975 and w2071;
w2073 <= not w2066 and not w2072;
w2074 <= not b(6) and not w2073;
w2075 <= not w1875 and not w1976;
w2076 <= not w1885 and w1918;
w2077 <= not w1914 and w2076;
w2078 <= not w1915 and not w1918;
w2079 <= not w2077 and not w2078;
w2080 <= w89 and not w2079;
w2081 <= not w1975 and w2080;
w2082 <= not w2075 and not w2081;
w2083 <= not b(5) and not w2082;
w2084 <= not w1884 and not w1976;
w2085 <= not w1893 and w1913;
w2086 <= not w1909 and w2085;
w2087 <= not w1910 and not w1913;
w2088 <= not w2086 and not w2087;
w2089 <= w89 and not w2088;
w2090 <= not w1975 and w2089;
w2091 <= not w2084 and not w2090;
w2092 <= not b(4) and not w2091;
w2093 <= not w1892 and not w1976;
w2094 <= not w1904 and w1908;
w2095 <= not w1903 and w2094;
w2096 <= not w1905 and not w1908;
w2097 <= not w2095 and not w2096;
w2098 <= w89 and not w2097;
w2099 <= not w1975 and w2098;
w2100 <= not w2093 and not w2099;
w2101 <= not b(3) and not w2100;
w2102 <= not w1897 and not w1976;
w2103 <= not w1900 and w1902;
w2104 <= not w1898 and w2103;
w2105 <= w89 and not w2104;
w2106 <= not w1903 and w2105;
w2107 <= not w1975 and w2106;
w2108 <= not w2102 and not w2107;
w2109 <= not b(2) and not w2108;
w2110 <= b(0) and not b(16);
w2111 <= w112 and w2110;
w2112 <= w332 and w2111;
w2113 <= w342 and w2112;
w2114 <= not w1975 and w2113;
w2115 <= a(48) and not w2114;
w2116 <= w14 and w1902;
w2117 <= w61 and w2116;
w2118 <= w255 and w2117;
w2119 <= not w1975 and w2118;
w2120 <= not w2115 and not w2119;
w2121 <= b(1) and not w2120;
w2122 <= not b(1) and not w2119;
w2123 <= not w2115 and w2122;
w2124 <= not w2121 and not w2123;
w2125 <= not a(47) and b(0);
w2126 <= not w2124 and not w2125;
w2127 <= not b(1) and not w2120;
w2128 <= not w2126 and not w2127;
w2129 <= b(2) and not w2107;
w2130 <= not w2102 and w2129;
w2131 <= not w2109 and not w2130;
w2132 <= not w2128 and w2131;
w2133 <= not w2109 and not w2132;
w2134 <= b(3) and not w2099;
w2135 <= not w2093 and w2134;
w2136 <= not w2101 and not w2135;
w2137 <= not w2133 and w2136;
w2138 <= not w2101 and not w2137;
w2139 <= b(4) and not w2090;
w2140 <= not w2084 and w2139;
w2141 <= not w2092 and not w2140;
w2142 <= not w2138 and w2141;
w2143 <= not w2092 and not w2142;
w2144 <= b(5) and not w2081;
w2145 <= not w2075 and w2144;
w2146 <= not w2083 and not w2145;
w2147 <= not w2143 and w2146;
w2148 <= not w2083 and not w2147;
w2149 <= b(6) and not w2072;
w2150 <= not w2066 and w2149;
w2151 <= not w2074 and not w2150;
w2152 <= not w2148 and w2151;
w2153 <= not w2074 and not w2152;
w2154 <= b(7) and not w2063;
w2155 <= not w2057 and w2154;
w2156 <= not w2065 and not w2155;
w2157 <= not w2153 and w2156;
w2158 <= not w2065 and not w2157;
w2159 <= b(8) and not w2054;
w2160 <= not w2048 and w2159;
w2161 <= not w2056 and not w2160;
w2162 <= not w2158 and w2161;
w2163 <= not w2056 and not w2162;
w2164 <= b(9) and not w2045;
w2165 <= not w2039 and w2164;
w2166 <= not w2047 and not w2165;
w2167 <= not w2163 and w2166;
w2168 <= not w2047 and not w2167;
w2169 <= b(10) and not w2036;
w2170 <= not w2030 and w2169;
w2171 <= not w2038 and not w2170;
w2172 <= not w2168 and w2171;
w2173 <= not w2038 and not w2172;
w2174 <= b(11) and not w2027;
w2175 <= not w2021 and w2174;
w2176 <= not w2029 and not w2175;
w2177 <= not w2173 and w2176;
w2178 <= not w2029 and not w2177;
w2179 <= b(12) and not w2018;
w2180 <= not w2012 and w2179;
w2181 <= not w2020 and not w2180;
w2182 <= not w2178 and w2181;
w2183 <= not w2020 and not w2182;
w2184 <= b(13) and not w2009;
w2185 <= not w2003 and w2184;
w2186 <= not w2011 and not w2185;
w2187 <= not w2183 and w2186;
w2188 <= not w2011 and not w2187;
w2189 <= b(14) and not w2000;
w2190 <= not w1994 and w2189;
w2191 <= not w2002 and not w2190;
w2192 <= not w2188 and w2191;
w2193 <= not w2002 and not w2192;
w2194 <= b(15) and not w1983;
w2195 <= not w1977 and w2194;
w2196 <= not w1993 and not w2195;
w2197 <= not w2193 and w2196;
w2198 <= not w1993 and not w2197;
w2199 <= b(16) and not w1985;
w2200 <= not w1990 and w2199;
w2201 <= not w1992 and not w2200;
w2202 <= not w2198 and w2201;
w2203 <= not w1992 and not w2202;
w2204 <= w218 and not w2203;
w2205 <= not w1984 and not w2204;
w2206 <= not w2002 and w2196;
w2207 <= not w2192 and w2206;
w2208 <= not w2193 and not w2196;
w2209 <= not w2207 and not w2208;
w2210 <= w218 and not w2209;
w2211 <= not w2203 and w2210;
w2212 <= not w2205 and not w2211;
w2213 <= not b(16) and not w2212;
w2214 <= not w2001 and not w2204;
w2215 <= not w2011 and w2191;
w2216 <= not w2187 and w2215;
w2217 <= not w2188 and not w2191;
w2218 <= not w2216 and not w2217;
w2219 <= w218 and not w2218;
w2220 <= not w2203 and w2219;
w2221 <= not w2214 and not w2220;
w2222 <= not b(15) and not w2221;
w2223 <= not w2010 and not w2204;
w2224 <= not w2020 and w2186;
w2225 <= not w2182 and w2224;
w2226 <= not w2183 and not w2186;
w2227 <= not w2225 and not w2226;
w2228 <= w218 and not w2227;
w2229 <= not w2203 and w2228;
w2230 <= not w2223 and not w2229;
w2231 <= not b(14) and not w2230;
w2232 <= not w2019 and not w2204;
w2233 <= not w2029 and w2181;
w2234 <= not w2177 and w2233;
w2235 <= not w2178 and not w2181;
w2236 <= not w2234 and not w2235;
w2237 <= w218 and not w2236;
w2238 <= not w2203 and w2237;
w2239 <= not w2232 and not w2238;
w2240 <= not b(13) and not w2239;
w2241 <= not w2028 and not w2204;
w2242 <= not w2038 and w2176;
w2243 <= not w2172 and w2242;
w2244 <= not w2173 and not w2176;
w2245 <= not w2243 and not w2244;
w2246 <= w218 and not w2245;
w2247 <= not w2203 and w2246;
w2248 <= not w2241 and not w2247;
w2249 <= not b(12) and not w2248;
w2250 <= not w2037 and not w2204;
w2251 <= not w2047 and w2171;
w2252 <= not w2167 and w2251;
w2253 <= not w2168 and not w2171;
w2254 <= not w2252 and not w2253;
w2255 <= w218 and not w2254;
w2256 <= not w2203 and w2255;
w2257 <= not w2250 and not w2256;
w2258 <= not b(11) and not w2257;
w2259 <= not w2046 and not w2204;
w2260 <= not w2056 and w2166;
w2261 <= not w2162 and w2260;
w2262 <= not w2163 and not w2166;
w2263 <= not w2261 and not w2262;
w2264 <= w218 and not w2263;
w2265 <= not w2203 and w2264;
w2266 <= not w2259 and not w2265;
w2267 <= not b(10) and not w2266;
w2268 <= not w2055 and not w2204;
w2269 <= not w2065 and w2161;
w2270 <= not w2157 and w2269;
w2271 <= not w2158 and not w2161;
w2272 <= not w2270 and not w2271;
w2273 <= w218 and not w2272;
w2274 <= not w2203 and w2273;
w2275 <= not w2268 and not w2274;
w2276 <= not b(9) and not w2275;
w2277 <= not w2064 and not w2204;
w2278 <= not w2074 and w2156;
w2279 <= not w2152 and w2278;
w2280 <= not w2153 and not w2156;
w2281 <= not w2279 and not w2280;
w2282 <= w218 and not w2281;
w2283 <= not w2203 and w2282;
w2284 <= not w2277 and not w2283;
w2285 <= not b(8) and not w2284;
w2286 <= not w2073 and not w2204;
w2287 <= not w2083 and w2151;
w2288 <= not w2147 and w2287;
w2289 <= not w2148 and not w2151;
w2290 <= not w2288 and not w2289;
w2291 <= w218 and not w2290;
w2292 <= not w2203 and w2291;
w2293 <= not w2286 and not w2292;
w2294 <= not b(7) and not w2293;
w2295 <= not w2082 and not w2204;
w2296 <= not w2092 and w2146;
w2297 <= not w2142 and w2296;
w2298 <= not w2143 and not w2146;
w2299 <= not w2297 and not w2298;
w2300 <= w218 and not w2299;
w2301 <= not w2203 and w2300;
w2302 <= not w2295 and not w2301;
w2303 <= not b(6) and not w2302;
w2304 <= not w2091 and not w2204;
w2305 <= not w2101 and w2141;
w2306 <= not w2137 and w2305;
w2307 <= not w2138 and not w2141;
w2308 <= not w2306 and not w2307;
w2309 <= w218 and not w2308;
w2310 <= not w2203 and w2309;
w2311 <= not w2304 and not w2310;
w2312 <= not b(5) and not w2311;
w2313 <= not w2100 and not w2204;
w2314 <= not w2109 and w2136;
w2315 <= not w2132 and w2314;
w2316 <= not w2133 and not w2136;
w2317 <= not w2315 and not w2316;
w2318 <= w218 and not w2317;
w2319 <= not w2203 and w2318;
w2320 <= not w2313 and not w2319;
w2321 <= not b(4) and not w2320;
w2322 <= not w2108 and not w2204;
w2323 <= not w2127 and w2131;
w2324 <= not w2126 and w2323;
w2325 <= not w2128 and not w2131;
w2326 <= not w2324 and not w2325;
w2327 <= w218 and not w2326;
w2328 <= not w2203 and w2327;
w2329 <= not w2322 and not w2328;
w2330 <= not b(3) and not w2329;
w2331 <= not w2120 and not w2204;
w2332 <= not w2123 and w2125;
w2333 <= not w2121 and w2332;
w2334 <= w218 and not w2333;
w2335 <= not w2126 and w2334;
w2336 <= not w2203 and w2335;
w2337 <= not w2331 and not w2336;
w2338 <= not b(2) and not w2337;
w2339 <= b(0) and not b(17);
w2340 <= w13 and w2339;
w2341 <= w52 and w2340;
w2342 <= w86 and w2341;
w2343 <= w84 and w2342;
w2344 <= w81 and w2343;
w2345 <= not w2203 and w2344;
w2346 <= a(47) and not w2345;
w2347 <= w112 and w2125;
w2348 <= w332 and w2347;
w2349 <= w342 and w2348;
w2350 <= not w2203 and w2349;
w2351 <= not w2346 and not w2350;
w2352 <= b(1) and not w2351;
w2353 <= not b(1) and not w2350;
w2354 <= not w2346 and w2353;
w2355 <= not w2352 and not w2354;
w2356 <= not a(46) and b(0);
w2357 <= not w2355 and not w2356;
w2358 <= not b(1) and not w2351;
w2359 <= not w2357 and not w2358;
w2360 <= b(2) and not w2336;
w2361 <= not w2331 and w2360;
w2362 <= not w2338 and not w2361;
w2363 <= not w2359 and w2362;
w2364 <= not w2338 and not w2363;
w2365 <= b(3) and not w2328;
w2366 <= not w2322 and w2365;
w2367 <= not w2330 and not w2366;
w2368 <= not w2364 and w2367;
w2369 <= not w2330 and not w2368;
w2370 <= b(4) and not w2319;
w2371 <= not w2313 and w2370;
w2372 <= not w2321 and not w2371;
w2373 <= not w2369 and w2372;
w2374 <= not w2321 and not w2373;
w2375 <= b(5) and not w2310;
w2376 <= not w2304 and w2375;
w2377 <= not w2312 and not w2376;
w2378 <= not w2374 and w2377;
w2379 <= not w2312 and not w2378;
w2380 <= b(6) and not w2301;
w2381 <= not w2295 and w2380;
w2382 <= not w2303 and not w2381;
w2383 <= not w2379 and w2382;
w2384 <= not w2303 and not w2383;
w2385 <= b(7) and not w2292;
w2386 <= not w2286 and w2385;
w2387 <= not w2294 and not w2386;
w2388 <= not w2384 and w2387;
w2389 <= not w2294 and not w2388;
w2390 <= b(8) and not w2283;
w2391 <= not w2277 and w2390;
w2392 <= not w2285 and not w2391;
w2393 <= not w2389 and w2392;
w2394 <= not w2285 and not w2393;
w2395 <= b(9) and not w2274;
w2396 <= not w2268 and w2395;
w2397 <= not w2276 and not w2396;
w2398 <= not w2394 and w2397;
w2399 <= not w2276 and not w2398;
w2400 <= b(10) and not w2265;
w2401 <= not w2259 and w2400;
w2402 <= not w2267 and not w2401;
w2403 <= not w2399 and w2402;
w2404 <= not w2267 and not w2403;
w2405 <= b(11) and not w2256;
w2406 <= not w2250 and w2405;
w2407 <= not w2258 and not w2406;
w2408 <= not w2404 and w2407;
w2409 <= not w2258 and not w2408;
w2410 <= b(12) and not w2247;
w2411 <= not w2241 and w2410;
w2412 <= not w2249 and not w2411;
w2413 <= not w2409 and w2412;
w2414 <= not w2249 and not w2413;
w2415 <= b(13) and not w2238;
w2416 <= not w2232 and w2415;
w2417 <= not w2240 and not w2416;
w2418 <= not w2414 and w2417;
w2419 <= not w2240 and not w2418;
w2420 <= b(14) and not w2229;
w2421 <= not w2223 and w2420;
w2422 <= not w2231 and not w2421;
w2423 <= not w2419 and w2422;
w2424 <= not w2231 and not w2423;
w2425 <= b(15) and not w2220;
w2426 <= not w2214 and w2425;
w2427 <= not w2222 and not w2426;
w2428 <= not w2424 and w2427;
w2429 <= not w2222 and not w2428;
w2430 <= b(16) and not w2211;
w2431 <= not w2205 and w2430;
w2432 <= not w2213 and not w2431;
w2433 <= not w2429 and w2432;
w2434 <= not w2213 and not w2433;
w2435 <= not w1991 and not w2204;
w2436 <= not w1993 and w2201;
w2437 <= not w2197 and w2436;
w2438 <= not w2198 and not w2201;
w2439 <= not w2437 and not w2438;
w2440 <= w2204 and not w2439;
w2441 <= not w2435 and not w2440;
w2442 <= not b(17) and not w2441;
w2443 <= b(17) and not w2435;
w2444 <= not w2440 and w2443;
w2445 <= w13 and w52;
w2446 <= w86 and w2445;
w2447 <= w84 and w2446;
w2448 <= w81 and w2447;
w2449 <= not w2444 and w2448;
w2450 <= not w2442 and w2449;
w2451 <= not w2434 and w2450;
w2452 <= w218 and not w2441;
w2453 <= not w2451 and not w2452;
w2454 <= not w2222 and w2432;
w2455 <= not w2428 and w2454;
w2456 <= not w2429 and not w2432;
w2457 <= not w2455 and not w2456;
w2458 <= not w2453 and not w2457;
w2459 <= not w2212 and not w2452;
w2460 <= not w2451 and w2459;
w2461 <= not w2458 and not w2460;
w2462 <= not w2213 and not w2444;
w2463 <= not w2442 and w2462;
w2464 <= not w2433 and w2463;
w2465 <= not w2442 and not w2444;
w2466 <= not w2434 and not w2465;
w2467 <= not w2464 and not w2466;
w2468 <= not w2453 and not w2467;
w2469 <= not w2441 and not w2452;
w2470 <= not w2451 and w2469;
w2471 <= not w2468 and not w2470;
w2472 <= not b(18) and not w2471;
w2473 <= not b(17) and not w2461;
w2474 <= not w2231 and w2427;
w2475 <= not w2423 and w2474;
w2476 <= not w2424 and not w2427;
w2477 <= not w2475 and not w2476;
w2478 <= not w2453 and not w2477;
w2479 <= not w2221 and not w2452;
w2480 <= not w2451 and w2479;
w2481 <= not w2478 and not w2480;
w2482 <= not b(16) and not w2481;
w2483 <= not w2240 and w2422;
w2484 <= not w2418 and w2483;
w2485 <= not w2419 and not w2422;
w2486 <= not w2484 and not w2485;
w2487 <= not w2453 and not w2486;
w2488 <= not w2230 and not w2452;
w2489 <= not w2451 and w2488;
w2490 <= not w2487 and not w2489;
w2491 <= not b(15) and not w2490;
w2492 <= not w2249 and w2417;
w2493 <= not w2413 and w2492;
w2494 <= not w2414 and not w2417;
w2495 <= not w2493 and not w2494;
w2496 <= not w2453 and not w2495;
w2497 <= not w2239 and not w2452;
w2498 <= not w2451 and w2497;
w2499 <= not w2496 and not w2498;
w2500 <= not b(14) and not w2499;
w2501 <= not w2258 and w2412;
w2502 <= not w2408 and w2501;
w2503 <= not w2409 and not w2412;
w2504 <= not w2502 and not w2503;
w2505 <= not w2453 and not w2504;
w2506 <= not w2248 and not w2452;
w2507 <= not w2451 and w2506;
w2508 <= not w2505 and not w2507;
w2509 <= not b(13) and not w2508;
w2510 <= not w2267 and w2407;
w2511 <= not w2403 and w2510;
w2512 <= not w2404 and not w2407;
w2513 <= not w2511 and not w2512;
w2514 <= not w2453 and not w2513;
w2515 <= not w2257 and not w2452;
w2516 <= not w2451 and w2515;
w2517 <= not w2514 and not w2516;
w2518 <= not b(12) and not w2517;
w2519 <= not w2276 and w2402;
w2520 <= not w2398 and w2519;
w2521 <= not w2399 and not w2402;
w2522 <= not w2520 and not w2521;
w2523 <= not w2453 and not w2522;
w2524 <= not w2266 and not w2452;
w2525 <= not w2451 and w2524;
w2526 <= not w2523 and not w2525;
w2527 <= not b(11) and not w2526;
w2528 <= not w2285 and w2397;
w2529 <= not w2393 and w2528;
w2530 <= not w2394 and not w2397;
w2531 <= not w2529 and not w2530;
w2532 <= not w2453 and not w2531;
w2533 <= not w2275 and not w2452;
w2534 <= not w2451 and w2533;
w2535 <= not w2532 and not w2534;
w2536 <= not b(10) and not w2535;
w2537 <= not w2294 and w2392;
w2538 <= not w2388 and w2537;
w2539 <= not w2389 and not w2392;
w2540 <= not w2538 and not w2539;
w2541 <= not w2453 and not w2540;
w2542 <= not w2284 and not w2452;
w2543 <= not w2451 and w2542;
w2544 <= not w2541 and not w2543;
w2545 <= not b(9) and not w2544;
w2546 <= not w2303 and w2387;
w2547 <= not w2383 and w2546;
w2548 <= not w2384 and not w2387;
w2549 <= not w2547 and not w2548;
w2550 <= not w2453 and not w2549;
w2551 <= not w2293 and not w2452;
w2552 <= not w2451 and w2551;
w2553 <= not w2550 and not w2552;
w2554 <= not b(8) and not w2553;
w2555 <= not w2312 and w2382;
w2556 <= not w2378 and w2555;
w2557 <= not w2379 and not w2382;
w2558 <= not w2556 and not w2557;
w2559 <= not w2453 and not w2558;
w2560 <= not w2302 and not w2452;
w2561 <= not w2451 and w2560;
w2562 <= not w2559 and not w2561;
w2563 <= not b(7) and not w2562;
w2564 <= not w2321 and w2377;
w2565 <= not w2373 and w2564;
w2566 <= not w2374 and not w2377;
w2567 <= not w2565 and not w2566;
w2568 <= not w2453 and not w2567;
w2569 <= not w2311 and not w2452;
w2570 <= not w2451 and w2569;
w2571 <= not w2568 and not w2570;
w2572 <= not b(6) and not w2571;
w2573 <= not w2330 and w2372;
w2574 <= not w2368 and w2573;
w2575 <= not w2369 and not w2372;
w2576 <= not w2574 and not w2575;
w2577 <= not w2453 and not w2576;
w2578 <= not w2320 and not w2452;
w2579 <= not w2451 and w2578;
w2580 <= not w2577 and not w2579;
w2581 <= not b(5) and not w2580;
w2582 <= not w2338 and w2367;
w2583 <= not w2363 and w2582;
w2584 <= not w2364 and not w2367;
w2585 <= not w2583 and not w2584;
w2586 <= not w2453 and not w2585;
w2587 <= not w2329 and not w2452;
w2588 <= not w2451 and w2587;
w2589 <= not w2586 and not w2588;
w2590 <= not b(4) and not w2589;
w2591 <= not w2358 and w2362;
w2592 <= not w2357 and w2591;
w2593 <= not w2359 and not w2362;
w2594 <= not w2592 and not w2593;
w2595 <= not w2453 and not w2594;
w2596 <= not w2337 and not w2452;
w2597 <= not w2451 and w2596;
w2598 <= not w2595 and not w2597;
w2599 <= not b(3) and not w2598;
w2600 <= not w2354 and w2356;
w2601 <= not w2352 and w2600;
w2602 <= not w2357 and not w2601;
w2603 <= not w2453 and w2602;
w2604 <= not w2351 and not w2452;
w2605 <= not w2451 and w2604;
w2606 <= not w2603 and not w2605;
w2607 <= not b(2) and not w2606;
w2608 <= b(0) and not w2453;
w2609 <= a(46) and not w2608;
w2610 <= w2356 and not w2453;
w2611 <= not w2609 and not w2610;
w2612 <= b(1) and not w2611;
w2613 <= not b(1) and not w2610;
w2614 <= not w2609 and w2613;
w2615 <= not w2612 and not w2614;
w2616 <= not a(45) and b(0);
w2617 <= not w2615 and not w2616;
w2618 <= not b(1) and not w2611;
w2619 <= not w2617 and not w2618;
w2620 <= b(2) and not w2605;
w2621 <= not w2603 and w2620;
w2622 <= not w2607 and not w2621;
w2623 <= not w2619 and w2622;
w2624 <= not w2607 and not w2623;
w2625 <= b(3) and not w2597;
w2626 <= not w2595 and w2625;
w2627 <= not w2599 and not w2626;
w2628 <= not w2624 and w2627;
w2629 <= not w2599 and not w2628;
w2630 <= b(4) and not w2588;
w2631 <= not w2586 and w2630;
w2632 <= not w2590 and not w2631;
w2633 <= not w2629 and w2632;
w2634 <= not w2590 and not w2633;
w2635 <= b(5) and not w2579;
w2636 <= not w2577 and w2635;
w2637 <= not w2581 and not w2636;
w2638 <= not w2634 and w2637;
w2639 <= not w2581 and not w2638;
w2640 <= b(6) and not w2570;
w2641 <= not w2568 and w2640;
w2642 <= not w2572 and not w2641;
w2643 <= not w2639 and w2642;
w2644 <= not w2572 and not w2643;
w2645 <= b(7) and not w2561;
w2646 <= not w2559 and w2645;
w2647 <= not w2563 and not w2646;
w2648 <= not w2644 and w2647;
w2649 <= not w2563 and not w2648;
w2650 <= b(8) and not w2552;
w2651 <= not w2550 and w2650;
w2652 <= not w2554 and not w2651;
w2653 <= not w2649 and w2652;
w2654 <= not w2554 and not w2653;
w2655 <= b(9) and not w2543;
w2656 <= not w2541 and w2655;
w2657 <= not w2545 and not w2656;
w2658 <= not w2654 and w2657;
w2659 <= not w2545 and not w2658;
w2660 <= b(10) and not w2534;
w2661 <= not w2532 and w2660;
w2662 <= not w2536 and not w2661;
w2663 <= not w2659 and w2662;
w2664 <= not w2536 and not w2663;
w2665 <= b(11) and not w2525;
w2666 <= not w2523 and w2665;
w2667 <= not w2527 and not w2666;
w2668 <= not w2664 and w2667;
w2669 <= not w2527 and not w2668;
w2670 <= b(12) and not w2516;
w2671 <= not w2514 and w2670;
w2672 <= not w2518 and not w2671;
w2673 <= not w2669 and w2672;
w2674 <= not w2518 and not w2673;
w2675 <= b(13) and not w2507;
w2676 <= not w2505 and w2675;
w2677 <= not w2509 and not w2676;
w2678 <= not w2674 and w2677;
w2679 <= not w2509 and not w2678;
w2680 <= b(14) and not w2498;
w2681 <= not w2496 and w2680;
w2682 <= not w2500 and not w2681;
w2683 <= not w2679 and w2682;
w2684 <= not w2500 and not w2683;
w2685 <= b(15) and not w2489;
w2686 <= not w2487 and w2685;
w2687 <= not w2491 and not w2686;
w2688 <= not w2684 and w2687;
w2689 <= not w2491 and not w2688;
w2690 <= b(16) and not w2480;
w2691 <= not w2478 and w2690;
w2692 <= not w2482 and not w2691;
w2693 <= not w2689 and w2692;
w2694 <= not w2482 and not w2693;
w2695 <= b(17) and not w2460;
w2696 <= not w2458 and w2695;
w2697 <= not w2473 and not w2696;
w2698 <= not w2694 and w2697;
w2699 <= not w2473 and not w2698;
w2700 <= b(18) and not w2470;
w2701 <= not w2468 and w2700;
w2702 <= not w2472 and not w2701;
w2703 <= not w2699 and w2702;
w2704 <= not w2472 and not w2703;
w2705 <= w109 and w111;
w2706 <= w120 and w2705;
w2707 <= w166 and w2706;
w2708 <= w151 and w2707;
w2709 <= not w2704 and w2708;
w2710 <= not w2461 and not w2709;
w2711 <= not w2482 and w2697;
w2712 <= not w2693 and w2711;
w2713 <= not w2694 and not w2697;
w2714 <= not w2712 and not w2713;
w2715 <= w2708 and not w2714;
w2716 <= not w2704 and w2715;
w2717 <= not w2710 and not w2716;
w2718 <= not w2471 and not w2709;
w2719 <= not w2473 and w2702;
w2720 <= not w2698 and w2719;
w2721 <= not w2699 and not w2702;
w2722 <= not w2720 and not w2721;
w2723 <= w2709 and not w2722;
w2724 <= not w2718 and not w2723;
w2725 <= not b(19) and not w2724;
w2726 <= not b(18) and not w2717;
w2727 <= not w2481 and not w2709;
w2728 <= not w2491 and w2692;
w2729 <= not w2688 and w2728;
w2730 <= not w2689 and not w2692;
w2731 <= not w2729 and not w2730;
w2732 <= w2708 and not w2731;
w2733 <= not w2704 and w2732;
w2734 <= not w2727 and not w2733;
w2735 <= not b(17) and not w2734;
w2736 <= not w2490 and not w2709;
w2737 <= not w2500 and w2687;
w2738 <= not w2683 and w2737;
w2739 <= not w2684 and not w2687;
w2740 <= not w2738 and not w2739;
w2741 <= w2708 and not w2740;
w2742 <= not w2704 and w2741;
w2743 <= not w2736 and not w2742;
w2744 <= not b(16) and not w2743;
w2745 <= not w2499 and not w2709;
w2746 <= not w2509 and w2682;
w2747 <= not w2678 and w2746;
w2748 <= not w2679 and not w2682;
w2749 <= not w2747 and not w2748;
w2750 <= w2708 and not w2749;
w2751 <= not w2704 and w2750;
w2752 <= not w2745 and not w2751;
w2753 <= not b(15) and not w2752;
w2754 <= not w2508 and not w2709;
w2755 <= not w2518 and w2677;
w2756 <= not w2673 and w2755;
w2757 <= not w2674 and not w2677;
w2758 <= not w2756 and not w2757;
w2759 <= w2708 and not w2758;
w2760 <= not w2704 and w2759;
w2761 <= not w2754 and not w2760;
w2762 <= not b(14) and not w2761;
w2763 <= not w2517 and not w2709;
w2764 <= not w2527 and w2672;
w2765 <= not w2668 and w2764;
w2766 <= not w2669 and not w2672;
w2767 <= not w2765 and not w2766;
w2768 <= w2708 and not w2767;
w2769 <= not w2704 and w2768;
w2770 <= not w2763 and not w2769;
w2771 <= not b(13) and not w2770;
w2772 <= not w2526 and not w2709;
w2773 <= not w2536 and w2667;
w2774 <= not w2663 and w2773;
w2775 <= not w2664 and not w2667;
w2776 <= not w2774 and not w2775;
w2777 <= w2708 and not w2776;
w2778 <= not w2704 and w2777;
w2779 <= not w2772 and not w2778;
w2780 <= not b(12) and not w2779;
w2781 <= not w2535 and not w2709;
w2782 <= not w2545 and w2662;
w2783 <= not w2658 and w2782;
w2784 <= not w2659 and not w2662;
w2785 <= not w2783 and not w2784;
w2786 <= w2708 and not w2785;
w2787 <= not w2704 and w2786;
w2788 <= not w2781 and not w2787;
w2789 <= not b(11) and not w2788;
w2790 <= not w2544 and not w2709;
w2791 <= not w2554 and w2657;
w2792 <= not w2653 and w2791;
w2793 <= not w2654 and not w2657;
w2794 <= not w2792 and not w2793;
w2795 <= w2708 and not w2794;
w2796 <= not w2704 and w2795;
w2797 <= not w2790 and not w2796;
w2798 <= not b(10) and not w2797;
w2799 <= not w2553 and not w2709;
w2800 <= not w2563 and w2652;
w2801 <= not w2648 and w2800;
w2802 <= not w2649 and not w2652;
w2803 <= not w2801 and not w2802;
w2804 <= w2708 and not w2803;
w2805 <= not w2704 and w2804;
w2806 <= not w2799 and not w2805;
w2807 <= not b(9) and not w2806;
w2808 <= not w2562 and not w2709;
w2809 <= not w2572 and w2647;
w2810 <= not w2643 and w2809;
w2811 <= not w2644 and not w2647;
w2812 <= not w2810 and not w2811;
w2813 <= w2708 and not w2812;
w2814 <= not w2704 and w2813;
w2815 <= not w2808 and not w2814;
w2816 <= not b(8) and not w2815;
w2817 <= not w2571 and not w2709;
w2818 <= not w2581 and w2642;
w2819 <= not w2638 and w2818;
w2820 <= not w2639 and not w2642;
w2821 <= not w2819 and not w2820;
w2822 <= w2708 and not w2821;
w2823 <= not w2704 and w2822;
w2824 <= not w2817 and not w2823;
w2825 <= not b(7) and not w2824;
w2826 <= not w2580 and not w2709;
w2827 <= not w2590 and w2637;
w2828 <= not w2633 and w2827;
w2829 <= not w2634 and not w2637;
w2830 <= not w2828 and not w2829;
w2831 <= w2708 and not w2830;
w2832 <= not w2704 and w2831;
w2833 <= not w2826 and not w2832;
w2834 <= not b(6) and not w2833;
w2835 <= not w2589 and not w2709;
w2836 <= not w2599 and w2632;
w2837 <= not w2628 and w2836;
w2838 <= not w2629 and not w2632;
w2839 <= not w2837 and not w2838;
w2840 <= w2708 and not w2839;
w2841 <= not w2704 and w2840;
w2842 <= not w2835 and not w2841;
w2843 <= not b(5) and not w2842;
w2844 <= not w2598 and not w2709;
w2845 <= not w2607 and w2627;
w2846 <= not w2623 and w2845;
w2847 <= not w2624 and not w2627;
w2848 <= not w2846 and not w2847;
w2849 <= w2708 and not w2848;
w2850 <= not w2704 and w2849;
w2851 <= not w2844 and not w2850;
w2852 <= not b(4) and not w2851;
w2853 <= not w2606 and not w2709;
w2854 <= not w2618 and w2622;
w2855 <= not w2617 and w2854;
w2856 <= not w2619 and not w2622;
w2857 <= not w2855 and not w2856;
w2858 <= w2708 and not w2857;
w2859 <= not w2704 and w2858;
w2860 <= not w2853 and not w2859;
w2861 <= not b(3) and not w2860;
w2862 <= not w2611 and not w2709;
w2863 <= not w2614 and w2616;
w2864 <= not w2612 and w2863;
w2865 <= w2708 and not w2864;
w2866 <= not w2617 and w2865;
w2867 <= not w2704 and w2866;
w2868 <= not w2862 and not w2867;
w2869 <= not b(2) and not w2868;
w2870 <= b(0) and not b(19);
w2871 <= w52 and w2870;
w2872 <= w86 and w2871;
w2873 <= w84 and w2872;
w2874 <= w81 and w2873;
w2875 <= not w2704 and w2874;
w2876 <= a(45) and not w2875;
w2877 <= w111 and w2616;
w2878 <= w109 and w2877;
w2879 <= w120 and w2878;
w2880 <= w166 and w2879;
w2881 <= w151 and w2880;
w2882 <= not w2704 and w2881;
w2883 <= not w2876 and not w2882;
w2884 <= b(1) and not w2883;
w2885 <= not b(1) and not w2882;
w2886 <= not w2876 and w2885;
w2887 <= not w2884 and not w2886;
w2888 <= not a(44) and b(0);
w2889 <= not w2887 and not w2888;
w2890 <= not b(1) and not w2883;
w2891 <= not w2889 and not w2890;
w2892 <= b(2) and not w2867;
w2893 <= not w2862 and w2892;
w2894 <= not w2869 and not w2893;
w2895 <= not w2891 and w2894;
w2896 <= not w2869 and not w2895;
w2897 <= b(3) and not w2859;
w2898 <= not w2853 and w2897;
w2899 <= not w2861 and not w2898;
w2900 <= not w2896 and w2899;
w2901 <= not w2861 and not w2900;
w2902 <= b(4) and not w2850;
w2903 <= not w2844 and w2902;
w2904 <= not w2852 and not w2903;
w2905 <= not w2901 and w2904;
w2906 <= not w2852 and not w2905;
w2907 <= b(5) and not w2841;
w2908 <= not w2835 and w2907;
w2909 <= not w2843 and not w2908;
w2910 <= not w2906 and w2909;
w2911 <= not w2843 and not w2910;
w2912 <= b(6) and not w2832;
w2913 <= not w2826 and w2912;
w2914 <= not w2834 and not w2913;
w2915 <= not w2911 and w2914;
w2916 <= not w2834 and not w2915;
w2917 <= b(7) and not w2823;
w2918 <= not w2817 and w2917;
w2919 <= not w2825 and not w2918;
w2920 <= not w2916 and w2919;
w2921 <= not w2825 and not w2920;
w2922 <= b(8) and not w2814;
w2923 <= not w2808 and w2922;
w2924 <= not w2816 and not w2923;
w2925 <= not w2921 and w2924;
w2926 <= not w2816 and not w2925;
w2927 <= b(9) and not w2805;
w2928 <= not w2799 and w2927;
w2929 <= not w2807 and not w2928;
w2930 <= not w2926 and w2929;
w2931 <= not w2807 and not w2930;
w2932 <= b(10) and not w2796;
w2933 <= not w2790 and w2932;
w2934 <= not w2798 and not w2933;
w2935 <= not w2931 and w2934;
w2936 <= not w2798 and not w2935;
w2937 <= b(11) and not w2787;
w2938 <= not w2781 and w2937;
w2939 <= not w2789 and not w2938;
w2940 <= not w2936 and w2939;
w2941 <= not w2789 and not w2940;
w2942 <= b(12) and not w2778;
w2943 <= not w2772 and w2942;
w2944 <= not w2780 and not w2943;
w2945 <= not w2941 and w2944;
w2946 <= not w2780 and not w2945;
w2947 <= b(13) and not w2769;
w2948 <= not w2763 and w2947;
w2949 <= not w2771 and not w2948;
w2950 <= not w2946 and w2949;
w2951 <= not w2771 and not w2950;
w2952 <= b(14) and not w2760;
w2953 <= not w2754 and w2952;
w2954 <= not w2762 and not w2953;
w2955 <= not w2951 and w2954;
w2956 <= not w2762 and not w2955;
w2957 <= b(15) and not w2751;
w2958 <= not w2745 and w2957;
w2959 <= not w2753 and not w2958;
w2960 <= not w2956 and w2959;
w2961 <= not w2753 and not w2960;
w2962 <= b(16) and not w2742;
w2963 <= not w2736 and w2962;
w2964 <= not w2744 and not w2963;
w2965 <= not w2961 and w2964;
w2966 <= not w2744 and not w2965;
w2967 <= b(17) and not w2733;
w2968 <= not w2727 and w2967;
w2969 <= not w2735 and not w2968;
w2970 <= not w2966 and w2969;
w2971 <= not w2735 and not w2970;
w2972 <= b(18) and not w2716;
w2973 <= not w2710 and w2972;
w2974 <= not w2726 and not w2973;
w2975 <= not w2971 and w2974;
w2976 <= not w2726 and not w2975;
w2977 <= b(19) and not w2718;
w2978 <= not w2723 and w2977;
w2979 <= not w2725 and not w2978;
w2980 <= not w2976 and w2979;
w2981 <= not w2725 and not w2980;
w2982 <= w63 and not w2981;
w2983 <= not w2717 and not w2982;
w2984 <= not w2735 and w2974;
w2985 <= not w2970 and w2984;
w2986 <= not w2971 and not w2974;
w2987 <= not w2985 and not w2986;
w2988 <= w63 and not w2987;
w2989 <= not w2981 and w2988;
w2990 <= not w2983 and not w2989;
w2991 <= not b(19) and not w2990;
w2992 <= not w2734 and not w2982;
w2993 <= not w2744 and w2969;
w2994 <= not w2965 and w2993;
w2995 <= not w2966 and not w2969;
w2996 <= not w2994 and not w2995;
w2997 <= w63 and not w2996;
w2998 <= not w2981 and w2997;
w2999 <= not w2992 and not w2998;
w3000 <= not b(18) and not w2999;
w3001 <= not w2743 and not w2982;
w3002 <= not w2753 and w2964;
w3003 <= not w2960 and w3002;
w3004 <= not w2961 and not w2964;
w3005 <= not w3003 and not w3004;
w3006 <= w63 and not w3005;
w3007 <= not w2981 and w3006;
w3008 <= not w3001 and not w3007;
w3009 <= not b(17) and not w3008;
w3010 <= not w2752 and not w2982;
w3011 <= not w2762 and w2959;
w3012 <= not w2955 and w3011;
w3013 <= not w2956 and not w2959;
w3014 <= not w3012 and not w3013;
w3015 <= w63 and not w3014;
w3016 <= not w2981 and w3015;
w3017 <= not w3010 and not w3016;
w3018 <= not b(16) and not w3017;
w3019 <= not w2761 and not w2982;
w3020 <= not w2771 and w2954;
w3021 <= not w2950 and w3020;
w3022 <= not w2951 and not w2954;
w3023 <= not w3021 and not w3022;
w3024 <= w63 and not w3023;
w3025 <= not w2981 and w3024;
w3026 <= not w3019 and not w3025;
w3027 <= not b(15) and not w3026;
w3028 <= not w2770 and not w2982;
w3029 <= not w2780 and w2949;
w3030 <= not w2945 and w3029;
w3031 <= not w2946 and not w2949;
w3032 <= not w3030 and not w3031;
w3033 <= w63 and not w3032;
w3034 <= not w2981 and w3033;
w3035 <= not w3028 and not w3034;
w3036 <= not b(14) and not w3035;
w3037 <= not w2779 and not w2982;
w3038 <= not w2789 and w2944;
w3039 <= not w2940 and w3038;
w3040 <= not w2941 and not w2944;
w3041 <= not w3039 and not w3040;
w3042 <= w63 and not w3041;
w3043 <= not w2981 and w3042;
w3044 <= not w3037 and not w3043;
w3045 <= not b(13) and not w3044;
w3046 <= not w2788 and not w2982;
w3047 <= not w2798 and w2939;
w3048 <= not w2935 and w3047;
w3049 <= not w2936 and not w2939;
w3050 <= not w3048 and not w3049;
w3051 <= w63 and not w3050;
w3052 <= not w2981 and w3051;
w3053 <= not w3046 and not w3052;
w3054 <= not b(12) and not w3053;
w3055 <= not w2797 and not w2982;
w3056 <= not w2807 and w2934;
w3057 <= not w2930 and w3056;
w3058 <= not w2931 and not w2934;
w3059 <= not w3057 and not w3058;
w3060 <= w63 and not w3059;
w3061 <= not w2981 and w3060;
w3062 <= not w3055 and not w3061;
w3063 <= not b(11) and not w3062;
w3064 <= not w2806 and not w2982;
w3065 <= not w2816 and w2929;
w3066 <= not w2925 and w3065;
w3067 <= not w2926 and not w2929;
w3068 <= not w3066 and not w3067;
w3069 <= w63 and not w3068;
w3070 <= not w2981 and w3069;
w3071 <= not w3064 and not w3070;
w3072 <= not b(10) and not w3071;
w3073 <= not w2815 and not w2982;
w3074 <= not w2825 and w2924;
w3075 <= not w2920 and w3074;
w3076 <= not w2921 and not w2924;
w3077 <= not w3075 and not w3076;
w3078 <= w63 and not w3077;
w3079 <= not w2981 and w3078;
w3080 <= not w3073 and not w3079;
w3081 <= not b(9) and not w3080;
w3082 <= not w2824 and not w2982;
w3083 <= not w2834 and w2919;
w3084 <= not w2915 and w3083;
w3085 <= not w2916 and not w2919;
w3086 <= not w3084 and not w3085;
w3087 <= w63 and not w3086;
w3088 <= not w2981 and w3087;
w3089 <= not w3082 and not w3088;
w3090 <= not b(8) and not w3089;
w3091 <= not w2833 and not w2982;
w3092 <= not w2843 and w2914;
w3093 <= not w2910 and w3092;
w3094 <= not w2911 and not w2914;
w3095 <= not w3093 and not w3094;
w3096 <= w63 and not w3095;
w3097 <= not w2981 and w3096;
w3098 <= not w3091 and not w3097;
w3099 <= not b(7) and not w3098;
w3100 <= not w2842 and not w2982;
w3101 <= not w2852 and w2909;
w3102 <= not w2905 and w3101;
w3103 <= not w2906 and not w2909;
w3104 <= not w3102 and not w3103;
w3105 <= w63 and not w3104;
w3106 <= not w2981 and w3105;
w3107 <= not w3100 and not w3106;
w3108 <= not b(6) and not w3107;
w3109 <= not w2851 and not w2982;
w3110 <= not w2861 and w2904;
w3111 <= not w2900 and w3110;
w3112 <= not w2901 and not w2904;
w3113 <= not w3111 and not w3112;
w3114 <= w63 and not w3113;
w3115 <= not w2981 and w3114;
w3116 <= not w3109 and not w3115;
w3117 <= not b(5) and not w3116;
w3118 <= not w2860 and not w2982;
w3119 <= not w2869 and w2899;
w3120 <= not w2895 and w3119;
w3121 <= not w2896 and not w2899;
w3122 <= not w3120 and not w3121;
w3123 <= w63 and not w3122;
w3124 <= not w2981 and w3123;
w3125 <= not w3118 and not w3124;
w3126 <= not b(4) and not w3125;
w3127 <= not w2868 and not w2982;
w3128 <= not w2890 and w2894;
w3129 <= not w2889 and w3128;
w3130 <= not w2891 and not w2894;
w3131 <= not w3129 and not w3130;
w3132 <= w63 and not w3131;
w3133 <= not w2981 and w3132;
w3134 <= not w3127 and not w3133;
w3135 <= not b(3) and not w3134;
w3136 <= not w2883 and not w2982;
w3137 <= not w2886 and w2888;
w3138 <= not w2884 and w3137;
w3139 <= w63 and not w3138;
w3140 <= not w2889 and w3139;
w3141 <= not w2981 and w3140;
w3142 <= not w3136 and not w3141;
w3143 <= not b(2) and not w3142;
w3144 <= b(0) and not b(20);
w3145 <= w109 and w3144;
w3146 <= w120 and w3145;
w3147 <= w166 and w3146;
w3148 <= w151 and w3147;
w3149 <= not w2981 and w3148;
w3150 <= a(44) and not w3149;
w3151 <= w52 and w2888;
w3152 <= w86 and w3151;
w3153 <= w84 and w3152;
w3154 <= w81 and w3153;
w3155 <= not w2981 and w3154;
w3156 <= not w3150 and not w3155;
w3157 <= b(1) and not w3156;
w3158 <= not b(1) and not w3155;
w3159 <= not w3150 and w3158;
w3160 <= not w3157 and not w3159;
w3161 <= not a(43) and b(0);
w3162 <= not w3160 and not w3161;
w3163 <= not b(1) and not w3156;
w3164 <= not w3162 and not w3163;
w3165 <= b(2) and not w3141;
w3166 <= not w3136 and w3165;
w3167 <= not w3143 and not w3166;
w3168 <= not w3164 and w3167;
w3169 <= not w3143 and not w3168;
w3170 <= b(3) and not w3133;
w3171 <= not w3127 and w3170;
w3172 <= not w3135 and not w3171;
w3173 <= not w3169 and w3172;
w3174 <= not w3135 and not w3173;
w3175 <= b(4) and not w3124;
w3176 <= not w3118 and w3175;
w3177 <= not w3126 and not w3176;
w3178 <= not w3174 and w3177;
w3179 <= not w3126 and not w3178;
w3180 <= b(5) and not w3115;
w3181 <= not w3109 and w3180;
w3182 <= not w3117 and not w3181;
w3183 <= not w3179 and w3182;
w3184 <= not w3117 and not w3183;
w3185 <= b(6) and not w3106;
w3186 <= not w3100 and w3185;
w3187 <= not w3108 and not w3186;
w3188 <= not w3184 and w3187;
w3189 <= not w3108 and not w3188;
w3190 <= b(7) and not w3097;
w3191 <= not w3091 and w3190;
w3192 <= not w3099 and not w3191;
w3193 <= not w3189 and w3192;
w3194 <= not w3099 and not w3193;
w3195 <= b(8) and not w3088;
w3196 <= not w3082 and w3195;
w3197 <= not w3090 and not w3196;
w3198 <= not w3194 and w3197;
w3199 <= not w3090 and not w3198;
w3200 <= b(9) and not w3079;
w3201 <= not w3073 and w3200;
w3202 <= not w3081 and not w3201;
w3203 <= not w3199 and w3202;
w3204 <= not w3081 and not w3203;
w3205 <= b(10) and not w3070;
w3206 <= not w3064 and w3205;
w3207 <= not w3072 and not w3206;
w3208 <= not w3204 and w3207;
w3209 <= not w3072 and not w3208;
w3210 <= b(11) and not w3061;
w3211 <= not w3055 and w3210;
w3212 <= not w3063 and not w3211;
w3213 <= not w3209 and w3212;
w3214 <= not w3063 and not w3213;
w3215 <= b(12) and not w3052;
w3216 <= not w3046 and w3215;
w3217 <= not w3054 and not w3216;
w3218 <= not w3214 and w3217;
w3219 <= not w3054 and not w3218;
w3220 <= b(13) and not w3043;
w3221 <= not w3037 and w3220;
w3222 <= not w3045 and not w3221;
w3223 <= not w3219 and w3222;
w3224 <= not w3045 and not w3223;
w3225 <= b(14) and not w3034;
w3226 <= not w3028 and w3225;
w3227 <= not w3036 and not w3226;
w3228 <= not w3224 and w3227;
w3229 <= not w3036 and not w3228;
w3230 <= b(15) and not w3025;
w3231 <= not w3019 and w3230;
w3232 <= not w3027 and not w3231;
w3233 <= not w3229 and w3232;
w3234 <= not w3027 and not w3233;
w3235 <= b(16) and not w3016;
w3236 <= not w3010 and w3235;
w3237 <= not w3018 and not w3236;
w3238 <= not w3234 and w3237;
w3239 <= not w3018 and not w3238;
w3240 <= b(17) and not w3007;
w3241 <= not w3001 and w3240;
w3242 <= not w3009 and not w3241;
w3243 <= not w3239 and w3242;
w3244 <= not w3009 and not w3243;
w3245 <= b(18) and not w2998;
w3246 <= not w2992 and w3245;
w3247 <= not w3000 and not w3246;
w3248 <= not w3244 and w3247;
w3249 <= not w3000 and not w3248;
w3250 <= b(19) and not w2989;
w3251 <= not w2983 and w3250;
w3252 <= not w2991 and not w3251;
w3253 <= not w3249 and w3252;
w3254 <= not w2991 and not w3253;
w3255 <= not w2724 and not w2982;
w3256 <= not w2726 and w2979;
w3257 <= not w2975 and w3256;
w3258 <= not w2976 and not w2979;
w3259 <= not w3257 and not w3258;
w3260 <= w2982 and not w3259;
w3261 <= not w3255 and not w3260;
w3262 <= not b(20) and not w3261;
w3263 <= b(20) and not w3255;
w3264 <= not w3260 and w3263;
w3265 <= w386 and not w3264;
w3266 <= not w3262 and w3265;
w3267 <= not w3254 and w3266;
w3268 <= w63 and not w3261;
w3269 <= not w3267 and not w3268;
w3270 <= not w3000 and w3252;
w3271 <= not w3248 and w3270;
w3272 <= not w3249 and not w3252;
w3273 <= not w3271 and not w3272;
w3274 <= not w3269 and not w3273;
w3275 <= not w2990 and not w3268;
w3276 <= not w3267 and w3275;
w3277 <= not w3274 and not w3276;
w3278 <= not w2991 and not w3264;
w3279 <= not w3262 and w3278;
w3280 <= not w3253 and w3279;
w3281 <= not w3262 and not w3264;
w3282 <= not w3254 and not w3281;
w3283 <= not w3280 and not w3282;
w3284 <= not w3269 and not w3283;
w3285 <= not w3261 and not w3268;
w3286 <= not w3267 and w3285;
w3287 <= not w3284 and not w3286;
w3288 <= not b(21) and not w3287;
w3289 <= not b(20) and not w3277;
w3290 <= not w3009 and w3247;
w3291 <= not w3243 and w3290;
w3292 <= not w3244 and not w3247;
w3293 <= not w3291 and not w3292;
w3294 <= not w3269 and not w3293;
w3295 <= not w2999 and not w3268;
w3296 <= not w3267 and w3295;
w3297 <= not w3294 and not w3296;
w3298 <= not b(19) and not w3297;
w3299 <= not w3018 and w3242;
w3300 <= not w3238 and w3299;
w3301 <= not w3239 and not w3242;
w3302 <= not w3300 and not w3301;
w3303 <= not w3269 and not w3302;
w3304 <= not w3008 and not w3268;
w3305 <= not w3267 and w3304;
w3306 <= not w3303 and not w3305;
w3307 <= not b(18) and not w3306;
w3308 <= not w3027 and w3237;
w3309 <= not w3233 and w3308;
w3310 <= not w3234 and not w3237;
w3311 <= not w3309 and not w3310;
w3312 <= not w3269 and not w3311;
w3313 <= not w3017 and not w3268;
w3314 <= not w3267 and w3313;
w3315 <= not w3312 and not w3314;
w3316 <= not b(17) and not w3315;
w3317 <= not w3036 and w3232;
w3318 <= not w3228 and w3317;
w3319 <= not w3229 and not w3232;
w3320 <= not w3318 and not w3319;
w3321 <= not w3269 and not w3320;
w3322 <= not w3026 and not w3268;
w3323 <= not w3267 and w3322;
w3324 <= not w3321 and not w3323;
w3325 <= not b(16) and not w3324;
w3326 <= not w3045 and w3227;
w3327 <= not w3223 and w3326;
w3328 <= not w3224 and not w3227;
w3329 <= not w3327 and not w3328;
w3330 <= not w3269 and not w3329;
w3331 <= not w3035 and not w3268;
w3332 <= not w3267 and w3331;
w3333 <= not w3330 and not w3332;
w3334 <= not b(15) and not w3333;
w3335 <= not w3054 and w3222;
w3336 <= not w3218 and w3335;
w3337 <= not w3219 and not w3222;
w3338 <= not w3336 and not w3337;
w3339 <= not w3269 and not w3338;
w3340 <= not w3044 and not w3268;
w3341 <= not w3267 and w3340;
w3342 <= not w3339 and not w3341;
w3343 <= not b(14) and not w3342;
w3344 <= not w3063 and w3217;
w3345 <= not w3213 and w3344;
w3346 <= not w3214 and not w3217;
w3347 <= not w3345 and not w3346;
w3348 <= not w3269 and not w3347;
w3349 <= not w3053 and not w3268;
w3350 <= not w3267 and w3349;
w3351 <= not w3348 and not w3350;
w3352 <= not b(13) and not w3351;
w3353 <= not w3072 and w3212;
w3354 <= not w3208 and w3353;
w3355 <= not w3209 and not w3212;
w3356 <= not w3354 and not w3355;
w3357 <= not w3269 and not w3356;
w3358 <= not w3062 and not w3268;
w3359 <= not w3267 and w3358;
w3360 <= not w3357 and not w3359;
w3361 <= not b(12) and not w3360;
w3362 <= not w3081 and w3207;
w3363 <= not w3203 and w3362;
w3364 <= not w3204 and not w3207;
w3365 <= not w3363 and not w3364;
w3366 <= not w3269 and not w3365;
w3367 <= not w3071 and not w3268;
w3368 <= not w3267 and w3367;
w3369 <= not w3366 and not w3368;
w3370 <= not b(11) and not w3369;
w3371 <= not w3090 and w3202;
w3372 <= not w3198 and w3371;
w3373 <= not w3199 and not w3202;
w3374 <= not w3372 and not w3373;
w3375 <= not w3269 and not w3374;
w3376 <= not w3080 and not w3268;
w3377 <= not w3267 and w3376;
w3378 <= not w3375 and not w3377;
w3379 <= not b(10) and not w3378;
w3380 <= not w3099 and w3197;
w3381 <= not w3193 and w3380;
w3382 <= not w3194 and not w3197;
w3383 <= not w3381 and not w3382;
w3384 <= not w3269 and not w3383;
w3385 <= not w3089 and not w3268;
w3386 <= not w3267 and w3385;
w3387 <= not w3384 and not w3386;
w3388 <= not b(9) and not w3387;
w3389 <= not w3108 and w3192;
w3390 <= not w3188 and w3389;
w3391 <= not w3189 and not w3192;
w3392 <= not w3390 and not w3391;
w3393 <= not w3269 and not w3392;
w3394 <= not w3098 and not w3268;
w3395 <= not w3267 and w3394;
w3396 <= not w3393 and not w3395;
w3397 <= not b(8) and not w3396;
w3398 <= not w3117 and w3187;
w3399 <= not w3183 and w3398;
w3400 <= not w3184 and not w3187;
w3401 <= not w3399 and not w3400;
w3402 <= not w3269 and not w3401;
w3403 <= not w3107 and not w3268;
w3404 <= not w3267 and w3403;
w3405 <= not w3402 and not w3404;
w3406 <= not b(7) and not w3405;
w3407 <= not w3126 and w3182;
w3408 <= not w3178 and w3407;
w3409 <= not w3179 and not w3182;
w3410 <= not w3408 and not w3409;
w3411 <= not w3269 and not w3410;
w3412 <= not w3116 and not w3268;
w3413 <= not w3267 and w3412;
w3414 <= not w3411 and not w3413;
w3415 <= not b(6) and not w3414;
w3416 <= not w3135 and w3177;
w3417 <= not w3173 and w3416;
w3418 <= not w3174 and not w3177;
w3419 <= not w3417 and not w3418;
w3420 <= not w3269 and not w3419;
w3421 <= not w3125 and not w3268;
w3422 <= not w3267 and w3421;
w3423 <= not w3420 and not w3422;
w3424 <= not b(5) and not w3423;
w3425 <= not w3143 and w3172;
w3426 <= not w3168 and w3425;
w3427 <= not w3169 and not w3172;
w3428 <= not w3426 and not w3427;
w3429 <= not w3269 and not w3428;
w3430 <= not w3134 and not w3268;
w3431 <= not w3267 and w3430;
w3432 <= not w3429 and not w3431;
w3433 <= not b(4) and not w3432;
w3434 <= not w3163 and w3167;
w3435 <= not w3162 and w3434;
w3436 <= not w3164 and not w3167;
w3437 <= not w3435 and not w3436;
w3438 <= not w3269 and not w3437;
w3439 <= not w3142 and not w3268;
w3440 <= not w3267 and w3439;
w3441 <= not w3438 and not w3440;
w3442 <= not b(3) and not w3441;
w3443 <= not w3159 and w3161;
w3444 <= not w3157 and w3443;
w3445 <= not w3162 and not w3444;
w3446 <= not w3269 and w3445;
w3447 <= not w3156 and not w3268;
w3448 <= not w3267 and w3447;
w3449 <= not w3446 and not w3448;
w3450 <= not b(2) and not w3449;
w3451 <= b(0) and not w3269;
w3452 <= a(43) and not w3451;
w3453 <= w3161 and not w3269;
w3454 <= not w3452 and not w3453;
w3455 <= b(1) and not w3454;
w3456 <= not b(1) and not w3453;
w3457 <= not w3452 and w3456;
w3458 <= not w3455 and not w3457;
w3459 <= not a(42) and b(0);
w3460 <= not w3458 and not w3459;
w3461 <= not b(1) and not w3454;
w3462 <= not w3460 and not w3461;
w3463 <= b(2) and not w3448;
w3464 <= not w3446 and w3463;
w3465 <= not w3450 and not w3464;
w3466 <= not w3462 and w3465;
w3467 <= not w3450 and not w3466;
w3468 <= b(3) and not w3440;
w3469 <= not w3438 and w3468;
w3470 <= not w3442 and not w3469;
w3471 <= not w3467 and w3470;
w3472 <= not w3442 and not w3471;
w3473 <= b(4) and not w3431;
w3474 <= not w3429 and w3473;
w3475 <= not w3433 and not w3474;
w3476 <= not w3472 and w3475;
w3477 <= not w3433 and not w3476;
w3478 <= b(5) and not w3422;
w3479 <= not w3420 and w3478;
w3480 <= not w3424 and not w3479;
w3481 <= not w3477 and w3480;
w3482 <= not w3424 and not w3481;
w3483 <= b(6) and not w3413;
w3484 <= not w3411 and w3483;
w3485 <= not w3415 and not w3484;
w3486 <= not w3482 and w3485;
w3487 <= not w3415 and not w3486;
w3488 <= b(7) and not w3404;
w3489 <= not w3402 and w3488;
w3490 <= not w3406 and not w3489;
w3491 <= not w3487 and w3490;
w3492 <= not w3406 and not w3491;
w3493 <= b(8) and not w3395;
w3494 <= not w3393 and w3493;
w3495 <= not w3397 and not w3494;
w3496 <= not w3492 and w3495;
w3497 <= not w3397 and not w3496;
w3498 <= b(9) and not w3386;
w3499 <= not w3384 and w3498;
w3500 <= not w3388 and not w3499;
w3501 <= not w3497 and w3500;
w3502 <= not w3388 and not w3501;
w3503 <= b(10) and not w3377;
w3504 <= not w3375 and w3503;
w3505 <= not w3379 and not w3504;
w3506 <= not w3502 and w3505;
w3507 <= not w3379 and not w3506;
w3508 <= b(11) and not w3368;
w3509 <= not w3366 and w3508;
w3510 <= not w3370 and not w3509;
w3511 <= not w3507 and w3510;
w3512 <= not w3370 and not w3511;
w3513 <= b(12) and not w3359;
w3514 <= not w3357 and w3513;
w3515 <= not w3361 and not w3514;
w3516 <= not w3512 and w3515;
w3517 <= not w3361 and not w3516;
w3518 <= b(13) and not w3350;
w3519 <= not w3348 and w3518;
w3520 <= not w3352 and not w3519;
w3521 <= not w3517 and w3520;
w3522 <= not w3352 and not w3521;
w3523 <= b(14) and not w3341;
w3524 <= not w3339 and w3523;
w3525 <= not w3343 and not w3524;
w3526 <= not w3522 and w3525;
w3527 <= not w3343 and not w3526;
w3528 <= b(15) and not w3332;
w3529 <= not w3330 and w3528;
w3530 <= not w3334 and not w3529;
w3531 <= not w3527 and w3530;
w3532 <= not w3334 and not w3531;
w3533 <= b(16) and not w3323;
w3534 <= not w3321 and w3533;
w3535 <= not w3325 and not w3534;
w3536 <= not w3532 and w3535;
w3537 <= not w3325 and not w3536;
w3538 <= b(17) and not w3314;
w3539 <= not w3312 and w3538;
w3540 <= not w3316 and not w3539;
w3541 <= not w3537 and w3540;
w3542 <= not w3316 and not w3541;
w3543 <= b(18) and not w3305;
w3544 <= not w3303 and w3543;
w3545 <= not w3307 and not w3544;
w3546 <= not w3542 and w3545;
w3547 <= not w3307 and not w3546;
w3548 <= b(19) and not w3296;
w3549 <= not w3294 and w3548;
w3550 <= not w3298 and not w3549;
w3551 <= not w3547 and w3550;
w3552 <= not w3298 and not w3551;
w3553 <= b(20) and not w3276;
w3554 <= not w3274 and w3553;
w3555 <= not w3289 and not w3554;
w3556 <= not w3552 and w3555;
w3557 <= not w3289 and not w3556;
w3558 <= b(21) and not w3286;
w3559 <= not w3284 and w3558;
w3560 <= not w3288 and not w3559;
w3561 <= not w3557 and w3560;
w3562 <= not w3288 and not w3561;
w3563 <= w49 and w51;
w3564 <= w60 and w3563;
w3565 <= w46 and w3564;
w3566 <= w31 and w3565;
w3567 <= not w3562 and w3566;
w3568 <= not w3277 and not w3567;
w3569 <= not w3298 and w3555;
w3570 <= not w3551 and w3569;
w3571 <= not w3552 and not w3555;
w3572 <= not w3570 and not w3571;
w3573 <= w3566 and not w3572;
w3574 <= not w3562 and w3573;
w3575 <= not w3568 and not w3574;
w3576 <= not w3287 and not w3567;
w3577 <= not w3289 and w3560;
w3578 <= not w3556 and w3577;
w3579 <= not w3557 and not w3560;
w3580 <= not w3578 and not w3579;
w3581 <= w3567 and not w3580;
w3582 <= not w3576 and not w3581;
w3583 <= not b(22) and not w3582;
w3584 <= not b(21) and not w3575;
w3585 <= not w3297 and not w3567;
w3586 <= not w3307 and w3550;
w3587 <= not w3546 and w3586;
w3588 <= not w3547 and not w3550;
w3589 <= not w3587 and not w3588;
w3590 <= w3566 and not w3589;
w3591 <= not w3562 and w3590;
w3592 <= not w3585 and not w3591;
w3593 <= not b(20) and not w3592;
w3594 <= not w3306 and not w3567;
w3595 <= not w3316 and w3545;
w3596 <= not w3541 and w3595;
w3597 <= not w3542 and not w3545;
w3598 <= not w3596 and not w3597;
w3599 <= w3566 and not w3598;
w3600 <= not w3562 and w3599;
w3601 <= not w3594 and not w3600;
w3602 <= not b(19) and not w3601;
w3603 <= not w3315 and not w3567;
w3604 <= not w3325 and w3540;
w3605 <= not w3536 and w3604;
w3606 <= not w3537 and not w3540;
w3607 <= not w3605 and not w3606;
w3608 <= w3566 and not w3607;
w3609 <= not w3562 and w3608;
w3610 <= not w3603 and not w3609;
w3611 <= not b(18) and not w3610;
w3612 <= not w3324 and not w3567;
w3613 <= not w3334 and w3535;
w3614 <= not w3531 and w3613;
w3615 <= not w3532 and not w3535;
w3616 <= not w3614 and not w3615;
w3617 <= w3566 and not w3616;
w3618 <= not w3562 and w3617;
w3619 <= not w3612 and not w3618;
w3620 <= not b(17) and not w3619;
w3621 <= not w3333 and not w3567;
w3622 <= not w3343 and w3530;
w3623 <= not w3526 and w3622;
w3624 <= not w3527 and not w3530;
w3625 <= not w3623 and not w3624;
w3626 <= w3566 and not w3625;
w3627 <= not w3562 and w3626;
w3628 <= not w3621 and not w3627;
w3629 <= not b(16) and not w3628;
w3630 <= not w3342 and not w3567;
w3631 <= not w3352 and w3525;
w3632 <= not w3521 and w3631;
w3633 <= not w3522 and not w3525;
w3634 <= not w3632 and not w3633;
w3635 <= w3566 and not w3634;
w3636 <= not w3562 and w3635;
w3637 <= not w3630 and not w3636;
w3638 <= not b(15) and not w3637;
w3639 <= not w3351 and not w3567;
w3640 <= not w3361 and w3520;
w3641 <= not w3516 and w3640;
w3642 <= not w3517 and not w3520;
w3643 <= not w3641 and not w3642;
w3644 <= w3566 and not w3643;
w3645 <= not w3562 and w3644;
w3646 <= not w3639 and not w3645;
w3647 <= not b(14) and not w3646;
w3648 <= not w3360 and not w3567;
w3649 <= not w3370 and w3515;
w3650 <= not w3511 and w3649;
w3651 <= not w3512 and not w3515;
w3652 <= not w3650 and not w3651;
w3653 <= w3566 and not w3652;
w3654 <= not w3562 and w3653;
w3655 <= not w3648 and not w3654;
w3656 <= not b(13) and not w3655;
w3657 <= not w3369 and not w3567;
w3658 <= not w3379 and w3510;
w3659 <= not w3506 and w3658;
w3660 <= not w3507 and not w3510;
w3661 <= not w3659 and not w3660;
w3662 <= w3566 and not w3661;
w3663 <= not w3562 and w3662;
w3664 <= not w3657 and not w3663;
w3665 <= not b(12) and not w3664;
w3666 <= not w3378 and not w3567;
w3667 <= not w3388 and w3505;
w3668 <= not w3501 and w3667;
w3669 <= not w3502 and not w3505;
w3670 <= not w3668 and not w3669;
w3671 <= w3566 and not w3670;
w3672 <= not w3562 and w3671;
w3673 <= not w3666 and not w3672;
w3674 <= not b(11) and not w3673;
w3675 <= not w3387 and not w3567;
w3676 <= not w3397 and w3500;
w3677 <= not w3496 and w3676;
w3678 <= not w3497 and not w3500;
w3679 <= not w3677 and not w3678;
w3680 <= w3566 and not w3679;
w3681 <= not w3562 and w3680;
w3682 <= not w3675 and not w3681;
w3683 <= not b(10) and not w3682;
w3684 <= not w3396 and not w3567;
w3685 <= not w3406 and w3495;
w3686 <= not w3491 and w3685;
w3687 <= not w3492 and not w3495;
w3688 <= not w3686 and not w3687;
w3689 <= w3566 and not w3688;
w3690 <= not w3562 and w3689;
w3691 <= not w3684 and not w3690;
w3692 <= not b(9) and not w3691;
w3693 <= not w3405 and not w3567;
w3694 <= not w3415 and w3490;
w3695 <= not w3486 and w3694;
w3696 <= not w3487 and not w3490;
w3697 <= not w3695 and not w3696;
w3698 <= w3566 and not w3697;
w3699 <= not w3562 and w3698;
w3700 <= not w3693 and not w3699;
w3701 <= not b(8) and not w3700;
w3702 <= not w3414 and not w3567;
w3703 <= not w3424 and w3485;
w3704 <= not w3481 and w3703;
w3705 <= not w3482 and not w3485;
w3706 <= not w3704 and not w3705;
w3707 <= w3566 and not w3706;
w3708 <= not w3562 and w3707;
w3709 <= not w3702 and not w3708;
w3710 <= not b(7) and not w3709;
w3711 <= not w3423 and not w3567;
w3712 <= not w3433 and w3480;
w3713 <= not w3476 and w3712;
w3714 <= not w3477 and not w3480;
w3715 <= not w3713 and not w3714;
w3716 <= w3566 and not w3715;
w3717 <= not w3562 and w3716;
w3718 <= not w3711 and not w3717;
w3719 <= not b(6) and not w3718;
w3720 <= not w3432 and not w3567;
w3721 <= not w3442 and w3475;
w3722 <= not w3471 and w3721;
w3723 <= not w3472 and not w3475;
w3724 <= not w3722 and not w3723;
w3725 <= w3566 and not w3724;
w3726 <= not w3562 and w3725;
w3727 <= not w3720 and not w3726;
w3728 <= not b(5) and not w3727;
w3729 <= not w3441 and not w3567;
w3730 <= not w3450 and w3470;
w3731 <= not w3466 and w3730;
w3732 <= not w3467 and not w3470;
w3733 <= not w3731 and not w3732;
w3734 <= w3566 and not w3733;
w3735 <= not w3562 and w3734;
w3736 <= not w3729 and not w3735;
w3737 <= not b(4) and not w3736;
w3738 <= not w3449 and not w3567;
w3739 <= not w3461 and w3465;
w3740 <= not w3460 and w3739;
w3741 <= not w3462 and not w3465;
w3742 <= not w3740 and not w3741;
w3743 <= w3566 and not w3742;
w3744 <= not w3562 and w3743;
w3745 <= not w3738 and not w3744;
w3746 <= not b(3) and not w3745;
w3747 <= not w3454 and not w3567;
w3748 <= not w3457 and w3459;
w3749 <= not w3455 and w3748;
w3750 <= w3566 and not w3749;
w3751 <= not w3460 and w3750;
w3752 <= not w3562 and w3751;
w3753 <= not w3747 and not w3752;
w3754 <= not b(2) and not w3753;
w3755 <= b(0) and not b(22);
w3756 <= w108 and w3755;
w3757 <= w119 and w3756;
w3758 <= w331 and w3757;
w3759 <= w341 and w3758;
w3760 <= w338 and w3759;
w3761 <= not w3562 and w3760;
w3762 <= a(42) and not w3761;
w3763 <= w51 and w3459;
w3764 <= w49 and w3763;
w3765 <= w60 and w3764;
w3766 <= w46 and w3765;
w3767 <= w31 and w3766;
w3768 <= not w3562 and w3767;
w3769 <= not w3762 and not w3768;
w3770 <= b(1) and not w3769;
w3771 <= not b(1) and not w3768;
w3772 <= not w3762 and w3771;
w3773 <= not w3770 and not w3772;
w3774 <= not a(41) and b(0);
w3775 <= not w3773 and not w3774;
w3776 <= not b(1) and not w3769;
w3777 <= not w3775 and not w3776;
w3778 <= b(2) and not w3752;
w3779 <= not w3747 and w3778;
w3780 <= not w3754 and not w3779;
w3781 <= not w3777 and w3780;
w3782 <= not w3754 and not w3781;
w3783 <= b(3) and not w3744;
w3784 <= not w3738 and w3783;
w3785 <= not w3746 and not w3784;
w3786 <= not w3782 and w3785;
w3787 <= not w3746 and not w3786;
w3788 <= b(4) and not w3735;
w3789 <= not w3729 and w3788;
w3790 <= not w3737 and not w3789;
w3791 <= not w3787 and w3790;
w3792 <= not w3737 and not w3791;
w3793 <= b(5) and not w3726;
w3794 <= not w3720 and w3793;
w3795 <= not w3728 and not w3794;
w3796 <= not w3792 and w3795;
w3797 <= not w3728 and not w3796;
w3798 <= b(6) and not w3717;
w3799 <= not w3711 and w3798;
w3800 <= not w3719 and not w3799;
w3801 <= not w3797 and w3800;
w3802 <= not w3719 and not w3801;
w3803 <= b(7) and not w3708;
w3804 <= not w3702 and w3803;
w3805 <= not w3710 and not w3804;
w3806 <= not w3802 and w3805;
w3807 <= not w3710 and not w3806;
w3808 <= b(8) and not w3699;
w3809 <= not w3693 and w3808;
w3810 <= not w3701 and not w3809;
w3811 <= not w3807 and w3810;
w3812 <= not w3701 and not w3811;
w3813 <= b(9) and not w3690;
w3814 <= not w3684 and w3813;
w3815 <= not w3692 and not w3814;
w3816 <= not w3812 and w3815;
w3817 <= not w3692 and not w3816;
w3818 <= b(10) and not w3681;
w3819 <= not w3675 and w3818;
w3820 <= not w3683 and not w3819;
w3821 <= not w3817 and w3820;
w3822 <= not w3683 and not w3821;
w3823 <= b(11) and not w3672;
w3824 <= not w3666 and w3823;
w3825 <= not w3674 and not w3824;
w3826 <= not w3822 and w3825;
w3827 <= not w3674 and not w3826;
w3828 <= b(12) and not w3663;
w3829 <= not w3657 and w3828;
w3830 <= not w3665 and not w3829;
w3831 <= not w3827 and w3830;
w3832 <= not w3665 and not w3831;
w3833 <= b(13) and not w3654;
w3834 <= not w3648 and w3833;
w3835 <= not w3656 and not w3834;
w3836 <= not w3832 and w3835;
w3837 <= not w3656 and not w3836;
w3838 <= b(14) and not w3645;
w3839 <= not w3639 and w3838;
w3840 <= not w3647 and not w3839;
w3841 <= not w3837 and w3840;
w3842 <= not w3647 and not w3841;
w3843 <= b(15) and not w3636;
w3844 <= not w3630 and w3843;
w3845 <= not w3638 and not w3844;
w3846 <= not w3842 and w3845;
w3847 <= not w3638 and not w3846;
w3848 <= b(16) and not w3627;
w3849 <= not w3621 and w3848;
w3850 <= not w3629 and not w3849;
w3851 <= not w3847 and w3850;
w3852 <= not w3629 and not w3851;
w3853 <= b(17) and not w3618;
w3854 <= not w3612 and w3853;
w3855 <= not w3620 and not w3854;
w3856 <= not w3852 and w3855;
w3857 <= not w3620 and not w3856;
w3858 <= b(18) and not w3609;
w3859 <= not w3603 and w3858;
w3860 <= not w3611 and not w3859;
w3861 <= not w3857 and w3860;
w3862 <= not w3611 and not w3861;
w3863 <= b(19) and not w3600;
w3864 <= not w3594 and w3863;
w3865 <= not w3602 and not w3864;
w3866 <= not w3862 and w3865;
w3867 <= not w3602 and not w3866;
w3868 <= b(20) and not w3591;
w3869 <= not w3585 and w3868;
w3870 <= not w3593 and not w3869;
w3871 <= not w3867 and w3870;
w3872 <= not w3593 and not w3871;
w3873 <= b(21) and not w3574;
w3874 <= not w3568 and w3873;
w3875 <= not w3584 and not w3874;
w3876 <= not w3872 and w3875;
w3877 <= not w3584 and not w3876;
w3878 <= b(22) and not w3576;
w3879 <= not w3581 and w3878;
w3880 <= not w3583 and not w3879;
w3881 <= not w3877 and w3880;
w3882 <= not w3583 and not w3881;
w3883 <= w108 and w119;
w3884 <= w331 and w3883;
w3885 <= w341 and w3884;
w3886 <= w338 and w3885;
w3887 <= not w3882 and w3886;
w3888 <= not w3575 and not w3887;
w3889 <= not w3593 and w3875;
w3890 <= not w3871 and w3889;
w3891 <= not w3872 and not w3875;
w3892 <= not w3890 and not w3891;
w3893 <= w3886 and not w3892;
w3894 <= not w3882 and w3893;
w3895 <= not w3888 and not w3894;
w3896 <= not b(22) and not w3895;
w3897 <= not w3592 and not w3887;
w3898 <= not w3602 and w3870;
w3899 <= not w3866 and w3898;
w3900 <= not w3867 and not w3870;
w3901 <= not w3899 and not w3900;
w3902 <= w3886 and not w3901;
w3903 <= not w3882 and w3902;
w3904 <= not w3897 and not w3903;
w3905 <= not b(21) and not w3904;
w3906 <= not w3601 and not w3887;
w3907 <= not w3611 and w3865;
w3908 <= not w3861 and w3907;
w3909 <= not w3862 and not w3865;
w3910 <= not w3908 and not w3909;
w3911 <= w3886 and not w3910;
w3912 <= not w3882 and w3911;
w3913 <= not w3906 and not w3912;
w3914 <= not b(20) and not w3913;
w3915 <= not w3610 and not w3887;
w3916 <= not w3620 and w3860;
w3917 <= not w3856 and w3916;
w3918 <= not w3857 and not w3860;
w3919 <= not w3917 and not w3918;
w3920 <= w3886 and not w3919;
w3921 <= not w3882 and w3920;
w3922 <= not w3915 and not w3921;
w3923 <= not b(19) and not w3922;
w3924 <= not w3619 and not w3887;
w3925 <= not w3629 and w3855;
w3926 <= not w3851 and w3925;
w3927 <= not w3852 and not w3855;
w3928 <= not w3926 and not w3927;
w3929 <= w3886 and not w3928;
w3930 <= not w3882 and w3929;
w3931 <= not w3924 and not w3930;
w3932 <= not b(18) and not w3931;
w3933 <= not w3628 and not w3887;
w3934 <= not w3638 and w3850;
w3935 <= not w3846 and w3934;
w3936 <= not w3847 and not w3850;
w3937 <= not w3935 and not w3936;
w3938 <= w3886 and not w3937;
w3939 <= not w3882 and w3938;
w3940 <= not w3933 and not w3939;
w3941 <= not b(17) and not w3940;
w3942 <= not w3637 and not w3887;
w3943 <= not w3647 and w3845;
w3944 <= not w3841 and w3943;
w3945 <= not w3842 and not w3845;
w3946 <= not w3944 and not w3945;
w3947 <= w3886 and not w3946;
w3948 <= not w3882 and w3947;
w3949 <= not w3942 and not w3948;
w3950 <= not b(16) and not w3949;
w3951 <= not w3646 and not w3887;
w3952 <= not w3656 and w3840;
w3953 <= not w3836 and w3952;
w3954 <= not w3837 and not w3840;
w3955 <= not w3953 and not w3954;
w3956 <= w3886 and not w3955;
w3957 <= not w3882 and w3956;
w3958 <= not w3951 and not w3957;
w3959 <= not b(15) and not w3958;
w3960 <= not w3655 and not w3887;
w3961 <= not w3665 and w3835;
w3962 <= not w3831 and w3961;
w3963 <= not w3832 and not w3835;
w3964 <= not w3962 and not w3963;
w3965 <= w3886 and not w3964;
w3966 <= not w3882 and w3965;
w3967 <= not w3960 and not w3966;
w3968 <= not b(14) and not w3967;
w3969 <= not w3664 and not w3887;
w3970 <= not w3674 and w3830;
w3971 <= not w3826 and w3970;
w3972 <= not w3827 and not w3830;
w3973 <= not w3971 and not w3972;
w3974 <= w3886 and not w3973;
w3975 <= not w3882 and w3974;
w3976 <= not w3969 and not w3975;
w3977 <= not b(13) and not w3976;
w3978 <= not w3673 and not w3887;
w3979 <= not w3683 and w3825;
w3980 <= not w3821 and w3979;
w3981 <= not w3822 and not w3825;
w3982 <= not w3980 and not w3981;
w3983 <= w3886 and not w3982;
w3984 <= not w3882 and w3983;
w3985 <= not w3978 and not w3984;
w3986 <= not b(12) and not w3985;
w3987 <= not w3682 and not w3887;
w3988 <= not w3692 and w3820;
w3989 <= not w3816 and w3988;
w3990 <= not w3817 and not w3820;
w3991 <= not w3989 and not w3990;
w3992 <= w3886 and not w3991;
w3993 <= not w3882 and w3992;
w3994 <= not w3987 and not w3993;
w3995 <= not b(11) and not w3994;
w3996 <= not w3691 and not w3887;
w3997 <= not w3701 and w3815;
w3998 <= not w3811 and w3997;
w3999 <= not w3812 and not w3815;
w4000 <= not w3998 and not w3999;
w4001 <= w3886 and not w4000;
w4002 <= not w3882 and w4001;
w4003 <= not w3996 and not w4002;
w4004 <= not b(10) and not w4003;
w4005 <= not w3700 and not w3887;
w4006 <= not w3710 and w3810;
w4007 <= not w3806 and w4006;
w4008 <= not w3807 and not w3810;
w4009 <= not w4007 and not w4008;
w4010 <= w3886 and not w4009;
w4011 <= not w3882 and w4010;
w4012 <= not w4005 and not w4011;
w4013 <= not b(9) and not w4012;
w4014 <= not w3709 and not w3887;
w4015 <= not w3719 and w3805;
w4016 <= not w3801 and w4015;
w4017 <= not w3802 and not w3805;
w4018 <= not w4016 and not w4017;
w4019 <= w3886 and not w4018;
w4020 <= not w3882 and w4019;
w4021 <= not w4014 and not w4020;
w4022 <= not b(8) and not w4021;
w4023 <= not w3718 and not w3887;
w4024 <= not w3728 and w3800;
w4025 <= not w3796 and w4024;
w4026 <= not w3797 and not w3800;
w4027 <= not w4025 and not w4026;
w4028 <= w3886 and not w4027;
w4029 <= not w3882 and w4028;
w4030 <= not w4023 and not w4029;
w4031 <= not b(7) and not w4030;
w4032 <= not w3727 and not w3887;
w4033 <= not w3737 and w3795;
w4034 <= not w3791 and w4033;
w4035 <= not w3792 and not w3795;
w4036 <= not w4034 and not w4035;
w4037 <= w3886 and not w4036;
w4038 <= not w3882 and w4037;
w4039 <= not w4032 and not w4038;
w4040 <= not b(6) and not w4039;
w4041 <= not w3736 and not w3887;
w4042 <= not w3746 and w3790;
w4043 <= not w3786 and w4042;
w4044 <= not w3787 and not w3790;
w4045 <= not w4043 and not w4044;
w4046 <= w3886 and not w4045;
w4047 <= not w3882 and w4046;
w4048 <= not w4041 and not w4047;
w4049 <= not b(5) and not w4048;
w4050 <= not w3745 and not w3887;
w4051 <= not w3754 and w3785;
w4052 <= not w3781 and w4051;
w4053 <= not w3782 and not w3785;
w4054 <= not w4052 and not w4053;
w4055 <= w3886 and not w4054;
w4056 <= not w3882 and w4055;
w4057 <= not w4050 and not w4056;
w4058 <= not b(4) and not w4057;
w4059 <= not w3753 and not w3887;
w4060 <= not w3776 and w3780;
w4061 <= not w3775 and w4060;
w4062 <= not w3777 and not w3780;
w4063 <= not w4061 and not w4062;
w4064 <= w3886 and not w4063;
w4065 <= not w3882 and w4064;
w4066 <= not w4059 and not w4065;
w4067 <= not b(3) and not w4066;
w4068 <= not w3769 and not w3887;
w4069 <= not w3772 and w3774;
w4070 <= not w3770 and w4069;
w4071 <= w3886 and not w4070;
w4072 <= not w3775 and w4071;
w4073 <= not w3882 and w4072;
w4074 <= not w4068 and not w4073;
w4075 <= not b(2) and not w4074;
w4076 <= b(0) and not b(23);
w4077 <= w49 and w4076;
w4078 <= w60 and w4077;
w4079 <= w46 and w4078;
w4080 <= w31 and w4079;
w4081 <= not w3882 and w4080;
w4082 <= a(41) and not w4081;
w4083 <= w108 and w3774;
w4084 <= w119 and w4083;
w4085 <= w331 and w4084;
w4086 <= w341 and w4085;
w4087 <= w338 and w4086;
w4088 <= not w3882 and w4087;
w4089 <= not w4082 and not w4088;
w4090 <= b(1) and not w4089;
w4091 <= not b(1) and not w4088;
w4092 <= not w4082 and w4091;
w4093 <= not w4090 and not w4092;
w4094 <= not a(40) and b(0);
w4095 <= not w4093 and not w4094;
w4096 <= not b(1) and not w4089;
w4097 <= not w4095 and not w4096;
w4098 <= b(2) and not w4073;
w4099 <= not w4068 and w4098;
w4100 <= not w4075 and not w4099;
w4101 <= not w4097 and w4100;
w4102 <= not w4075 and not w4101;
w4103 <= b(3) and not w4065;
w4104 <= not w4059 and w4103;
w4105 <= not w4067 and not w4104;
w4106 <= not w4102 and w4105;
w4107 <= not w4067 and not w4106;
w4108 <= b(4) and not w4056;
w4109 <= not w4050 and w4108;
w4110 <= not w4058 and not w4109;
w4111 <= not w4107 and w4110;
w4112 <= not w4058 and not w4111;
w4113 <= b(5) and not w4047;
w4114 <= not w4041 and w4113;
w4115 <= not w4049 and not w4114;
w4116 <= not w4112 and w4115;
w4117 <= not w4049 and not w4116;
w4118 <= b(6) and not w4038;
w4119 <= not w4032 and w4118;
w4120 <= not w4040 and not w4119;
w4121 <= not w4117 and w4120;
w4122 <= not w4040 and not w4121;
w4123 <= b(7) and not w4029;
w4124 <= not w4023 and w4123;
w4125 <= not w4031 and not w4124;
w4126 <= not w4122 and w4125;
w4127 <= not w4031 and not w4126;
w4128 <= b(8) and not w4020;
w4129 <= not w4014 and w4128;
w4130 <= not w4022 and not w4129;
w4131 <= not w4127 and w4130;
w4132 <= not w4022 and not w4131;
w4133 <= b(9) and not w4011;
w4134 <= not w4005 and w4133;
w4135 <= not w4013 and not w4134;
w4136 <= not w4132 and w4135;
w4137 <= not w4013 and not w4136;
w4138 <= b(10) and not w4002;
w4139 <= not w3996 and w4138;
w4140 <= not w4004 and not w4139;
w4141 <= not w4137 and w4140;
w4142 <= not w4004 and not w4141;
w4143 <= b(11) and not w3993;
w4144 <= not w3987 and w4143;
w4145 <= not w3995 and not w4144;
w4146 <= not w4142 and w4145;
w4147 <= not w3995 and not w4146;
w4148 <= b(12) and not w3984;
w4149 <= not w3978 and w4148;
w4150 <= not w3986 and not w4149;
w4151 <= not w4147 and w4150;
w4152 <= not w3986 and not w4151;
w4153 <= b(13) and not w3975;
w4154 <= not w3969 and w4153;
w4155 <= not w3977 and not w4154;
w4156 <= not w4152 and w4155;
w4157 <= not w3977 and not w4156;
w4158 <= b(14) and not w3966;
w4159 <= not w3960 and w4158;
w4160 <= not w3968 and not w4159;
w4161 <= not w4157 and w4160;
w4162 <= not w3968 and not w4161;
w4163 <= b(15) and not w3957;
w4164 <= not w3951 and w4163;
w4165 <= not w3959 and not w4164;
w4166 <= not w4162 and w4165;
w4167 <= not w3959 and not w4166;
w4168 <= b(16) and not w3948;
w4169 <= not w3942 and w4168;
w4170 <= not w3950 and not w4169;
w4171 <= not w4167 and w4170;
w4172 <= not w3950 and not w4171;
w4173 <= b(17) and not w3939;
w4174 <= not w3933 and w4173;
w4175 <= not w3941 and not w4174;
w4176 <= not w4172 and w4175;
w4177 <= not w3941 and not w4176;
w4178 <= b(18) and not w3930;
w4179 <= not w3924 and w4178;
w4180 <= not w3932 and not w4179;
w4181 <= not w4177 and w4180;
w4182 <= not w3932 and not w4181;
w4183 <= b(19) and not w3921;
w4184 <= not w3915 and w4183;
w4185 <= not w3923 and not w4184;
w4186 <= not w4182 and w4185;
w4187 <= not w3923 and not w4186;
w4188 <= b(20) and not w3912;
w4189 <= not w3906 and w4188;
w4190 <= not w3914 and not w4189;
w4191 <= not w4187 and w4190;
w4192 <= not w3914 and not w4191;
w4193 <= b(21) and not w3903;
w4194 <= not w3897 and w4193;
w4195 <= not w3905 and not w4194;
w4196 <= not w4192 and w4195;
w4197 <= not w3905 and not w4196;
w4198 <= b(22) and not w3894;
w4199 <= not w3888 and w4198;
w4200 <= not w3896 and not w4199;
w4201 <= not w4197 and w4200;
w4202 <= not w3896 and not w4201;
w4203 <= not w3582 and not w3887;
w4204 <= not w3584 and w3880;
w4205 <= not w3876 and w4204;
w4206 <= not w3877 and not w3880;
w4207 <= not w4205 and not w4206;
w4208 <= w3887 and not w4207;
w4209 <= not w4203 and not w4208;
w4210 <= not b(23) and not w4209;
w4211 <= b(23) and not w4203;
w4212 <= not w4208 and w4211;
w4213 <= w84 and w86;
w4214 <= w81 and w4213;
w4215 <= not w4212 and w4214;
w4216 <= not w4210 and w4215;
w4217 <= not w4202 and w4216;
w4218 <= w3886 and not w4209;
w4219 <= not w4217 and not w4218;
w4220 <= not w3905 and w4200;
w4221 <= not w4196 and w4220;
w4222 <= not w4197 and not w4200;
w4223 <= not w4221 and not w4222;
w4224 <= not w4219 and not w4223;
w4225 <= not w3895 and not w4218;
w4226 <= not w4217 and w4225;
w4227 <= not w4224 and not w4226;
w4228 <= not w3896 and not w4212;
w4229 <= not w4210 and w4228;
w4230 <= not w4201 and w4229;
w4231 <= not w4210 and not w4212;
w4232 <= not w4202 and not w4231;
w4233 <= not w4230 and not w4232;
w4234 <= not w4219 and not w4233;
w4235 <= not w4209 and not w4218;
w4236 <= not w4217 and w4235;
w4237 <= not w4234 and not w4236;
w4238 <= not b(24) and not w4237;
w4239 <= not b(23) and not w4227;
w4240 <= not w3914 and w4195;
w4241 <= not w4191 and w4240;
w4242 <= not w4192 and not w4195;
w4243 <= not w4241 and not w4242;
w4244 <= not w4219 and not w4243;
w4245 <= not w3904 and not w4218;
w4246 <= not w4217 and w4245;
w4247 <= not w4244 and not w4246;
w4248 <= not b(22) and not w4247;
w4249 <= not w3923 and w4190;
w4250 <= not w4186 and w4249;
w4251 <= not w4187 and not w4190;
w4252 <= not w4250 and not w4251;
w4253 <= not w4219 and not w4252;
w4254 <= not w3913 and not w4218;
w4255 <= not w4217 and w4254;
w4256 <= not w4253 and not w4255;
w4257 <= not b(21) and not w4256;
w4258 <= not w3932 and w4185;
w4259 <= not w4181 and w4258;
w4260 <= not w4182 and not w4185;
w4261 <= not w4259 and not w4260;
w4262 <= not w4219 and not w4261;
w4263 <= not w3922 and not w4218;
w4264 <= not w4217 and w4263;
w4265 <= not w4262 and not w4264;
w4266 <= not b(20) and not w4265;
w4267 <= not w3941 and w4180;
w4268 <= not w4176 and w4267;
w4269 <= not w4177 and not w4180;
w4270 <= not w4268 and not w4269;
w4271 <= not w4219 and not w4270;
w4272 <= not w3931 and not w4218;
w4273 <= not w4217 and w4272;
w4274 <= not w4271 and not w4273;
w4275 <= not b(19) and not w4274;
w4276 <= not w3950 and w4175;
w4277 <= not w4171 and w4276;
w4278 <= not w4172 and not w4175;
w4279 <= not w4277 and not w4278;
w4280 <= not w4219 and not w4279;
w4281 <= not w3940 and not w4218;
w4282 <= not w4217 and w4281;
w4283 <= not w4280 and not w4282;
w4284 <= not b(18) and not w4283;
w4285 <= not w3959 and w4170;
w4286 <= not w4166 and w4285;
w4287 <= not w4167 and not w4170;
w4288 <= not w4286 and not w4287;
w4289 <= not w4219 and not w4288;
w4290 <= not w3949 and not w4218;
w4291 <= not w4217 and w4290;
w4292 <= not w4289 and not w4291;
w4293 <= not b(17) and not w4292;
w4294 <= not w3968 and w4165;
w4295 <= not w4161 and w4294;
w4296 <= not w4162 and not w4165;
w4297 <= not w4295 and not w4296;
w4298 <= not w4219 and not w4297;
w4299 <= not w3958 and not w4218;
w4300 <= not w4217 and w4299;
w4301 <= not w4298 and not w4300;
w4302 <= not b(16) and not w4301;
w4303 <= not w3977 and w4160;
w4304 <= not w4156 and w4303;
w4305 <= not w4157 and not w4160;
w4306 <= not w4304 and not w4305;
w4307 <= not w4219 and not w4306;
w4308 <= not w3967 and not w4218;
w4309 <= not w4217 and w4308;
w4310 <= not w4307 and not w4309;
w4311 <= not b(15) and not w4310;
w4312 <= not w3986 and w4155;
w4313 <= not w4151 and w4312;
w4314 <= not w4152 and not w4155;
w4315 <= not w4313 and not w4314;
w4316 <= not w4219 and not w4315;
w4317 <= not w3976 and not w4218;
w4318 <= not w4217 and w4317;
w4319 <= not w4316 and not w4318;
w4320 <= not b(14) and not w4319;
w4321 <= not w3995 and w4150;
w4322 <= not w4146 and w4321;
w4323 <= not w4147 and not w4150;
w4324 <= not w4322 and not w4323;
w4325 <= not w4219 and not w4324;
w4326 <= not w3985 and not w4218;
w4327 <= not w4217 and w4326;
w4328 <= not w4325 and not w4327;
w4329 <= not b(13) and not w4328;
w4330 <= not w4004 and w4145;
w4331 <= not w4141 and w4330;
w4332 <= not w4142 and not w4145;
w4333 <= not w4331 and not w4332;
w4334 <= not w4219 and not w4333;
w4335 <= not w3994 and not w4218;
w4336 <= not w4217 and w4335;
w4337 <= not w4334 and not w4336;
w4338 <= not b(12) and not w4337;
w4339 <= not w4013 and w4140;
w4340 <= not w4136 and w4339;
w4341 <= not w4137 and not w4140;
w4342 <= not w4340 and not w4341;
w4343 <= not w4219 and not w4342;
w4344 <= not w4003 and not w4218;
w4345 <= not w4217 and w4344;
w4346 <= not w4343 and not w4345;
w4347 <= not b(11) and not w4346;
w4348 <= not w4022 and w4135;
w4349 <= not w4131 and w4348;
w4350 <= not w4132 and not w4135;
w4351 <= not w4349 and not w4350;
w4352 <= not w4219 and not w4351;
w4353 <= not w4012 and not w4218;
w4354 <= not w4217 and w4353;
w4355 <= not w4352 and not w4354;
w4356 <= not b(10) and not w4355;
w4357 <= not w4031 and w4130;
w4358 <= not w4126 and w4357;
w4359 <= not w4127 and not w4130;
w4360 <= not w4358 and not w4359;
w4361 <= not w4219 and not w4360;
w4362 <= not w4021 and not w4218;
w4363 <= not w4217 and w4362;
w4364 <= not w4361 and not w4363;
w4365 <= not b(9) and not w4364;
w4366 <= not w4040 and w4125;
w4367 <= not w4121 and w4366;
w4368 <= not w4122 and not w4125;
w4369 <= not w4367 and not w4368;
w4370 <= not w4219 and not w4369;
w4371 <= not w4030 and not w4218;
w4372 <= not w4217 and w4371;
w4373 <= not w4370 and not w4372;
w4374 <= not b(8) and not w4373;
w4375 <= not w4049 and w4120;
w4376 <= not w4116 and w4375;
w4377 <= not w4117 and not w4120;
w4378 <= not w4376 and not w4377;
w4379 <= not w4219 and not w4378;
w4380 <= not w4039 and not w4218;
w4381 <= not w4217 and w4380;
w4382 <= not w4379 and not w4381;
w4383 <= not b(7) and not w4382;
w4384 <= not w4058 and w4115;
w4385 <= not w4111 and w4384;
w4386 <= not w4112 and not w4115;
w4387 <= not w4385 and not w4386;
w4388 <= not w4219 and not w4387;
w4389 <= not w4048 and not w4218;
w4390 <= not w4217 and w4389;
w4391 <= not w4388 and not w4390;
w4392 <= not b(6) and not w4391;
w4393 <= not w4067 and w4110;
w4394 <= not w4106 and w4393;
w4395 <= not w4107 and not w4110;
w4396 <= not w4394 and not w4395;
w4397 <= not w4219 and not w4396;
w4398 <= not w4057 and not w4218;
w4399 <= not w4217 and w4398;
w4400 <= not w4397 and not w4399;
w4401 <= not b(5) and not w4400;
w4402 <= not w4075 and w4105;
w4403 <= not w4101 and w4402;
w4404 <= not w4102 and not w4105;
w4405 <= not w4403 and not w4404;
w4406 <= not w4219 and not w4405;
w4407 <= not w4066 and not w4218;
w4408 <= not w4217 and w4407;
w4409 <= not w4406 and not w4408;
w4410 <= not b(4) and not w4409;
w4411 <= not w4096 and w4100;
w4412 <= not w4095 and w4411;
w4413 <= not w4097 and not w4100;
w4414 <= not w4412 and not w4413;
w4415 <= not w4219 and not w4414;
w4416 <= not w4074 and not w4218;
w4417 <= not w4217 and w4416;
w4418 <= not w4415 and not w4417;
w4419 <= not b(3) and not w4418;
w4420 <= not w4092 and w4094;
w4421 <= not w4090 and w4420;
w4422 <= not w4095 and not w4421;
w4423 <= not w4219 and w4422;
w4424 <= not w4089 and not w4218;
w4425 <= not w4217 and w4424;
w4426 <= not w4423 and not w4425;
w4427 <= not b(2) and not w4426;
w4428 <= b(0) and not w4219;
w4429 <= a(40) and not w4428;
w4430 <= w4094 and not w4219;
w4431 <= not w4429 and not w4430;
w4432 <= b(1) and not w4431;
w4433 <= not b(1) and not w4430;
w4434 <= not w4429 and w4433;
w4435 <= not w4432 and not w4434;
w4436 <= not a(39) and b(0);
w4437 <= not w4435 and not w4436;
w4438 <= not b(1) and not w4431;
w4439 <= not w4437 and not w4438;
w4440 <= b(2) and not w4425;
w4441 <= not w4423 and w4440;
w4442 <= not w4427 and not w4441;
w4443 <= not w4439 and w4442;
w4444 <= not w4427 and not w4443;
w4445 <= b(3) and not w4417;
w4446 <= not w4415 and w4445;
w4447 <= not w4419 and not w4446;
w4448 <= not w4444 and w4447;
w4449 <= not w4419 and not w4448;
w4450 <= b(4) and not w4408;
w4451 <= not w4406 and w4450;
w4452 <= not w4410 and not w4451;
w4453 <= not w4449 and w4452;
w4454 <= not w4410 and not w4453;
w4455 <= b(5) and not w4399;
w4456 <= not w4397 and w4455;
w4457 <= not w4401 and not w4456;
w4458 <= not w4454 and w4457;
w4459 <= not w4401 and not w4458;
w4460 <= b(6) and not w4390;
w4461 <= not w4388 and w4460;
w4462 <= not w4392 and not w4461;
w4463 <= not w4459 and w4462;
w4464 <= not w4392 and not w4463;
w4465 <= b(7) and not w4381;
w4466 <= not w4379 and w4465;
w4467 <= not w4383 and not w4466;
w4468 <= not w4464 and w4467;
w4469 <= not w4383 and not w4468;
w4470 <= b(8) and not w4372;
w4471 <= not w4370 and w4470;
w4472 <= not w4374 and not w4471;
w4473 <= not w4469 and w4472;
w4474 <= not w4374 and not w4473;
w4475 <= b(9) and not w4363;
w4476 <= not w4361 and w4475;
w4477 <= not w4365 and not w4476;
w4478 <= not w4474 and w4477;
w4479 <= not w4365 and not w4478;
w4480 <= b(10) and not w4354;
w4481 <= not w4352 and w4480;
w4482 <= not w4356 and not w4481;
w4483 <= not w4479 and w4482;
w4484 <= not w4356 and not w4483;
w4485 <= b(11) and not w4345;
w4486 <= not w4343 and w4485;
w4487 <= not w4347 and not w4486;
w4488 <= not w4484 and w4487;
w4489 <= not w4347 and not w4488;
w4490 <= b(12) and not w4336;
w4491 <= not w4334 and w4490;
w4492 <= not w4338 and not w4491;
w4493 <= not w4489 and w4492;
w4494 <= not w4338 and not w4493;
w4495 <= b(13) and not w4327;
w4496 <= not w4325 and w4495;
w4497 <= not w4329 and not w4496;
w4498 <= not w4494 and w4497;
w4499 <= not w4329 and not w4498;
w4500 <= b(14) and not w4318;
w4501 <= not w4316 and w4500;
w4502 <= not w4320 and not w4501;
w4503 <= not w4499 and w4502;
w4504 <= not w4320 and not w4503;
w4505 <= b(15) and not w4309;
w4506 <= not w4307 and w4505;
w4507 <= not w4311 and not w4506;
w4508 <= not w4504 and w4507;
w4509 <= not w4311 and not w4508;
w4510 <= b(16) and not w4300;
w4511 <= not w4298 and w4510;
w4512 <= not w4302 and not w4511;
w4513 <= not w4509 and w4512;
w4514 <= not w4302 and not w4513;
w4515 <= b(17) and not w4291;
w4516 <= not w4289 and w4515;
w4517 <= not w4293 and not w4516;
w4518 <= not w4514 and w4517;
w4519 <= not w4293 and not w4518;
w4520 <= b(18) and not w4282;
w4521 <= not w4280 and w4520;
w4522 <= not w4284 and not w4521;
w4523 <= not w4519 and w4522;
w4524 <= not w4284 and not w4523;
w4525 <= b(19) and not w4273;
w4526 <= not w4271 and w4525;
w4527 <= not w4275 and not w4526;
w4528 <= not w4524 and w4527;
w4529 <= not w4275 and not w4528;
w4530 <= b(20) and not w4264;
w4531 <= not w4262 and w4530;
w4532 <= not w4266 and not w4531;
w4533 <= not w4529 and w4532;
w4534 <= not w4266 and not w4533;
w4535 <= b(21) and not w4255;
w4536 <= not w4253 and w4535;
w4537 <= not w4257 and not w4536;
w4538 <= not w4534 and w4537;
w4539 <= not w4257 and not w4538;
w4540 <= b(22) and not w4246;
w4541 <= not w4244 and w4540;
w4542 <= not w4248 and not w4541;
w4543 <= not w4539 and w4542;
w4544 <= not w4248 and not w4543;
w4545 <= b(23) and not w4226;
w4546 <= not w4224 and w4545;
w4547 <= not w4239 and not w4546;
w4548 <= not w4544 and w4547;
w4549 <= not w4239 and not w4548;
w4550 <= b(24) and not w4236;
w4551 <= not w4234 and w4550;
w4552 <= not w4238 and not w4551;
w4553 <= not w4549 and w4552;
w4554 <= not w4238 and not w4553;
w4555 <= w120 and w166;
w4556 <= w151 and w4555;
w4557 <= not w4554 and w4556;
w4558 <= not w4227 and not w4557;
w4559 <= not w4248 and w4547;
w4560 <= not w4543 and w4559;
w4561 <= not w4544 and not w4547;
w4562 <= not w4560 and not w4561;
w4563 <= w4556 and not w4562;
w4564 <= not w4554 and w4563;
w4565 <= not w4558 and not w4564;
w4566 <= not w4237 and not w4557;
w4567 <= not w4239 and w4552;
w4568 <= not w4548 and w4567;
w4569 <= not w4549 and not w4552;
w4570 <= not w4568 and not w4569;
w4571 <= w4557 and not w4570;
w4572 <= not w4566 and not w4571;
w4573 <= not b(25) and not w4572;
w4574 <= not b(24) and not w4565;
w4575 <= not w4247 and not w4557;
w4576 <= not w4257 and w4542;
w4577 <= not w4538 and w4576;
w4578 <= not w4539 and not w4542;
w4579 <= not w4577 and not w4578;
w4580 <= w4556 and not w4579;
w4581 <= not w4554 and w4580;
w4582 <= not w4575 and not w4581;
w4583 <= not b(23) and not w4582;
w4584 <= not w4256 and not w4557;
w4585 <= not w4266 and w4537;
w4586 <= not w4533 and w4585;
w4587 <= not w4534 and not w4537;
w4588 <= not w4586 and not w4587;
w4589 <= w4556 and not w4588;
w4590 <= not w4554 and w4589;
w4591 <= not w4584 and not w4590;
w4592 <= not b(22) and not w4591;
w4593 <= not w4265 and not w4557;
w4594 <= not w4275 and w4532;
w4595 <= not w4528 and w4594;
w4596 <= not w4529 and not w4532;
w4597 <= not w4595 and not w4596;
w4598 <= w4556 and not w4597;
w4599 <= not w4554 and w4598;
w4600 <= not w4593 and not w4599;
w4601 <= not b(21) and not w4600;
w4602 <= not w4274 and not w4557;
w4603 <= not w4284 and w4527;
w4604 <= not w4523 and w4603;
w4605 <= not w4524 and not w4527;
w4606 <= not w4604 and not w4605;
w4607 <= w4556 and not w4606;
w4608 <= not w4554 and w4607;
w4609 <= not w4602 and not w4608;
w4610 <= not b(20) and not w4609;
w4611 <= not w4283 and not w4557;
w4612 <= not w4293 and w4522;
w4613 <= not w4518 and w4612;
w4614 <= not w4519 and not w4522;
w4615 <= not w4613 and not w4614;
w4616 <= w4556 and not w4615;
w4617 <= not w4554 and w4616;
w4618 <= not w4611 and not w4617;
w4619 <= not b(19) and not w4618;
w4620 <= not w4292 and not w4557;
w4621 <= not w4302 and w4517;
w4622 <= not w4513 and w4621;
w4623 <= not w4514 and not w4517;
w4624 <= not w4622 and not w4623;
w4625 <= w4556 and not w4624;
w4626 <= not w4554 and w4625;
w4627 <= not w4620 and not w4626;
w4628 <= not b(18) and not w4627;
w4629 <= not w4301 and not w4557;
w4630 <= not w4311 and w4512;
w4631 <= not w4508 and w4630;
w4632 <= not w4509 and not w4512;
w4633 <= not w4631 and not w4632;
w4634 <= w4556 and not w4633;
w4635 <= not w4554 and w4634;
w4636 <= not w4629 and not w4635;
w4637 <= not b(17) and not w4636;
w4638 <= not w4310 and not w4557;
w4639 <= not w4320 and w4507;
w4640 <= not w4503 and w4639;
w4641 <= not w4504 and not w4507;
w4642 <= not w4640 and not w4641;
w4643 <= w4556 and not w4642;
w4644 <= not w4554 and w4643;
w4645 <= not w4638 and not w4644;
w4646 <= not b(16) and not w4645;
w4647 <= not w4319 and not w4557;
w4648 <= not w4329 and w4502;
w4649 <= not w4498 and w4648;
w4650 <= not w4499 and not w4502;
w4651 <= not w4649 and not w4650;
w4652 <= w4556 and not w4651;
w4653 <= not w4554 and w4652;
w4654 <= not w4647 and not w4653;
w4655 <= not b(15) and not w4654;
w4656 <= not w4328 and not w4557;
w4657 <= not w4338 and w4497;
w4658 <= not w4493 and w4657;
w4659 <= not w4494 and not w4497;
w4660 <= not w4658 and not w4659;
w4661 <= w4556 and not w4660;
w4662 <= not w4554 and w4661;
w4663 <= not w4656 and not w4662;
w4664 <= not b(14) and not w4663;
w4665 <= not w4337 and not w4557;
w4666 <= not w4347 and w4492;
w4667 <= not w4488 and w4666;
w4668 <= not w4489 and not w4492;
w4669 <= not w4667 and not w4668;
w4670 <= w4556 and not w4669;
w4671 <= not w4554 and w4670;
w4672 <= not w4665 and not w4671;
w4673 <= not b(13) and not w4672;
w4674 <= not w4346 and not w4557;
w4675 <= not w4356 and w4487;
w4676 <= not w4483 and w4675;
w4677 <= not w4484 and not w4487;
w4678 <= not w4676 and not w4677;
w4679 <= w4556 and not w4678;
w4680 <= not w4554 and w4679;
w4681 <= not w4674 and not w4680;
w4682 <= not b(12) and not w4681;
w4683 <= not w4355 and not w4557;
w4684 <= not w4365 and w4482;
w4685 <= not w4478 and w4684;
w4686 <= not w4479 and not w4482;
w4687 <= not w4685 and not w4686;
w4688 <= w4556 and not w4687;
w4689 <= not w4554 and w4688;
w4690 <= not w4683 and not w4689;
w4691 <= not b(11) and not w4690;
w4692 <= not w4364 and not w4557;
w4693 <= not w4374 and w4477;
w4694 <= not w4473 and w4693;
w4695 <= not w4474 and not w4477;
w4696 <= not w4694 and not w4695;
w4697 <= w4556 and not w4696;
w4698 <= not w4554 and w4697;
w4699 <= not w4692 and not w4698;
w4700 <= not b(10) and not w4699;
w4701 <= not w4373 and not w4557;
w4702 <= not w4383 and w4472;
w4703 <= not w4468 and w4702;
w4704 <= not w4469 and not w4472;
w4705 <= not w4703 and not w4704;
w4706 <= w4556 and not w4705;
w4707 <= not w4554 and w4706;
w4708 <= not w4701 and not w4707;
w4709 <= not b(9) and not w4708;
w4710 <= not w4382 and not w4557;
w4711 <= not w4392 and w4467;
w4712 <= not w4463 and w4711;
w4713 <= not w4464 and not w4467;
w4714 <= not w4712 and not w4713;
w4715 <= w4556 and not w4714;
w4716 <= not w4554 and w4715;
w4717 <= not w4710 and not w4716;
w4718 <= not b(8) and not w4717;
w4719 <= not w4391 and not w4557;
w4720 <= not w4401 and w4462;
w4721 <= not w4458 and w4720;
w4722 <= not w4459 and not w4462;
w4723 <= not w4721 and not w4722;
w4724 <= w4556 and not w4723;
w4725 <= not w4554 and w4724;
w4726 <= not w4719 and not w4725;
w4727 <= not b(7) and not w4726;
w4728 <= not w4400 and not w4557;
w4729 <= not w4410 and w4457;
w4730 <= not w4453 and w4729;
w4731 <= not w4454 and not w4457;
w4732 <= not w4730 and not w4731;
w4733 <= w4556 and not w4732;
w4734 <= not w4554 and w4733;
w4735 <= not w4728 and not w4734;
w4736 <= not b(6) and not w4735;
w4737 <= not w4409 and not w4557;
w4738 <= not w4419 and w4452;
w4739 <= not w4448 and w4738;
w4740 <= not w4449 and not w4452;
w4741 <= not w4739 and not w4740;
w4742 <= w4556 and not w4741;
w4743 <= not w4554 and w4742;
w4744 <= not w4737 and not w4743;
w4745 <= not b(5) and not w4744;
w4746 <= not w4418 and not w4557;
w4747 <= not w4427 and w4447;
w4748 <= not w4443 and w4747;
w4749 <= not w4444 and not w4447;
w4750 <= not w4748 and not w4749;
w4751 <= w4556 and not w4750;
w4752 <= not w4554 and w4751;
w4753 <= not w4746 and not w4752;
w4754 <= not b(4) and not w4753;
w4755 <= not w4426 and not w4557;
w4756 <= not w4438 and w4442;
w4757 <= not w4437 and w4756;
w4758 <= not w4439 and not w4442;
w4759 <= not w4757 and not w4758;
w4760 <= w4556 and not w4759;
w4761 <= not w4554 and w4760;
w4762 <= not w4755 and not w4761;
w4763 <= not b(3) and not w4762;
w4764 <= not w4431 and not w4557;
w4765 <= not w4434 and w4436;
w4766 <= not w4432 and w4765;
w4767 <= w4556 and not w4766;
w4768 <= not w4437 and w4767;
w4769 <= not w4554 and w4768;
w4770 <= not w4764 and not w4769;
w4771 <= not b(2) and not w4770;
w4772 <= b(0) and not b(25);
w4773 <= w48 and w4772;
w4774 <= w59 and w4773;
w4775 <= w84 and w4774;
w4776 <= w81 and w4775;
w4777 <= not w4554 and w4776;
w4778 <= a(39) and not w4777;
w4779 <= w119 and w4436;
w4780 <= w331 and w4779;
w4781 <= w341 and w4780;
w4782 <= w338 and w4781;
w4783 <= not w4554 and w4782;
w4784 <= not w4778 and not w4783;
w4785 <= b(1) and not w4784;
w4786 <= not b(1) and not w4783;
w4787 <= not w4778 and w4786;
w4788 <= not w4785 and not w4787;
w4789 <= not a(38) and b(0);
w4790 <= not w4788 and not w4789;
w4791 <= not b(1) and not w4784;
w4792 <= not w4790 and not w4791;
w4793 <= b(2) and not w4769;
w4794 <= not w4764 and w4793;
w4795 <= not w4771 and not w4794;
w4796 <= not w4792 and w4795;
w4797 <= not w4771 and not w4796;
w4798 <= b(3) and not w4761;
w4799 <= not w4755 and w4798;
w4800 <= not w4763 and not w4799;
w4801 <= not w4797 and w4800;
w4802 <= not w4763 and not w4801;
w4803 <= b(4) and not w4752;
w4804 <= not w4746 and w4803;
w4805 <= not w4754 and not w4804;
w4806 <= not w4802 and w4805;
w4807 <= not w4754 and not w4806;
w4808 <= b(5) and not w4743;
w4809 <= not w4737 and w4808;
w4810 <= not w4745 and not w4809;
w4811 <= not w4807 and w4810;
w4812 <= not w4745 and not w4811;
w4813 <= b(6) and not w4734;
w4814 <= not w4728 and w4813;
w4815 <= not w4736 and not w4814;
w4816 <= not w4812 and w4815;
w4817 <= not w4736 and not w4816;
w4818 <= b(7) and not w4725;
w4819 <= not w4719 and w4818;
w4820 <= not w4727 and not w4819;
w4821 <= not w4817 and w4820;
w4822 <= not w4727 and not w4821;
w4823 <= b(8) and not w4716;
w4824 <= not w4710 and w4823;
w4825 <= not w4718 and not w4824;
w4826 <= not w4822 and w4825;
w4827 <= not w4718 and not w4826;
w4828 <= b(9) and not w4707;
w4829 <= not w4701 and w4828;
w4830 <= not w4709 and not w4829;
w4831 <= not w4827 and w4830;
w4832 <= not w4709 and not w4831;
w4833 <= b(10) and not w4698;
w4834 <= not w4692 and w4833;
w4835 <= not w4700 and not w4834;
w4836 <= not w4832 and w4835;
w4837 <= not w4700 and not w4836;
w4838 <= b(11) and not w4689;
w4839 <= not w4683 and w4838;
w4840 <= not w4691 and not w4839;
w4841 <= not w4837 and w4840;
w4842 <= not w4691 and not w4841;
w4843 <= b(12) and not w4680;
w4844 <= not w4674 and w4843;
w4845 <= not w4682 and not w4844;
w4846 <= not w4842 and w4845;
w4847 <= not w4682 and not w4846;
w4848 <= b(13) and not w4671;
w4849 <= not w4665 and w4848;
w4850 <= not w4673 and not w4849;
w4851 <= not w4847 and w4850;
w4852 <= not w4673 and not w4851;
w4853 <= b(14) and not w4662;
w4854 <= not w4656 and w4853;
w4855 <= not w4664 and not w4854;
w4856 <= not w4852 and w4855;
w4857 <= not w4664 and not w4856;
w4858 <= b(15) and not w4653;
w4859 <= not w4647 and w4858;
w4860 <= not w4655 and not w4859;
w4861 <= not w4857 and w4860;
w4862 <= not w4655 and not w4861;
w4863 <= b(16) and not w4644;
w4864 <= not w4638 and w4863;
w4865 <= not w4646 and not w4864;
w4866 <= not w4862 and w4865;
w4867 <= not w4646 and not w4866;
w4868 <= b(17) and not w4635;
w4869 <= not w4629 and w4868;
w4870 <= not w4637 and not w4869;
w4871 <= not w4867 and w4870;
w4872 <= not w4637 and not w4871;
w4873 <= b(18) and not w4626;
w4874 <= not w4620 and w4873;
w4875 <= not w4628 and not w4874;
w4876 <= not w4872 and w4875;
w4877 <= not w4628 and not w4876;
w4878 <= b(19) and not w4617;
w4879 <= not w4611 and w4878;
w4880 <= not w4619 and not w4879;
w4881 <= not w4877 and w4880;
w4882 <= not w4619 and not w4881;
w4883 <= b(20) and not w4608;
w4884 <= not w4602 and w4883;
w4885 <= not w4610 and not w4884;
w4886 <= not w4882 and w4885;
w4887 <= not w4610 and not w4886;
w4888 <= b(21) and not w4599;
w4889 <= not w4593 and w4888;
w4890 <= not w4601 and not w4889;
w4891 <= not w4887 and w4890;
w4892 <= not w4601 and not w4891;
w4893 <= b(22) and not w4590;
w4894 <= not w4584 and w4893;
w4895 <= not w4592 and not w4894;
w4896 <= not w4892 and w4895;
w4897 <= not w4592 and not w4896;
w4898 <= b(23) and not w4581;
w4899 <= not w4575 and w4898;
w4900 <= not w4583 and not w4899;
w4901 <= not w4897 and w4900;
w4902 <= not w4583 and not w4901;
w4903 <= b(24) and not w4564;
w4904 <= not w4558 and w4903;
w4905 <= not w4574 and not w4904;
w4906 <= not w4902 and w4905;
w4907 <= not w4574 and not w4906;
w4908 <= b(25) and not w4566;
w4909 <= not w4571 and w4908;
w4910 <= not w4573 and not w4909;
w4911 <= not w4907 and w4910;
w4912 <= not w4573 and not w4911;
w4913 <= w48 and w59;
w4914 <= w84 and w4913;
w4915 <= w81 and w4914;
w4916 <= not w4912 and w4915;
w4917 <= not w4565 and not w4916;
w4918 <= not w4583 and w4905;
w4919 <= not w4901 and w4918;
w4920 <= not w4902 and not w4905;
w4921 <= not w4919 and not w4920;
w4922 <= w4915 and not w4921;
w4923 <= not w4912 and w4922;
w4924 <= not w4917 and not w4923;
w4925 <= not b(25) and not w4924;
w4926 <= not w4582 and not w4916;
w4927 <= not w4592 and w4900;
w4928 <= not w4896 and w4927;
w4929 <= not w4897 and not w4900;
w4930 <= not w4928 and not w4929;
w4931 <= w4915 and not w4930;
w4932 <= not w4912 and w4931;
w4933 <= not w4926 and not w4932;
w4934 <= not b(24) and not w4933;
w4935 <= not w4591 and not w4916;
w4936 <= not w4601 and w4895;
w4937 <= not w4891 and w4936;
w4938 <= not w4892 and not w4895;
w4939 <= not w4937 and not w4938;
w4940 <= w4915 and not w4939;
w4941 <= not w4912 and w4940;
w4942 <= not w4935 and not w4941;
w4943 <= not b(23) and not w4942;
w4944 <= not w4600 and not w4916;
w4945 <= not w4610 and w4890;
w4946 <= not w4886 and w4945;
w4947 <= not w4887 and not w4890;
w4948 <= not w4946 and not w4947;
w4949 <= w4915 and not w4948;
w4950 <= not w4912 and w4949;
w4951 <= not w4944 and not w4950;
w4952 <= not b(22) and not w4951;
w4953 <= not w4609 and not w4916;
w4954 <= not w4619 and w4885;
w4955 <= not w4881 and w4954;
w4956 <= not w4882 and not w4885;
w4957 <= not w4955 and not w4956;
w4958 <= w4915 and not w4957;
w4959 <= not w4912 and w4958;
w4960 <= not w4953 and not w4959;
w4961 <= not b(21) and not w4960;
w4962 <= not w4618 and not w4916;
w4963 <= not w4628 and w4880;
w4964 <= not w4876 and w4963;
w4965 <= not w4877 and not w4880;
w4966 <= not w4964 and not w4965;
w4967 <= w4915 and not w4966;
w4968 <= not w4912 and w4967;
w4969 <= not w4962 and not w4968;
w4970 <= not b(20) and not w4969;
w4971 <= not w4627 and not w4916;
w4972 <= not w4637 and w4875;
w4973 <= not w4871 and w4972;
w4974 <= not w4872 and not w4875;
w4975 <= not w4973 and not w4974;
w4976 <= w4915 and not w4975;
w4977 <= not w4912 and w4976;
w4978 <= not w4971 and not w4977;
w4979 <= not b(19) and not w4978;
w4980 <= not w4636 and not w4916;
w4981 <= not w4646 and w4870;
w4982 <= not w4866 and w4981;
w4983 <= not w4867 and not w4870;
w4984 <= not w4982 and not w4983;
w4985 <= w4915 and not w4984;
w4986 <= not w4912 and w4985;
w4987 <= not w4980 and not w4986;
w4988 <= not b(18) and not w4987;
w4989 <= not w4645 and not w4916;
w4990 <= not w4655 and w4865;
w4991 <= not w4861 and w4990;
w4992 <= not w4862 and not w4865;
w4993 <= not w4991 and not w4992;
w4994 <= w4915 and not w4993;
w4995 <= not w4912 and w4994;
w4996 <= not w4989 and not w4995;
w4997 <= not b(17) and not w4996;
w4998 <= not w4654 and not w4916;
w4999 <= not w4664 and w4860;
w5000 <= not w4856 and w4999;
w5001 <= not w4857 and not w4860;
w5002 <= not w5000 and not w5001;
w5003 <= w4915 and not w5002;
w5004 <= not w4912 and w5003;
w5005 <= not w4998 and not w5004;
w5006 <= not b(16) and not w5005;
w5007 <= not w4663 and not w4916;
w5008 <= not w4673 and w4855;
w5009 <= not w4851 and w5008;
w5010 <= not w4852 and not w4855;
w5011 <= not w5009 and not w5010;
w5012 <= w4915 and not w5011;
w5013 <= not w4912 and w5012;
w5014 <= not w5007 and not w5013;
w5015 <= not b(15) and not w5014;
w5016 <= not w4672 and not w4916;
w5017 <= not w4682 and w4850;
w5018 <= not w4846 and w5017;
w5019 <= not w4847 and not w4850;
w5020 <= not w5018 and not w5019;
w5021 <= w4915 and not w5020;
w5022 <= not w4912 and w5021;
w5023 <= not w5016 and not w5022;
w5024 <= not b(14) and not w5023;
w5025 <= not w4681 and not w4916;
w5026 <= not w4691 and w4845;
w5027 <= not w4841 and w5026;
w5028 <= not w4842 and not w4845;
w5029 <= not w5027 and not w5028;
w5030 <= w4915 and not w5029;
w5031 <= not w4912 and w5030;
w5032 <= not w5025 and not w5031;
w5033 <= not b(13) and not w5032;
w5034 <= not w4690 and not w4916;
w5035 <= not w4700 and w4840;
w5036 <= not w4836 and w5035;
w5037 <= not w4837 and not w4840;
w5038 <= not w5036 and not w5037;
w5039 <= w4915 and not w5038;
w5040 <= not w4912 and w5039;
w5041 <= not w5034 and not w5040;
w5042 <= not b(12) and not w5041;
w5043 <= not w4699 and not w4916;
w5044 <= not w4709 and w4835;
w5045 <= not w4831 and w5044;
w5046 <= not w4832 and not w4835;
w5047 <= not w5045 and not w5046;
w5048 <= w4915 and not w5047;
w5049 <= not w4912 and w5048;
w5050 <= not w5043 and not w5049;
w5051 <= not b(11) and not w5050;
w5052 <= not w4708 and not w4916;
w5053 <= not w4718 and w4830;
w5054 <= not w4826 and w5053;
w5055 <= not w4827 and not w4830;
w5056 <= not w5054 and not w5055;
w5057 <= w4915 and not w5056;
w5058 <= not w4912 and w5057;
w5059 <= not w5052 and not w5058;
w5060 <= not b(10) and not w5059;
w5061 <= not w4717 and not w4916;
w5062 <= not w4727 and w4825;
w5063 <= not w4821 and w5062;
w5064 <= not w4822 and not w4825;
w5065 <= not w5063 and not w5064;
w5066 <= w4915 and not w5065;
w5067 <= not w4912 and w5066;
w5068 <= not w5061 and not w5067;
w5069 <= not b(9) and not w5068;
w5070 <= not w4726 and not w4916;
w5071 <= not w4736 and w4820;
w5072 <= not w4816 and w5071;
w5073 <= not w4817 and not w4820;
w5074 <= not w5072 and not w5073;
w5075 <= w4915 and not w5074;
w5076 <= not w4912 and w5075;
w5077 <= not w5070 and not w5076;
w5078 <= not b(8) and not w5077;
w5079 <= not w4735 and not w4916;
w5080 <= not w4745 and w4815;
w5081 <= not w4811 and w5080;
w5082 <= not w4812 and not w4815;
w5083 <= not w5081 and not w5082;
w5084 <= w4915 and not w5083;
w5085 <= not w4912 and w5084;
w5086 <= not w5079 and not w5085;
w5087 <= not b(7) and not w5086;
w5088 <= not w4744 and not w4916;
w5089 <= not w4754 and w4810;
w5090 <= not w4806 and w5089;
w5091 <= not w4807 and not w4810;
w5092 <= not w5090 and not w5091;
w5093 <= w4915 and not w5092;
w5094 <= not w4912 and w5093;
w5095 <= not w5088 and not w5094;
w5096 <= not b(6) and not w5095;
w5097 <= not w4753 and not w4916;
w5098 <= not w4763 and w4805;
w5099 <= not w4801 and w5098;
w5100 <= not w4802 and not w4805;
w5101 <= not w5099 and not w5100;
w5102 <= w4915 and not w5101;
w5103 <= not w4912 and w5102;
w5104 <= not w5097 and not w5103;
w5105 <= not b(5) and not w5104;
w5106 <= not w4762 and not w4916;
w5107 <= not w4771 and w4800;
w5108 <= not w4796 and w5107;
w5109 <= not w4797 and not w4800;
w5110 <= not w5108 and not w5109;
w5111 <= w4915 and not w5110;
w5112 <= not w4912 and w5111;
w5113 <= not w5106 and not w5112;
w5114 <= not b(4) and not w5113;
w5115 <= not w4770 and not w4916;
w5116 <= not w4791 and w4795;
w5117 <= not w4790 and w5116;
w5118 <= not w4792 and not w4795;
w5119 <= not w5117 and not w5118;
w5120 <= w4915 and not w5119;
w5121 <= not w4912 and w5120;
w5122 <= not w5115 and not w5121;
w5123 <= not b(3) and not w5122;
w5124 <= not w4784 and not w4916;
w5125 <= not w4787 and w4789;
w5126 <= not w4785 and w5125;
w5127 <= w4915 and not w5126;
w5128 <= not w4790 and w5127;
w5129 <= not w4912 and w5128;
w5130 <= not w5124 and not w5129;
w5131 <= not b(2) and not w5130;
w5132 <= b(0) and not b(26);
w5133 <= w118 and w5132;
w5134 <= w116 and w5133;
w5135 <= w166 and w5134;
w5136 <= w151 and w5135;
w5137 <= not w4912 and w5136;
w5138 <= a(38) and not w5137;
w5139 <= w48 and w4789;
w5140 <= w59 and w5139;
w5141 <= w84 and w5140;
w5142 <= w81 and w5141;
w5143 <= not w4912 and w5142;
w5144 <= not w5138 and not w5143;
w5145 <= b(1) and not w5144;
w5146 <= not b(1) and not w5143;
w5147 <= not w5138 and w5146;
w5148 <= not w5145 and not w5147;
w5149 <= not a(37) and b(0);
w5150 <= not w5148 and not w5149;
w5151 <= not b(1) and not w5144;
w5152 <= not w5150 and not w5151;
w5153 <= b(2) and not w5129;
w5154 <= not w5124 and w5153;
w5155 <= not w5131 and not w5154;
w5156 <= not w5152 and w5155;
w5157 <= not w5131 and not w5156;
w5158 <= b(3) and not w5121;
w5159 <= not w5115 and w5158;
w5160 <= not w5123 and not w5159;
w5161 <= not w5157 and w5160;
w5162 <= not w5123 and not w5161;
w5163 <= b(4) and not w5112;
w5164 <= not w5106 and w5163;
w5165 <= not w5114 and not w5164;
w5166 <= not w5162 and w5165;
w5167 <= not w5114 and not w5166;
w5168 <= b(5) and not w5103;
w5169 <= not w5097 and w5168;
w5170 <= not w5105 and not w5169;
w5171 <= not w5167 and w5170;
w5172 <= not w5105 and not w5171;
w5173 <= b(6) and not w5094;
w5174 <= not w5088 and w5173;
w5175 <= not w5096 and not w5174;
w5176 <= not w5172 and w5175;
w5177 <= not w5096 and not w5176;
w5178 <= b(7) and not w5085;
w5179 <= not w5079 and w5178;
w5180 <= not w5087 and not w5179;
w5181 <= not w5177 and w5180;
w5182 <= not w5087 and not w5181;
w5183 <= b(8) and not w5076;
w5184 <= not w5070 and w5183;
w5185 <= not w5078 and not w5184;
w5186 <= not w5182 and w5185;
w5187 <= not w5078 and not w5186;
w5188 <= b(9) and not w5067;
w5189 <= not w5061 and w5188;
w5190 <= not w5069 and not w5189;
w5191 <= not w5187 and w5190;
w5192 <= not w5069 and not w5191;
w5193 <= b(10) and not w5058;
w5194 <= not w5052 and w5193;
w5195 <= not w5060 and not w5194;
w5196 <= not w5192 and w5195;
w5197 <= not w5060 and not w5196;
w5198 <= b(11) and not w5049;
w5199 <= not w5043 and w5198;
w5200 <= not w5051 and not w5199;
w5201 <= not w5197 and w5200;
w5202 <= not w5051 and not w5201;
w5203 <= b(12) and not w5040;
w5204 <= not w5034 and w5203;
w5205 <= not w5042 and not w5204;
w5206 <= not w5202 and w5205;
w5207 <= not w5042 and not w5206;
w5208 <= b(13) and not w5031;
w5209 <= not w5025 and w5208;
w5210 <= not w5033 and not w5209;
w5211 <= not w5207 and w5210;
w5212 <= not w5033 and not w5211;
w5213 <= b(14) and not w5022;
w5214 <= not w5016 and w5213;
w5215 <= not w5024 and not w5214;
w5216 <= not w5212 and w5215;
w5217 <= not w5024 and not w5216;
w5218 <= b(15) and not w5013;
w5219 <= not w5007 and w5218;
w5220 <= not w5015 and not w5219;
w5221 <= not w5217 and w5220;
w5222 <= not w5015 and not w5221;
w5223 <= b(16) and not w5004;
w5224 <= not w4998 and w5223;
w5225 <= not w5006 and not w5224;
w5226 <= not w5222 and w5225;
w5227 <= not w5006 and not w5226;
w5228 <= b(17) and not w4995;
w5229 <= not w4989 and w5228;
w5230 <= not w4997 and not w5229;
w5231 <= not w5227 and w5230;
w5232 <= not w4997 and not w5231;
w5233 <= b(18) and not w4986;
w5234 <= not w4980 and w5233;
w5235 <= not w4988 and not w5234;
w5236 <= not w5232 and w5235;
w5237 <= not w4988 and not w5236;
w5238 <= b(19) and not w4977;
w5239 <= not w4971 and w5238;
w5240 <= not w4979 and not w5239;
w5241 <= not w5237 and w5240;
w5242 <= not w4979 and not w5241;
w5243 <= b(20) and not w4968;
w5244 <= not w4962 and w5243;
w5245 <= not w4970 and not w5244;
w5246 <= not w5242 and w5245;
w5247 <= not w4970 and not w5246;
w5248 <= b(21) and not w4959;
w5249 <= not w4953 and w5248;
w5250 <= not w4961 and not w5249;
w5251 <= not w5247 and w5250;
w5252 <= not w4961 and not w5251;
w5253 <= b(22) and not w4950;
w5254 <= not w4944 and w5253;
w5255 <= not w4952 and not w5254;
w5256 <= not w5252 and w5255;
w5257 <= not w4952 and not w5256;
w5258 <= b(23) and not w4941;
w5259 <= not w4935 and w5258;
w5260 <= not w4943 and not w5259;
w5261 <= not w5257 and w5260;
w5262 <= not w4943 and not w5261;
w5263 <= b(24) and not w4932;
w5264 <= not w4926 and w5263;
w5265 <= not w4934 and not w5264;
w5266 <= not w5262 and w5265;
w5267 <= not w4934 and not w5266;
w5268 <= b(25) and not w4923;
w5269 <= not w4917 and w5268;
w5270 <= not w4925 and not w5269;
w5271 <= not w5267 and w5270;
w5272 <= not w4925 and not w5271;
w5273 <= not w4572 and not w4916;
w5274 <= not w4574 and w4910;
w5275 <= not w4906 and w5274;
w5276 <= not w4907 and not w4910;
w5277 <= not w5275 and not w5276;
w5278 <= w4916 and not w5277;
w5279 <= not w5273 and not w5278;
w5280 <= not b(26) and not w5279;
w5281 <= b(26) and not w5273;
w5282 <= not w5278 and w5281;
w5283 <= w116 and w118;
w5284 <= w166 and w5283;
w5285 <= w151 and w5284;
w5286 <= not w5282 and w5285;
w5287 <= not w5280 and w5286;
w5288 <= not w5272 and w5287;
w5289 <= w4915 and not w5279;
w5290 <= not w5288 and not w5289;
w5291 <= not w4934 and w5270;
w5292 <= not w5266 and w5291;
w5293 <= not w5267 and not w5270;
w5294 <= not w5292 and not w5293;
w5295 <= not w5290 and not w5294;
w5296 <= not w4924 and not w5289;
w5297 <= not w5288 and w5296;
w5298 <= not w5295 and not w5297;
w5299 <= not w4925 and not w5282;
w5300 <= not w5280 and w5299;
w5301 <= not w5271 and w5300;
w5302 <= not w5280 and not w5282;
w5303 <= not w5272 and not w5302;
w5304 <= not w5301 and not w5303;
w5305 <= not w5290 and not w5304;
w5306 <= not w5279 and not w5289;
w5307 <= not w5288 and w5306;
w5308 <= not w5305 and not w5307;
w5309 <= not b(27) and not w5308;
w5310 <= not b(26) and not w5298;
w5311 <= not w4943 and w5265;
w5312 <= not w5261 and w5311;
w5313 <= not w5262 and not w5265;
w5314 <= not w5312 and not w5313;
w5315 <= not w5290 and not w5314;
w5316 <= not w4933 and not w5289;
w5317 <= not w5288 and w5316;
w5318 <= not w5315 and not w5317;
w5319 <= not b(25) and not w5318;
w5320 <= not w4952 and w5260;
w5321 <= not w5256 and w5320;
w5322 <= not w5257 and not w5260;
w5323 <= not w5321 and not w5322;
w5324 <= not w5290 and not w5323;
w5325 <= not w4942 and not w5289;
w5326 <= not w5288 and w5325;
w5327 <= not w5324 and not w5326;
w5328 <= not b(24) and not w5327;
w5329 <= not w4961 and w5255;
w5330 <= not w5251 and w5329;
w5331 <= not w5252 and not w5255;
w5332 <= not w5330 and not w5331;
w5333 <= not w5290 and not w5332;
w5334 <= not w4951 and not w5289;
w5335 <= not w5288 and w5334;
w5336 <= not w5333 and not w5335;
w5337 <= not b(23) and not w5336;
w5338 <= not w4970 and w5250;
w5339 <= not w5246 and w5338;
w5340 <= not w5247 and not w5250;
w5341 <= not w5339 and not w5340;
w5342 <= not w5290 and not w5341;
w5343 <= not w4960 and not w5289;
w5344 <= not w5288 and w5343;
w5345 <= not w5342 and not w5344;
w5346 <= not b(22) and not w5345;
w5347 <= not w4979 and w5245;
w5348 <= not w5241 and w5347;
w5349 <= not w5242 and not w5245;
w5350 <= not w5348 and not w5349;
w5351 <= not w5290 and not w5350;
w5352 <= not w4969 and not w5289;
w5353 <= not w5288 and w5352;
w5354 <= not w5351 and not w5353;
w5355 <= not b(21) and not w5354;
w5356 <= not w4988 and w5240;
w5357 <= not w5236 and w5356;
w5358 <= not w5237 and not w5240;
w5359 <= not w5357 and not w5358;
w5360 <= not w5290 and not w5359;
w5361 <= not w4978 and not w5289;
w5362 <= not w5288 and w5361;
w5363 <= not w5360 and not w5362;
w5364 <= not b(20) and not w5363;
w5365 <= not w4997 and w5235;
w5366 <= not w5231 and w5365;
w5367 <= not w5232 and not w5235;
w5368 <= not w5366 and not w5367;
w5369 <= not w5290 and not w5368;
w5370 <= not w4987 and not w5289;
w5371 <= not w5288 and w5370;
w5372 <= not w5369 and not w5371;
w5373 <= not b(19) and not w5372;
w5374 <= not w5006 and w5230;
w5375 <= not w5226 and w5374;
w5376 <= not w5227 and not w5230;
w5377 <= not w5375 and not w5376;
w5378 <= not w5290 and not w5377;
w5379 <= not w4996 and not w5289;
w5380 <= not w5288 and w5379;
w5381 <= not w5378 and not w5380;
w5382 <= not b(18) and not w5381;
w5383 <= not w5015 and w5225;
w5384 <= not w5221 and w5383;
w5385 <= not w5222 and not w5225;
w5386 <= not w5384 and not w5385;
w5387 <= not w5290 and not w5386;
w5388 <= not w5005 and not w5289;
w5389 <= not w5288 and w5388;
w5390 <= not w5387 and not w5389;
w5391 <= not b(17) and not w5390;
w5392 <= not w5024 and w5220;
w5393 <= not w5216 and w5392;
w5394 <= not w5217 and not w5220;
w5395 <= not w5393 and not w5394;
w5396 <= not w5290 and not w5395;
w5397 <= not w5014 and not w5289;
w5398 <= not w5288 and w5397;
w5399 <= not w5396 and not w5398;
w5400 <= not b(16) and not w5399;
w5401 <= not w5033 and w5215;
w5402 <= not w5211 and w5401;
w5403 <= not w5212 and not w5215;
w5404 <= not w5402 and not w5403;
w5405 <= not w5290 and not w5404;
w5406 <= not w5023 and not w5289;
w5407 <= not w5288 and w5406;
w5408 <= not w5405 and not w5407;
w5409 <= not b(15) and not w5408;
w5410 <= not w5042 and w5210;
w5411 <= not w5206 and w5410;
w5412 <= not w5207 and not w5210;
w5413 <= not w5411 and not w5412;
w5414 <= not w5290 and not w5413;
w5415 <= not w5032 and not w5289;
w5416 <= not w5288 and w5415;
w5417 <= not w5414 and not w5416;
w5418 <= not b(14) and not w5417;
w5419 <= not w5051 and w5205;
w5420 <= not w5201 and w5419;
w5421 <= not w5202 and not w5205;
w5422 <= not w5420 and not w5421;
w5423 <= not w5290 and not w5422;
w5424 <= not w5041 and not w5289;
w5425 <= not w5288 and w5424;
w5426 <= not w5423 and not w5425;
w5427 <= not b(13) and not w5426;
w5428 <= not w5060 and w5200;
w5429 <= not w5196 and w5428;
w5430 <= not w5197 and not w5200;
w5431 <= not w5429 and not w5430;
w5432 <= not w5290 and not w5431;
w5433 <= not w5050 and not w5289;
w5434 <= not w5288 and w5433;
w5435 <= not w5432 and not w5434;
w5436 <= not b(12) and not w5435;
w5437 <= not w5069 and w5195;
w5438 <= not w5191 and w5437;
w5439 <= not w5192 and not w5195;
w5440 <= not w5438 and not w5439;
w5441 <= not w5290 and not w5440;
w5442 <= not w5059 and not w5289;
w5443 <= not w5288 and w5442;
w5444 <= not w5441 and not w5443;
w5445 <= not b(11) and not w5444;
w5446 <= not w5078 and w5190;
w5447 <= not w5186 and w5446;
w5448 <= not w5187 and not w5190;
w5449 <= not w5447 and not w5448;
w5450 <= not w5290 and not w5449;
w5451 <= not w5068 and not w5289;
w5452 <= not w5288 and w5451;
w5453 <= not w5450 and not w5452;
w5454 <= not b(10) and not w5453;
w5455 <= not w5087 and w5185;
w5456 <= not w5181 and w5455;
w5457 <= not w5182 and not w5185;
w5458 <= not w5456 and not w5457;
w5459 <= not w5290 and not w5458;
w5460 <= not w5077 and not w5289;
w5461 <= not w5288 and w5460;
w5462 <= not w5459 and not w5461;
w5463 <= not b(9) and not w5462;
w5464 <= not w5096 and w5180;
w5465 <= not w5176 and w5464;
w5466 <= not w5177 and not w5180;
w5467 <= not w5465 and not w5466;
w5468 <= not w5290 and not w5467;
w5469 <= not w5086 and not w5289;
w5470 <= not w5288 and w5469;
w5471 <= not w5468 and not w5470;
w5472 <= not b(8) and not w5471;
w5473 <= not w5105 and w5175;
w5474 <= not w5171 and w5473;
w5475 <= not w5172 and not w5175;
w5476 <= not w5474 and not w5475;
w5477 <= not w5290 and not w5476;
w5478 <= not w5095 and not w5289;
w5479 <= not w5288 and w5478;
w5480 <= not w5477 and not w5479;
w5481 <= not b(7) and not w5480;
w5482 <= not w5114 and w5170;
w5483 <= not w5166 and w5482;
w5484 <= not w5167 and not w5170;
w5485 <= not w5483 and not w5484;
w5486 <= not w5290 and not w5485;
w5487 <= not w5104 and not w5289;
w5488 <= not w5288 and w5487;
w5489 <= not w5486 and not w5488;
w5490 <= not b(6) and not w5489;
w5491 <= not w5123 and w5165;
w5492 <= not w5161 and w5491;
w5493 <= not w5162 and not w5165;
w5494 <= not w5492 and not w5493;
w5495 <= not w5290 and not w5494;
w5496 <= not w5113 and not w5289;
w5497 <= not w5288 and w5496;
w5498 <= not w5495 and not w5497;
w5499 <= not b(5) and not w5498;
w5500 <= not w5131 and w5160;
w5501 <= not w5156 and w5500;
w5502 <= not w5157 and not w5160;
w5503 <= not w5501 and not w5502;
w5504 <= not w5290 and not w5503;
w5505 <= not w5122 and not w5289;
w5506 <= not w5288 and w5505;
w5507 <= not w5504 and not w5506;
w5508 <= not b(4) and not w5507;
w5509 <= not w5151 and w5155;
w5510 <= not w5150 and w5509;
w5511 <= not w5152 and not w5155;
w5512 <= not w5510 and not w5511;
w5513 <= not w5290 and not w5512;
w5514 <= not w5130 and not w5289;
w5515 <= not w5288 and w5514;
w5516 <= not w5513 and not w5515;
w5517 <= not b(3) and not w5516;
w5518 <= not w5147 and w5149;
w5519 <= not w5145 and w5518;
w5520 <= not w5150 and not w5519;
w5521 <= not w5290 and w5520;
w5522 <= not w5144 and not w5289;
w5523 <= not w5288 and w5522;
w5524 <= not w5521 and not w5523;
w5525 <= not b(2) and not w5524;
w5526 <= b(0) and not w5290;
w5527 <= a(37) and not w5526;
w5528 <= w5149 and not w5290;
w5529 <= not w5527 and not w5528;
w5530 <= b(1) and not w5529;
w5531 <= not b(1) and not w5528;
w5532 <= not w5527 and w5531;
w5533 <= not w5530 and not w5532;
w5534 <= not a(36) and b(0);
w5535 <= not w5533 and not w5534;
w5536 <= not b(1) and not w5529;
w5537 <= not w5535 and not w5536;
w5538 <= b(2) and not w5523;
w5539 <= not w5521 and w5538;
w5540 <= not w5525 and not w5539;
w5541 <= not w5537 and w5540;
w5542 <= not w5525 and not w5541;
w5543 <= b(3) and not w5515;
w5544 <= not w5513 and w5543;
w5545 <= not w5517 and not w5544;
w5546 <= not w5542 and w5545;
w5547 <= not w5517 and not w5546;
w5548 <= b(4) and not w5506;
w5549 <= not w5504 and w5548;
w5550 <= not w5508 and not w5549;
w5551 <= not w5547 and w5550;
w5552 <= not w5508 and not w5551;
w5553 <= b(5) and not w5497;
w5554 <= not w5495 and w5553;
w5555 <= not w5499 and not w5554;
w5556 <= not w5552 and w5555;
w5557 <= not w5499 and not w5556;
w5558 <= b(6) and not w5488;
w5559 <= not w5486 and w5558;
w5560 <= not w5490 and not w5559;
w5561 <= not w5557 and w5560;
w5562 <= not w5490 and not w5561;
w5563 <= b(7) and not w5479;
w5564 <= not w5477 and w5563;
w5565 <= not w5481 and not w5564;
w5566 <= not w5562 and w5565;
w5567 <= not w5481 and not w5566;
w5568 <= b(8) and not w5470;
w5569 <= not w5468 and w5568;
w5570 <= not w5472 and not w5569;
w5571 <= not w5567 and w5570;
w5572 <= not w5472 and not w5571;
w5573 <= b(9) and not w5461;
w5574 <= not w5459 and w5573;
w5575 <= not w5463 and not w5574;
w5576 <= not w5572 and w5575;
w5577 <= not w5463 and not w5576;
w5578 <= b(10) and not w5452;
w5579 <= not w5450 and w5578;
w5580 <= not w5454 and not w5579;
w5581 <= not w5577 and w5580;
w5582 <= not w5454 and not w5581;
w5583 <= b(11) and not w5443;
w5584 <= not w5441 and w5583;
w5585 <= not w5445 and not w5584;
w5586 <= not w5582 and w5585;
w5587 <= not w5445 and not w5586;
w5588 <= b(12) and not w5434;
w5589 <= not w5432 and w5588;
w5590 <= not w5436 and not w5589;
w5591 <= not w5587 and w5590;
w5592 <= not w5436 and not w5591;
w5593 <= b(13) and not w5425;
w5594 <= not w5423 and w5593;
w5595 <= not w5427 and not w5594;
w5596 <= not w5592 and w5595;
w5597 <= not w5427 and not w5596;
w5598 <= b(14) and not w5416;
w5599 <= not w5414 and w5598;
w5600 <= not w5418 and not w5599;
w5601 <= not w5597 and w5600;
w5602 <= not w5418 and not w5601;
w5603 <= b(15) and not w5407;
w5604 <= not w5405 and w5603;
w5605 <= not w5409 and not w5604;
w5606 <= not w5602 and w5605;
w5607 <= not w5409 and not w5606;
w5608 <= b(16) and not w5398;
w5609 <= not w5396 and w5608;
w5610 <= not w5400 and not w5609;
w5611 <= not w5607 and w5610;
w5612 <= not w5400 and not w5611;
w5613 <= b(17) and not w5389;
w5614 <= not w5387 and w5613;
w5615 <= not w5391 and not w5614;
w5616 <= not w5612 and w5615;
w5617 <= not w5391 and not w5616;
w5618 <= b(18) and not w5380;
w5619 <= not w5378 and w5618;
w5620 <= not w5382 and not w5619;
w5621 <= not w5617 and w5620;
w5622 <= not w5382 and not w5621;
w5623 <= b(19) and not w5371;
w5624 <= not w5369 and w5623;
w5625 <= not w5373 and not w5624;
w5626 <= not w5622 and w5625;
w5627 <= not w5373 and not w5626;
w5628 <= b(20) and not w5362;
w5629 <= not w5360 and w5628;
w5630 <= not w5364 and not w5629;
w5631 <= not w5627 and w5630;
w5632 <= not w5364 and not w5631;
w5633 <= b(21) and not w5353;
w5634 <= not w5351 and w5633;
w5635 <= not w5355 and not w5634;
w5636 <= not w5632 and w5635;
w5637 <= not w5355 and not w5636;
w5638 <= b(22) and not w5344;
w5639 <= not w5342 and w5638;
w5640 <= not w5346 and not w5639;
w5641 <= not w5637 and w5640;
w5642 <= not w5346 and not w5641;
w5643 <= b(23) and not w5335;
w5644 <= not w5333 and w5643;
w5645 <= not w5337 and not w5644;
w5646 <= not w5642 and w5645;
w5647 <= not w5337 and not w5646;
w5648 <= b(24) and not w5326;
w5649 <= not w5324 and w5648;
w5650 <= not w5328 and not w5649;
w5651 <= not w5647 and w5650;
w5652 <= not w5328 and not w5651;
w5653 <= b(25) and not w5317;
w5654 <= not w5315 and w5653;
w5655 <= not w5319 and not w5654;
w5656 <= not w5652 and w5655;
w5657 <= not w5319 and not w5656;
w5658 <= b(26) and not w5297;
w5659 <= not w5295 and w5658;
w5660 <= not w5310 and not w5659;
w5661 <= not w5657 and w5660;
w5662 <= not w5310 and not w5661;
w5663 <= b(27) and not w5307;
w5664 <= not w5305 and w5663;
w5665 <= not w5309 and not w5664;
w5666 <= not w5662 and w5665;
w5667 <= not w5309 and not w5666;
w5668 <= w46 and w60;
w5669 <= w31 and w5668;
w5670 <= not w5667 and w5669;
w5671 <= not w5298 and not w5670;
w5672 <= not w5319 and w5660;
w5673 <= not w5656 and w5672;
w5674 <= not w5657 and not w5660;
w5675 <= not w5673 and not w5674;
w5676 <= w5669 and not w5675;
w5677 <= not w5667 and w5676;
w5678 <= not w5671 and not w5677;
w5679 <= not w5308 and not w5670;
w5680 <= not w5310 and w5665;
w5681 <= not w5661 and w5680;
w5682 <= not w5662 and not w5665;
w5683 <= not w5681 and not w5682;
w5684 <= w5670 and not w5683;
w5685 <= not w5679 and not w5684;
w5686 <= not b(28) and not w5685;
w5687 <= not b(27) and not w5678;
w5688 <= not w5318 and not w5670;
w5689 <= not w5328 and w5655;
w5690 <= not w5651 and w5689;
w5691 <= not w5652 and not w5655;
w5692 <= not w5690 and not w5691;
w5693 <= w5669 and not w5692;
w5694 <= not w5667 and w5693;
w5695 <= not w5688 and not w5694;
w5696 <= not b(26) and not w5695;
w5697 <= not w5327 and not w5670;
w5698 <= not w5337 and w5650;
w5699 <= not w5646 and w5698;
w5700 <= not w5647 and not w5650;
w5701 <= not w5699 and not w5700;
w5702 <= w5669 and not w5701;
w5703 <= not w5667 and w5702;
w5704 <= not w5697 and not w5703;
w5705 <= not b(25) and not w5704;
w5706 <= not w5336 and not w5670;
w5707 <= not w5346 and w5645;
w5708 <= not w5641 and w5707;
w5709 <= not w5642 and not w5645;
w5710 <= not w5708 and not w5709;
w5711 <= w5669 and not w5710;
w5712 <= not w5667 and w5711;
w5713 <= not w5706 and not w5712;
w5714 <= not b(24) and not w5713;
w5715 <= not w5345 and not w5670;
w5716 <= not w5355 and w5640;
w5717 <= not w5636 and w5716;
w5718 <= not w5637 and not w5640;
w5719 <= not w5717 and not w5718;
w5720 <= w5669 and not w5719;
w5721 <= not w5667 and w5720;
w5722 <= not w5715 and not w5721;
w5723 <= not b(23) and not w5722;
w5724 <= not w5354 and not w5670;
w5725 <= not w5364 and w5635;
w5726 <= not w5631 and w5725;
w5727 <= not w5632 and not w5635;
w5728 <= not w5726 and not w5727;
w5729 <= w5669 and not w5728;
w5730 <= not w5667 and w5729;
w5731 <= not w5724 and not w5730;
w5732 <= not b(22) and not w5731;
w5733 <= not w5363 and not w5670;
w5734 <= not w5373 and w5630;
w5735 <= not w5626 and w5734;
w5736 <= not w5627 and not w5630;
w5737 <= not w5735 and not w5736;
w5738 <= w5669 and not w5737;
w5739 <= not w5667 and w5738;
w5740 <= not w5733 and not w5739;
w5741 <= not b(21) and not w5740;
w5742 <= not w5372 and not w5670;
w5743 <= not w5382 and w5625;
w5744 <= not w5621 and w5743;
w5745 <= not w5622 and not w5625;
w5746 <= not w5744 and not w5745;
w5747 <= w5669 and not w5746;
w5748 <= not w5667 and w5747;
w5749 <= not w5742 and not w5748;
w5750 <= not b(20) and not w5749;
w5751 <= not w5381 and not w5670;
w5752 <= not w5391 and w5620;
w5753 <= not w5616 and w5752;
w5754 <= not w5617 and not w5620;
w5755 <= not w5753 and not w5754;
w5756 <= w5669 and not w5755;
w5757 <= not w5667 and w5756;
w5758 <= not w5751 and not w5757;
w5759 <= not b(19) and not w5758;
w5760 <= not w5390 and not w5670;
w5761 <= not w5400 and w5615;
w5762 <= not w5611 and w5761;
w5763 <= not w5612 and not w5615;
w5764 <= not w5762 and not w5763;
w5765 <= w5669 and not w5764;
w5766 <= not w5667 and w5765;
w5767 <= not w5760 and not w5766;
w5768 <= not b(18) and not w5767;
w5769 <= not w5399 and not w5670;
w5770 <= not w5409 and w5610;
w5771 <= not w5606 and w5770;
w5772 <= not w5607 and not w5610;
w5773 <= not w5771 and not w5772;
w5774 <= w5669 and not w5773;
w5775 <= not w5667 and w5774;
w5776 <= not w5769 and not w5775;
w5777 <= not b(17) and not w5776;
w5778 <= not w5408 and not w5670;
w5779 <= not w5418 and w5605;
w5780 <= not w5601 and w5779;
w5781 <= not w5602 and not w5605;
w5782 <= not w5780 and not w5781;
w5783 <= w5669 and not w5782;
w5784 <= not w5667 and w5783;
w5785 <= not w5778 and not w5784;
w5786 <= not b(16) and not w5785;
w5787 <= not w5417 and not w5670;
w5788 <= not w5427 and w5600;
w5789 <= not w5596 and w5788;
w5790 <= not w5597 and not w5600;
w5791 <= not w5789 and not w5790;
w5792 <= w5669 and not w5791;
w5793 <= not w5667 and w5792;
w5794 <= not w5787 and not w5793;
w5795 <= not b(15) and not w5794;
w5796 <= not w5426 and not w5670;
w5797 <= not w5436 and w5595;
w5798 <= not w5591 and w5797;
w5799 <= not w5592 and not w5595;
w5800 <= not w5798 and not w5799;
w5801 <= w5669 and not w5800;
w5802 <= not w5667 and w5801;
w5803 <= not w5796 and not w5802;
w5804 <= not b(14) and not w5803;
w5805 <= not w5435 and not w5670;
w5806 <= not w5445 and w5590;
w5807 <= not w5586 and w5806;
w5808 <= not w5587 and not w5590;
w5809 <= not w5807 and not w5808;
w5810 <= w5669 and not w5809;
w5811 <= not w5667 and w5810;
w5812 <= not w5805 and not w5811;
w5813 <= not b(13) and not w5812;
w5814 <= not w5444 and not w5670;
w5815 <= not w5454 and w5585;
w5816 <= not w5581 and w5815;
w5817 <= not w5582 and not w5585;
w5818 <= not w5816 and not w5817;
w5819 <= w5669 and not w5818;
w5820 <= not w5667 and w5819;
w5821 <= not w5814 and not w5820;
w5822 <= not b(12) and not w5821;
w5823 <= not w5453 and not w5670;
w5824 <= not w5463 and w5580;
w5825 <= not w5576 and w5824;
w5826 <= not w5577 and not w5580;
w5827 <= not w5825 and not w5826;
w5828 <= w5669 and not w5827;
w5829 <= not w5667 and w5828;
w5830 <= not w5823 and not w5829;
w5831 <= not b(11) and not w5830;
w5832 <= not w5462 and not w5670;
w5833 <= not w5472 and w5575;
w5834 <= not w5571 and w5833;
w5835 <= not w5572 and not w5575;
w5836 <= not w5834 and not w5835;
w5837 <= w5669 and not w5836;
w5838 <= not w5667 and w5837;
w5839 <= not w5832 and not w5838;
w5840 <= not b(10) and not w5839;
w5841 <= not w5471 and not w5670;
w5842 <= not w5481 and w5570;
w5843 <= not w5566 and w5842;
w5844 <= not w5567 and not w5570;
w5845 <= not w5843 and not w5844;
w5846 <= w5669 and not w5845;
w5847 <= not w5667 and w5846;
w5848 <= not w5841 and not w5847;
w5849 <= not b(9) and not w5848;
w5850 <= not w5480 and not w5670;
w5851 <= not w5490 and w5565;
w5852 <= not w5561 and w5851;
w5853 <= not w5562 and not w5565;
w5854 <= not w5852 and not w5853;
w5855 <= w5669 and not w5854;
w5856 <= not w5667 and w5855;
w5857 <= not w5850 and not w5856;
w5858 <= not b(8) and not w5857;
w5859 <= not w5489 and not w5670;
w5860 <= not w5499 and w5560;
w5861 <= not w5556 and w5860;
w5862 <= not w5557 and not w5560;
w5863 <= not w5861 and not w5862;
w5864 <= w5669 and not w5863;
w5865 <= not w5667 and w5864;
w5866 <= not w5859 and not w5865;
w5867 <= not b(7) and not w5866;
w5868 <= not w5498 and not w5670;
w5869 <= not w5508 and w5555;
w5870 <= not w5551 and w5869;
w5871 <= not w5552 and not w5555;
w5872 <= not w5870 and not w5871;
w5873 <= w5669 and not w5872;
w5874 <= not w5667 and w5873;
w5875 <= not w5868 and not w5874;
w5876 <= not b(6) and not w5875;
w5877 <= not w5507 and not w5670;
w5878 <= not w5517 and w5550;
w5879 <= not w5546 and w5878;
w5880 <= not w5547 and not w5550;
w5881 <= not w5879 and not w5880;
w5882 <= w5669 and not w5881;
w5883 <= not w5667 and w5882;
w5884 <= not w5877 and not w5883;
w5885 <= not b(5) and not w5884;
w5886 <= not w5516 and not w5670;
w5887 <= not w5525 and w5545;
w5888 <= not w5541 and w5887;
w5889 <= not w5542 and not w5545;
w5890 <= not w5888 and not w5889;
w5891 <= w5669 and not w5890;
w5892 <= not w5667 and w5891;
w5893 <= not w5886 and not w5892;
w5894 <= not b(4) and not w5893;
w5895 <= not w5524 and not w5670;
w5896 <= not w5536 and w5540;
w5897 <= not w5535 and w5896;
w5898 <= not w5537 and not w5540;
w5899 <= not w5897 and not w5898;
w5900 <= w5669 and not w5899;
w5901 <= not w5667 and w5900;
w5902 <= not w5895 and not w5901;
w5903 <= not b(3) and not w5902;
w5904 <= not w5529 and not w5670;
w5905 <= not w5532 and w5534;
w5906 <= not w5530 and w5905;
w5907 <= w5669 and not w5906;
w5908 <= not w5535 and w5907;
w5909 <= not w5667 and w5908;
w5910 <= not w5904 and not w5909;
w5911 <= not b(2) and not w5910;
w5912 <= b(0) and not b(28);
w5913 <= w116 and w5912;
w5914 <= w166 and w5913;
w5915 <= w151 and w5914;
w5916 <= not w5667 and w5915;
w5917 <= a(36) and not w5916;
w5918 <= w59 and w5534;
w5919 <= w84 and w5918;
w5920 <= w81 and w5919;
w5921 <= not w5667 and w5920;
w5922 <= not w5917 and not w5921;
w5923 <= b(1) and not w5922;
w5924 <= not b(1) and not w5921;
w5925 <= not w5917 and w5924;
w5926 <= not w5923 and not w5925;
w5927 <= not a(35) and b(0);
w5928 <= not w5926 and not w5927;
w5929 <= not b(1) and not w5922;
w5930 <= not w5928 and not w5929;
w5931 <= b(2) and not w5909;
w5932 <= not w5904 and w5931;
w5933 <= not w5911 and not w5932;
w5934 <= not w5930 and w5933;
w5935 <= not w5911 and not w5934;
w5936 <= b(3) and not w5901;
w5937 <= not w5895 and w5936;
w5938 <= not w5903 and not w5937;
w5939 <= not w5935 and w5938;
w5940 <= not w5903 and not w5939;
w5941 <= b(4) and not w5892;
w5942 <= not w5886 and w5941;
w5943 <= not w5894 and not w5942;
w5944 <= not w5940 and w5943;
w5945 <= not w5894 and not w5944;
w5946 <= b(5) and not w5883;
w5947 <= not w5877 and w5946;
w5948 <= not w5885 and not w5947;
w5949 <= not w5945 and w5948;
w5950 <= not w5885 and not w5949;
w5951 <= b(6) and not w5874;
w5952 <= not w5868 and w5951;
w5953 <= not w5876 and not w5952;
w5954 <= not w5950 and w5953;
w5955 <= not w5876 and not w5954;
w5956 <= b(7) and not w5865;
w5957 <= not w5859 and w5956;
w5958 <= not w5867 and not w5957;
w5959 <= not w5955 and w5958;
w5960 <= not w5867 and not w5959;
w5961 <= b(8) and not w5856;
w5962 <= not w5850 and w5961;
w5963 <= not w5858 and not w5962;
w5964 <= not w5960 and w5963;
w5965 <= not w5858 and not w5964;
w5966 <= b(9) and not w5847;
w5967 <= not w5841 and w5966;
w5968 <= not w5849 and not w5967;
w5969 <= not w5965 and w5968;
w5970 <= not w5849 and not w5969;
w5971 <= b(10) and not w5838;
w5972 <= not w5832 and w5971;
w5973 <= not w5840 and not w5972;
w5974 <= not w5970 and w5973;
w5975 <= not w5840 and not w5974;
w5976 <= b(11) and not w5829;
w5977 <= not w5823 and w5976;
w5978 <= not w5831 and not w5977;
w5979 <= not w5975 and w5978;
w5980 <= not w5831 and not w5979;
w5981 <= b(12) and not w5820;
w5982 <= not w5814 and w5981;
w5983 <= not w5822 and not w5982;
w5984 <= not w5980 and w5983;
w5985 <= not w5822 and not w5984;
w5986 <= b(13) and not w5811;
w5987 <= not w5805 and w5986;
w5988 <= not w5813 and not w5987;
w5989 <= not w5985 and w5988;
w5990 <= not w5813 and not w5989;
w5991 <= b(14) and not w5802;
w5992 <= not w5796 and w5991;
w5993 <= not w5804 and not w5992;
w5994 <= not w5990 and w5993;
w5995 <= not w5804 and not w5994;
w5996 <= b(15) and not w5793;
w5997 <= not w5787 and w5996;
w5998 <= not w5795 and not w5997;
w5999 <= not w5995 and w5998;
w6000 <= not w5795 and not w5999;
w6001 <= b(16) and not w5784;
w6002 <= not w5778 and w6001;
w6003 <= not w5786 and not w6002;
w6004 <= not w6000 and w6003;
w6005 <= not w5786 and not w6004;
w6006 <= b(17) and not w5775;
w6007 <= not w5769 and w6006;
w6008 <= not w5777 and not w6007;
w6009 <= not w6005 and w6008;
w6010 <= not w5777 and not w6009;
w6011 <= b(18) and not w5766;
w6012 <= not w5760 and w6011;
w6013 <= not w5768 and not w6012;
w6014 <= not w6010 and w6013;
w6015 <= not w5768 and not w6014;
w6016 <= b(19) and not w5757;
w6017 <= not w5751 and w6016;
w6018 <= not w5759 and not w6017;
w6019 <= not w6015 and w6018;
w6020 <= not w5759 and not w6019;
w6021 <= b(20) and not w5748;
w6022 <= not w5742 and w6021;
w6023 <= not w5750 and not w6022;
w6024 <= not w6020 and w6023;
w6025 <= not w5750 and not w6024;
w6026 <= b(21) and not w5739;
w6027 <= not w5733 and w6026;
w6028 <= not w5741 and not w6027;
w6029 <= not w6025 and w6028;
w6030 <= not w5741 and not w6029;
w6031 <= b(22) and not w5730;
w6032 <= not w5724 and w6031;
w6033 <= not w5732 and not w6032;
w6034 <= not w6030 and w6033;
w6035 <= not w5732 and not w6034;
w6036 <= b(23) and not w5721;
w6037 <= not w5715 and w6036;
w6038 <= not w5723 and not w6037;
w6039 <= not w6035 and w6038;
w6040 <= not w5723 and not w6039;
w6041 <= b(24) and not w5712;
w6042 <= not w5706 and w6041;
w6043 <= not w5714 and not w6042;
w6044 <= not w6040 and w6043;
w6045 <= not w5714 and not w6044;
w6046 <= b(25) and not w5703;
w6047 <= not w5697 and w6046;
w6048 <= not w5705 and not w6047;
w6049 <= not w6045 and w6048;
w6050 <= not w5705 and not w6049;
w6051 <= b(26) and not w5694;
w6052 <= not w5688 and w6051;
w6053 <= not w5696 and not w6052;
w6054 <= not w6050 and w6053;
w6055 <= not w5696 and not w6054;
w6056 <= b(27) and not w5677;
w6057 <= not w5671 and w6056;
w6058 <= not w5687 and not w6057;
w6059 <= not w6055 and w6058;
w6060 <= not w5687 and not w6059;
w6061 <= b(28) and not w5679;
w6062 <= not w5684 and w6061;
w6063 <= not w5686 and not w6062;
w6064 <= not w6060 and w6063;
w6065 <= not w5686 and not w6064;
w6066 <= w331 and w341;
w6067 <= w338 and w6066;
w6068 <= not w6065 and w6067;
w6069 <= not w5678 and not w6068;
w6070 <= not w5696 and w6058;
w6071 <= not w6054 and w6070;
w6072 <= not w6055 and not w6058;
w6073 <= not w6071 and not w6072;
w6074 <= w6067 and not w6073;
w6075 <= not w6065 and w6074;
w6076 <= not w6069 and not w6075;
w6077 <= not b(28) and not w6076;
w6078 <= not w5695 and not w6068;
w6079 <= not w5705 and w6053;
w6080 <= not w6049 and w6079;
w6081 <= not w6050 and not w6053;
w6082 <= not w6080 and not w6081;
w6083 <= w6067 and not w6082;
w6084 <= not w6065 and w6083;
w6085 <= not w6078 and not w6084;
w6086 <= not b(27) and not w6085;
w6087 <= not w5704 and not w6068;
w6088 <= not w5714 and w6048;
w6089 <= not w6044 and w6088;
w6090 <= not w6045 and not w6048;
w6091 <= not w6089 and not w6090;
w6092 <= w6067 and not w6091;
w6093 <= not w6065 and w6092;
w6094 <= not w6087 and not w6093;
w6095 <= not b(26) and not w6094;
w6096 <= not w5713 and not w6068;
w6097 <= not w5723 and w6043;
w6098 <= not w6039 and w6097;
w6099 <= not w6040 and not w6043;
w6100 <= not w6098 and not w6099;
w6101 <= w6067 and not w6100;
w6102 <= not w6065 and w6101;
w6103 <= not w6096 and not w6102;
w6104 <= not b(25) and not w6103;
w6105 <= not w5722 and not w6068;
w6106 <= not w5732 and w6038;
w6107 <= not w6034 and w6106;
w6108 <= not w6035 and not w6038;
w6109 <= not w6107 and not w6108;
w6110 <= w6067 and not w6109;
w6111 <= not w6065 and w6110;
w6112 <= not w6105 and not w6111;
w6113 <= not b(24) and not w6112;
w6114 <= not w5731 and not w6068;
w6115 <= not w5741 and w6033;
w6116 <= not w6029 and w6115;
w6117 <= not w6030 and not w6033;
w6118 <= not w6116 and not w6117;
w6119 <= w6067 and not w6118;
w6120 <= not w6065 and w6119;
w6121 <= not w6114 and not w6120;
w6122 <= not b(23) and not w6121;
w6123 <= not w5740 and not w6068;
w6124 <= not w5750 and w6028;
w6125 <= not w6024 and w6124;
w6126 <= not w6025 and not w6028;
w6127 <= not w6125 and not w6126;
w6128 <= w6067 and not w6127;
w6129 <= not w6065 and w6128;
w6130 <= not w6123 and not w6129;
w6131 <= not b(22) and not w6130;
w6132 <= not w5749 and not w6068;
w6133 <= not w5759 and w6023;
w6134 <= not w6019 and w6133;
w6135 <= not w6020 and not w6023;
w6136 <= not w6134 and not w6135;
w6137 <= w6067 and not w6136;
w6138 <= not w6065 and w6137;
w6139 <= not w6132 and not w6138;
w6140 <= not b(21) and not w6139;
w6141 <= not w5758 and not w6068;
w6142 <= not w5768 and w6018;
w6143 <= not w6014 and w6142;
w6144 <= not w6015 and not w6018;
w6145 <= not w6143 and not w6144;
w6146 <= w6067 and not w6145;
w6147 <= not w6065 and w6146;
w6148 <= not w6141 and not w6147;
w6149 <= not b(20) and not w6148;
w6150 <= not w5767 and not w6068;
w6151 <= not w5777 and w6013;
w6152 <= not w6009 and w6151;
w6153 <= not w6010 and not w6013;
w6154 <= not w6152 and not w6153;
w6155 <= w6067 and not w6154;
w6156 <= not w6065 and w6155;
w6157 <= not w6150 and not w6156;
w6158 <= not b(19) and not w6157;
w6159 <= not w5776 and not w6068;
w6160 <= not w5786 and w6008;
w6161 <= not w6004 and w6160;
w6162 <= not w6005 and not w6008;
w6163 <= not w6161 and not w6162;
w6164 <= w6067 and not w6163;
w6165 <= not w6065 and w6164;
w6166 <= not w6159 and not w6165;
w6167 <= not b(18) and not w6166;
w6168 <= not w5785 and not w6068;
w6169 <= not w5795 and w6003;
w6170 <= not w5999 and w6169;
w6171 <= not w6000 and not w6003;
w6172 <= not w6170 and not w6171;
w6173 <= w6067 and not w6172;
w6174 <= not w6065 and w6173;
w6175 <= not w6168 and not w6174;
w6176 <= not b(17) and not w6175;
w6177 <= not w5794 and not w6068;
w6178 <= not w5804 and w5998;
w6179 <= not w5994 and w6178;
w6180 <= not w5995 and not w5998;
w6181 <= not w6179 and not w6180;
w6182 <= w6067 and not w6181;
w6183 <= not w6065 and w6182;
w6184 <= not w6177 and not w6183;
w6185 <= not b(16) and not w6184;
w6186 <= not w5803 and not w6068;
w6187 <= not w5813 and w5993;
w6188 <= not w5989 and w6187;
w6189 <= not w5990 and not w5993;
w6190 <= not w6188 and not w6189;
w6191 <= w6067 and not w6190;
w6192 <= not w6065 and w6191;
w6193 <= not w6186 and not w6192;
w6194 <= not b(15) and not w6193;
w6195 <= not w5812 and not w6068;
w6196 <= not w5822 and w5988;
w6197 <= not w5984 and w6196;
w6198 <= not w5985 and not w5988;
w6199 <= not w6197 and not w6198;
w6200 <= w6067 and not w6199;
w6201 <= not w6065 and w6200;
w6202 <= not w6195 and not w6201;
w6203 <= not b(14) and not w6202;
w6204 <= not w5821 and not w6068;
w6205 <= not w5831 and w5983;
w6206 <= not w5979 and w6205;
w6207 <= not w5980 and not w5983;
w6208 <= not w6206 and not w6207;
w6209 <= w6067 and not w6208;
w6210 <= not w6065 and w6209;
w6211 <= not w6204 and not w6210;
w6212 <= not b(13) and not w6211;
w6213 <= not w5830 and not w6068;
w6214 <= not w5840 and w5978;
w6215 <= not w5974 and w6214;
w6216 <= not w5975 and not w5978;
w6217 <= not w6215 and not w6216;
w6218 <= w6067 and not w6217;
w6219 <= not w6065 and w6218;
w6220 <= not w6213 and not w6219;
w6221 <= not b(12) and not w6220;
w6222 <= not w5839 and not w6068;
w6223 <= not w5849 and w5973;
w6224 <= not w5969 and w6223;
w6225 <= not w5970 and not w5973;
w6226 <= not w6224 and not w6225;
w6227 <= w6067 and not w6226;
w6228 <= not w6065 and w6227;
w6229 <= not w6222 and not w6228;
w6230 <= not b(11) and not w6229;
w6231 <= not w5848 and not w6068;
w6232 <= not w5858 and w5968;
w6233 <= not w5964 and w6232;
w6234 <= not w5965 and not w5968;
w6235 <= not w6233 and not w6234;
w6236 <= w6067 and not w6235;
w6237 <= not w6065 and w6236;
w6238 <= not w6231 and not w6237;
w6239 <= not b(10) and not w6238;
w6240 <= not w5857 and not w6068;
w6241 <= not w5867 and w5963;
w6242 <= not w5959 and w6241;
w6243 <= not w5960 and not w5963;
w6244 <= not w6242 and not w6243;
w6245 <= w6067 and not w6244;
w6246 <= not w6065 and w6245;
w6247 <= not w6240 and not w6246;
w6248 <= not b(9) and not w6247;
w6249 <= not w5866 and not w6068;
w6250 <= not w5876 and w5958;
w6251 <= not w5954 and w6250;
w6252 <= not w5955 and not w5958;
w6253 <= not w6251 and not w6252;
w6254 <= w6067 and not w6253;
w6255 <= not w6065 and w6254;
w6256 <= not w6249 and not w6255;
w6257 <= not b(8) and not w6256;
w6258 <= not w5875 and not w6068;
w6259 <= not w5885 and w5953;
w6260 <= not w5949 and w6259;
w6261 <= not w5950 and not w5953;
w6262 <= not w6260 and not w6261;
w6263 <= w6067 and not w6262;
w6264 <= not w6065 and w6263;
w6265 <= not w6258 and not w6264;
w6266 <= not b(7) and not w6265;
w6267 <= not w5884 and not w6068;
w6268 <= not w5894 and w5948;
w6269 <= not w5944 and w6268;
w6270 <= not w5945 and not w5948;
w6271 <= not w6269 and not w6270;
w6272 <= w6067 and not w6271;
w6273 <= not w6065 and w6272;
w6274 <= not w6267 and not w6273;
w6275 <= not b(6) and not w6274;
w6276 <= not w5893 and not w6068;
w6277 <= not w5903 and w5943;
w6278 <= not w5939 and w6277;
w6279 <= not w5940 and not w5943;
w6280 <= not w6278 and not w6279;
w6281 <= w6067 and not w6280;
w6282 <= not w6065 and w6281;
w6283 <= not w6276 and not w6282;
w6284 <= not b(5) and not w6283;
w6285 <= not w5902 and not w6068;
w6286 <= not w5911 and w5938;
w6287 <= not w5934 and w6286;
w6288 <= not w5935 and not w5938;
w6289 <= not w6287 and not w6288;
w6290 <= w6067 and not w6289;
w6291 <= not w6065 and w6290;
w6292 <= not w6285 and not w6291;
w6293 <= not b(4) and not w6292;
w6294 <= not w5910 and not w6068;
w6295 <= not w5929 and w5933;
w6296 <= not w5928 and w6295;
w6297 <= not w5930 and not w5933;
w6298 <= not w6296 and not w6297;
w6299 <= w6067 and not w6298;
w6300 <= not w6065 and w6299;
w6301 <= not w6294 and not w6300;
w6302 <= not b(3) and not w6301;
w6303 <= not w5922 and not w6068;
w6304 <= not w5925 and w5927;
w6305 <= not w5923 and w6304;
w6306 <= w6067 and not w6305;
w6307 <= not w5928 and w6306;
w6308 <= not w6065 and w6307;
w6309 <= not w6303 and not w6308;
w6310 <= not b(2) and not w6309;
w6311 <= b(0) and not b(29);
w6312 <= w58 and w6311;
w6313 <= w56 and w6312;
w6314 <= w46 and w6313;
w6315 <= w31 and w6314;
w6316 <= not w6065 and w6315;
w6317 <= a(35) and not w6316;
w6318 <= w116 and w5927;
w6319 <= w166 and w6318;
w6320 <= w151 and w6319;
w6321 <= not w6065 and w6320;
w6322 <= not w6317 and not w6321;
w6323 <= b(1) and not w6322;
w6324 <= not b(1) and not w6321;
w6325 <= not w6317 and w6324;
w6326 <= not w6323 and not w6325;
w6327 <= not a(34) and b(0);
w6328 <= not w6326 and not w6327;
w6329 <= not b(1) and not w6322;
w6330 <= not w6328 and not w6329;
w6331 <= b(2) and not w6308;
w6332 <= not w6303 and w6331;
w6333 <= not w6310 and not w6332;
w6334 <= not w6330 and w6333;
w6335 <= not w6310 and not w6334;
w6336 <= b(3) and not w6300;
w6337 <= not w6294 and w6336;
w6338 <= not w6302 and not w6337;
w6339 <= not w6335 and w6338;
w6340 <= not w6302 and not w6339;
w6341 <= b(4) and not w6291;
w6342 <= not w6285 and w6341;
w6343 <= not w6293 and not w6342;
w6344 <= not w6340 and w6343;
w6345 <= not w6293 and not w6344;
w6346 <= b(5) and not w6282;
w6347 <= not w6276 and w6346;
w6348 <= not w6284 and not w6347;
w6349 <= not w6345 and w6348;
w6350 <= not w6284 and not w6349;
w6351 <= b(6) and not w6273;
w6352 <= not w6267 and w6351;
w6353 <= not w6275 and not w6352;
w6354 <= not w6350 and w6353;
w6355 <= not w6275 and not w6354;
w6356 <= b(7) and not w6264;
w6357 <= not w6258 and w6356;
w6358 <= not w6266 and not w6357;
w6359 <= not w6355 and w6358;
w6360 <= not w6266 and not w6359;
w6361 <= b(8) and not w6255;
w6362 <= not w6249 and w6361;
w6363 <= not w6257 and not w6362;
w6364 <= not w6360 and w6363;
w6365 <= not w6257 and not w6364;
w6366 <= b(9) and not w6246;
w6367 <= not w6240 and w6366;
w6368 <= not w6248 and not w6367;
w6369 <= not w6365 and w6368;
w6370 <= not w6248 and not w6369;
w6371 <= b(10) and not w6237;
w6372 <= not w6231 and w6371;
w6373 <= not w6239 and not w6372;
w6374 <= not w6370 and w6373;
w6375 <= not w6239 and not w6374;
w6376 <= b(11) and not w6228;
w6377 <= not w6222 and w6376;
w6378 <= not w6230 and not w6377;
w6379 <= not w6375 and w6378;
w6380 <= not w6230 and not w6379;
w6381 <= b(12) and not w6219;
w6382 <= not w6213 and w6381;
w6383 <= not w6221 and not w6382;
w6384 <= not w6380 and w6383;
w6385 <= not w6221 and not w6384;
w6386 <= b(13) and not w6210;
w6387 <= not w6204 and w6386;
w6388 <= not w6212 and not w6387;
w6389 <= not w6385 and w6388;
w6390 <= not w6212 and not w6389;
w6391 <= b(14) and not w6201;
w6392 <= not w6195 and w6391;
w6393 <= not w6203 and not w6392;
w6394 <= not w6390 and w6393;
w6395 <= not w6203 and not w6394;
w6396 <= b(15) and not w6192;
w6397 <= not w6186 and w6396;
w6398 <= not w6194 and not w6397;
w6399 <= not w6395 and w6398;
w6400 <= not w6194 and not w6399;
w6401 <= b(16) and not w6183;
w6402 <= not w6177 and w6401;
w6403 <= not w6185 and not w6402;
w6404 <= not w6400 and w6403;
w6405 <= not w6185 and not w6404;
w6406 <= b(17) and not w6174;
w6407 <= not w6168 and w6406;
w6408 <= not w6176 and not w6407;
w6409 <= not w6405 and w6408;
w6410 <= not w6176 and not w6409;
w6411 <= b(18) and not w6165;
w6412 <= not w6159 and w6411;
w6413 <= not w6167 and not w6412;
w6414 <= not w6410 and w6413;
w6415 <= not w6167 and not w6414;
w6416 <= b(19) and not w6156;
w6417 <= not w6150 and w6416;
w6418 <= not w6158 and not w6417;
w6419 <= not w6415 and w6418;
w6420 <= not w6158 and not w6419;
w6421 <= b(20) and not w6147;
w6422 <= not w6141 and w6421;
w6423 <= not w6149 and not w6422;
w6424 <= not w6420 and w6423;
w6425 <= not w6149 and not w6424;
w6426 <= b(21) and not w6138;
w6427 <= not w6132 and w6426;
w6428 <= not w6140 and not w6427;
w6429 <= not w6425 and w6428;
w6430 <= not w6140 and not w6429;
w6431 <= b(22) and not w6129;
w6432 <= not w6123 and w6431;
w6433 <= not w6131 and not w6432;
w6434 <= not w6430 and w6433;
w6435 <= not w6131 and not w6434;
w6436 <= b(23) and not w6120;
w6437 <= not w6114 and w6436;
w6438 <= not w6122 and not w6437;
w6439 <= not w6435 and w6438;
w6440 <= not w6122 and not w6439;
w6441 <= b(24) and not w6111;
w6442 <= not w6105 and w6441;
w6443 <= not w6113 and not w6442;
w6444 <= not w6440 and w6443;
w6445 <= not w6113 and not w6444;
w6446 <= b(25) and not w6102;
w6447 <= not w6096 and w6446;
w6448 <= not w6104 and not w6447;
w6449 <= not w6445 and w6448;
w6450 <= not w6104 and not w6449;
w6451 <= b(26) and not w6093;
w6452 <= not w6087 and w6451;
w6453 <= not w6095 and not w6452;
w6454 <= not w6450 and w6453;
w6455 <= not w6095 and not w6454;
w6456 <= b(27) and not w6084;
w6457 <= not w6078 and w6456;
w6458 <= not w6086 and not w6457;
w6459 <= not w6455 and w6458;
w6460 <= not w6086 and not w6459;
w6461 <= b(28) and not w6075;
w6462 <= not w6069 and w6461;
w6463 <= not w6077 and not w6462;
w6464 <= not w6460 and w6463;
w6465 <= not w6077 and not w6464;
w6466 <= not w5685 and not w6068;
w6467 <= not w5687 and w6063;
w6468 <= not w6059 and w6467;
w6469 <= not w6060 and not w6063;
w6470 <= not w6468 and not w6469;
w6471 <= w6068 and not w6470;
w6472 <= not w6466 and not w6471;
w6473 <= not b(29) and not w6472;
w6474 <= b(29) and not w6466;
w6475 <= not w6471 and w6474;
w6476 <= w56 and w58;
w6477 <= w46 and w6476;
w6478 <= w31 and w6477;
w6479 <= not w6475 and w6478;
w6480 <= not w6473 and w6479;
w6481 <= not w6465 and w6480;
w6482 <= w6067 and not w6472;
w6483 <= not w6481 and not w6482;
w6484 <= not w6086 and w6463;
w6485 <= not w6459 and w6484;
w6486 <= not w6460 and not w6463;
w6487 <= not w6485 and not w6486;
w6488 <= not w6483 and not w6487;
w6489 <= not w6076 and not w6482;
w6490 <= not w6481 and w6489;
w6491 <= not w6488 and not w6490;
w6492 <= not w6077 and not w6475;
w6493 <= not w6473 and w6492;
w6494 <= not w6464 and w6493;
w6495 <= not w6473 and not w6475;
w6496 <= not w6465 and not w6495;
w6497 <= not w6494 and not w6496;
w6498 <= not w6483 and not w6497;
w6499 <= not w6472 and not w6482;
w6500 <= not w6481 and w6499;
w6501 <= not w6498 and not w6500;
w6502 <= not b(30) and not w6501;
w6503 <= not b(29) and not w6491;
w6504 <= not w6095 and w6458;
w6505 <= not w6454 and w6504;
w6506 <= not w6455 and not w6458;
w6507 <= not w6505 and not w6506;
w6508 <= not w6483 and not w6507;
w6509 <= not w6085 and not w6482;
w6510 <= not w6481 and w6509;
w6511 <= not w6508 and not w6510;
w6512 <= not b(28) and not w6511;
w6513 <= not w6104 and w6453;
w6514 <= not w6449 and w6513;
w6515 <= not w6450 and not w6453;
w6516 <= not w6514 and not w6515;
w6517 <= not w6483 and not w6516;
w6518 <= not w6094 and not w6482;
w6519 <= not w6481 and w6518;
w6520 <= not w6517 and not w6519;
w6521 <= not b(27) and not w6520;
w6522 <= not w6113 and w6448;
w6523 <= not w6444 and w6522;
w6524 <= not w6445 and not w6448;
w6525 <= not w6523 and not w6524;
w6526 <= not w6483 and not w6525;
w6527 <= not w6103 and not w6482;
w6528 <= not w6481 and w6527;
w6529 <= not w6526 and not w6528;
w6530 <= not b(26) and not w6529;
w6531 <= not w6122 and w6443;
w6532 <= not w6439 and w6531;
w6533 <= not w6440 and not w6443;
w6534 <= not w6532 and not w6533;
w6535 <= not w6483 and not w6534;
w6536 <= not w6112 and not w6482;
w6537 <= not w6481 and w6536;
w6538 <= not w6535 and not w6537;
w6539 <= not b(25) and not w6538;
w6540 <= not w6131 and w6438;
w6541 <= not w6434 and w6540;
w6542 <= not w6435 and not w6438;
w6543 <= not w6541 and not w6542;
w6544 <= not w6483 and not w6543;
w6545 <= not w6121 and not w6482;
w6546 <= not w6481 and w6545;
w6547 <= not w6544 and not w6546;
w6548 <= not b(24) and not w6547;
w6549 <= not w6140 and w6433;
w6550 <= not w6429 and w6549;
w6551 <= not w6430 and not w6433;
w6552 <= not w6550 and not w6551;
w6553 <= not w6483 and not w6552;
w6554 <= not w6130 and not w6482;
w6555 <= not w6481 and w6554;
w6556 <= not w6553 and not w6555;
w6557 <= not b(23) and not w6556;
w6558 <= not w6149 and w6428;
w6559 <= not w6424 and w6558;
w6560 <= not w6425 and not w6428;
w6561 <= not w6559 and not w6560;
w6562 <= not w6483 and not w6561;
w6563 <= not w6139 and not w6482;
w6564 <= not w6481 and w6563;
w6565 <= not w6562 and not w6564;
w6566 <= not b(22) and not w6565;
w6567 <= not w6158 and w6423;
w6568 <= not w6419 and w6567;
w6569 <= not w6420 and not w6423;
w6570 <= not w6568 and not w6569;
w6571 <= not w6483 and not w6570;
w6572 <= not w6148 and not w6482;
w6573 <= not w6481 and w6572;
w6574 <= not w6571 and not w6573;
w6575 <= not b(21) and not w6574;
w6576 <= not w6167 and w6418;
w6577 <= not w6414 and w6576;
w6578 <= not w6415 and not w6418;
w6579 <= not w6577 and not w6578;
w6580 <= not w6483 and not w6579;
w6581 <= not w6157 and not w6482;
w6582 <= not w6481 and w6581;
w6583 <= not w6580 and not w6582;
w6584 <= not b(20) and not w6583;
w6585 <= not w6176 and w6413;
w6586 <= not w6409 and w6585;
w6587 <= not w6410 and not w6413;
w6588 <= not w6586 and not w6587;
w6589 <= not w6483 and not w6588;
w6590 <= not w6166 and not w6482;
w6591 <= not w6481 and w6590;
w6592 <= not w6589 and not w6591;
w6593 <= not b(19) and not w6592;
w6594 <= not w6185 and w6408;
w6595 <= not w6404 and w6594;
w6596 <= not w6405 and not w6408;
w6597 <= not w6595 and not w6596;
w6598 <= not w6483 and not w6597;
w6599 <= not w6175 and not w6482;
w6600 <= not w6481 and w6599;
w6601 <= not w6598 and not w6600;
w6602 <= not b(18) and not w6601;
w6603 <= not w6194 and w6403;
w6604 <= not w6399 and w6603;
w6605 <= not w6400 and not w6403;
w6606 <= not w6604 and not w6605;
w6607 <= not w6483 and not w6606;
w6608 <= not w6184 and not w6482;
w6609 <= not w6481 and w6608;
w6610 <= not w6607 and not w6609;
w6611 <= not b(17) and not w6610;
w6612 <= not w6203 and w6398;
w6613 <= not w6394 and w6612;
w6614 <= not w6395 and not w6398;
w6615 <= not w6613 and not w6614;
w6616 <= not w6483 and not w6615;
w6617 <= not w6193 and not w6482;
w6618 <= not w6481 and w6617;
w6619 <= not w6616 and not w6618;
w6620 <= not b(16) and not w6619;
w6621 <= not w6212 and w6393;
w6622 <= not w6389 and w6621;
w6623 <= not w6390 and not w6393;
w6624 <= not w6622 and not w6623;
w6625 <= not w6483 and not w6624;
w6626 <= not w6202 and not w6482;
w6627 <= not w6481 and w6626;
w6628 <= not w6625 and not w6627;
w6629 <= not b(15) and not w6628;
w6630 <= not w6221 and w6388;
w6631 <= not w6384 and w6630;
w6632 <= not w6385 and not w6388;
w6633 <= not w6631 and not w6632;
w6634 <= not w6483 and not w6633;
w6635 <= not w6211 and not w6482;
w6636 <= not w6481 and w6635;
w6637 <= not w6634 and not w6636;
w6638 <= not b(14) and not w6637;
w6639 <= not w6230 and w6383;
w6640 <= not w6379 and w6639;
w6641 <= not w6380 and not w6383;
w6642 <= not w6640 and not w6641;
w6643 <= not w6483 and not w6642;
w6644 <= not w6220 and not w6482;
w6645 <= not w6481 and w6644;
w6646 <= not w6643 and not w6645;
w6647 <= not b(13) and not w6646;
w6648 <= not w6239 and w6378;
w6649 <= not w6374 and w6648;
w6650 <= not w6375 and not w6378;
w6651 <= not w6649 and not w6650;
w6652 <= not w6483 and not w6651;
w6653 <= not w6229 and not w6482;
w6654 <= not w6481 and w6653;
w6655 <= not w6652 and not w6654;
w6656 <= not b(12) and not w6655;
w6657 <= not w6248 and w6373;
w6658 <= not w6369 and w6657;
w6659 <= not w6370 and not w6373;
w6660 <= not w6658 and not w6659;
w6661 <= not w6483 and not w6660;
w6662 <= not w6238 and not w6482;
w6663 <= not w6481 and w6662;
w6664 <= not w6661 and not w6663;
w6665 <= not b(11) and not w6664;
w6666 <= not w6257 and w6368;
w6667 <= not w6364 and w6666;
w6668 <= not w6365 and not w6368;
w6669 <= not w6667 and not w6668;
w6670 <= not w6483 and not w6669;
w6671 <= not w6247 and not w6482;
w6672 <= not w6481 and w6671;
w6673 <= not w6670 and not w6672;
w6674 <= not b(10) and not w6673;
w6675 <= not w6266 and w6363;
w6676 <= not w6359 and w6675;
w6677 <= not w6360 and not w6363;
w6678 <= not w6676 and not w6677;
w6679 <= not w6483 and not w6678;
w6680 <= not w6256 and not w6482;
w6681 <= not w6481 and w6680;
w6682 <= not w6679 and not w6681;
w6683 <= not b(9) and not w6682;
w6684 <= not w6275 and w6358;
w6685 <= not w6354 and w6684;
w6686 <= not w6355 and not w6358;
w6687 <= not w6685 and not w6686;
w6688 <= not w6483 and not w6687;
w6689 <= not w6265 and not w6482;
w6690 <= not w6481 and w6689;
w6691 <= not w6688 and not w6690;
w6692 <= not b(8) and not w6691;
w6693 <= not w6284 and w6353;
w6694 <= not w6349 and w6693;
w6695 <= not w6350 and not w6353;
w6696 <= not w6694 and not w6695;
w6697 <= not w6483 and not w6696;
w6698 <= not w6274 and not w6482;
w6699 <= not w6481 and w6698;
w6700 <= not w6697 and not w6699;
w6701 <= not b(7) and not w6700;
w6702 <= not w6293 and w6348;
w6703 <= not w6344 and w6702;
w6704 <= not w6345 and not w6348;
w6705 <= not w6703 and not w6704;
w6706 <= not w6483 and not w6705;
w6707 <= not w6283 and not w6482;
w6708 <= not w6481 and w6707;
w6709 <= not w6706 and not w6708;
w6710 <= not b(6) and not w6709;
w6711 <= not w6302 and w6343;
w6712 <= not w6339 and w6711;
w6713 <= not w6340 and not w6343;
w6714 <= not w6712 and not w6713;
w6715 <= not w6483 and not w6714;
w6716 <= not w6292 and not w6482;
w6717 <= not w6481 and w6716;
w6718 <= not w6715 and not w6717;
w6719 <= not b(5) and not w6718;
w6720 <= not w6310 and w6338;
w6721 <= not w6334 and w6720;
w6722 <= not w6335 and not w6338;
w6723 <= not w6721 and not w6722;
w6724 <= not w6483 and not w6723;
w6725 <= not w6301 and not w6482;
w6726 <= not w6481 and w6725;
w6727 <= not w6724 and not w6726;
w6728 <= not b(4) and not w6727;
w6729 <= not w6329 and w6333;
w6730 <= not w6328 and w6729;
w6731 <= not w6330 and not w6333;
w6732 <= not w6730 and not w6731;
w6733 <= not w6483 and not w6732;
w6734 <= not w6309 and not w6482;
w6735 <= not w6481 and w6734;
w6736 <= not w6733 and not w6735;
w6737 <= not b(3) and not w6736;
w6738 <= not w6325 and w6327;
w6739 <= not w6323 and w6738;
w6740 <= not w6328 and not w6739;
w6741 <= not w6483 and w6740;
w6742 <= not w6322 and not w6482;
w6743 <= not w6481 and w6742;
w6744 <= not w6741 and not w6743;
w6745 <= not b(2) and not w6744;
w6746 <= b(0) and not w6483;
w6747 <= a(34) and not w6746;
w6748 <= w6327 and not w6483;
w6749 <= not w6747 and not w6748;
w6750 <= b(1) and not w6749;
w6751 <= not b(1) and not w6748;
w6752 <= not w6747 and w6751;
w6753 <= not w6750 and not w6752;
w6754 <= not a(33) and b(0);
w6755 <= not w6753 and not w6754;
w6756 <= not b(1) and not w6749;
w6757 <= not w6755 and not w6756;
w6758 <= b(2) and not w6743;
w6759 <= not w6741 and w6758;
w6760 <= not w6745 and not w6759;
w6761 <= not w6757 and w6760;
w6762 <= not w6745 and not w6761;
w6763 <= b(3) and not w6735;
w6764 <= not w6733 and w6763;
w6765 <= not w6737 and not w6764;
w6766 <= not w6762 and w6765;
w6767 <= not w6737 and not w6766;
w6768 <= b(4) and not w6726;
w6769 <= not w6724 and w6768;
w6770 <= not w6728 and not w6769;
w6771 <= not w6767 and w6770;
w6772 <= not w6728 and not w6771;
w6773 <= b(5) and not w6717;
w6774 <= not w6715 and w6773;
w6775 <= not w6719 and not w6774;
w6776 <= not w6772 and w6775;
w6777 <= not w6719 and not w6776;
w6778 <= b(6) and not w6708;
w6779 <= not w6706 and w6778;
w6780 <= not w6710 and not w6779;
w6781 <= not w6777 and w6780;
w6782 <= not w6710 and not w6781;
w6783 <= b(7) and not w6699;
w6784 <= not w6697 and w6783;
w6785 <= not w6701 and not w6784;
w6786 <= not w6782 and w6785;
w6787 <= not w6701 and not w6786;
w6788 <= b(8) and not w6690;
w6789 <= not w6688 and w6788;
w6790 <= not w6692 and not w6789;
w6791 <= not w6787 and w6790;
w6792 <= not w6692 and not w6791;
w6793 <= b(9) and not w6681;
w6794 <= not w6679 and w6793;
w6795 <= not w6683 and not w6794;
w6796 <= not w6792 and w6795;
w6797 <= not w6683 and not w6796;
w6798 <= b(10) and not w6672;
w6799 <= not w6670 and w6798;
w6800 <= not w6674 and not w6799;
w6801 <= not w6797 and w6800;
w6802 <= not w6674 and not w6801;
w6803 <= b(11) and not w6663;
w6804 <= not w6661 and w6803;
w6805 <= not w6665 and not w6804;
w6806 <= not w6802 and w6805;
w6807 <= not w6665 and not w6806;
w6808 <= b(12) and not w6654;
w6809 <= not w6652 and w6808;
w6810 <= not w6656 and not w6809;
w6811 <= not w6807 and w6810;
w6812 <= not w6656 and not w6811;
w6813 <= b(13) and not w6645;
w6814 <= not w6643 and w6813;
w6815 <= not w6647 and not w6814;
w6816 <= not w6812 and w6815;
w6817 <= not w6647 and not w6816;
w6818 <= b(14) and not w6636;
w6819 <= not w6634 and w6818;
w6820 <= not w6638 and not w6819;
w6821 <= not w6817 and w6820;
w6822 <= not w6638 and not w6821;
w6823 <= b(15) and not w6627;
w6824 <= not w6625 and w6823;
w6825 <= not w6629 and not w6824;
w6826 <= not w6822 and w6825;
w6827 <= not w6629 and not w6826;
w6828 <= b(16) and not w6618;
w6829 <= not w6616 and w6828;
w6830 <= not w6620 and not w6829;
w6831 <= not w6827 and w6830;
w6832 <= not w6620 and not w6831;
w6833 <= b(17) and not w6609;
w6834 <= not w6607 and w6833;
w6835 <= not w6611 and not w6834;
w6836 <= not w6832 and w6835;
w6837 <= not w6611 and not w6836;
w6838 <= b(18) and not w6600;
w6839 <= not w6598 and w6838;
w6840 <= not w6602 and not w6839;
w6841 <= not w6837 and w6840;
w6842 <= not w6602 and not w6841;
w6843 <= b(19) and not w6591;
w6844 <= not w6589 and w6843;
w6845 <= not w6593 and not w6844;
w6846 <= not w6842 and w6845;
w6847 <= not w6593 and not w6846;
w6848 <= b(20) and not w6582;
w6849 <= not w6580 and w6848;
w6850 <= not w6584 and not w6849;
w6851 <= not w6847 and w6850;
w6852 <= not w6584 and not w6851;
w6853 <= b(21) and not w6573;
w6854 <= not w6571 and w6853;
w6855 <= not w6575 and not w6854;
w6856 <= not w6852 and w6855;
w6857 <= not w6575 and not w6856;
w6858 <= b(22) and not w6564;
w6859 <= not w6562 and w6858;
w6860 <= not w6566 and not w6859;
w6861 <= not w6857 and w6860;
w6862 <= not w6566 and not w6861;
w6863 <= b(23) and not w6555;
w6864 <= not w6553 and w6863;
w6865 <= not w6557 and not w6864;
w6866 <= not w6862 and w6865;
w6867 <= not w6557 and not w6866;
w6868 <= b(24) and not w6546;
w6869 <= not w6544 and w6868;
w6870 <= not w6548 and not w6869;
w6871 <= not w6867 and w6870;
w6872 <= not w6548 and not w6871;
w6873 <= b(25) and not w6537;
w6874 <= not w6535 and w6873;
w6875 <= not w6539 and not w6874;
w6876 <= not w6872 and w6875;
w6877 <= not w6539 and not w6876;
w6878 <= b(26) and not w6528;
w6879 <= not w6526 and w6878;
w6880 <= not w6530 and not w6879;
w6881 <= not w6877 and w6880;
w6882 <= not w6530 and not w6881;
w6883 <= b(27) and not w6519;
w6884 <= not w6517 and w6883;
w6885 <= not w6521 and not w6884;
w6886 <= not w6882 and w6885;
w6887 <= not w6521 and not w6886;
w6888 <= b(28) and not w6510;
w6889 <= not w6508 and w6888;
w6890 <= not w6512 and not w6889;
w6891 <= not w6887 and w6890;
w6892 <= not w6512 and not w6891;
w6893 <= b(29) and not w6490;
w6894 <= not w6488 and w6893;
w6895 <= not w6503 and not w6894;
w6896 <= not w6892 and w6895;
w6897 <= not w6503 and not w6896;
w6898 <= b(30) and not w6500;
w6899 <= not w6498 and w6898;
w6900 <= not w6502 and not w6899;
w6901 <= not w6897 and w6900;
w6902 <= not w6502 and not w6901;
w6903 <= w115 and w157;
w6904 <= w341 and w6903;
w6905 <= w338 and w6904;
w6906 <= not w6902 and w6905;
w6907 <= not w6491 and not w6906;
w6908 <= not w6512 and w6895;
w6909 <= not w6891 and w6908;
w6910 <= not w6892 and not w6895;
w6911 <= not w6909 and not w6910;
w6912 <= w6905 and not w6911;
w6913 <= not w6902 and w6912;
w6914 <= not w6907 and not w6913;
w6915 <= not w6501 and not w6906;
w6916 <= not w6503 and w6900;
w6917 <= not w6896 and w6916;
w6918 <= not w6897 and not w6900;
w6919 <= not w6917 and not w6918;
w6920 <= w6906 and not w6919;
w6921 <= not w6915 and not w6920;
w6922 <= not b(31) and not w6921;
w6923 <= not b(30) and not w6914;
w6924 <= not w6511 and not w6906;
w6925 <= not w6521 and w6890;
w6926 <= not w6886 and w6925;
w6927 <= not w6887 and not w6890;
w6928 <= not w6926 and not w6927;
w6929 <= w6905 and not w6928;
w6930 <= not w6902 and w6929;
w6931 <= not w6924 and not w6930;
w6932 <= not b(29) and not w6931;
w6933 <= not w6520 and not w6906;
w6934 <= not w6530 and w6885;
w6935 <= not w6881 and w6934;
w6936 <= not w6882 and not w6885;
w6937 <= not w6935 and not w6936;
w6938 <= w6905 and not w6937;
w6939 <= not w6902 and w6938;
w6940 <= not w6933 and not w6939;
w6941 <= not b(28) and not w6940;
w6942 <= not w6529 and not w6906;
w6943 <= not w6539 and w6880;
w6944 <= not w6876 and w6943;
w6945 <= not w6877 and not w6880;
w6946 <= not w6944 and not w6945;
w6947 <= w6905 and not w6946;
w6948 <= not w6902 and w6947;
w6949 <= not w6942 and not w6948;
w6950 <= not b(27) and not w6949;
w6951 <= not w6538 and not w6906;
w6952 <= not w6548 and w6875;
w6953 <= not w6871 and w6952;
w6954 <= not w6872 and not w6875;
w6955 <= not w6953 and not w6954;
w6956 <= w6905 and not w6955;
w6957 <= not w6902 and w6956;
w6958 <= not w6951 and not w6957;
w6959 <= not b(26) and not w6958;
w6960 <= not w6547 and not w6906;
w6961 <= not w6557 and w6870;
w6962 <= not w6866 and w6961;
w6963 <= not w6867 and not w6870;
w6964 <= not w6962 and not w6963;
w6965 <= w6905 and not w6964;
w6966 <= not w6902 and w6965;
w6967 <= not w6960 and not w6966;
w6968 <= not b(25) and not w6967;
w6969 <= not w6556 and not w6906;
w6970 <= not w6566 and w6865;
w6971 <= not w6861 and w6970;
w6972 <= not w6862 and not w6865;
w6973 <= not w6971 and not w6972;
w6974 <= w6905 and not w6973;
w6975 <= not w6902 and w6974;
w6976 <= not w6969 and not w6975;
w6977 <= not b(24) and not w6976;
w6978 <= not w6565 and not w6906;
w6979 <= not w6575 and w6860;
w6980 <= not w6856 and w6979;
w6981 <= not w6857 and not w6860;
w6982 <= not w6980 and not w6981;
w6983 <= w6905 and not w6982;
w6984 <= not w6902 and w6983;
w6985 <= not w6978 and not w6984;
w6986 <= not b(23) and not w6985;
w6987 <= not w6574 and not w6906;
w6988 <= not w6584 and w6855;
w6989 <= not w6851 and w6988;
w6990 <= not w6852 and not w6855;
w6991 <= not w6989 and not w6990;
w6992 <= w6905 and not w6991;
w6993 <= not w6902 and w6992;
w6994 <= not w6987 and not w6993;
w6995 <= not b(22) and not w6994;
w6996 <= not w6583 and not w6906;
w6997 <= not w6593 and w6850;
w6998 <= not w6846 and w6997;
w6999 <= not w6847 and not w6850;
w7000 <= not w6998 and not w6999;
w7001 <= w6905 and not w7000;
w7002 <= not w6902 and w7001;
w7003 <= not w6996 and not w7002;
w7004 <= not b(21) and not w7003;
w7005 <= not w6592 and not w6906;
w7006 <= not w6602 and w6845;
w7007 <= not w6841 and w7006;
w7008 <= not w6842 and not w6845;
w7009 <= not w7007 and not w7008;
w7010 <= w6905 and not w7009;
w7011 <= not w6902 and w7010;
w7012 <= not w7005 and not w7011;
w7013 <= not b(20) and not w7012;
w7014 <= not w6601 and not w6906;
w7015 <= not w6611 and w6840;
w7016 <= not w6836 and w7015;
w7017 <= not w6837 and not w6840;
w7018 <= not w7016 and not w7017;
w7019 <= w6905 and not w7018;
w7020 <= not w6902 and w7019;
w7021 <= not w7014 and not w7020;
w7022 <= not b(19) and not w7021;
w7023 <= not w6610 and not w6906;
w7024 <= not w6620 and w6835;
w7025 <= not w6831 and w7024;
w7026 <= not w6832 and not w6835;
w7027 <= not w7025 and not w7026;
w7028 <= w6905 and not w7027;
w7029 <= not w6902 and w7028;
w7030 <= not w7023 and not w7029;
w7031 <= not b(18) and not w7030;
w7032 <= not w6619 and not w6906;
w7033 <= not w6629 and w6830;
w7034 <= not w6826 and w7033;
w7035 <= not w6827 and not w6830;
w7036 <= not w7034 and not w7035;
w7037 <= w6905 and not w7036;
w7038 <= not w6902 and w7037;
w7039 <= not w7032 and not w7038;
w7040 <= not b(17) and not w7039;
w7041 <= not w6628 and not w6906;
w7042 <= not w6638 and w6825;
w7043 <= not w6821 and w7042;
w7044 <= not w6822 and not w6825;
w7045 <= not w7043 and not w7044;
w7046 <= w6905 and not w7045;
w7047 <= not w6902 and w7046;
w7048 <= not w7041 and not w7047;
w7049 <= not b(16) and not w7048;
w7050 <= not w6637 and not w6906;
w7051 <= not w6647 and w6820;
w7052 <= not w6816 and w7051;
w7053 <= not w6817 and not w6820;
w7054 <= not w7052 and not w7053;
w7055 <= w6905 and not w7054;
w7056 <= not w6902 and w7055;
w7057 <= not w7050 and not w7056;
w7058 <= not b(15) and not w7057;
w7059 <= not w6646 and not w6906;
w7060 <= not w6656 and w6815;
w7061 <= not w6811 and w7060;
w7062 <= not w6812 and not w6815;
w7063 <= not w7061 and not w7062;
w7064 <= w6905 and not w7063;
w7065 <= not w6902 and w7064;
w7066 <= not w7059 and not w7065;
w7067 <= not b(14) and not w7066;
w7068 <= not w6655 and not w6906;
w7069 <= not w6665 and w6810;
w7070 <= not w6806 and w7069;
w7071 <= not w6807 and not w6810;
w7072 <= not w7070 and not w7071;
w7073 <= w6905 and not w7072;
w7074 <= not w6902 and w7073;
w7075 <= not w7068 and not w7074;
w7076 <= not b(13) and not w7075;
w7077 <= not w6664 and not w6906;
w7078 <= not w6674 and w6805;
w7079 <= not w6801 and w7078;
w7080 <= not w6802 and not w6805;
w7081 <= not w7079 and not w7080;
w7082 <= w6905 and not w7081;
w7083 <= not w6902 and w7082;
w7084 <= not w7077 and not w7083;
w7085 <= not b(12) and not w7084;
w7086 <= not w6673 and not w6906;
w7087 <= not w6683 and w6800;
w7088 <= not w6796 and w7087;
w7089 <= not w6797 and not w6800;
w7090 <= not w7088 and not w7089;
w7091 <= w6905 and not w7090;
w7092 <= not w6902 and w7091;
w7093 <= not w7086 and not w7092;
w7094 <= not b(11) and not w7093;
w7095 <= not w6682 and not w6906;
w7096 <= not w6692 and w6795;
w7097 <= not w6791 and w7096;
w7098 <= not w6792 and not w6795;
w7099 <= not w7097 and not w7098;
w7100 <= w6905 and not w7099;
w7101 <= not w6902 and w7100;
w7102 <= not w7095 and not w7101;
w7103 <= not b(10) and not w7102;
w7104 <= not w6691 and not w6906;
w7105 <= not w6701 and w6790;
w7106 <= not w6786 and w7105;
w7107 <= not w6787 and not w6790;
w7108 <= not w7106 and not w7107;
w7109 <= w6905 and not w7108;
w7110 <= not w6902 and w7109;
w7111 <= not w7104 and not w7110;
w7112 <= not b(9) and not w7111;
w7113 <= not w6700 and not w6906;
w7114 <= not w6710 and w6785;
w7115 <= not w6781 and w7114;
w7116 <= not w6782 and not w6785;
w7117 <= not w7115 and not w7116;
w7118 <= w6905 and not w7117;
w7119 <= not w6902 and w7118;
w7120 <= not w7113 and not w7119;
w7121 <= not b(8) and not w7120;
w7122 <= not w6709 and not w6906;
w7123 <= not w6719 and w6780;
w7124 <= not w6776 and w7123;
w7125 <= not w6777 and not w6780;
w7126 <= not w7124 and not w7125;
w7127 <= w6905 and not w7126;
w7128 <= not w6902 and w7127;
w7129 <= not w7122 and not w7128;
w7130 <= not b(7) and not w7129;
w7131 <= not w6718 and not w6906;
w7132 <= not w6728 and w6775;
w7133 <= not w6771 and w7132;
w7134 <= not w6772 and not w6775;
w7135 <= not w7133 and not w7134;
w7136 <= w6905 and not w7135;
w7137 <= not w6902 and w7136;
w7138 <= not w7131 and not w7137;
w7139 <= not b(6) and not w7138;
w7140 <= not w6727 and not w6906;
w7141 <= not w6737 and w6770;
w7142 <= not w6766 and w7141;
w7143 <= not w6767 and not w6770;
w7144 <= not w7142 and not w7143;
w7145 <= w6905 and not w7144;
w7146 <= not w6902 and w7145;
w7147 <= not w7140 and not w7146;
w7148 <= not b(5) and not w7147;
w7149 <= not w6736 and not w6906;
w7150 <= not w6745 and w6765;
w7151 <= not w6761 and w7150;
w7152 <= not w6762 and not w6765;
w7153 <= not w7151 and not w7152;
w7154 <= w6905 and not w7153;
w7155 <= not w6902 and w7154;
w7156 <= not w7149 and not w7155;
w7157 <= not b(4) and not w7156;
w7158 <= not w6744 and not w6906;
w7159 <= not w6756 and w6760;
w7160 <= not w6755 and w7159;
w7161 <= not w6757 and not w6760;
w7162 <= not w7160 and not w7161;
w7163 <= w6905 and not w7162;
w7164 <= not w6902 and w7163;
w7165 <= not w7158 and not w7164;
w7166 <= not b(3) and not w7165;
w7167 <= not w6749 and not w6906;
w7168 <= not w6752 and w6754;
w7169 <= not w6750 and w7168;
w7170 <= w6905 and not w7169;
w7171 <= not w6755 and w7170;
w7172 <= not w6902 and w7171;
w7173 <= not w7167 and not w7172;
w7174 <= not b(2) and not w7173;
w7175 <= b(0) and not b(31);
w7176 <= w56 and w7175;
w7177 <= w46 and w7176;
w7178 <= w31 and w7177;
w7179 <= not w6902 and w7178;
w7180 <= a(33) and not w7179;
w7181 <= w115 and w6754;
w7182 <= w157 and w7181;
w7183 <= w341 and w7182;
w7184 <= w338 and w7183;
w7185 <= not w6902 and w7184;
w7186 <= not w7180 and not w7185;
w7187 <= b(1) and not w7186;
w7188 <= not b(1) and not w7185;
w7189 <= not w7180 and w7188;
w7190 <= not w7187 and not w7189;
w7191 <= not a(32) and b(0);
w7192 <= not w7190 and not w7191;
w7193 <= not b(1) and not w7186;
w7194 <= not w7192 and not w7193;
w7195 <= b(2) and not w7172;
w7196 <= not w7167 and w7195;
w7197 <= not w7174 and not w7196;
w7198 <= not w7194 and w7197;
w7199 <= not w7174 and not w7198;
w7200 <= b(3) and not w7164;
w7201 <= not w7158 and w7200;
w7202 <= not w7166 and not w7201;
w7203 <= not w7199 and w7202;
w7204 <= not w7166 and not w7203;
w7205 <= b(4) and not w7155;
w7206 <= not w7149 and w7205;
w7207 <= not w7157 and not w7206;
w7208 <= not w7204 and w7207;
w7209 <= not w7157 and not w7208;
w7210 <= b(5) and not w7146;
w7211 <= not w7140 and w7210;
w7212 <= not w7148 and not w7211;
w7213 <= not w7209 and w7212;
w7214 <= not w7148 and not w7213;
w7215 <= b(6) and not w7137;
w7216 <= not w7131 and w7215;
w7217 <= not w7139 and not w7216;
w7218 <= not w7214 and w7217;
w7219 <= not w7139 and not w7218;
w7220 <= b(7) and not w7128;
w7221 <= not w7122 and w7220;
w7222 <= not w7130 and not w7221;
w7223 <= not w7219 and w7222;
w7224 <= not w7130 and not w7223;
w7225 <= b(8) and not w7119;
w7226 <= not w7113 and w7225;
w7227 <= not w7121 and not w7226;
w7228 <= not w7224 and w7227;
w7229 <= not w7121 and not w7228;
w7230 <= b(9) and not w7110;
w7231 <= not w7104 and w7230;
w7232 <= not w7112 and not w7231;
w7233 <= not w7229 and w7232;
w7234 <= not w7112 and not w7233;
w7235 <= b(10) and not w7101;
w7236 <= not w7095 and w7235;
w7237 <= not w7103 and not w7236;
w7238 <= not w7234 and w7237;
w7239 <= not w7103 and not w7238;
w7240 <= b(11) and not w7092;
w7241 <= not w7086 and w7240;
w7242 <= not w7094 and not w7241;
w7243 <= not w7239 and w7242;
w7244 <= not w7094 and not w7243;
w7245 <= b(12) and not w7083;
w7246 <= not w7077 and w7245;
w7247 <= not w7085 and not w7246;
w7248 <= not w7244 and w7247;
w7249 <= not w7085 and not w7248;
w7250 <= b(13) and not w7074;
w7251 <= not w7068 and w7250;
w7252 <= not w7076 and not w7251;
w7253 <= not w7249 and w7252;
w7254 <= not w7076 and not w7253;
w7255 <= b(14) and not w7065;
w7256 <= not w7059 and w7255;
w7257 <= not w7067 and not w7256;
w7258 <= not w7254 and w7257;
w7259 <= not w7067 and not w7258;
w7260 <= b(15) and not w7056;
w7261 <= not w7050 and w7260;
w7262 <= not w7058 and not w7261;
w7263 <= not w7259 and w7262;
w7264 <= not w7058 and not w7263;
w7265 <= b(16) and not w7047;
w7266 <= not w7041 and w7265;
w7267 <= not w7049 and not w7266;
w7268 <= not w7264 and w7267;
w7269 <= not w7049 and not w7268;
w7270 <= b(17) and not w7038;
w7271 <= not w7032 and w7270;
w7272 <= not w7040 and not w7271;
w7273 <= not w7269 and w7272;
w7274 <= not w7040 and not w7273;
w7275 <= b(18) and not w7029;
w7276 <= not w7023 and w7275;
w7277 <= not w7031 and not w7276;
w7278 <= not w7274 and w7277;
w7279 <= not w7031 and not w7278;
w7280 <= b(19) and not w7020;
w7281 <= not w7014 and w7280;
w7282 <= not w7022 and not w7281;
w7283 <= not w7279 and w7282;
w7284 <= not w7022 and not w7283;
w7285 <= b(20) and not w7011;
w7286 <= not w7005 and w7285;
w7287 <= not w7013 and not w7286;
w7288 <= not w7284 and w7287;
w7289 <= not w7013 and not w7288;
w7290 <= b(21) and not w7002;
w7291 <= not w6996 and w7290;
w7292 <= not w7004 and not w7291;
w7293 <= not w7289 and w7292;
w7294 <= not w7004 and not w7293;
w7295 <= b(22) and not w6993;
w7296 <= not w6987 and w7295;
w7297 <= not w6995 and not w7296;
w7298 <= not w7294 and w7297;
w7299 <= not w6995 and not w7298;
w7300 <= b(23) and not w6984;
w7301 <= not w6978 and w7300;
w7302 <= not w6986 and not w7301;
w7303 <= not w7299 and w7302;
w7304 <= not w6986 and not w7303;
w7305 <= b(24) and not w6975;
w7306 <= not w6969 and w7305;
w7307 <= not w6977 and not w7306;
w7308 <= not w7304 and w7307;
w7309 <= not w6977 and not w7308;
w7310 <= b(25) and not w6966;
w7311 <= not w6960 and w7310;
w7312 <= not w6968 and not w7311;
w7313 <= not w7309 and w7312;
w7314 <= not w6968 and not w7313;
w7315 <= b(26) and not w6957;
w7316 <= not w6951 and w7315;
w7317 <= not w6959 and not w7316;
w7318 <= not w7314 and w7317;
w7319 <= not w6959 and not w7318;
w7320 <= b(27) and not w6948;
w7321 <= not w6942 and w7320;
w7322 <= not w6950 and not w7321;
w7323 <= not w7319 and w7322;
w7324 <= not w6950 and not w7323;
w7325 <= b(28) and not w6939;
w7326 <= not w6933 and w7325;
w7327 <= not w6941 and not w7326;
w7328 <= not w7324 and w7327;
w7329 <= not w6941 and not w7328;
w7330 <= b(29) and not w6930;
w7331 <= not w6924 and w7330;
w7332 <= not w6932 and not w7331;
w7333 <= not w7329 and w7332;
w7334 <= not w6932 and not w7333;
w7335 <= b(30) and not w6913;
w7336 <= not w6907 and w7335;
w7337 <= not w6923 and not w7336;
w7338 <= not w7334 and w7337;
w7339 <= not w6923 and not w7338;
w7340 <= b(31) and not w6915;
w7341 <= not w6920 and w7340;
w7342 <= not w6922 and not w7341;
w7343 <= not w7339 and w7342;
w7344 <= not w6922 and not w7343;
w7345 <= w175 and not w7344;
w7346 <= not w6914 and not w7345;
w7347 <= not w6932 and w7337;
w7348 <= not w7333 and w7347;
w7349 <= not w7334 and not w7337;
w7350 <= not w7348 and not w7349;
w7351 <= w175 and not w7350;
w7352 <= not w7344 and w7351;
w7353 <= not w7346 and not w7352;
w7354 <= not b(31) and not w7353;
w7355 <= not w6931 and not w7345;
w7356 <= not w6941 and w7332;
w7357 <= not w7328 and w7356;
w7358 <= not w7329 and not w7332;
w7359 <= not w7357 and not w7358;
w7360 <= w175 and not w7359;
w7361 <= not w7344 and w7360;
w7362 <= not w7355 and not w7361;
w7363 <= not b(30) and not w7362;
w7364 <= not w6940 and not w7345;
w7365 <= not w6950 and w7327;
w7366 <= not w7323 and w7365;
w7367 <= not w7324 and not w7327;
w7368 <= not w7366 and not w7367;
w7369 <= w175 and not w7368;
w7370 <= not w7344 and w7369;
w7371 <= not w7364 and not w7370;
w7372 <= not b(29) and not w7371;
w7373 <= not w6949 and not w7345;
w7374 <= not w6959 and w7322;
w7375 <= not w7318 and w7374;
w7376 <= not w7319 and not w7322;
w7377 <= not w7375 and not w7376;
w7378 <= w175 and not w7377;
w7379 <= not w7344 and w7378;
w7380 <= not w7373 and not w7379;
w7381 <= not b(28) and not w7380;
w7382 <= not w6958 and not w7345;
w7383 <= not w6968 and w7317;
w7384 <= not w7313 and w7383;
w7385 <= not w7314 and not w7317;
w7386 <= not w7384 and not w7385;
w7387 <= w175 and not w7386;
w7388 <= not w7344 and w7387;
w7389 <= not w7382 and not w7388;
w7390 <= not b(27) and not w7389;
w7391 <= not w6967 and not w7345;
w7392 <= not w6977 and w7312;
w7393 <= not w7308 and w7392;
w7394 <= not w7309 and not w7312;
w7395 <= not w7393 and not w7394;
w7396 <= w175 and not w7395;
w7397 <= not w7344 and w7396;
w7398 <= not w7391 and not w7397;
w7399 <= not b(26) and not w7398;
w7400 <= not w6976 and not w7345;
w7401 <= not w6986 and w7307;
w7402 <= not w7303 and w7401;
w7403 <= not w7304 and not w7307;
w7404 <= not w7402 and not w7403;
w7405 <= w175 and not w7404;
w7406 <= not w7344 and w7405;
w7407 <= not w7400 and not w7406;
w7408 <= not b(25) and not w7407;
w7409 <= not w6985 and not w7345;
w7410 <= not w6995 and w7302;
w7411 <= not w7298 and w7410;
w7412 <= not w7299 and not w7302;
w7413 <= not w7411 and not w7412;
w7414 <= w175 and not w7413;
w7415 <= not w7344 and w7414;
w7416 <= not w7409 and not w7415;
w7417 <= not b(24) and not w7416;
w7418 <= not w6994 and not w7345;
w7419 <= not w7004 and w7297;
w7420 <= not w7293 and w7419;
w7421 <= not w7294 and not w7297;
w7422 <= not w7420 and not w7421;
w7423 <= w175 and not w7422;
w7424 <= not w7344 and w7423;
w7425 <= not w7418 and not w7424;
w7426 <= not b(23) and not w7425;
w7427 <= not w7003 and not w7345;
w7428 <= not w7013 and w7292;
w7429 <= not w7288 and w7428;
w7430 <= not w7289 and not w7292;
w7431 <= not w7429 and not w7430;
w7432 <= w175 and not w7431;
w7433 <= not w7344 and w7432;
w7434 <= not w7427 and not w7433;
w7435 <= not b(22) and not w7434;
w7436 <= not w7012 and not w7345;
w7437 <= not w7022 and w7287;
w7438 <= not w7283 and w7437;
w7439 <= not w7284 and not w7287;
w7440 <= not w7438 and not w7439;
w7441 <= w175 and not w7440;
w7442 <= not w7344 and w7441;
w7443 <= not w7436 and not w7442;
w7444 <= not b(21) and not w7443;
w7445 <= not w7021 and not w7345;
w7446 <= not w7031 and w7282;
w7447 <= not w7278 and w7446;
w7448 <= not w7279 and not w7282;
w7449 <= not w7447 and not w7448;
w7450 <= w175 and not w7449;
w7451 <= not w7344 and w7450;
w7452 <= not w7445 and not w7451;
w7453 <= not b(20) and not w7452;
w7454 <= not w7030 and not w7345;
w7455 <= not w7040 and w7277;
w7456 <= not w7273 and w7455;
w7457 <= not w7274 and not w7277;
w7458 <= not w7456 and not w7457;
w7459 <= w175 and not w7458;
w7460 <= not w7344 and w7459;
w7461 <= not w7454 and not w7460;
w7462 <= not b(19) and not w7461;
w7463 <= not w7039 and not w7345;
w7464 <= not w7049 and w7272;
w7465 <= not w7268 and w7464;
w7466 <= not w7269 and not w7272;
w7467 <= not w7465 and not w7466;
w7468 <= w175 and not w7467;
w7469 <= not w7344 and w7468;
w7470 <= not w7463 and not w7469;
w7471 <= not b(18) and not w7470;
w7472 <= not w7048 and not w7345;
w7473 <= not w7058 and w7267;
w7474 <= not w7263 and w7473;
w7475 <= not w7264 and not w7267;
w7476 <= not w7474 and not w7475;
w7477 <= w175 and not w7476;
w7478 <= not w7344 and w7477;
w7479 <= not w7472 and not w7478;
w7480 <= not b(17) and not w7479;
w7481 <= not w7057 and not w7345;
w7482 <= not w7067 and w7262;
w7483 <= not w7258 and w7482;
w7484 <= not w7259 and not w7262;
w7485 <= not w7483 and not w7484;
w7486 <= w175 and not w7485;
w7487 <= not w7344 and w7486;
w7488 <= not w7481 and not w7487;
w7489 <= not b(16) and not w7488;
w7490 <= not w7066 and not w7345;
w7491 <= not w7076 and w7257;
w7492 <= not w7253 and w7491;
w7493 <= not w7254 and not w7257;
w7494 <= not w7492 and not w7493;
w7495 <= w175 and not w7494;
w7496 <= not w7344 and w7495;
w7497 <= not w7490 and not w7496;
w7498 <= not b(15) and not w7497;
w7499 <= not w7075 and not w7345;
w7500 <= not w7085 and w7252;
w7501 <= not w7248 and w7500;
w7502 <= not w7249 and not w7252;
w7503 <= not w7501 and not w7502;
w7504 <= w175 and not w7503;
w7505 <= not w7344 and w7504;
w7506 <= not w7499 and not w7505;
w7507 <= not b(14) and not w7506;
w7508 <= not w7084 and not w7345;
w7509 <= not w7094 and w7247;
w7510 <= not w7243 and w7509;
w7511 <= not w7244 and not w7247;
w7512 <= not w7510 and not w7511;
w7513 <= w175 and not w7512;
w7514 <= not w7344 and w7513;
w7515 <= not w7508 and not w7514;
w7516 <= not b(13) and not w7515;
w7517 <= not w7093 and not w7345;
w7518 <= not w7103 and w7242;
w7519 <= not w7238 and w7518;
w7520 <= not w7239 and not w7242;
w7521 <= not w7519 and not w7520;
w7522 <= w175 and not w7521;
w7523 <= not w7344 and w7522;
w7524 <= not w7517 and not w7523;
w7525 <= not b(12) and not w7524;
w7526 <= not w7102 and not w7345;
w7527 <= not w7112 and w7237;
w7528 <= not w7233 and w7527;
w7529 <= not w7234 and not w7237;
w7530 <= not w7528 and not w7529;
w7531 <= w175 and not w7530;
w7532 <= not w7344 and w7531;
w7533 <= not w7526 and not w7532;
w7534 <= not b(11) and not w7533;
w7535 <= not w7111 and not w7345;
w7536 <= not w7121 and w7232;
w7537 <= not w7228 and w7536;
w7538 <= not w7229 and not w7232;
w7539 <= not w7537 and not w7538;
w7540 <= w175 and not w7539;
w7541 <= not w7344 and w7540;
w7542 <= not w7535 and not w7541;
w7543 <= not b(10) and not w7542;
w7544 <= not w7120 and not w7345;
w7545 <= not w7130 and w7227;
w7546 <= not w7223 and w7545;
w7547 <= not w7224 and not w7227;
w7548 <= not w7546 and not w7547;
w7549 <= w175 and not w7548;
w7550 <= not w7344 and w7549;
w7551 <= not w7544 and not w7550;
w7552 <= not b(9) and not w7551;
w7553 <= not w7129 and not w7345;
w7554 <= not w7139 and w7222;
w7555 <= not w7218 and w7554;
w7556 <= not w7219 and not w7222;
w7557 <= not w7555 and not w7556;
w7558 <= w175 and not w7557;
w7559 <= not w7344 and w7558;
w7560 <= not w7553 and not w7559;
w7561 <= not b(8) and not w7560;
w7562 <= not w7138 and not w7345;
w7563 <= not w7148 and w7217;
w7564 <= not w7213 and w7563;
w7565 <= not w7214 and not w7217;
w7566 <= not w7564 and not w7565;
w7567 <= w175 and not w7566;
w7568 <= not w7344 and w7567;
w7569 <= not w7562 and not w7568;
w7570 <= not b(7) and not w7569;
w7571 <= not w7147 and not w7345;
w7572 <= not w7157 and w7212;
w7573 <= not w7208 and w7572;
w7574 <= not w7209 and not w7212;
w7575 <= not w7573 and not w7574;
w7576 <= w175 and not w7575;
w7577 <= not w7344 and w7576;
w7578 <= not w7571 and not w7577;
w7579 <= not b(6) and not w7578;
w7580 <= not w7156 and not w7345;
w7581 <= not w7166 and w7207;
w7582 <= not w7203 and w7581;
w7583 <= not w7204 and not w7207;
w7584 <= not w7582 and not w7583;
w7585 <= w175 and not w7584;
w7586 <= not w7344 and w7585;
w7587 <= not w7580 and not w7586;
w7588 <= not b(5) and not w7587;
w7589 <= not w7165 and not w7345;
w7590 <= not w7174 and w7202;
w7591 <= not w7198 and w7590;
w7592 <= not w7199 and not w7202;
w7593 <= not w7591 and not w7592;
w7594 <= w175 and not w7593;
w7595 <= not w7344 and w7594;
w7596 <= not w7589 and not w7595;
w7597 <= not b(4) and not w7596;
w7598 <= not w7173 and not w7345;
w7599 <= not w7193 and w7197;
w7600 <= not w7192 and w7599;
w7601 <= not w7194 and not w7197;
w7602 <= not w7600 and not w7601;
w7603 <= w175 and not w7602;
w7604 <= not w7344 and w7603;
w7605 <= not w7598 and not w7604;
w7606 <= not b(3) and not w7605;
w7607 <= not w7186 and not w7345;
w7608 <= not w7189 and w7191;
w7609 <= not w7187 and w7608;
w7610 <= w175 and not w7609;
w7611 <= not w7192 and w7610;
w7612 <= not w7344 and w7611;
w7613 <= not w7607 and not w7612;
w7614 <= not b(2) and not w7613;
w7615 <= b(0) and not b(32);
w7616 <= w157 and w7615;
w7617 <= w341 and w7616;
w7618 <= w338 and w7617;
w7619 <= not w7344 and w7618;
w7620 <= a(32) and not w7619;
w7621 <= w56 and w7191;
w7622 <= w46 and w7621;
w7623 <= w31 and w7622;
w7624 <= not w7344 and w7623;
w7625 <= not w7620 and not w7624;
w7626 <= b(1) and not w7625;
w7627 <= not b(1) and not w7624;
w7628 <= not w7620 and w7627;
w7629 <= not w7626 and not w7628;
w7630 <= not a(31) and b(0);
w7631 <= not w7629 and not w7630;
w7632 <= not b(1) and not w7625;
w7633 <= not w7631 and not w7632;
w7634 <= b(2) and not w7612;
w7635 <= not w7607 and w7634;
w7636 <= not w7614 and not w7635;
w7637 <= not w7633 and w7636;
w7638 <= not w7614 and not w7637;
w7639 <= b(3) and not w7604;
w7640 <= not w7598 and w7639;
w7641 <= not w7606 and not w7640;
w7642 <= not w7638 and w7641;
w7643 <= not w7606 and not w7642;
w7644 <= b(4) and not w7595;
w7645 <= not w7589 and w7644;
w7646 <= not w7597 and not w7645;
w7647 <= not w7643 and w7646;
w7648 <= not w7597 and not w7647;
w7649 <= b(5) and not w7586;
w7650 <= not w7580 and w7649;
w7651 <= not w7588 and not w7650;
w7652 <= not w7648 and w7651;
w7653 <= not w7588 and not w7652;
w7654 <= b(6) and not w7577;
w7655 <= not w7571 and w7654;
w7656 <= not w7579 and not w7655;
w7657 <= not w7653 and w7656;
w7658 <= not w7579 and not w7657;
w7659 <= b(7) and not w7568;
w7660 <= not w7562 and w7659;
w7661 <= not w7570 and not w7660;
w7662 <= not w7658 and w7661;
w7663 <= not w7570 and not w7662;
w7664 <= b(8) and not w7559;
w7665 <= not w7553 and w7664;
w7666 <= not w7561 and not w7665;
w7667 <= not w7663 and w7666;
w7668 <= not w7561 and not w7667;
w7669 <= b(9) and not w7550;
w7670 <= not w7544 and w7669;
w7671 <= not w7552 and not w7670;
w7672 <= not w7668 and w7671;
w7673 <= not w7552 and not w7672;
w7674 <= b(10) and not w7541;
w7675 <= not w7535 and w7674;
w7676 <= not w7543 and not w7675;
w7677 <= not w7673 and w7676;
w7678 <= not w7543 and not w7677;
w7679 <= b(11) and not w7532;
w7680 <= not w7526 and w7679;
w7681 <= not w7534 and not w7680;
w7682 <= not w7678 and w7681;
w7683 <= not w7534 and not w7682;
w7684 <= b(12) and not w7523;
w7685 <= not w7517 and w7684;
w7686 <= not w7525 and not w7685;
w7687 <= not w7683 and w7686;
w7688 <= not w7525 and not w7687;
w7689 <= b(13) and not w7514;
w7690 <= not w7508 and w7689;
w7691 <= not w7516 and not w7690;
w7692 <= not w7688 and w7691;
w7693 <= not w7516 and not w7692;
w7694 <= b(14) and not w7505;
w7695 <= not w7499 and w7694;
w7696 <= not w7507 and not w7695;
w7697 <= not w7693 and w7696;
w7698 <= not w7507 and not w7697;
w7699 <= b(15) and not w7496;
w7700 <= not w7490 and w7699;
w7701 <= not w7498 and not w7700;
w7702 <= not w7698 and w7701;
w7703 <= not w7498 and not w7702;
w7704 <= b(16) and not w7487;
w7705 <= not w7481 and w7704;
w7706 <= not w7489 and not w7705;
w7707 <= not w7703 and w7706;
w7708 <= not w7489 and not w7707;
w7709 <= b(17) and not w7478;
w7710 <= not w7472 and w7709;
w7711 <= not w7480 and not w7710;
w7712 <= not w7708 and w7711;
w7713 <= not w7480 and not w7712;
w7714 <= b(18) and not w7469;
w7715 <= not w7463 and w7714;
w7716 <= not w7471 and not w7715;
w7717 <= not w7713 and w7716;
w7718 <= not w7471 and not w7717;
w7719 <= b(19) and not w7460;
w7720 <= not w7454 and w7719;
w7721 <= not w7462 and not w7720;
w7722 <= not w7718 and w7721;
w7723 <= not w7462 and not w7722;
w7724 <= b(20) and not w7451;
w7725 <= not w7445 and w7724;
w7726 <= not w7453 and not w7725;
w7727 <= not w7723 and w7726;
w7728 <= not w7453 and not w7727;
w7729 <= b(21) and not w7442;
w7730 <= not w7436 and w7729;
w7731 <= not w7444 and not w7730;
w7732 <= not w7728 and w7731;
w7733 <= not w7444 and not w7732;
w7734 <= b(22) and not w7433;
w7735 <= not w7427 and w7734;
w7736 <= not w7435 and not w7735;
w7737 <= not w7733 and w7736;
w7738 <= not w7435 and not w7737;
w7739 <= b(23) and not w7424;
w7740 <= not w7418 and w7739;
w7741 <= not w7426 and not w7740;
w7742 <= not w7738 and w7741;
w7743 <= not w7426 and not w7742;
w7744 <= b(24) and not w7415;
w7745 <= not w7409 and w7744;
w7746 <= not w7417 and not w7745;
w7747 <= not w7743 and w7746;
w7748 <= not w7417 and not w7747;
w7749 <= b(25) and not w7406;
w7750 <= not w7400 and w7749;
w7751 <= not w7408 and not w7750;
w7752 <= not w7748 and w7751;
w7753 <= not w7408 and not w7752;
w7754 <= b(26) and not w7397;
w7755 <= not w7391 and w7754;
w7756 <= not w7399 and not w7755;
w7757 <= not w7753 and w7756;
w7758 <= not w7399 and not w7757;
w7759 <= b(27) and not w7388;
w7760 <= not w7382 and w7759;
w7761 <= not w7390 and not w7760;
w7762 <= not w7758 and w7761;
w7763 <= not w7390 and not w7762;
w7764 <= b(28) and not w7379;
w7765 <= not w7373 and w7764;
w7766 <= not w7381 and not w7765;
w7767 <= not w7763 and w7766;
w7768 <= not w7381 and not w7767;
w7769 <= b(29) and not w7370;
w7770 <= not w7364 and w7769;
w7771 <= not w7372 and not w7770;
w7772 <= not w7768 and w7771;
w7773 <= not w7372 and not w7772;
w7774 <= b(30) and not w7361;
w7775 <= not w7355 and w7774;
w7776 <= not w7363 and not w7775;
w7777 <= not w7773 and w7776;
w7778 <= not w7363 and not w7777;
w7779 <= b(31) and not w7352;
w7780 <= not w7346 and w7779;
w7781 <= not w7354 and not w7780;
w7782 <= not w7778 and w7781;
w7783 <= not w7354 and not w7782;
w7784 <= not w6921 and not w7345;
w7785 <= not w6923 and w7342;
w7786 <= not w7338 and w7785;
w7787 <= not w7339 and not w7342;
w7788 <= not w7786 and not w7787;
w7789 <= w7345 and not w7788;
w7790 <= not w7784 and not w7789;
w7791 <= not b(32) and not w7790;
w7792 <= b(32) and not w7784;
w7793 <= not w7789 and w7792;
w7794 <= w167 and not w7793;
w7795 <= not w7791 and w7794;
w7796 <= not w7783 and w7795;
w7797 <= w175 and not w7790;
w7798 <= not w7796 and not w7797;
w7799 <= not w7363 and w7781;
w7800 <= not w7777 and w7799;
w7801 <= not w7778 and not w7781;
w7802 <= not w7800 and not w7801;
w7803 <= not w7798 and not w7802;
w7804 <= not w7353 and not w7797;
w7805 <= not w7796 and w7804;
w7806 <= not w7803 and not w7805;
w7807 <= not w7354 and not w7793;
w7808 <= not w7791 and w7807;
w7809 <= not w7782 and w7808;
w7810 <= not w7791 and not w7793;
w7811 <= not w7783 and not w7810;
w7812 <= not w7809 and not w7811;
w7813 <= not w7798 and not w7812;
w7814 <= not w7790 and not w7797;
w7815 <= not w7796 and w7814;
w7816 <= not w7813 and not w7815;
w7817 <= not b(33) and not w7816;
w7818 <= not b(32) and not w7806;
w7819 <= not w7372 and w7776;
w7820 <= not w7772 and w7819;
w7821 <= not w7773 and not w7776;
w7822 <= not w7820 and not w7821;
w7823 <= not w7798 and not w7822;
w7824 <= not w7362 and not w7797;
w7825 <= not w7796 and w7824;
w7826 <= not w7823 and not w7825;
w7827 <= not b(31) and not w7826;
w7828 <= not w7381 and w7771;
w7829 <= not w7767 and w7828;
w7830 <= not w7768 and not w7771;
w7831 <= not w7829 and not w7830;
w7832 <= not w7798 and not w7831;
w7833 <= not w7371 and not w7797;
w7834 <= not w7796 and w7833;
w7835 <= not w7832 and not w7834;
w7836 <= not b(30) and not w7835;
w7837 <= not w7390 and w7766;
w7838 <= not w7762 and w7837;
w7839 <= not w7763 and not w7766;
w7840 <= not w7838 and not w7839;
w7841 <= not w7798 and not w7840;
w7842 <= not w7380 and not w7797;
w7843 <= not w7796 and w7842;
w7844 <= not w7841 and not w7843;
w7845 <= not b(29) and not w7844;
w7846 <= not w7399 and w7761;
w7847 <= not w7757 and w7846;
w7848 <= not w7758 and not w7761;
w7849 <= not w7847 and not w7848;
w7850 <= not w7798 and not w7849;
w7851 <= not w7389 and not w7797;
w7852 <= not w7796 and w7851;
w7853 <= not w7850 and not w7852;
w7854 <= not b(28) and not w7853;
w7855 <= not w7408 and w7756;
w7856 <= not w7752 and w7855;
w7857 <= not w7753 and not w7756;
w7858 <= not w7856 and not w7857;
w7859 <= not w7798 and not w7858;
w7860 <= not w7398 and not w7797;
w7861 <= not w7796 and w7860;
w7862 <= not w7859 and not w7861;
w7863 <= not b(27) and not w7862;
w7864 <= not w7417 and w7751;
w7865 <= not w7747 and w7864;
w7866 <= not w7748 and not w7751;
w7867 <= not w7865 and not w7866;
w7868 <= not w7798 and not w7867;
w7869 <= not w7407 and not w7797;
w7870 <= not w7796 and w7869;
w7871 <= not w7868 and not w7870;
w7872 <= not b(26) and not w7871;
w7873 <= not w7426 and w7746;
w7874 <= not w7742 and w7873;
w7875 <= not w7743 and not w7746;
w7876 <= not w7874 and not w7875;
w7877 <= not w7798 and not w7876;
w7878 <= not w7416 and not w7797;
w7879 <= not w7796 and w7878;
w7880 <= not w7877 and not w7879;
w7881 <= not b(25) and not w7880;
w7882 <= not w7435 and w7741;
w7883 <= not w7737 and w7882;
w7884 <= not w7738 and not w7741;
w7885 <= not w7883 and not w7884;
w7886 <= not w7798 and not w7885;
w7887 <= not w7425 and not w7797;
w7888 <= not w7796 and w7887;
w7889 <= not w7886 and not w7888;
w7890 <= not b(24) and not w7889;
w7891 <= not w7444 and w7736;
w7892 <= not w7732 and w7891;
w7893 <= not w7733 and not w7736;
w7894 <= not w7892 and not w7893;
w7895 <= not w7798 and not w7894;
w7896 <= not w7434 and not w7797;
w7897 <= not w7796 and w7896;
w7898 <= not w7895 and not w7897;
w7899 <= not b(23) and not w7898;
w7900 <= not w7453 and w7731;
w7901 <= not w7727 and w7900;
w7902 <= not w7728 and not w7731;
w7903 <= not w7901 and not w7902;
w7904 <= not w7798 and not w7903;
w7905 <= not w7443 and not w7797;
w7906 <= not w7796 and w7905;
w7907 <= not w7904 and not w7906;
w7908 <= not b(22) and not w7907;
w7909 <= not w7462 and w7726;
w7910 <= not w7722 and w7909;
w7911 <= not w7723 and not w7726;
w7912 <= not w7910 and not w7911;
w7913 <= not w7798 and not w7912;
w7914 <= not w7452 and not w7797;
w7915 <= not w7796 and w7914;
w7916 <= not w7913 and not w7915;
w7917 <= not b(21) and not w7916;
w7918 <= not w7471 and w7721;
w7919 <= not w7717 and w7918;
w7920 <= not w7718 and not w7721;
w7921 <= not w7919 and not w7920;
w7922 <= not w7798 and not w7921;
w7923 <= not w7461 and not w7797;
w7924 <= not w7796 and w7923;
w7925 <= not w7922 and not w7924;
w7926 <= not b(20) and not w7925;
w7927 <= not w7480 and w7716;
w7928 <= not w7712 and w7927;
w7929 <= not w7713 and not w7716;
w7930 <= not w7928 and not w7929;
w7931 <= not w7798 and not w7930;
w7932 <= not w7470 and not w7797;
w7933 <= not w7796 and w7932;
w7934 <= not w7931 and not w7933;
w7935 <= not b(19) and not w7934;
w7936 <= not w7489 and w7711;
w7937 <= not w7707 and w7936;
w7938 <= not w7708 and not w7711;
w7939 <= not w7937 and not w7938;
w7940 <= not w7798 and not w7939;
w7941 <= not w7479 and not w7797;
w7942 <= not w7796 and w7941;
w7943 <= not w7940 and not w7942;
w7944 <= not b(18) and not w7943;
w7945 <= not w7498 and w7706;
w7946 <= not w7702 and w7945;
w7947 <= not w7703 and not w7706;
w7948 <= not w7946 and not w7947;
w7949 <= not w7798 and not w7948;
w7950 <= not w7488 and not w7797;
w7951 <= not w7796 and w7950;
w7952 <= not w7949 and not w7951;
w7953 <= not b(17) and not w7952;
w7954 <= not w7507 and w7701;
w7955 <= not w7697 and w7954;
w7956 <= not w7698 and not w7701;
w7957 <= not w7955 and not w7956;
w7958 <= not w7798 and not w7957;
w7959 <= not w7497 and not w7797;
w7960 <= not w7796 and w7959;
w7961 <= not w7958 and not w7960;
w7962 <= not b(16) and not w7961;
w7963 <= not w7516 and w7696;
w7964 <= not w7692 and w7963;
w7965 <= not w7693 and not w7696;
w7966 <= not w7964 and not w7965;
w7967 <= not w7798 and not w7966;
w7968 <= not w7506 and not w7797;
w7969 <= not w7796 and w7968;
w7970 <= not w7967 and not w7969;
w7971 <= not b(15) and not w7970;
w7972 <= not w7525 and w7691;
w7973 <= not w7687 and w7972;
w7974 <= not w7688 and not w7691;
w7975 <= not w7973 and not w7974;
w7976 <= not w7798 and not w7975;
w7977 <= not w7515 and not w7797;
w7978 <= not w7796 and w7977;
w7979 <= not w7976 and not w7978;
w7980 <= not b(14) and not w7979;
w7981 <= not w7534 and w7686;
w7982 <= not w7682 and w7981;
w7983 <= not w7683 and not w7686;
w7984 <= not w7982 and not w7983;
w7985 <= not w7798 and not w7984;
w7986 <= not w7524 and not w7797;
w7987 <= not w7796 and w7986;
w7988 <= not w7985 and not w7987;
w7989 <= not b(13) and not w7988;
w7990 <= not w7543 and w7681;
w7991 <= not w7677 and w7990;
w7992 <= not w7678 and not w7681;
w7993 <= not w7991 and not w7992;
w7994 <= not w7798 and not w7993;
w7995 <= not w7533 and not w7797;
w7996 <= not w7796 and w7995;
w7997 <= not w7994 and not w7996;
w7998 <= not b(12) and not w7997;
w7999 <= not w7552 and w7676;
w8000 <= not w7672 and w7999;
w8001 <= not w7673 and not w7676;
w8002 <= not w8000 and not w8001;
w8003 <= not w7798 and not w8002;
w8004 <= not w7542 and not w7797;
w8005 <= not w7796 and w8004;
w8006 <= not w8003 and not w8005;
w8007 <= not b(11) and not w8006;
w8008 <= not w7561 and w7671;
w8009 <= not w7667 and w8008;
w8010 <= not w7668 and not w7671;
w8011 <= not w8009 and not w8010;
w8012 <= not w7798 and not w8011;
w8013 <= not w7551 and not w7797;
w8014 <= not w7796 and w8013;
w8015 <= not w8012 and not w8014;
w8016 <= not b(10) and not w8015;
w8017 <= not w7570 and w7666;
w8018 <= not w7662 and w8017;
w8019 <= not w7663 and not w7666;
w8020 <= not w8018 and not w8019;
w8021 <= not w7798 and not w8020;
w8022 <= not w7560 and not w7797;
w8023 <= not w7796 and w8022;
w8024 <= not w8021 and not w8023;
w8025 <= not b(9) and not w8024;
w8026 <= not w7579 and w7661;
w8027 <= not w7657 and w8026;
w8028 <= not w7658 and not w7661;
w8029 <= not w8027 and not w8028;
w8030 <= not w7798 and not w8029;
w8031 <= not w7569 and not w7797;
w8032 <= not w7796 and w8031;
w8033 <= not w8030 and not w8032;
w8034 <= not b(8) and not w8033;
w8035 <= not w7588 and w7656;
w8036 <= not w7652 and w8035;
w8037 <= not w7653 and not w7656;
w8038 <= not w8036 and not w8037;
w8039 <= not w7798 and not w8038;
w8040 <= not w7578 and not w7797;
w8041 <= not w7796 and w8040;
w8042 <= not w8039 and not w8041;
w8043 <= not b(7) and not w8042;
w8044 <= not w7597 and w7651;
w8045 <= not w7647 and w8044;
w8046 <= not w7648 and not w7651;
w8047 <= not w8045 and not w8046;
w8048 <= not w7798 and not w8047;
w8049 <= not w7587 and not w7797;
w8050 <= not w7796 and w8049;
w8051 <= not w8048 and not w8050;
w8052 <= not b(6) and not w8051;
w8053 <= not w7606 and w7646;
w8054 <= not w7642 and w8053;
w8055 <= not w7643 and not w7646;
w8056 <= not w8054 and not w8055;
w8057 <= not w7798 and not w8056;
w8058 <= not w7596 and not w7797;
w8059 <= not w7796 and w8058;
w8060 <= not w8057 and not w8059;
w8061 <= not b(5) and not w8060;
w8062 <= not w7614 and w7641;
w8063 <= not w7637 and w8062;
w8064 <= not w7638 and not w7641;
w8065 <= not w8063 and not w8064;
w8066 <= not w7798 and not w8065;
w8067 <= not w7605 and not w7797;
w8068 <= not w7796 and w8067;
w8069 <= not w8066 and not w8068;
w8070 <= not b(4) and not w8069;
w8071 <= not w7632 and w7636;
w8072 <= not w7631 and w8071;
w8073 <= not w7633 and not w7636;
w8074 <= not w8072 and not w8073;
w8075 <= not w7798 and not w8074;
w8076 <= not w7613 and not w7797;
w8077 <= not w7796 and w8076;
w8078 <= not w8075 and not w8077;
w8079 <= not b(3) and not w8078;
w8080 <= not w7628 and w7630;
w8081 <= not w7626 and w8080;
w8082 <= not w7631 and not w8081;
w8083 <= not w7798 and w8082;
w8084 <= not w7625 and not w7797;
w8085 <= not w7796 and w8084;
w8086 <= not w8083 and not w8085;
w8087 <= not b(2) and not w8086;
w8088 <= b(0) and not w7798;
w8089 <= a(31) and not w8088;
w8090 <= w7630 and not w7798;
w8091 <= not w8089 and not w8090;
w8092 <= b(1) and not w8091;
w8093 <= not b(1) and not w8090;
w8094 <= not w8089 and w8093;
w8095 <= not w8092 and not w8094;
w8096 <= not a(30) and b(0);
w8097 <= not w8095 and not w8096;
w8098 <= not b(1) and not w8091;
w8099 <= not w8097 and not w8098;
w8100 <= b(2) and not w8085;
w8101 <= not w8083 and w8100;
w8102 <= not w8087 and not w8101;
w8103 <= not w8099 and w8102;
w8104 <= not w8087 and not w8103;
w8105 <= b(3) and not w8077;
w8106 <= not w8075 and w8105;
w8107 <= not w8079 and not w8106;
w8108 <= not w8104 and w8107;
w8109 <= not w8079 and not w8108;
w8110 <= b(4) and not w8068;
w8111 <= not w8066 and w8110;
w8112 <= not w8070 and not w8111;
w8113 <= not w8109 and w8112;
w8114 <= not w8070 and not w8113;
w8115 <= b(5) and not w8059;
w8116 <= not w8057 and w8115;
w8117 <= not w8061 and not w8116;
w8118 <= not w8114 and w8117;
w8119 <= not w8061 and not w8118;
w8120 <= b(6) and not w8050;
w8121 <= not w8048 and w8120;
w8122 <= not w8052 and not w8121;
w8123 <= not w8119 and w8122;
w8124 <= not w8052 and not w8123;
w8125 <= b(7) and not w8041;
w8126 <= not w8039 and w8125;
w8127 <= not w8043 and not w8126;
w8128 <= not w8124 and w8127;
w8129 <= not w8043 and not w8128;
w8130 <= b(8) and not w8032;
w8131 <= not w8030 and w8130;
w8132 <= not w8034 and not w8131;
w8133 <= not w8129 and w8132;
w8134 <= not w8034 and not w8133;
w8135 <= b(9) and not w8023;
w8136 <= not w8021 and w8135;
w8137 <= not w8025 and not w8136;
w8138 <= not w8134 and w8137;
w8139 <= not w8025 and not w8138;
w8140 <= b(10) and not w8014;
w8141 <= not w8012 and w8140;
w8142 <= not w8016 and not w8141;
w8143 <= not w8139 and w8142;
w8144 <= not w8016 and not w8143;
w8145 <= b(11) and not w8005;
w8146 <= not w8003 and w8145;
w8147 <= not w8007 and not w8146;
w8148 <= not w8144 and w8147;
w8149 <= not w8007 and not w8148;
w8150 <= b(12) and not w7996;
w8151 <= not w7994 and w8150;
w8152 <= not w7998 and not w8151;
w8153 <= not w8149 and w8152;
w8154 <= not w7998 and not w8153;
w8155 <= b(13) and not w7987;
w8156 <= not w7985 and w8155;
w8157 <= not w7989 and not w8156;
w8158 <= not w8154 and w8157;
w8159 <= not w7989 and not w8158;
w8160 <= b(14) and not w7978;
w8161 <= not w7976 and w8160;
w8162 <= not w7980 and not w8161;
w8163 <= not w8159 and w8162;
w8164 <= not w7980 and not w8163;
w8165 <= b(15) and not w7969;
w8166 <= not w7967 and w8165;
w8167 <= not w7971 and not w8166;
w8168 <= not w8164 and w8167;
w8169 <= not w7971 and not w8168;
w8170 <= b(16) and not w7960;
w8171 <= not w7958 and w8170;
w8172 <= not w7962 and not w8171;
w8173 <= not w8169 and w8172;
w8174 <= not w7962 and not w8173;
w8175 <= b(17) and not w7951;
w8176 <= not w7949 and w8175;
w8177 <= not w7953 and not w8176;
w8178 <= not w8174 and w8177;
w8179 <= not w7953 and not w8178;
w8180 <= b(18) and not w7942;
w8181 <= not w7940 and w8180;
w8182 <= not w7944 and not w8181;
w8183 <= not w8179 and w8182;
w8184 <= not w7944 and not w8183;
w8185 <= b(19) and not w7933;
w8186 <= not w7931 and w8185;
w8187 <= not w7935 and not w8186;
w8188 <= not w8184 and w8187;
w8189 <= not w7935 and not w8188;
w8190 <= b(20) and not w7924;
w8191 <= not w7922 and w8190;
w8192 <= not w7926 and not w8191;
w8193 <= not w8189 and w8192;
w8194 <= not w7926 and not w8193;
w8195 <= b(21) and not w7915;
w8196 <= not w7913 and w8195;
w8197 <= not w7917 and not w8196;
w8198 <= not w8194 and w8197;
w8199 <= not w7917 and not w8198;
w8200 <= b(22) and not w7906;
w8201 <= not w7904 and w8200;
w8202 <= not w7908 and not w8201;
w8203 <= not w8199 and w8202;
w8204 <= not w7908 and not w8203;
w8205 <= b(23) and not w7897;
w8206 <= not w7895 and w8205;
w8207 <= not w7899 and not w8206;
w8208 <= not w8204 and w8207;
w8209 <= not w7899 and not w8208;
w8210 <= b(24) and not w7888;
w8211 <= not w7886 and w8210;
w8212 <= not w7890 and not w8211;
w8213 <= not w8209 and w8212;
w8214 <= not w7890 and not w8213;
w8215 <= b(25) and not w7879;
w8216 <= not w7877 and w8215;
w8217 <= not w7881 and not w8216;
w8218 <= not w8214 and w8217;
w8219 <= not w7881 and not w8218;
w8220 <= b(26) and not w7870;
w8221 <= not w7868 and w8220;
w8222 <= not w7872 and not w8221;
w8223 <= not w8219 and w8222;
w8224 <= not w7872 and not w8223;
w8225 <= b(27) and not w7861;
w8226 <= not w7859 and w8225;
w8227 <= not w7863 and not w8226;
w8228 <= not w8224 and w8227;
w8229 <= not w7863 and not w8228;
w8230 <= b(28) and not w7852;
w8231 <= not w7850 and w8230;
w8232 <= not w7854 and not w8231;
w8233 <= not w8229 and w8232;
w8234 <= not w7854 and not w8233;
w8235 <= b(29) and not w7843;
w8236 <= not w7841 and w8235;
w8237 <= not w7845 and not w8236;
w8238 <= not w8234 and w8237;
w8239 <= not w7845 and not w8238;
w8240 <= b(30) and not w7834;
w8241 <= not w7832 and w8240;
w8242 <= not w7836 and not w8241;
w8243 <= not w8239 and w8242;
w8244 <= not w7836 and not w8243;
w8245 <= b(31) and not w7825;
w8246 <= not w7823 and w8245;
w8247 <= not w7827 and not w8246;
w8248 <= not w8244 and w8247;
w8249 <= not w7827 and not w8248;
w8250 <= b(32) and not w7805;
w8251 <= not w7803 and w8250;
w8252 <= not w7818 and not w8251;
w8253 <= not w8249 and w8252;
w8254 <= not w7818 and not w8253;
w8255 <= b(33) and not w7815;
w8256 <= not w7813 and w8255;
w8257 <= not w7817 and not w8256;
w8258 <= not w8254 and w8257;
w8259 <= not w7817 and not w8258;
w8260 <= w37 and w55;
w8261 <= w83 and w8260;
w8262 <= w81 and w8261;
w8263 <= not w8259 and w8262;
w8264 <= not w7806 and not w8263;
w8265 <= not w7827 and w8252;
w8266 <= not w8248 and w8265;
w8267 <= not w8249 and not w8252;
w8268 <= not w8266 and not w8267;
w8269 <= w8262 and not w8268;
w8270 <= not w8259 and w8269;
w8271 <= not w8264 and not w8270;
w8272 <= not w7816 and not w8263;
w8273 <= not w7818 and w8257;
w8274 <= not w8253 and w8273;
w8275 <= not w8254 and not w8257;
w8276 <= not w8274 and not w8275;
w8277 <= w8263 and not w8276;
w8278 <= not w8272 and not w8277;
w8279 <= not b(34) and not w8278;
w8280 <= not b(33) and not w8271;
w8281 <= not w7826 and not w8263;
w8282 <= not w7836 and w8247;
w8283 <= not w8243 and w8282;
w8284 <= not w8244 and not w8247;
w8285 <= not w8283 and not w8284;
w8286 <= w8262 and not w8285;
w8287 <= not w8259 and w8286;
w8288 <= not w8281 and not w8287;
w8289 <= not b(32) and not w8288;
w8290 <= not w7835 and not w8263;
w8291 <= not w7845 and w8242;
w8292 <= not w8238 and w8291;
w8293 <= not w8239 and not w8242;
w8294 <= not w8292 and not w8293;
w8295 <= w8262 and not w8294;
w8296 <= not w8259 and w8295;
w8297 <= not w8290 and not w8296;
w8298 <= not b(31) and not w8297;
w8299 <= not w7844 and not w8263;
w8300 <= not w7854 and w8237;
w8301 <= not w8233 and w8300;
w8302 <= not w8234 and not w8237;
w8303 <= not w8301 and not w8302;
w8304 <= w8262 and not w8303;
w8305 <= not w8259 and w8304;
w8306 <= not w8299 and not w8305;
w8307 <= not b(30) and not w8306;
w8308 <= not w7853 and not w8263;
w8309 <= not w7863 and w8232;
w8310 <= not w8228 and w8309;
w8311 <= not w8229 and not w8232;
w8312 <= not w8310 and not w8311;
w8313 <= w8262 and not w8312;
w8314 <= not w8259 and w8313;
w8315 <= not w8308 and not w8314;
w8316 <= not b(29) and not w8315;
w8317 <= not w7862 and not w8263;
w8318 <= not w7872 and w8227;
w8319 <= not w8223 and w8318;
w8320 <= not w8224 and not w8227;
w8321 <= not w8319 and not w8320;
w8322 <= w8262 and not w8321;
w8323 <= not w8259 and w8322;
w8324 <= not w8317 and not w8323;
w8325 <= not b(28) and not w8324;
w8326 <= not w7871 and not w8263;
w8327 <= not w7881 and w8222;
w8328 <= not w8218 and w8327;
w8329 <= not w8219 and not w8222;
w8330 <= not w8328 and not w8329;
w8331 <= w8262 and not w8330;
w8332 <= not w8259 and w8331;
w8333 <= not w8326 and not w8332;
w8334 <= not b(27) and not w8333;
w8335 <= not w7880 and not w8263;
w8336 <= not w7890 and w8217;
w8337 <= not w8213 and w8336;
w8338 <= not w8214 and not w8217;
w8339 <= not w8337 and not w8338;
w8340 <= w8262 and not w8339;
w8341 <= not w8259 and w8340;
w8342 <= not w8335 and not w8341;
w8343 <= not b(26) and not w8342;
w8344 <= not w7889 and not w8263;
w8345 <= not w7899 and w8212;
w8346 <= not w8208 and w8345;
w8347 <= not w8209 and not w8212;
w8348 <= not w8346 and not w8347;
w8349 <= w8262 and not w8348;
w8350 <= not w8259 and w8349;
w8351 <= not w8344 and not w8350;
w8352 <= not b(25) and not w8351;
w8353 <= not w7898 and not w8263;
w8354 <= not w7908 and w8207;
w8355 <= not w8203 and w8354;
w8356 <= not w8204 and not w8207;
w8357 <= not w8355 and not w8356;
w8358 <= w8262 and not w8357;
w8359 <= not w8259 and w8358;
w8360 <= not w8353 and not w8359;
w8361 <= not b(24) and not w8360;
w8362 <= not w7907 and not w8263;
w8363 <= not w7917 and w8202;
w8364 <= not w8198 and w8363;
w8365 <= not w8199 and not w8202;
w8366 <= not w8364 and not w8365;
w8367 <= w8262 and not w8366;
w8368 <= not w8259 and w8367;
w8369 <= not w8362 and not w8368;
w8370 <= not b(23) and not w8369;
w8371 <= not w7916 and not w8263;
w8372 <= not w7926 and w8197;
w8373 <= not w8193 and w8372;
w8374 <= not w8194 and not w8197;
w8375 <= not w8373 and not w8374;
w8376 <= w8262 and not w8375;
w8377 <= not w8259 and w8376;
w8378 <= not w8371 and not w8377;
w8379 <= not b(22) and not w8378;
w8380 <= not w7925 and not w8263;
w8381 <= not w7935 and w8192;
w8382 <= not w8188 and w8381;
w8383 <= not w8189 and not w8192;
w8384 <= not w8382 and not w8383;
w8385 <= w8262 and not w8384;
w8386 <= not w8259 and w8385;
w8387 <= not w8380 and not w8386;
w8388 <= not b(21) and not w8387;
w8389 <= not w7934 and not w8263;
w8390 <= not w7944 and w8187;
w8391 <= not w8183 and w8390;
w8392 <= not w8184 and not w8187;
w8393 <= not w8391 and not w8392;
w8394 <= w8262 and not w8393;
w8395 <= not w8259 and w8394;
w8396 <= not w8389 and not w8395;
w8397 <= not b(20) and not w8396;
w8398 <= not w7943 and not w8263;
w8399 <= not w7953 and w8182;
w8400 <= not w8178 and w8399;
w8401 <= not w8179 and not w8182;
w8402 <= not w8400 and not w8401;
w8403 <= w8262 and not w8402;
w8404 <= not w8259 and w8403;
w8405 <= not w8398 and not w8404;
w8406 <= not b(19) and not w8405;
w8407 <= not w7952 and not w8263;
w8408 <= not w7962 and w8177;
w8409 <= not w8173 and w8408;
w8410 <= not w8174 and not w8177;
w8411 <= not w8409 and not w8410;
w8412 <= w8262 and not w8411;
w8413 <= not w8259 and w8412;
w8414 <= not w8407 and not w8413;
w8415 <= not b(18) and not w8414;
w8416 <= not w7961 and not w8263;
w8417 <= not w7971 and w8172;
w8418 <= not w8168 and w8417;
w8419 <= not w8169 and not w8172;
w8420 <= not w8418 and not w8419;
w8421 <= w8262 and not w8420;
w8422 <= not w8259 and w8421;
w8423 <= not w8416 and not w8422;
w8424 <= not b(17) and not w8423;
w8425 <= not w7970 and not w8263;
w8426 <= not w7980 and w8167;
w8427 <= not w8163 and w8426;
w8428 <= not w8164 and not w8167;
w8429 <= not w8427 and not w8428;
w8430 <= w8262 and not w8429;
w8431 <= not w8259 and w8430;
w8432 <= not w8425 and not w8431;
w8433 <= not b(16) and not w8432;
w8434 <= not w7979 and not w8263;
w8435 <= not w7989 and w8162;
w8436 <= not w8158 and w8435;
w8437 <= not w8159 and not w8162;
w8438 <= not w8436 and not w8437;
w8439 <= w8262 and not w8438;
w8440 <= not w8259 and w8439;
w8441 <= not w8434 and not w8440;
w8442 <= not b(15) and not w8441;
w8443 <= not w7988 and not w8263;
w8444 <= not w7998 and w8157;
w8445 <= not w8153 and w8444;
w8446 <= not w8154 and not w8157;
w8447 <= not w8445 and not w8446;
w8448 <= w8262 and not w8447;
w8449 <= not w8259 and w8448;
w8450 <= not w8443 and not w8449;
w8451 <= not b(14) and not w8450;
w8452 <= not w7997 and not w8263;
w8453 <= not w8007 and w8152;
w8454 <= not w8148 and w8453;
w8455 <= not w8149 and not w8152;
w8456 <= not w8454 and not w8455;
w8457 <= w8262 and not w8456;
w8458 <= not w8259 and w8457;
w8459 <= not w8452 and not w8458;
w8460 <= not b(13) and not w8459;
w8461 <= not w8006 and not w8263;
w8462 <= not w8016 and w8147;
w8463 <= not w8143 and w8462;
w8464 <= not w8144 and not w8147;
w8465 <= not w8463 and not w8464;
w8466 <= w8262 and not w8465;
w8467 <= not w8259 and w8466;
w8468 <= not w8461 and not w8467;
w8469 <= not b(12) and not w8468;
w8470 <= not w8015 and not w8263;
w8471 <= not w8025 and w8142;
w8472 <= not w8138 and w8471;
w8473 <= not w8139 and not w8142;
w8474 <= not w8472 and not w8473;
w8475 <= w8262 and not w8474;
w8476 <= not w8259 and w8475;
w8477 <= not w8470 and not w8476;
w8478 <= not b(11) and not w8477;
w8479 <= not w8024 and not w8263;
w8480 <= not w8034 and w8137;
w8481 <= not w8133 and w8480;
w8482 <= not w8134 and not w8137;
w8483 <= not w8481 and not w8482;
w8484 <= w8262 and not w8483;
w8485 <= not w8259 and w8484;
w8486 <= not w8479 and not w8485;
w8487 <= not b(10) and not w8486;
w8488 <= not w8033 and not w8263;
w8489 <= not w8043 and w8132;
w8490 <= not w8128 and w8489;
w8491 <= not w8129 and not w8132;
w8492 <= not w8490 and not w8491;
w8493 <= w8262 and not w8492;
w8494 <= not w8259 and w8493;
w8495 <= not w8488 and not w8494;
w8496 <= not b(9) and not w8495;
w8497 <= not w8042 and not w8263;
w8498 <= not w8052 and w8127;
w8499 <= not w8123 and w8498;
w8500 <= not w8124 and not w8127;
w8501 <= not w8499 and not w8500;
w8502 <= w8262 and not w8501;
w8503 <= not w8259 and w8502;
w8504 <= not w8497 and not w8503;
w8505 <= not b(8) and not w8504;
w8506 <= not w8051 and not w8263;
w8507 <= not w8061 and w8122;
w8508 <= not w8118 and w8507;
w8509 <= not w8119 and not w8122;
w8510 <= not w8508 and not w8509;
w8511 <= w8262 and not w8510;
w8512 <= not w8259 and w8511;
w8513 <= not w8506 and not w8512;
w8514 <= not b(7) and not w8513;
w8515 <= not w8060 and not w8263;
w8516 <= not w8070 and w8117;
w8517 <= not w8113 and w8516;
w8518 <= not w8114 and not w8117;
w8519 <= not w8517 and not w8518;
w8520 <= w8262 and not w8519;
w8521 <= not w8259 and w8520;
w8522 <= not w8515 and not w8521;
w8523 <= not b(6) and not w8522;
w8524 <= not w8069 and not w8263;
w8525 <= not w8079 and w8112;
w8526 <= not w8108 and w8525;
w8527 <= not w8109 and not w8112;
w8528 <= not w8526 and not w8527;
w8529 <= w8262 and not w8528;
w8530 <= not w8259 and w8529;
w8531 <= not w8524 and not w8530;
w8532 <= not b(5) and not w8531;
w8533 <= not w8078 and not w8263;
w8534 <= not w8087 and w8107;
w8535 <= not w8103 and w8534;
w8536 <= not w8104 and not w8107;
w8537 <= not w8535 and not w8536;
w8538 <= w8262 and not w8537;
w8539 <= not w8259 and w8538;
w8540 <= not w8533 and not w8539;
w8541 <= not b(4) and not w8540;
w8542 <= not w8086 and not w8263;
w8543 <= not w8098 and w8102;
w8544 <= not w8097 and w8543;
w8545 <= not w8099 and not w8102;
w8546 <= not w8544 and not w8545;
w8547 <= w8262 and not w8546;
w8548 <= not w8259 and w8547;
w8549 <= not w8542 and not w8548;
w8550 <= not b(3) and not w8549;
w8551 <= not w8091 and not w8263;
w8552 <= not w8094 and w8096;
w8553 <= not w8092 and w8552;
w8554 <= w8262 and not w8553;
w8555 <= not w8097 and w8554;
w8556 <= not w8259 and w8555;
w8557 <= not w8551 and not w8556;
w8558 <= not b(2) and not w8557;
w8559 <= b(0) and not b(34);
w8560 <= w156 and w8559;
w8561 <= w154 and w8560;
w8562 <= w165 and w8561;
w8563 <= w151 and w8562;
w8564 <= not w8259 and w8563;
w8565 <= a(30) and not w8564;
w8566 <= w55 and w8096;
w8567 <= w37 and w8566;
w8568 <= w83 and w8567;
w8569 <= w81 and w8568;
w8570 <= not w8259 and w8569;
w8571 <= not w8565 and not w8570;
w8572 <= b(1) and not w8571;
w8573 <= not b(1) and not w8570;
w8574 <= not w8565 and w8573;
w8575 <= not w8572 and not w8574;
w8576 <= not a(29) and b(0);
w8577 <= not w8575 and not w8576;
w8578 <= not b(1) and not w8571;
w8579 <= not w8577 and not w8578;
w8580 <= b(2) and not w8556;
w8581 <= not w8551 and w8580;
w8582 <= not w8558 and not w8581;
w8583 <= not w8579 and w8582;
w8584 <= not w8558 and not w8583;
w8585 <= b(3) and not w8548;
w8586 <= not w8542 and w8585;
w8587 <= not w8550 and not w8586;
w8588 <= not w8584 and w8587;
w8589 <= not w8550 and not w8588;
w8590 <= b(4) and not w8539;
w8591 <= not w8533 and w8590;
w8592 <= not w8541 and not w8591;
w8593 <= not w8589 and w8592;
w8594 <= not w8541 and not w8593;
w8595 <= b(5) and not w8530;
w8596 <= not w8524 and w8595;
w8597 <= not w8532 and not w8596;
w8598 <= not w8594 and w8597;
w8599 <= not w8532 and not w8598;
w8600 <= b(6) and not w8521;
w8601 <= not w8515 and w8600;
w8602 <= not w8523 and not w8601;
w8603 <= not w8599 and w8602;
w8604 <= not w8523 and not w8603;
w8605 <= b(7) and not w8512;
w8606 <= not w8506 and w8605;
w8607 <= not w8514 and not w8606;
w8608 <= not w8604 and w8607;
w8609 <= not w8514 and not w8608;
w8610 <= b(8) and not w8503;
w8611 <= not w8497 and w8610;
w8612 <= not w8505 and not w8611;
w8613 <= not w8609 and w8612;
w8614 <= not w8505 and not w8613;
w8615 <= b(9) and not w8494;
w8616 <= not w8488 and w8615;
w8617 <= not w8496 and not w8616;
w8618 <= not w8614 and w8617;
w8619 <= not w8496 and not w8618;
w8620 <= b(10) and not w8485;
w8621 <= not w8479 and w8620;
w8622 <= not w8487 and not w8621;
w8623 <= not w8619 and w8622;
w8624 <= not w8487 and not w8623;
w8625 <= b(11) and not w8476;
w8626 <= not w8470 and w8625;
w8627 <= not w8478 and not w8626;
w8628 <= not w8624 and w8627;
w8629 <= not w8478 and not w8628;
w8630 <= b(12) and not w8467;
w8631 <= not w8461 and w8630;
w8632 <= not w8469 and not w8631;
w8633 <= not w8629 and w8632;
w8634 <= not w8469 and not w8633;
w8635 <= b(13) and not w8458;
w8636 <= not w8452 and w8635;
w8637 <= not w8460 and not w8636;
w8638 <= not w8634 and w8637;
w8639 <= not w8460 and not w8638;
w8640 <= b(14) and not w8449;
w8641 <= not w8443 and w8640;
w8642 <= not w8451 and not w8641;
w8643 <= not w8639 and w8642;
w8644 <= not w8451 and not w8643;
w8645 <= b(15) and not w8440;
w8646 <= not w8434 and w8645;
w8647 <= not w8442 and not w8646;
w8648 <= not w8644 and w8647;
w8649 <= not w8442 and not w8648;
w8650 <= b(16) and not w8431;
w8651 <= not w8425 and w8650;
w8652 <= not w8433 and not w8651;
w8653 <= not w8649 and w8652;
w8654 <= not w8433 and not w8653;
w8655 <= b(17) and not w8422;
w8656 <= not w8416 and w8655;
w8657 <= not w8424 and not w8656;
w8658 <= not w8654 and w8657;
w8659 <= not w8424 and not w8658;
w8660 <= b(18) and not w8413;
w8661 <= not w8407 and w8660;
w8662 <= not w8415 and not w8661;
w8663 <= not w8659 and w8662;
w8664 <= not w8415 and not w8663;
w8665 <= b(19) and not w8404;
w8666 <= not w8398 and w8665;
w8667 <= not w8406 and not w8666;
w8668 <= not w8664 and w8667;
w8669 <= not w8406 and not w8668;
w8670 <= b(20) and not w8395;
w8671 <= not w8389 and w8670;
w8672 <= not w8397 and not w8671;
w8673 <= not w8669 and w8672;
w8674 <= not w8397 and not w8673;
w8675 <= b(21) and not w8386;
w8676 <= not w8380 and w8675;
w8677 <= not w8388 and not w8676;
w8678 <= not w8674 and w8677;
w8679 <= not w8388 and not w8678;
w8680 <= b(22) and not w8377;
w8681 <= not w8371 and w8680;
w8682 <= not w8379 and not w8681;
w8683 <= not w8679 and w8682;
w8684 <= not w8379 and not w8683;
w8685 <= b(23) and not w8368;
w8686 <= not w8362 and w8685;
w8687 <= not w8370 and not w8686;
w8688 <= not w8684 and w8687;
w8689 <= not w8370 and not w8688;
w8690 <= b(24) and not w8359;
w8691 <= not w8353 and w8690;
w8692 <= not w8361 and not w8691;
w8693 <= not w8689 and w8692;
w8694 <= not w8361 and not w8693;
w8695 <= b(25) and not w8350;
w8696 <= not w8344 and w8695;
w8697 <= not w8352 and not w8696;
w8698 <= not w8694 and w8697;
w8699 <= not w8352 and not w8698;
w8700 <= b(26) and not w8341;
w8701 <= not w8335 and w8700;
w8702 <= not w8343 and not w8701;
w8703 <= not w8699 and w8702;
w8704 <= not w8343 and not w8703;
w8705 <= b(27) and not w8332;
w8706 <= not w8326 and w8705;
w8707 <= not w8334 and not w8706;
w8708 <= not w8704 and w8707;
w8709 <= not w8334 and not w8708;
w8710 <= b(28) and not w8323;
w8711 <= not w8317 and w8710;
w8712 <= not w8325 and not w8711;
w8713 <= not w8709 and w8712;
w8714 <= not w8325 and not w8713;
w8715 <= b(29) and not w8314;
w8716 <= not w8308 and w8715;
w8717 <= not w8316 and not w8716;
w8718 <= not w8714 and w8717;
w8719 <= not w8316 and not w8718;
w8720 <= b(30) and not w8305;
w8721 <= not w8299 and w8720;
w8722 <= not w8307 and not w8721;
w8723 <= not w8719 and w8722;
w8724 <= not w8307 and not w8723;
w8725 <= b(31) and not w8296;
w8726 <= not w8290 and w8725;
w8727 <= not w8298 and not w8726;
w8728 <= not w8724 and w8727;
w8729 <= not w8298 and not w8728;
w8730 <= b(32) and not w8287;
w8731 <= not w8281 and w8730;
w8732 <= not w8289 and not w8731;
w8733 <= not w8729 and w8732;
w8734 <= not w8289 and not w8733;
w8735 <= b(33) and not w8270;
w8736 <= not w8264 and w8735;
w8737 <= not w8280 and not w8736;
w8738 <= not w8734 and w8737;
w8739 <= not w8280 and not w8738;
w8740 <= b(34) and not w8272;
w8741 <= not w8277 and w8740;
w8742 <= not w8279 and not w8741;
w8743 <= not w8739 and w8742;
w8744 <= not w8279 and not w8743;
w8745 <= w154 and w156;
w8746 <= w165 and w8745;
w8747 <= w151 and w8746;
w8748 <= not w8744 and w8747;
w8749 <= not w8271 and not w8748;
w8750 <= not w8289 and w8737;
w8751 <= not w8733 and w8750;
w8752 <= not w8734 and not w8737;
w8753 <= not w8751 and not w8752;
w8754 <= w8747 and not w8753;
w8755 <= not w8744 and w8754;
w8756 <= not w8749 and not w8755;
w8757 <= not b(34) and not w8756;
w8758 <= not w8288 and not w8748;
w8759 <= not w8298 and w8732;
w8760 <= not w8728 and w8759;
w8761 <= not w8729 and not w8732;
w8762 <= not w8760 and not w8761;
w8763 <= w8747 and not w8762;
w8764 <= not w8744 and w8763;
w8765 <= not w8758 and not w8764;
w8766 <= not b(33) and not w8765;
w8767 <= not w8297 and not w8748;
w8768 <= not w8307 and w8727;
w8769 <= not w8723 and w8768;
w8770 <= not w8724 and not w8727;
w8771 <= not w8769 and not w8770;
w8772 <= w8747 and not w8771;
w8773 <= not w8744 and w8772;
w8774 <= not w8767 and not w8773;
w8775 <= not b(32) and not w8774;
w8776 <= not w8306 and not w8748;
w8777 <= not w8316 and w8722;
w8778 <= not w8718 and w8777;
w8779 <= not w8719 and not w8722;
w8780 <= not w8778 and not w8779;
w8781 <= w8747 and not w8780;
w8782 <= not w8744 and w8781;
w8783 <= not w8776 and not w8782;
w8784 <= not b(31) and not w8783;
w8785 <= not w8315 and not w8748;
w8786 <= not w8325 and w8717;
w8787 <= not w8713 and w8786;
w8788 <= not w8714 and not w8717;
w8789 <= not w8787 and not w8788;
w8790 <= w8747 and not w8789;
w8791 <= not w8744 and w8790;
w8792 <= not w8785 and not w8791;
w8793 <= not b(30) and not w8792;
w8794 <= not w8324 and not w8748;
w8795 <= not w8334 and w8712;
w8796 <= not w8708 and w8795;
w8797 <= not w8709 and not w8712;
w8798 <= not w8796 and not w8797;
w8799 <= w8747 and not w8798;
w8800 <= not w8744 and w8799;
w8801 <= not w8794 and not w8800;
w8802 <= not b(29) and not w8801;
w8803 <= not w8333 and not w8748;
w8804 <= not w8343 and w8707;
w8805 <= not w8703 and w8804;
w8806 <= not w8704 and not w8707;
w8807 <= not w8805 and not w8806;
w8808 <= w8747 and not w8807;
w8809 <= not w8744 and w8808;
w8810 <= not w8803 and not w8809;
w8811 <= not b(28) and not w8810;
w8812 <= not w8342 and not w8748;
w8813 <= not w8352 and w8702;
w8814 <= not w8698 and w8813;
w8815 <= not w8699 and not w8702;
w8816 <= not w8814 and not w8815;
w8817 <= w8747 and not w8816;
w8818 <= not w8744 and w8817;
w8819 <= not w8812 and not w8818;
w8820 <= not b(27) and not w8819;
w8821 <= not w8351 and not w8748;
w8822 <= not w8361 and w8697;
w8823 <= not w8693 and w8822;
w8824 <= not w8694 and not w8697;
w8825 <= not w8823 and not w8824;
w8826 <= w8747 and not w8825;
w8827 <= not w8744 and w8826;
w8828 <= not w8821 and not w8827;
w8829 <= not b(26) and not w8828;
w8830 <= not w8360 and not w8748;
w8831 <= not w8370 and w8692;
w8832 <= not w8688 and w8831;
w8833 <= not w8689 and not w8692;
w8834 <= not w8832 and not w8833;
w8835 <= w8747 and not w8834;
w8836 <= not w8744 and w8835;
w8837 <= not w8830 and not w8836;
w8838 <= not b(25) and not w8837;
w8839 <= not w8369 and not w8748;
w8840 <= not w8379 and w8687;
w8841 <= not w8683 and w8840;
w8842 <= not w8684 and not w8687;
w8843 <= not w8841 and not w8842;
w8844 <= w8747 and not w8843;
w8845 <= not w8744 and w8844;
w8846 <= not w8839 and not w8845;
w8847 <= not b(24) and not w8846;
w8848 <= not w8378 and not w8748;
w8849 <= not w8388 and w8682;
w8850 <= not w8678 and w8849;
w8851 <= not w8679 and not w8682;
w8852 <= not w8850 and not w8851;
w8853 <= w8747 and not w8852;
w8854 <= not w8744 and w8853;
w8855 <= not w8848 and not w8854;
w8856 <= not b(23) and not w8855;
w8857 <= not w8387 and not w8748;
w8858 <= not w8397 and w8677;
w8859 <= not w8673 and w8858;
w8860 <= not w8674 and not w8677;
w8861 <= not w8859 and not w8860;
w8862 <= w8747 and not w8861;
w8863 <= not w8744 and w8862;
w8864 <= not w8857 and not w8863;
w8865 <= not b(22) and not w8864;
w8866 <= not w8396 and not w8748;
w8867 <= not w8406 and w8672;
w8868 <= not w8668 and w8867;
w8869 <= not w8669 and not w8672;
w8870 <= not w8868 and not w8869;
w8871 <= w8747 and not w8870;
w8872 <= not w8744 and w8871;
w8873 <= not w8866 and not w8872;
w8874 <= not b(21) and not w8873;
w8875 <= not w8405 and not w8748;
w8876 <= not w8415 and w8667;
w8877 <= not w8663 and w8876;
w8878 <= not w8664 and not w8667;
w8879 <= not w8877 and not w8878;
w8880 <= w8747 and not w8879;
w8881 <= not w8744 and w8880;
w8882 <= not w8875 and not w8881;
w8883 <= not b(20) and not w8882;
w8884 <= not w8414 and not w8748;
w8885 <= not w8424 and w8662;
w8886 <= not w8658 and w8885;
w8887 <= not w8659 and not w8662;
w8888 <= not w8886 and not w8887;
w8889 <= w8747 and not w8888;
w8890 <= not w8744 and w8889;
w8891 <= not w8884 and not w8890;
w8892 <= not b(19) and not w8891;
w8893 <= not w8423 and not w8748;
w8894 <= not w8433 and w8657;
w8895 <= not w8653 and w8894;
w8896 <= not w8654 and not w8657;
w8897 <= not w8895 and not w8896;
w8898 <= w8747 and not w8897;
w8899 <= not w8744 and w8898;
w8900 <= not w8893 and not w8899;
w8901 <= not b(18) and not w8900;
w8902 <= not w8432 and not w8748;
w8903 <= not w8442 and w8652;
w8904 <= not w8648 and w8903;
w8905 <= not w8649 and not w8652;
w8906 <= not w8904 and not w8905;
w8907 <= w8747 and not w8906;
w8908 <= not w8744 and w8907;
w8909 <= not w8902 and not w8908;
w8910 <= not b(17) and not w8909;
w8911 <= not w8441 and not w8748;
w8912 <= not w8451 and w8647;
w8913 <= not w8643 and w8912;
w8914 <= not w8644 and not w8647;
w8915 <= not w8913 and not w8914;
w8916 <= w8747 and not w8915;
w8917 <= not w8744 and w8916;
w8918 <= not w8911 and not w8917;
w8919 <= not b(16) and not w8918;
w8920 <= not w8450 and not w8748;
w8921 <= not w8460 and w8642;
w8922 <= not w8638 and w8921;
w8923 <= not w8639 and not w8642;
w8924 <= not w8922 and not w8923;
w8925 <= w8747 and not w8924;
w8926 <= not w8744 and w8925;
w8927 <= not w8920 and not w8926;
w8928 <= not b(15) and not w8927;
w8929 <= not w8459 and not w8748;
w8930 <= not w8469 and w8637;
w8931 <= not w8633 and w8930;
w8932 <= not w8634 and not w8637;
w8933 <= not w8931 and not w8932;
w8934 <= w8747 and not w8933;
w8935 <= not w8744 and w8934;
w8936 <= not w8929 and not w8935;
w8937 <= not b(14) and not w8936;
w8938 <= not w8468 and not w8748;
w8939 <= not w8478 and w8632;
w8940 <= not w8628 and w8939;
w8941 <= not w8629 and not w8632;
w8942 <= not w8940 and not w8941;
w8943 <= w8747 and not w8942;
w8944 <= not w8744 and w8943;
w8945 <= not w8938 and not w8944;
w8946 <= not b(13) and not w8945;
w8947 <= not w8477 and not w8748;
w8948 <= not w8487 and w8627;
w8949 <= not w8623 and w8948;
w8950 <= not w8624 and not w8627;
w8951 <= not w8949 and not w8950;
w8952 <= w8747 and not w8951;
w8953 <= not w8744 and w8952;
w8954 <= not w8947 and not w8953;
w8955 <= not b(12) and not w8954;
w8956 <= not w8486 and not w8748;
w8957 <= not w8496 and w8622;
w8958 <= not w8618 and w8957;
w8959 <= not w8619 and not w8622;
w8960 <= not w8958 and not w8959;
w8961 <= w8747 and not w8960;
w8962 <= not w8744 and w8961;
w8963 <= not w8956 and not w8962;
w8964 <= not b(11) and not w8963;
w8965 <= not w8495 and not w8748;
w8966 <= not w8505 and w8617;
w8967 <= not w8613 and w8966;
w8968 <= not w8614 and not w8617;
w8969 <= not w8967 and not w8968;
w8970 <= w8747 and not w8969;
w8971 <= not w8744 and w8970;
w8972 <= not w8965 and not w8971;
w8973 <= not b(10) and not w8972;
w8974 <= not w8504 and not w8748;
w8975 <= not w8514 and w8612;
w8976 <= not w8608 and w8975;
w8977 <= not w8609 and not w8612;
w8978 <= not w8976 and not w8977;
w8979 <= w8747 and not w8978;
w8980 <= not w8744 and w8979;
w8981 <= not w8974 and not w8980;
w8982 <= not b(9) and not w8981;
w8983 <= not w8513 and not w8748;
w8984 <= not w8523 and w8607;
w8985 <= not w8603 and w8984;
w8986 <= not w8604 and not w8607;
w8987 <= not w8985 and not w8986;
w8988 <= w8747 and not w8987;
w8989 <= not w8744 and w8988;
w8990 <= not w8983 and not w8989;
w8991 <= not b(8) and not w8990;
w8992 <= not w8522 and not w8748;
w8993 <= not w8532 and w8602;
w8994 <= not w8598 and w8993;
w8995 <= not w8599 and not w8602;
w8996 <= not w8994 and not w8995;
w8997 <= w8747 and not w8996;
w8998 <= not w8744 and w8997;
w8999 <= not w8992 and not w8998;
w9000 <= not b(7) and not w8999;
w9001 <= not w8531 and not w8748;
w9002 <= not w8541 and w8597;
w9003 <= not w8593 and w9002;
w9004 <= not w8594 and not w8597;
w9005 <= not w9003 and not w9004;
w9006 <= w8747 and not w9005;
w9007 <= not w8744 and w9006;
w9008 <= not w9001 and not w9007;
w9009 <= not b(6) and not w9008;
w9010 <= not w8540 and not w8748;
w9011 <= not w8550 and w8592;
w9012 <= not w8588 and w9011;
w9013 <= not w8589 and not w8592;
w9014 <= not w9012 and not w9013;
w9015 <= w8747 and not w9014;
w9016 <= not w8744 and w9015;
w9017 <= not w9010 and not w9016;
w9018 <= not b(5) and not w9017;
w9019 <= not w8549 and not w8748;
w9020 <= not w8558 and w8587;
w9021 <= not w8583 and w9020;
w9022 <= not w8584 and not w8587;
w9023 <= not w9021 and not w9022;
w9024 <= w8747 and not w9023;
w9025 <= not w8744 and w9024;
w9026 <= not w9019 and not w9025;
w9027 <= not b(4) and not w9026;
w9028 <= not w8557 and not w8748;
w9029 <= not w8578 and w8582;
w9030 <= not w8577 and w9029;
w9031 <= not w8579 and not w8582;
w9032 <= not w9030 and not w9031;
w9033 <= w8747 and not w9032;
w9034 <= not w8744 and w9033;
w9035 <= not w9028 and not w9034;
w9036 <= not b(3) and not w9035;
w9037 <= not w8571 and not w8748;
w9038 <= not w8574 and w8576;
w9039 <= not w8572 and w9038;
w9040 <= w8747 and not w9039;
w9041 <= not w8577 and w9040;
w9042 <= not w8744 and w9041;
w9043 <= not w9037 and not w9042;
w9044 <= not b(2) and not w9043;
w9045 <= b(0) and not b(35);
w9046 <= w37 and w9045;
w9047 <= w83 and w9046;
w9048 <= w81 and w9047;
w9049 <= not w8744 and w9048;
w9050 <= a(29) and not w9049;
w9051 <= w156 and w8576;
w9052 <= w154 and w9051;
w9053 <= w165 and w9052;
w9054 <= w151 and w9053;
w9055 <= not w8744 and w9054;
w9056 <= not w9050 and not w9055;
w9057 <= b(1) and not w9056;
w9058 <= not b(1) and not w9055;
w9059 <= not w9050 and w9058;
w9060 <= not w9057 and not w9059;
w9061 <= not a(28) and b(0);
w9062 <= not w9060 and not w9061;
w9063 <= not b(1) and not w9056;
w9064 <= not w9062 and not w9063;
w9065 <= b(2) and not w9042;
w9066 <= not w9037 and w9065;
w9067 <= not w9044 and not w9066;
w9068 <= not w9064 and w9067;
w9069 <= not w9044 and not w9068;
w9070 <= b(3) and not w9034;
w9071 <= not w9028 and w9070;
w9072 <= not w9036 and not w9071;
w9073 <= not w9069 and w9072;
w9074 <= not w9036 and not w9073;
w9075 <= b(4) and not w9025;
w9076 <= not w9019 and w9075;
w9077 <= not w9027 and not w9076;
w9078 <= not w9074 and w9077;
w9079 <= not w9027 and not w9078;
w9080 <= b(5) and not w9016;
w9081 <= not w9010 and w9080;
w9082 <= not w9018 and not w9081;
w9083 <= not w9079 and w9082;
w9084 <= not w9018 and not w9083;
w9085 <= b(6) and not w9007;
w9086 <= not w9001 and w9085;
w9087 <= not w9009 and not w9086;
w9088 <= not w9084 and w9087;
w9089 <= not w9009 and not w9088;
w9090 <= b(7) and not w8998;
w9091 <= not w8992 and w9090;
w9092 <= not w9000 and not w9091;
w9093 <= not w9089 and w9092;
w9094 <= not w9000 and not w9093;
w9095 <= b(8) and not w8989;
w9096 <= not w8983 and w9095;
w9097 <= not w8991 and not w9096;
w9098 <= not w9094 and w9097;
w9099 <= not w8991 and not w9098;
w9100 <= b(9) and not w8980;
w9101 <= not w8974 and w9100;
w9102 <= not w8982 and not w9101;
w9103 <= not w9099 and w9102;
w9104 <= not w8982 and not w9103;
w9105 <= b(10) and not w8971;
w9106 <= not w8965 and w9105;
w9107 <= not w8973 and not w9106;
w9108 <= not w9104 and w9107;
w9109 <= not w8973 and not w9108;
w9110 <= b(11) and not w8962;
w9111 <= not w8956 and w9110;
w9112 <= not w8964 and not w9111;
w9113 <= not w9109 and w9112;
w9114 <= not w8964 and not w9113;
w9115 <= b(12) and not w8953;
w9116 <= not w8947 and w9115;
w9117 <= not w8955 and not w9116;
w9118 <= not w9114 and w9117;
w9119 <= not w8955 and not w9118;
w9120 <= b(13) and not w8944;
w9121 <= not w8938 and w9120;
w9122 <= not w8946 and not w9121;
w9123 <= not w9119 and w9122;
w9124 <= not w8946 and not w9123;
w9125 <= b(14) and not w8935;
w9126 <= not w8929 and w9125;
w9127 <= not w8937 and not w9126;
w9128 <= not w9124 and w9127;
w9129 <= not w8937 and not w9128;
w9130 <= b(15) and not w8926;
w9131 <= not w8920 and w9130;
w9132 <= not w8928 and not w9131;
w9133 <= not w9129 and w9132;
w9134 <= not w8928 and not w9133;
w9135 <= b(16) and not w8917;
w9136 <= not w8911 and w9135;
w9137 <= not w8919 and not w9136;
w9138 <= not w9134 and w9137;
w9139 <= not w8919 and not w9138;
w9140 <= b(17) and not w8908;
w9141 <= not w8902 and w9140;
w9142 <= not w8910 and not w9141;
w9143 <= not w9139 and w9142;
w9144 <= not w8910 and not w9143;
w9145 <= b(18) and not w8899;
w9146 <= not w8893 and w9145;
w9147 <= not w8901 and not w9146;
w9148 <= not w9144 and w9147;
w9149 <= not w8901 and not w9148;
w9150 <= b(19) and not w8890;
w9151 <= not w8884 and w9150;
w9152 <= not w8892 and not w9151;
w9153 <= not w9149 and w9152;
w9154 <= not w8892 and not w9153;
w9155 <= b(20) and not w8881;
w9156 <= not w8875 and w9155;
w9157 <= not w8883 and not w9156;
w9158 <= not w9154 and w9157;
w9159 <= not w8883 and not w9158;
w9160 <= b(21) and not w8872;
w9161 <= not w8866 and w9160;
w9162 <= not w8874 and not w9161;
w9163 <= not w9159 and w9162;
w9164 <= not w8874 and not w9163;
w9165 <= b(22) and not w8863;
w9166 <= not w8857 and w9165;
w9167 <= not w8865 and not w9166;
w9168 <= not w9164 and w9167;
w9169 <= not w8865 and not w9168;
w9170 <= b(23) and not w8854;
w9171 <= not w8848 and w9170;
w9172 <= not w8856 and not w9171;
w9173 <= not w9169 and w9172;
w9174 <= not w8856 and not w9173;
w9175 <= b(24) and not w8845;
w9176 <= not w8839 and w9175;
w9177 <= not w8847 and not w9176;
w9178 <= not w9174 and w9177;
w9179 <= not w8847 and not w9178;
w9180 <= b(25) and not w8836;
w9181 <= not w8830 and w9180;
w9182 <= not w8838 and not w9181;
w9183 <= not w9179 and w9182;
w9184 <= not w8838 and not w9183;
w9185 <= b(26) and not w8827;
w9186 <= not w8821 and w9185;
w9187 <= not w8829 and not w9186;
w9188 <= not w9184 and w9187;
w9189 <= not w8829 and not w9188;
w9190 <= b(27) and not w8818;
w9191 <= not w8812 and w9190;
w9192 <= not w8820 and not w9191;
w9193 <= not w9189 and w9192;
w9194 <= not w8820 and not w9193;
w9195 <= b(28) and not w8809;
w9196 <= not w8803 and w9195;
w9197 <= not w8811 and not w9196;
w9198 <= not w9194 and w9197;
w9199 <= not w8811 and not w9198;
w9200 <= b(29) and not w8800;
w9201 <= not w8794 and w9200;
w9202 <= not w8802 and not w9201;
w9203 <= not w9199 and w9202;
w9204 <= not w8802 and not w9203;
w9205 <= b(30) and not w8791;
w9206 <= not w8785 and w9205;
w9207 <= not w8793 and not w9206;
w9208 <= not w9204 and w9207;
w9209 <= not w8793 and not w9208;
w9210 <= b(31) and not w8782;
w9211 <= not w8776 and w9210;
w9212 <= not w8784 and not w9211;
w9213 <= not w9209 and w9212;
w9214 <= not w8784 and not w9213;
w9215 <= b(32) and not w8773;
w9216 <= not w8767 and w9215;
w9217 <= not w8775 and not w9216;
w9218 <= not w9214 and w9217;
w9219 <= not w8775 and not w9218;
w9220 <= b(33) and not w8764;
w9221 <= not w8758 and w9220;
w9222 <= not w8766 and not w9221;
w9223 <= not w9219 and w9222;
w9224 <= not w8766 and not w9223;
w9225 <= b(34) and not w8755;
w9226 <= not w8749 and w9225;
w9227 <= not w8757 and not w9226;
w9228 <= not w9224 and w9227;
w9229 <= not w8757 and not w9228;
w9230 <= not w8278 and not w8748;
w9231 <= not w8280 and w8742;
w9232 <= not w8738 and w9231;
w9233 <= not w8739 and not w8742;
w9234 <= not w9232 and not w9233;
w9235 <= w8748 and not w9234;
w9236 <= not w9230 and not w9235;
w9237 <= not b(35) and not w9236;
w9238 <= b(35) and not w9230;
w9239 <= not w9235 and w9238;
w9240 <= w255 and not w9239;
w9241 <= not w9237 and w9240;
w9242 <= not w9229 and w9241;
w9243 <= w8747 and not w9236;
w9244 <= not w9242 and not w9243;
w9245 <= not w8766 and w9227;
w9246 <= not w9223 and w9245;
w9247 <= not w9224 and not w9227;
w9248 <= not w9246 and not w9247;
w9249 <= not w9244 and not w9248;
w9250 <= not w8756 and not w9243;
w9251 <= not w9242 and w9250;
w9252 <= not w9249 and not w9251;
w9253 <= not w8757 and not w9239;
w9254 <= not w9237 and w9253;
w9255 <= not w9228 and w9254;
w9256 <= not w9237 and not w9239;
w9257 <= not w9229 and not w9256;
w9258 <= not w9255 and not w9257;
w9259 <= not w9244 and not w9258;
w9260 <= not w9236 and not w9243;
w9261 <= not w9242 and w9260;
w9262 <= not w9259 and not w9261;
w9263 <= not b(36) and not w9262;
w9264 <= not b(35) and not w9252;
w9265 <= not w8775 and w9222;
w9266 <= not w9218 and w9265;
w9267 <= not w9219 and not w9222;
w9268 <= not w9266 and not w9267;
w9269 <= not w9244 and not w9268;
w9270 <= not w8765 and not w9243;
w9271 <= not w9242 and w9270;
w9272 <= not w9269 and not w9271;
w9273 <= not b(34) and not w9272;
w9274 <= not w8784 and w9217;
w9275 <= not w9213 and w9274;
w9276 <= not w9214 and not w9217;
w9277 <= not w9275 and not w9276;
w9278 <= not w9244 and not w9277;
w9279 <= not w8774 and not w9243;
w9280 <= not w9242 and w9279;
w9281 <= not w9278 and not w9280;
w9282 <= not b(33) and not w9281;
w9283 <= not w8793 and w9212;
w9284 <= not w9208 and w9283;
w9285 <= not w9209 and not w9212;
w9286 <= not w9284 and not w9285;
w9287 <= not w9244 and not w9286;
w9288 <= not w8783 and not w9243;
w9289 <= not w9242 and w9288;
w9290 <= not w9287 and not w9289;
w9291 <= not b(32) and not w9290;
w9292 <= not w8802 and w9207;
w9293 <= not w9203 and w9292;
w9294 <= not w9204 and not w9207;
w9295 <= not w9293 and not w9294;
w9296 <= not w9244 and not w9295;
w9297 <= not w8792 and not w9243;
w9298 <= not w9242 and w9297;
w9299 <= not w9296 and not w9298;
w9300 <= not b(31) and not w9299;
w9301 <= not w8811 and w9202;
w9302 <= not w9198 and w9301;
w9303 <= not w9199 and not w9202;
w9304 <= not w9302 and not w9303;
w9305 <= not w9244 and not w9304;
w9306 <= not w8801 and not w9243;
w9307 <= not w9242 and w9306;
w9308 <= not w9305 and not w9307;
w9309 <= not b(30) and not w9308;
w9310 <= not w8820 and w9197;
w9311 <= not w9193 and w9310;
w9312 <= not w9194 and not w9197;
w9313 <= not w9311 and not w9312;
w9314 <= not w9244 and not w9313;
w9315 <= not w8810 and not w9243;
w9316 <= not w9242 and w9315;
w9317 <= not w9314 and not w9316;
w9318 <= not b(29) and not w9317;
w9319 <= not w8829 and w9192;
w9320 <= not w9188 and w9319;
w9321 <= not w9189 and not w9192;
w9322 <= not w9320 and not w9321;
w9323 <= not w9244 and not w9322;
w9324 <= not w8819 and not w9243;
w9325 <= not w9242 and w9324;
w9326 <= not w9323 and not w9325;
w9327 <= not b(28) and not w9326;
w9328 <= not w8838 and w9187;
w9329 <= not w9183 and w9328;
w9330 <= not w9184 and not w9187;
w9331 <= not w9329 and not w9330;
w9332 <= not w9244 and not w9331;
w9333 <= not w8828 and not w9243;
w9334 <= not w9242 and w9333;
w9335 <= not w9332 and not w9334;
w9336 <= not b(27) and not w9335;
w9337 <= not w8847 and w9182;
w9338 <= not w9178 and w9337;
w9339 <= not w9179 and not w9182;
w9340 <= not w9338 and not w9339;
w9341 <= not w9244 and not w9340;
w9342 <= not w8837 and not w9243;
w9343 <= not w9242 and w9342;
w9344 <= not w9341 and not w9343;
w9345 <= not b(26) and not w9344;
w9346 <= not w8856 and w9177;
w9347 <= not w9173 and w9346;
w9348 <= not w9174 and not w9177;
w9349 <= not w9347 and not w9348;
w9350 <= not w9244 and not w9349;
w9351 <= not w8846 and not w9243;
w9352 <= not w9242 and w9351;
w9353 <= not w9350 and not w9352;
w9354 <= not b(25) and not w9353;
w9355 <= not w8865 and w9172;
w9356 <= not w9168 and w9355;
w9357 <= not w9169 and not w9172;
w9358 <= not w9356 and not w9357;
w9359 <= not w9244 and not w9358;
w9360 <= not w8855 and not w9243;
w9361 <= not w9242 and w9360;
w9362 <= not w9359 and not w9361;
w9363 <= not b(24) and not w9362;
w9364 <= not w8874 and w9167;
w9365 <= not w9163 and w9364;
w9366 <= not w9164 and not w9167;
w9367 <= not w9365 and not w9366;
w9368 <= not w9244 and not w9367;
w9369 <= not w8864 and not w9243;
w9370 <= not w9242 and w9369;
w9371 <= not w9368 and not w9370;
w9372 <= not b(23) and not w9371;
w9373 <= not w8883 and w9162;
w9374 <= not w9158 and w9373;
w9375 <= not w9159 and not w9162;
w9376 <= not w9374 and not w9375;
w9377 <= not w9244 and not w9376;
w9378 <= not w8873 and not w9243;
w9379 <= not w9242 and w9378;
w9380 <= not w9377 and not w9379;
w9381 <= not b(22) and not w9380;
w9382 <= not w8892 and w9157;
w9383 <= not w9153 and w9382;
w9384 <= not w9154 and not w9157;
w9385 <= not w9383 and not w9384;
w9386 <= not w9244 and not w9385;
w9387 <= not w8882 and not w9243;
w9388 <= not w9242 and w9387;
w9389 <= not w9386 and not w9388;
w9390 <= not b(21) and not w9389;
w9391 <= not w8901 and w9152;
w9392 <= not w9148 and w9391;
w9393 <= not w9149 and not w9152;
w9394 <= not w9392 and not w9393;
w9395 <= not w9244 and not w9394;
w9396 <= not w8891 and not w9243;
w9397 <= not w9242 and w9396;
w9398 <= not w9395 and not w9397;
w9399 <= not b(20) and not w9398;
w9400 <= not w8910 and w9147;
w9401 <= not w9143 and w9400;
w9402 <= not w9144 and not w9147;
w9403 <= not w9401 and not w9402;
w9404 <= not w9244 and not w9403;
w9405 <= not w8900 and not w9243;
w9406 <= not w9242 and w9405;
w9407 <= not w9404 and not w9406;
w9408 <= not b(19) and not w9407;
w9409 <= not w8919 and w9142;
w9410 <= not w9138 and w9409;
w9411 <= not w9139 and not w9142;
w9412 <= not w9410 and not w9411;
w9413 <= not w9244 and not w9412;
w9414 <= not w8909 and not w9243;
w9415 <= not w9242 and w9414;
w9416 <= not w9413 and not w9415;
w9417 <= not b(18) and not w9416;
w9418 <= not w8928 and w9137;
w9419 <= not w9133 and w9418;
w9420 <= not w9134 and not w9137;
w9421 <= not w9419 and not w9420;
w9422 <= not w9244 and not w9421;
w9423 <= not w8918 and not w9243;
w9424 <= not w9242 and w9423;
w9425 <= not w9422 and not w9424;
w9426 <= not b(17) and not w9425;
w9427 <= not w8937 and w9132;
w9428 <= not w9128 and w9427;
w9429 <= not w9129 and not w9132;
w9430 <= not w9428 and not w9429;
w9431 <= not w9244 and not w9430;
w9432 <= not w8927 and not w9243;
w9433 <= not w9242 and w9432;
w9434 <= not w9431 and not w9433;
w9435 <= not b(16) and not w9434;
w9436 <= not w8946 and w9127;
w9437 <= not w9123 and w9436;
w9438 <= not w9124 and not w9127;
w9439 <= not w9437 and not w9438;
w9440 <= not w9244 and not w9439;
w9441 <= not w8936 and not w9243;
w9442 <= not w9242 and w9441;
w9443 <= not w9440 and not w9442;
w9444 <= not b(15) and not w9443;
w9445 <= not w8955 and w9122;
w9446 <= not w9118 and w9445;
w9447 <= not w9119 and not w9122;
w9448 <= not w9446 and not w9447;
w9449 <= not w9244 and not w9448;
w9450 <= not w8945 and not w9243;
w9451 <= not w9242 and w9450;
w9452 <= not w9449 and not w9451;
w9453 <= not b(14) and not w9452;
w9454 <= not w8964 and w9117;
w9455 <= not w9113 and w9454;
w9456 <= not w9114 and not w9117;
w9457 <= not w9455 and not w9456;
w9458 <= not w9244 and not w9457;
w9459 <= not w8954 and not w9243;
w9460 <= not w9242 and w9459;
w9461 <= not w9458 and not w9460;
w9462 <= not b(13) and not w9461;
w9463 <= not w8973 and w9112;
w9464 <= not w9108 and w9463;
w9465 <= not w9109 and not w9112;
w9466 <= not w9464 and not w9465;
w9467 <= not w9244 and not w9466;
w9468 <= not w8963 and not w9243;
w9469 <= not w9242 and w9468;
w9470 <= not w9467 and not w9469;
w9471 <= not b(12) and not w9470;
w9472 <= not w8982 and w9107;
w9473 <= not w9103 and w9472;
w9474 <= not w9104 and not w9107;
w9475 <= not w9473 and not w9474;
w9476 <= not w9244 and not w9475;
w9477 <= not w8972 and not w9243;
w9478 <= not w9242 and w9477;
w9479 <= not w9476 and not w9478;
w9480 <= not b(11) and not w9479;
w9481 <= not w8991 and w9102;
w9482 <= not w9098 and w9481;
w9483 <= not w9099 and not w9102;
w9484 <= not w9482 and not w9483;
w9485 <= not w9244 and not w9484;
w9486 <= not w8981 and not w9243;
w9487 <= not w9242 and w9486;
w9488 <= not w9485 and not w9487;
w9489 <= not b(10) and not w9488;
w9490 <= not w9000 and w9097;
w9491 <= not w9093 and w9490;
w9492 <= not w9094 and not w9097;
w9493 <= not w9491 and not w9492;
w9494 <= not w9244 and not w9493;
w9495 <= not w8990 and not w9243;
w9496 <= not w9242 and w9495;
w9497 <= not w9494 and not w9496;
w9498 <= not b(9) and not w9497;
w9499 <= not w9009 and w9092;
w9500 <= not w9088 and w9499;
w9501 <= not w9089 and not w9092;
w9502 <= not w9500 and not w9501;
w9503 <= not w9244 and not w9502;
w9504 <= not w8999 and not w9243;
w9505 <= not w9242 and w9504;
w9506 <= not w9503 and not w9505;
w9507 <= not b(8) and not w9506;
w9508 <= not w9018 and w9087;
w9509 <= not w9083 and w9508;
w9510 <= not w9084 and not w9087;
w9511 <= not w9509 and not w9510;
w9512 <= not w9244 and not w9511;
w9513 <= not w9008 and not w9243;
w9514 <= not w9242 and w9513;
w9515 <= not w9512 and not w9514;
w9516 <= not b(7) and not w9515;
w9517 <= not w9027 and w9082;
w9518 <= not w9078 and w9517;
w9519 <= not w9079 and not w9082;
w9520 <= not w9518 and not w9519;
w9521 <= not w9244 and not w9520;
w9522 <= not w9017 and not w9243;
w9523 <= not w9242 and w9522;
w9524 <= not w9521 and not w9523;
w9525 <= not b(6) and not w9524;
w9526 <= not w9036 and w9077;
w9527 <= not w9073 and w9526;
w9528 <= not w9074 and not w9077;
w9529 <= not w9527 and not w9528;
w9530 <= not w9244 and not w9529;
w9531 <= not w9026 and not w9243;
w9532 <= not w9242 and w9531;
w9533 <= not w9530 and not w9532;
w9534 <= not b(5) and not w9533;
w9535 <= not w9044 and w9072;
w9536 <= not w9068 and w9535;
w9537 <= not w9069 and not w9072;
w9538 <= not w9536 and not w9537;
w9539 <= not w9244 and not w9538;
w9540 <= not w9035 and not w9243;
w9541 <= not w9242 and w9540;
w9542 <= not w9539 and not w9541;
w9543 <= not b(4) and not w9542;
w9544 <= not w9063 and w9067;
w9545 <= not w9062 and w9544;
w9546 <= not w9064 and not w9067;
w9547 <= not w9545 and not w9546;
w9548 <= not w9244 and not w9547;
w9549 <= not w9043 and not w9243;
w9550 <= not w9242 and w9549;
w9551 <= not w9548 and not w9550;
w9552 <= not b(3) and not w9551;
w9553 <= not w9059 and w9061;
w9554 <= not w9057 and w9553;
w9555 <= not w9062 and not w9554;
w9556 <= not w9244 and w9555;
w9557 <= not w9056 and not w9243;
w9558 <= not w9242 and w9557;
w9559 <= not w9556 and not w9558;
w9560 <= not b(2) and not w9559;
w9561 <= b(0) and not w9244;
w9562 <= a(28) and not w9561;
w9563 <= w9061 and not w9244;
w9564 <= not w9562 and not w9563;
w9565 <= b(1) and not w9564;
w9566 <= not b(1) and not w9563;
w9567 <= not w9562 and w9566;
w9568 <= not w9565 and not w9567;
w9569 <= not a(27) and b(0);
w9570 <= not w9568 and not w9569;
w9571 <= not b(1) and not w9564;
w9572 <= not w9570 and not w9571;
w9573 <= b(2) and not w9558;
w9574 <= not w9556 and w9573;
w9575 <= not w9560 and not w9574;
w9576 <= not w9572 and w9575;
w9577 <= not w9560 and not w9576;
w9578 <= b(3) and not w9550;
w9579 <= not w9548 and w9578;
w9580 <= not w9552 and not w9579;
w9581 <= not w9577 and w9580;
w9582 <= not w9552 and not w9581;
w9583 <= b(4) and not w9541;
w9584 <= not w9539 and w9583;
w9585 <= not w9543 and not w9584;
w9586 <= not w9582 and w9585;
w9587 <= not w9543 and not w9586;
w9588 <= b(5) and not w9532;
w9589 <= not w9530 and w9588;
w9590 <= not w9534 and not w9589;
w9591 <= not w9587 and w9590;
w9592 <= not w9534 and not w9591;
w9593 <= b(6) and not w9523;
w9594 <= not w9521 and w9593;
w9595 <= not w9525 and not w9594;
w9596 <= not w9592 and w9595;
w9597 <= not w9525 and not w9596;
w9598 <= b(7) and not w9514;
w9599 <= not w9512 and w9598;
w9600 <= not w9516 and not w9599;
w9601 <= not w9597 and w9600;
w9602 <= not w9516 and not w9601;
w9603 <= b(8) and not w9505;
w9604 <= not w9503 and w9603;
w9605 <= not w9507 and not w9604;
w9606 <= not w9602 and w9605;
w9607 <= not w9507 and not w9606;
w9608 <= b(9) and not w9496;
w9609 <= not w9494 and w9608;
w9610 <= not w9498 and not w9609;
w9611 <= not w9607 and w9610;
w9612 <= not w9498 and not w9611;
w9613 <= b(10) and not w9487;
w9614 <= not w9485 and w9613;
w9615 <= not w9489 and not w9614;
w9616 <= not w9612 and w9615;
w9617 <= not w9489 and not w9616;
w9618 <= b(11) and not w9478;
w9619 <= not w9476 and w9618;
w9620 <= not w9480 and not w9619;
w9621 <= not w9617 and w9620;
w9622 <= not w9480 and not w9621;
w9623 <= b(12) and not w9469;
w9624 <= not w9467 and w9623;
w9625 <= not w9471 and not w9624;
w9626 <= not w9622 and w9625;
w9627 <= not w9471 and not w9626;
w9628 <= b(13) and not w9460;
w9629 <= not w9458 and w9628;
w9630 <= not w9462 and not w9629;
w9631 <= not w9627 and w9630;
w9632 <= not w9462 and not w9631;
w9633 <= b(14) and not w9451;
w9634 <= not w9449 and w9633;
w9635 <= not w9453 and not w9634;
w9636 <= not w9632 and w9635;
w9637 <= not w9453 and not w9636;
w9638 <= b(15) and not w9442;
w9639 <= not w9440 and w9638;
w9640 <= not w9444 and not w9639;
w9641 <= not w9637 and w9640;
w9642 <= not w9444 and not w9641;
w9643 <= b(16) and not w9433;
w9644 <= not w9431 and w9643;
w9645 <= not w9435 and not w9644;
w9646 <= not w9642 and w9645;
w9647 <= not w9435 and not w9646;
w9648 <= b(17) and not w9424;
w9649 <= not w9422 and w9648;
w9650 <= not w9426 and not w9649;
w9651 <= not w9647 and w9650;
w9652 <= not w9426 and not w9651;
w9653 <= b(18) and not w9415;
w9654 <= not w9413 and w9653;
w9655 <= not w9417 and not w9654;
w9656 <= not w9652 and w9655;
w9657 <= not w9417 and not w9656;
w9658 <= b(19) and not w9406;
w9659 <= not w9404 and w9658;
w9660 <= not w9408 and not w9659;
w9661 <= not w9657 and w9660;
w9662 <= not w9408 and not w9661;
w9663 <= b(20) and not w9397;
w9664 <= not w9395 and w9663;
w9665 <= not w9399 and not w9664;
w9666 <= not w9662 and w9665;
w9667 <= not w9399 and not w9666;
w9668 <= b(21) and not w9388;
w9669 <= not w9386 and w9668;
w9670 <= not w9390 and not w9669;
w9671 <= not w9667 and w9670;
w9672 <= not w9390 and not w9671;
w9673 <= b(22) and not w9379;
w9674 <= not w9377 and w9673;
w9675 <= not w9381 and not w9674;
w9676 <= not w9672 and w9675;
w9677 <= not w9381 and not w9676;
w9678 <= b(23) and not w9370;
w9679 <= not w9368 and w9678;
w9680 <= not w9372 and not w9679;
w9681 <= not w9677 and w9680;
w9682 <= not w9372 and not w9681;
w9683 <= b(24) and not w9361;
w9684 <= not w9359 and w9683;
w9685 <= not w9363 and not w9684;
w9686 <= not w9682 and w9685;
w9687 <= not w9363 and not w9686;
w9688 <= b(25) and not w9352;
w9689 <= not w9350 and w9688;
w9690 <= not w9354 and not w9689;
w9691 <= not w9687 and w9690;
w9692 <= not w9354 and not w9691;
w9693 <= b(26) and not w9343;
w9694 <= not w9341 and w9693;
w9695 <= not w9345 and not w9694;
w9696 <= not w9692 and w9695;
w9697 <= not w9345 and not w9696;
w9698 <= b(27) and not w9334;
w9699 <= not w9332 and w9698;
w9700 <= not w9336 and not w9699;
w9701 <= not w9697 and w9700;
w9702 <= not w9336 and not w9701;
w9703 <= b(28) and not w9325;
w9704 <= not w9323 and w9703;
w9705 <= not w9327 and not w9704;
w9706 <= not w9702 and w9705;
w9707 <= not w9327 and not w9706;
w9708 <= b(29) and not w9316;
w9709 <= not w9314 and w9708;
w9710 <= not w9318 and not w9709;
w9711 <= not w9707 and w9710;
w9712 <= not w9318 and not w9711;
w9713 <= b(30) and not w9307;
w9714 <= not w9305 and w9713;
w9715 <= not w9309 and not w9714;
w9716 <= not w9712 and w9715;
w9717 <= not w9309 and not w9716;
w9718 <= b(31) and not w9298;
w9719 <= not w9296 and w9718;
w9720 <= not w9300 and not w9719;
w9721 <= not w9717 and w9720;
w9722 <= not w9300 and not w9721;
w9723 <= b(32) and not w9289;
w9724 <= not w9287 and w9723;
w9725 <= not w9291 and not w9724;
w9726 <= not w9722 and w9725;
w9727 <= not w9291 and not w9726;
w9728 <= b(33) and not w9280;
w9729 <= not w9278 and w9728;
w9730 <= not w9282 and not w9729;
w9731 <= not w9727 and w9730;
w9732 <= not w9282 and not w9731;
w9733 <= b(34) and not w9271;
w9734 <= not w9269 and w9733;
w9735 <= not w9273 and not w9734;
w9736 <= not w9732 and w9735;
w9737 <= not w9273 and not w9736;
w9738 <= b(35) and not w9251;
w9739 <= not w9249 and w9738;
w9740 <= not w9264 and not w9739;
w9741 <= not w9737 and w9740;
w9742 <= not w9264 and not w9741;
w9743 <= b(36) and not w9261;
w9744 <= not w9259 and w9743;
w9745 <= not w9263 and not w9744;
w9746 <= not w9742 and w9745;
w9747 <= not w9263 and not w9746;
w9748 <= w342 and not w9747;
w9749 <= not w9252 and not w9748;
w9750 <= not w9273 and w9740;
w9751 <= not w9736 and w9750;
w9752 <= not w9737 and not w9740;
w9753 <= not w9751 and not w9752;
w9754 <= w342 and not w9753;
w9755 <= not w9747 and w9754;
w9756 <= not w9749 and not w9755;
w9757 <= not w9262 and not w9748;
w9758 <= not w9264 and w9745;
w9759 <= not w9741 and w9758;
w9760 <= not w9742 and not w9745;
w9761 <= not w9759 and not w9760;
w9762 <= w9748 and not w9761;
w9763 <= not w9757 and not w9762;
w9764 <= not b(37) and not w9763;
w9765 <= not b(36) and not w9756;
w9766 <= not w9272 and not w9748;
w9767 <= not w9282 and w9735;
w9768 <= not w9731 and w9767;
w9769 <= not w9732 and not w9735;
w9770 <= not w9768 and not w9769;
w9771 <= w342 and not w9770;
w9772 <= not w9747 and w9771;
w9773 <= not w9766 and not w9772;
w9774 <= not b(35) and not w9773;
w9775 <= not w9281 and not w9748;
w9776 <= not w9291 and w9730;
w9777 <= not w9726 and w9776;
w9778 <= not w9727 and not w9730;
w9779 <= not w9777 and not w9778;
w9780 <= w342 and not w9779;
w9781 <= not w9747 and w9780;
w9782 <= not w9775 and not w9781;
w9783 <= not b(34) and not w9782;
w9784 <= not w9290 and not w9748;
w9785 <= not w9300 and w9725;
w9786 <= not w9721 and w9785;
w9787 <= not w9722 and not w9725;
w9788 <= not w9786 and not w9787;
w9789 <= w342 and not w9788;
w9790 <= not w9747 and w9789;
w9791 <= not w9784 and not w9790;
w9792 <= not b(33) and not w9791;
w9793 <= not w9299 and not w9748;
w9794 <= not w9309 and w9720;
w9795 <= not w9716 and w9794;
w9796 <= not w9717 and not w9720;
w9797 <= not w9795 and not w9796;
w9798 <= w342 and not w9797;
w9799 <= not w9747 and w9798;
w9800 <= not w9793 and not w9799;
w9801 <= not b(32) and not w9800;
w9802 <= not w9308 and not w9748;
w9803 <= not w9318 and w9715;
w9804 <= not w9711 and w9803;
w9805 <= not w9712 and not w9715;
w9806 <= not w9804 and not w9805;
w9807 <= w342 and not w9806;
w9808 <= not w9747 and w9807;
w9809 <= not w9802 and not w9808;
w9810 <= not b(31) and not w9809;
w9811 <= not w9317 and not w9748;
w9812 <= not w9327 and w9710;
w9813 <= not w9706 and w9812;
w9814 <= not w9707 and not w9710;
w9815 <= not w9813 and not w9814;
w9816 <= w342 and not w9815;
w9817 <= not w9747 and w9816;
w9818 <= not w9811 and not w9817;
w9819 <= not b(30) and not w9818;
w9820 <= not w9326 and not w9748;
w9821 <= not w9336 and w9705;
w9822 <= not w9701 and w9821;
w9823 <= not w9702 and not w9705;
w9824 <= not w9822 and not w9823;
w9825 <= w342 and not w9824;
w9826 <= not w9747 and w9825;
w9827 <= not w9820 and not w9826;
w9828 <= not b(29) and not w9827;
w9829 <= not w9335 and not w9748;
w9830 <= not w9345 and w9700;
w9831 <= not w9696 and w9830;
w9832 <= not w9697 and not w9700;
w9833 <= not w9831 and not w9832;
w9834 <= w342 and not w9833;
w9835 <= not w9747 and w9834;
w9836 <= not w9829 and not w9835;
w9837 <= not b(28) and not w9836;
w9838 <= not w9344 and not w9748;
w9839 <= not w9354 and w9695;
w9840 <= not w9691 and w9839;
w9841 <= not w9692 and not w9695;
w9842 <= not w9840 and not w9841;
w9843 <= w342 and not w9842;
w9844 <= not w9747 and w9843;
w9845 <= not w9838 and not w9844;
w9846 <= not b(27) and not w9845;
w9847 <= not w9353 and not w9748;
w9848 <= not w9363 and w9690;
w9849 <= not w9686 and w9848;
w9850 <= not w9687 and not w9690;
w9851 <= not w9849 and not w9850;
w9852 <= w342 and not w9851;
w9853 <= not w9747 and w9852;
w9854 <= not w9847 and not w9853;
w9855 <= not b(26) and not w9854;
w9856 <= not w9362 and not w9748;
w9857 <= not w9372 and w9685;
w9858 <= not w9681 and w9857;
w9859 <= not w9682 and not w9685;
w9860 <= not w9858 and not w9859;
w9861 <= w342 and not w9860;
w9862 <= not w9747 and w9861;
w9863 <= not w9856 and not w9862;
w9864 <= not b(25) and not w9863;
w9865 <= not w9371 and not w9748;
w9866 <= not w9381 and w9680;
w9867 <= not w9676 and w9866;
w9868 <= not w9677 and not w9680;
w9869 <= not w9867 and not w9868;
w9870 <= w342 and not w9869;
w9871 <= not w9747 and w9870;
w9872 <= not w9865 and not w9871;
w9873 <= not b(24) and not w9872;
w9874 <= not w9380 and not w9748;
w9875 <= not w9390 and w9675;
w9876 <= not w9671 and w9875;
w9877 <= not w9672 and not w9675;
w9878 <= not w9876 and not w9877;
w9879 <= w342 and not w9878;
w9880 <= not w9747 and w9879;
w9881 <= not w9874 and not w9880;
w9882 <= not b(23) and not w9881;
w9883 <= not w9389 and not w9748;
w9884 <= not w9399 and w9670;
w9885 <= not w9666 and w9884;
w9886 <= not w9667 and not w9670;
w9887 <= not w9885 and not w9886;
w9888 <= w342 and not w9887;
w9889 <= not w9747 and w9888;
w9890 <= not w9883 and not w9889;
w9891 <= not b(22) and not w9890;
w9892 <= not w9398 and not w9748;
w9893 <= not w9408 and w9665;
w9894 <= not w9661 and w9893;
w9895 <= not w9662 and not w9665;
w9896 <= not w9894 and not w9895;
w9897 <= w342 and not w9896;
w9898 <= not w9747 and w9897;
w9899 <= not w9892 and not w9898;
w9900 <= not b(21) and not w9899;
w9901 <= not w9407 and not w9748;
w9902 <= not w9417 and w9660;
w9903 <= not w9656 and w9902;
w9904 <= not w9657 and not w9660;
w9905 <= not w9903 and not w9904;
w9906 <= w342 and not w9905;
w9907 <= not w9747 and w9906;
w9908 <= not w9901 and not w9907;
w9909 <= not b(20) and not w9908;
w9910 <= not w9416 and not w9748;
w9911 <= not w9426 and w9655;
w9912 <= not w9651 and w9911;
w9913 <= not w9652 and not w9655;
w9914 <= not w9912 and not w9913;
w9915 <= w342 and not w9914;
w9916 <= not w9747 and w9915;
w9917 <= not w9910 and not w9916;
w9918 <= not b(19) and not w9917;
w9919 <= not w9425 and not w9748;
w9920 <= not w9435 and w9650;
w9921 <= not w9646 and w9920;
w9922 <= not w9647 and not w9650;
w9923 <= not w9921 and not w9922;
w9924 <= w342 and not w9923;
w9925 <= not w9747 and w9924;
w9926 <= not w9919 and not w9925;
w9927 <= not b(18) and not w9926;
w9928 <= not w9434 and not w9748;
w9929 <= not w9444 and w9645;
w9930 <= not w9641 and w9929;
w9931 <= not w9642 and not w9645;
w9932 <= not w9930 and not w9931;
w9933 <= w342 and not w9932;
w9934 <= not w9747 and w9933;
w9935 <= not w9928 and not w9934;
w9936 <= not b(17) and not w9935;
w9937 <= not w9443 and not w9748;
w9938 <= not w9453 and w9640;
w9939 <= not w9636 and w9938;
w9940 <= not w9637 and not w9640;
w9941 <= not w9939 and not w9940;
w9942 <= w342 and not w9941;
w9943 <= not w9747 and w9942;
w9944 <= not w9937 and not w9943;
w9945 <= not b(16) and not w9944;
w9946 <= not w9452 and not w9748;
w9947 <= not w9462 and w9635;
w9948 <= not w9631 and w9947;
w9949 <= not w9632 and not w9635;
w9950 <= not w9948 and not w9949;
w9951 <= w342 and not w9950;
w9952 <= not w9747 and w9951;
w9953 <= not w9946 and not w9952;
w9954 <= not b(15) and not w9953;
w9955 <= not w9461 and not w9748;
w9956 <= not w9471 and w9630;
w9957 <= not w9626 and w9956;
w9958 <= not w9627 and not w9630;
w9959 <= not w9957 and not w9958;
w9960 <= w342 and not w9959;
w9961 <= not w9747 and w9960;
w9962 <= not w9955 and not w9961;
w9963 <= not b(14) and not w9962;
w9964 <= not w9470 and not w9748;
w9965 <= not w9480 and w9625;
w9966 <= not w9621 and w9965;
w9967 <= not w9622 and not w9625;
w9968 <= not w9966 and not w9967;
w9969 <= w342 and not w9968;
w9970 <= not w9747 and w9969;
w9971 <= not w9964 and not w9970;
w9972 <= not b(13) and not w9971;
w9973 <= not w9479 and not w9748;
w9974 <= not w9489 and w9620;
w9975 <= not w9616 and w9974;
w9976 <= not w9617 and not w9620;
w9977 <= not w9975 and not w9976;
w9978 <= w342 and not w9977;
w9979 <= not w9747 and w9978;
w9980 <= not w9973 and not w9979;
w9981 <= not b(12) and not w9980;
w9982 <= not w9488 and not w9748;
w9983 <= not w9498 and w9615;
w9984 <= not w9611 and w9983;
w9985 <= not w9612 and not w9615;
w9986 <= not w9984 and not w9985;
w9987 <= w342 and not w9986;
w9988 <= not w9747 and w9987;
w9989 <= not w9982 and not w9988;
w9990 <= not b(11) and not w9989;
w9991 <= not w9497 and not w9748;
w9992 <= not w9507 and w9610;
w9993 <= not w9606 and w9992;
w9994 <= not w9607 and not w9610;
w9995 <= not w9993 and not w9994;
w9996 <= w342 and not w9995;
w9997 <= not w9747 and w9996;
w9998 <= not w9991 and not w9997;
w9999 <= not b(10) and not w9998;
w10000 <= not w9506 and not w9748;
w10001 <= not w9516 and w9605;
w10002 <= not w9601 and w10001;
w10003 <= not w9602 and not w9605;
w10004 <= not w10002 and not w10003;
w10005 <= w342 and not w10004;
w10006 <= not w9747 and w10005;
w10007 <= not w10000 and not w10006;
w10008 <= not b(9) and not w10007;
w10009 <= not w9515 and not w9748;
w10010 <= not w9525 and w9600;
w10011 <= not w9596 and w10010;
w10012 <= not w9597 and not w9600;
w10013 <= not w10011 and not w10012;
w10014 <= w342 and not w10013;
w10015 <= not w9747 and w10014;
w10016 <= not w10009 and not w10015;
w10017 <= not b(8) and not w10016;
w10018 <= not w9524 and not w9748;
w10019 <= not w9534 and w9595;
w10020 <= not w9591 and w10019;
w10021 <= not w9592 and not w9595;
w10022 <= not w10020 and not w10021;
w10023 <= w342 and not w10022;
w10024 <= not w9747 and w10023;
w10025 <= not w10018 and not w10024;
w10026 <= not b(7) and not w10025;
w10027 <= not w9533 and not w9748;
w10028 <= not w9543 and w9590;
w10029 <= not w9586 and w10028;
w10030 <= not w9587 and not w9590;
w10031 <= not w10029 and not w10030;
w10032 <= w342 and not w10031;
w10033 <= not w9747 and w10032;
w10034 <= not w10027 and not w10033;
w10035 <= not b(6) and not w10034;
w10036 <= not w9542 and not w9748;
w10037 <= not w9552 and w9585;
w10038 <= not w9581 and w10037;
w10039 <= not w9582 and not w9585;
w10040 <= not w10038 and not w10039;
w10041 <= w342 and not w10040;
w10042 <= not w9747 and w10041;
w10043 <= not w10036 and not w10042;
w10044 <= not b(5) and not w10043;
w10045 <= not w9551 and not w9748;
w10046 <= not w9560 and w9580;
w10047 <= not w9576 and w10046;
w10048 <= not w9577 and not w9580;
w10049 <= not w10047 and not w10048;
w10050 <= w342 and not w10049;
w10051 <= not w9747 and w10050;
w10052 <= not w10045 and not w10051;
w10053 <= not b(4) and not w10052;
w10054 <= not w9559 and not w9748;
w10055 <= not w9571 and w9575;
w10056 <= not w9570 and w10055;
w10057 <= not w9572 and not w9575;
w10058 <= not w10056 and not w10057;
w10059 <= w342 and not w10058;
w10060 <= not w9747 and w10059;
w10061 <= not w10054 and not w10060;
w10062 <= not b(3) and not w10061;
w10063 <= not w9564 and not w9748;
w10064 <= not w9567 and w9569;
w10065 <= not w9565 and w10064;
w10066 <= w342 and not w10065;
w10067 <= not w9570 and w10066;
w10068 <= not w9747 and w10067;
w10069 <= not w10063 and not w10068;
w10070 <= not b(2) and not w10069;
w10071 <= b(0) and not b(37);
w10072 <= w36 and w10071;
w10073 <= w34 and w10072;
w10074 <= w45 and w10073;
w10075 <= w31 and w10074;
w10076 <= not w9747 and w10075;
w10077 <= a(27) and not w10076;
w10078 <= w154 and w9569;
w10079 <= w165 and w10078;
w10080 <= w151 and w10079;
w10081 <= not w9747 and w10080;
w10082 <= not w10077 and not w10081;
w10083 <= b(1) and not w10082;
w10084 <= not b(1) and not w10081;
w10085 <= not w10077 and w10084;
w10086 <= not w10083 and not w10085;
w10087 <= not a(26) and b(0);
w10088 <= not w10086 and not w10087;
w10089 <= not b(1) and not w10082;
w10090 <= not w10088 and not w10089;
w10091 <= b(2) and not w10068;
w10092 <= not w10063 and w10091;
w10093 <= not w10070 and not w10092;
w10094 <= not w10090 and w10093;
w10095 <= not w10070 and not w10094;
w10096 <= b(3) and not w10060;
w10097 <= not w10054 and w10096;
w10098 <= not w10062 and not w10097;
w10099 <= not w10095 and w10098;
w10100 <= not w10062 and not w10099;
w10101 <= b(4) and not w10051;
w10102 <= not w10045 and w10101;
w10103 <= not w10053 and not w10102;
w10104 <= not w10100 and w10103;
w10105 <= not w10053 and not w10104;
w10106 <= b(5) and not w10042;
w10107 <= not w10036 and w10106;
w10108 <= not w10044 and not w10107;
w10109 <= not w10105 and w10108;
w10110 <= not w10044 and not w10109;
w10111 <= b(6) and not w10033;
w10112 <= not w10027 and w10111;
w10113 <= not w10035 and not w10112;
w10114 <= not w10110 and w10113;
w10115 <= not w10035 and not w10114;
w10116 <= b(7) and not w10024;
w10117 <= not w10018 and w10116;
w10118 <= not w10026 and not w10117;
w10119 <= not w10115 and w10118;
w10120 <= not w10026 and not w10119;
w10121 <= b(8) and not w10015;
w10122 <= not w10009 and w10121;
w10123 <= not w10017 and not w10122;
w10124 <= not w10120 and w10123;
w10125 <= not w10017 and not w10124;
w10126 <= b(9) and not w10006;
w10127 <= not w10000 and w10126;
w10128 <= not w10008 and not w10127;
w10129 <= not w10125 and w10128;
w10130 <= not w10008 and not w10129;
w10131 <= b(10) and not w9997;
w10132 <= not w9991 and w10131;
w10133 <= not w9999 and not w10132;
w10134 <= not w10130 and w10133;
w10135 <= not w9999 and not w10134;
w10136 <= b(11) and not w9988;
w10137 <= not w9982 and w10136;
w10138 <= not w9990 and not w10137;
w10139 <= not w10135 and w10138;
w10140 <= not w9990 and not w10139;
w10141 <= b(12) and not w9979;
w10142 <= not w9973 and w10141;
w10143 <= not w9981 and not w10142;
w10144 <= not w10140 and w10143;
w10145 <= not w9981 and not w10144;
w10146 <= b(13) and not w9970;
w10147 <= not w9964 and w10146;
w10148 <= not w9972 and not w10147;
w10149 <= not w10145 and w10148;
w10150 <= not w9972 and not w10149;
w10151 <= b(14) and not w9961;
w10152 <= not w9955 and w10151;
w10153 <= not w9963 and not w10152;
w10154 <= not w10150 and w10153;
w10155 <= not w9963 and not w10154;
w10156 <= b(15) and not w9952;
w10157 <= not w9946 and w10156;
w10158 <= not w9954 and not w10157;
w10159 <= not w10155 and w10158;
w10160 <= not w9954 and not w10159;
w10161 <= b(16) and not w9943;
w10162 <= not w9937 and w10161;
w10163 <= not w9945 and not w10162;
w10164 <= not w10160 and w10163;
w10165 <= not w9945 and not w10164;
w10166 <= b(17) and not w9934;
w10167 <= not w9928 and w10166;
w10168 <= not w9936 and not w10167;
w10169 <= not w10165 and w10168;
w10170 <= not w9936 and not w10169;
w10171 <= b(18) and not w9925;
w10172 <= not w9919 and w10171;
w10173 <= not w9927 and not w10172;
w10174 <= not w10170 and w10173;
w10175 <= not w9927 and not w10174;
w10176 <= b(19) and not w9916;
w10177 <= not w9910 and w10176;
w10178 <= not w9918 and not w10177;
w10179 <= not w10175 and w10178;
w10180 <= not w9918 and not w10179;
w10181 <= b(20) and not w9907;
w10182 <= not w9901 and w10181;
w10183 <= not w9909 and not w10182;
w10184 <= not w10180 and w10183;
w10185 <= not w9909 and not w10184;
w10186 <= b(21) and not w9898;
w10187 <= not w9892 and w10186;
w10188 <= not w9900 and not w10187;
w10189 <= not w10185 and w10188;
w10190 <= not w9900 and not w10189;
w10191 <= b(22) and not w9889;
w10192 <= not w9883 and w10191;
w10193 <= not w9891 and not w10192;
w10194 <= not w10190 and w10193;
w10195 <= not w9891 and not w10194;
w10196 <= b(23) and not w9880;
w10197 <= not w9874 and w10196;
w10198 <= not w9882 and not w10197;
w10199 <= not w10195 and w10198;
w10200 <= not w9882 and not w10199;
w10201 <= b(24) and not w9871;
w10202 <= not w9865 and w10201;
w10203 <= not w9873 and not w10202;
w10204 <= not w10200 and w10203;
w10205 <= not w9873 and not w10204;
w10206 <= b(25) and not w9862;
w10207 <= not w9856 and w10206;
w10208 <= not w9864 and not w10207;
w10209 <= not w10205 and w10208;
w10210 <= not w9864 and not w10209;
w10211 <= b(26) and not w9853;
w10212 <= not w9847 and w10211;
w10213 <= not w9855 and not w10212;
w10214 <= not w10210 and w10213;
w10215 <= not w9855 and not w10214;
w10216 <= b(27) and not w9844;
w10217 <= not w9838 and w10216;
w10218 <= not w9846 and not w10217;
w10219 <= not w10215 and w10218;
w10220 <= not w9846 and not w10219;
w10221 <= b(28) and not w9835;
w10222 <= not w9829 and w10221;
w10223 <= not w9837 and not w10222;
w10224 <= not w10220 and w10223;
w10225 <= not w9837 and not w10224;
w10226 <= b(29) and not w9826;
w10227 <= not w9820 and w10226;
w10228 <= not w9828 and not w10227;
w10229 <= not w10225 and w10228;
w10230 <= not w9828 and not w10229;
w10231 <= b(30) and not w9817;
w10232 <= not w9811 and w10231;
w10233 <= not w9819 and not w10232;
w10234 <= not w10230 and w10233;
w10235 <= not w9819 and not w10234;
w10236 <= b(31) and not w9808;
w10237 <= not w9802 and w10236;
w10238 <= not w9810 and not w10237;
w10239 <= not w10235 and w10238;
w10240 <= not w9810 and not w10239;
w10241 <= b(32) and not w9799;
w10242 <= not w9793 and w10241;
w10243 <= not w9801 and not w10242;
w10244 <= not w10240 and w10243;
w10245 <= not w9801 and not w10244;
w10246 <= b(33) and not w9790;
w10247 <= not w9784 and w10246;
w10248 <= not w9792 and not w10247;
w10249 <= not w10245 and w10248;
w10250 <= not w9792 and not w10249;
w10251 <= b(34) and not w9781;
w10252 <= not w9775 and w10251;
w10253 <= not w9783 and not w10252;
w10254 <= not w10250 and w10253;
w10255 <= not w9783 and not w10254;
w10256 <= b(35) and not w9772;
w10257 <= not w9766 and w10256;
w10258 <= not w9774 and not w10257;
w10259 <= not w10255 and w10258;
w10260 <= not w9774 and not w10259;
w10261 <= b(36) and not w9755;
w10262 <= not w9749 and w10261;
w10263 <= not w9765 and not w10262;
w10264 <= not w10260 and w10263;
w10265 <= not w9765 and not w10264;
w10266 <= b(37) and not w9757;
w10267 <= not w9762 and w10266;
w10268 <= not w9764 and not w10267;
w10269 <= not w10265 and w10268;
w10270 <= not w9764 and not w10269;
w10271 <= w34 and w36;
w10272 <= w45 and w10271;
w10273 <= w31 and w10272;
w10274 <= not w10270 and w10273;
w10275 <= not w9756 and not w10274;
w10276 <= not w9774 and w10263;
w10277 <= not w10259 and w10276;
w10278 <= not w10260 and not w10263;
w10279 <= not w10277 and not w10278;
w10280 <= w10273 and not w10279;
w10281 <= not w10270 and w10280;
w10282 <= not w10275 and not w10281;
w10283 <= not b(37) and not w10282;
w10284 <= not w9773 and not w10274;
w10285 <= not w9783 and w10258;
w10286 <= not w10254 and w10285;
w10287 <= not w10255 and not w10258;
w10288 <= not w10286 and not w10287;
w10289 <= w10273 and not w10288;
w10290 <= not w10270 and w10289;
w10291 <= not w10284 and not w10290;
w10292 <= not b(36) and not w10291;
w10293 <= not w9782 and not w10274;
w10294 <= not w9792 and w10253;
w10295 <= not w10249 and w10294;
w10296 <= not w10250 and not w10253;
w10297 <= not w10295 and not w10296;
w10298 <= w10273 and not w10297;
w10299 <= not w10270 and w10298;
w10300 <= not w10293 and not w10299;
w10301 <= not b(35) and not w10300;
w10302 <= not w9791 and not w10274;
w10303 <= not w9801 and w10248;
w10304 <= not w10244 and w10303;
w10305 <= not w10245 and not w10248;
w10306 <= not w10304 and not w10305;
w10307 <= w10273 and not w10306;
w10308 <= not w10270 and w10307;
w10309 <= not w10302 and not w10308;
w10310 <= not b(34) and not w10309;
w10311 <= not w9800 and not w10274;
w10312 <= not w9810 and w10243;
w10313 <= not w10239 and w10312;
w10314 <= not w10240 and not w10243;
w10315 <= not w10313 and not w10314;
w10316 <= w10273 and not w10315;
w10317 <= not w10270 and w10316;
w10318 <= not w10311 and not w10317;
w10319 <= not b(33) and not w10318;
w10320 <= not w9809 and not w10274;
w10321 <= not w9819 and w10238;
w10322 <= not w10234 and w10321;
w10323 <= not w10235 and not w10238;
w10324 <= not w10322 and not w10323;
w10325 <= w10273 and not w10324;
w10326 <= not w10270 and w10325;
w10327 <= not w10320 and not w10326;
w10328 <= not b(32) and not w10327;
w10329 <= not w9818 and not w10274;
w10330 <= not w9828 and w10233;
w10331 <= not w10229 and w10330;
w10332 <= not w10230 and not w10233;
w10333 <= not w10331 and not w10332;
w10334 <= w10273 and not w10333;
w10335 <= not w10270 and w10334;
w10336 <= not w10329 and not w10335;
w10337 <= not b(31) and not w10336;
w10338 <= not w9827 and not w10274;
w10339 <= not w9837 and w10228;
w10340 <= not w10224 and w10339;
w10341 <= not w10225 and not w10228;
w10342 <= not w10340 and not w10341;
w10343 <= w10273 and not w10342;
w10344 <= not w10270 and w10343;
w10345 <= not w10338 and not w10344;
w10346 <= not b(30) and not w10345;
w10347 <= not w9836 and not w10274;
w10348 <= not w9846 and w10223;
w10349 <= not w10219 and w10348;
w10350 <= not w10220 and not w10223;
w10351 <= not w10349 and not w10350;
w10352 <= w10273 and not w10351;
w10353 <= not w10270 and w10352;
w10354 <= not w10347 and not w10353;
w10355 <= not b(29) and not w10354;
w10356 <= not w9845 and not w10274;
w10357 <= not w9855 and w10218;
w10358 <= not w10214 and w10357;
w10359 <= not w10215 and not w10218;
w10360 <= not w10358 and not w10359;
w10361 <= w10273 and not w10360;
w10362 <= not w10270 and w10361;
w10363 <= not w10356 and not w10362;
w10364 <= not b(28) and not w10363;
w10365 <= not w9854 and not w10274;
w10366 <= not w9864 and w10213;
w10367 <= not w10209 and w10366;
w10368 <= not w10210 and not w10213;
w10369 <= not w10367 and not w10368;
w10370 <= w10273 and not w10369;
w10371 <= not w10270 and w10370;
w10372 <= not w10365 and not w10371;
w10373 <= not b(27) and not w10372;
w10374 <= not w9863 and not w10274;
w10375 <= not w9873 and w10208;
w10376 <= not w10204 and w10375;
w10377 <= not w10205 and not w10208;
w10378 <= not w10376 and not w10377;
w10379 <= w10273 and not w10378;
w10380 <= not w10270 and w10379;
w10381 <= not w10374 and not w10380;
w10382 <= not b(26) and not w10381;
w10383 <= not w9872 and not w10274;
w10384 <= not w9882 and w10203;
w10385 <= not w10199 and w10384;
w10386 <= not w10200 and not w10203;
w10387 <= not w10385 and not w10386;
w10388 <= w10273 and not w10387;
w10389 <= not w10270 and w10388;
w10390 <= not w10383 and not w10389;
w10391 <= not b(25) and not w10390;
w10392 <= not w9881 and not w10274;
w10393 <= not w9891 and w10198;
w10394 <= not w10194 and w10393;
w10395 <= not w10195 and not w10198;
w10396 <= not w10394 and not w10395;
w10397 <= w10273 and not w10396;
w10398 <= not w10270 and w10397;
w10399 <= not w10392 and not w10398;
w10400 <= not b(24) and not w10399;
w10401 <= not w9890 and not w10274;
w10402 <= not w9900 and w10193;
w10403 <= not w10189 and w10402;
w10404 <= not w10190 and not w10193;
w10405 <= not w10403 and not w10404;
w10406 <= w10273 and not w10405;
w10407 <= not w10270 and w10406;
w10408 <= not w10401 and not w10407;
w10409 <= not b(23) and not w10408;
w10410 <= not w9899 and not w10274;
w10411 <= not w9909 and w10188;
w10412 <= not w10184 and w10411;
w10413 <= not w10185 and not w10188;
w10414 <= not w10412 and not w10413;
w10415 <= w10273 and not w10414;
w10416 <= not w10270 and w10415;
w10417 <= not w10410 and not w10416;
w10418 <= not b(22) and not w10417;
w10419 <= not w9908 and not w10274;
w10420 <= not w9918 and w10183;
w10421 <= not w10179 and w10420;
w10422 <= not w10180 and not w10183;
w10423 <= not w10421 and not w10422;
w10424 <= w10273 and not w10423;
w10425 <= not w10270 and w10424;
w10426 <= not w10419 and not w10425;
w10427 <= not b(21) and not w10426;
w10428 <= not w9917 and not w10274;
w10429 <= not w9927 and w10178;
w10430 <= not w10174 and w10429;
w10431 <= not w10175 and not w10178;
w10432 <= not w10430 and not w10431;
w10433 <= w10273 and not w10432;
w10434 <= not w10270 and w10433;
w10435 <= not w10428 and not w10434;
w10436 <= not b(20) and not w10435;
w10437 <= not w9926 and not w10274;
w10438 <= not w9936 and w10173;
w10439 <= not w10169 and w10438;
w10440 <= not w10170 and not w10173;
w10441 <= not w10439 and not w10440;
w10442 <= w10273 and not w10441;
w10443 <= not w10270 and w10442;
w10444 <= not w10437 and not w10443;
w10445 <= not b(19) and not w10444;
w10446 <= not w9935 and not w10274;
w10447 <= not w9945 and w10168;
w10448 <= not w10164 and w10447;
w10449 <= not w10165 and not w10168;
w10450 <= not w10448 and not w10449;
w10451 <= w10273 and not w10450;
w10452 <= not w10270 and w10451;
w10453 <= not w10446 and not w10452;
w10454 <= not b(18) and not w10453;
w10455 <= not w9944 and not w10274;
w10456 <= not w9954 and w10163;
w10457 <= not w10159 and w10456;
w10458 <= not w10160 and not w10163;
w10459 <= not w10457 and not w10458;
w10460 <= w10273 and not w10459;
w10461 <= not w10270 and w10460;
w10462 <= not w10455 and not w10461;
w10463 <= not b(17) and not w10462;
w10464 <= not w9953 and not w10274;
w10465 <= not w9963 and w10158;
w10466 <= not w10154 and w10465;
w10467 <= not w10155 and not w10158;
w10468 <= not w10466 and not w10467;
w10469 <= w10273 and not w10468;
w10470 <= not w10270 and w10469;
w10471 <= not w10464 and not w10470;
w10472 <= not b(16) and not w10471;
w10473 <= not w9962 and not w10274;
w10474 <= not w9972 and w10153;
w10475 <= not w10149 and w10474;
w10476 <= not w10150 and not w10153;
w10477 <= not w10475 and not w10476;
w10478 <= w10273 and not w10477;
w10479 <= not w10270 and w10478;
w10480 <= not w10473 and not w10479;
w10481 <= not b(15) and not w10480;
w10482 <= not w9971 and not w10274;
w10483 <= not w9981 and w10148;
w10484 <= not w10144 and w10483;
w10485 <= not w10145 and not w10148;
w10486 <= not w10484 and not w10485;
w10487 <= w10273 and not w10486;
w10488 <= not w10270 and w10487;
w10489 <= not w10482 and not w10488;
w10490 <= not b(14) and not w10489;
w10491 <= not w9980 and not w10274;
w10492 <= not w9990 and w10143;
w10493 <= not w10139 and w10492;
w10494 <= not w10140 and not w10143;
w10495 <= not w10493 and not w10494;
w10496 <= w10273 and not w10495;
w10497 <= not w10270 and w10496;
w10498 <= not w10491 and not w10497;
w10499 <= not b(13) and not w10498;
w10500 <= not w9989 and not w10274;
w10501 <= not w9999 and w10138;
w10502 <= not w10134 and w10501;
w10503 <= not w10135 and not w10138;
w10504 <= not w10502 and not w10503;
w10505 <= w10273 and not w10504;
w10506 <= not w10270 and w10505;
w10507 <= not w10500 and not w10506;
w10508 <= not b(12) and not w10507;
w10509 <= not w9998 and not w10274;
w10510 <= not w10008 and w10133;
w10511 <= not w10129 and w10510;
w10512 <= not w10130 and not w10133;
w10513 <= not w10511 and not w10512;
w10514 <= w10273 and not w10513;
w10515 <= not w10270 and w10514;
w10516 <= not w10509 and not w10515;
w10517 <= not b(11) and not w10516;
w10518 <= not w10007 and not w10274;
w10519 <= not w10017 and w10128;
w10520 <= not w10124 and w10519;
w10521 <= not w10125 and not w10128;
w10522 <= not w10520 and not w10521;
w10523 <= w10273 and not w10522;
w10524 <= not w10270 and w10523;
w10525 <= not w10518 and not w10524;
w10526 <= not b(10) and not w10525;
w10527 <= not w10016 and not w10274;
w10528 <= not w10026 and w10123;
w10529 <= not w10119 and w10528;
w10530 <= not w10120 and not w10123;
w10531 <= not w10529 and not w10530;
w10532 <= w10273 and not w10531;
w10533 <= not w10270 and w10532;
w10534 <= not w10527 and not w10533;
w10535 <= not b(9) and not w10534;
w10536 <= not w10025 and not w10274;
w10537 <= not w10035 and w10118;
w10538 <= not w10114 and w10537;
w10539 <= not w10115 and not w10118;
w10540 <= not w10538 and not w10539;
w10541 <= w10273 and not w10540;
w10542 <= not w10270 and w10541;
w10543 <= not w10536 and not w10542;
w10544 <= not b(8) and not w10543;
w10545 <= not w10034 and not w10274;
w10546 <= not w10044 and w10113;
w10547 <= not w10109 and w10546;
w10548 <= not w10110 and not w10113;
w10549 <= not w10547 and not w10548;
w10550 <= w10273 and not w10549;
w10551 <= not w10270 and w10550;
w10552 <= not w10545 and not w10551;
w10553 <= not b(7) and not w10552;
w10554 <= not w10043 and not w10274;
w10555 <= not w10053 and w10108;
w10556 <= not w10104 and w10555;
w10557 <= not w10105 and not w10108;
w10558 <= not w10556 and not w10557;
w10559 <= w10273 and not w10558;
w10560 <= not w10270 and w10559;
w10561 <= not w10554 and not w10560;
w10562 <= not b(6) and not w10561;
w10563 <= not w10052 and not w10274;
w10564 <= not w10062 and w10103;
w10565 <= not w10099 and w10564;
w10566 <= not w10100 and not w10103;
w10567 <= not w10565 and not w10566;
w10568 <= w10273 and not w10567;
w10569 <= not w10270 and w10568;
w10570 <= not w10563 and not w10569;
w10571 <= not b(5) and not w10570;
w10572 <= not w10061 and not w10274;
w10573 <= not w10070 and w10098;
w10574 <= not w10094 and w10573;
w10575 <= not w10095 and not w10098;
w10576 <= not w10574 and not w10575;
w10577 <= w10273 and not w10576;
w10578 <= not w10270 and w10577;
w10579 <= not w10572 and not w10578;
w10580 <= not b(4) and not w10579;
w10581 <= not w10069 and not w10274;
w10582 <= not w10089 and w10093;
w10583 <= not w10088 and w10582;
w10584 <= not w10090 and not w10093;
w10585 <= not w10583 and not w10584;
w10586 <= w10273 and not w10585;
w10587 <= not w10270 and w10586;
w10588 <= not w10581 and not w10587;
w10589 <= not b(3) and not w10588;
w10590 <= not w10082 and not w10274;
w10591 <= not w10085 and w10087;
w10592 <= not w10083 and w10591;
w10593 <= w10273 and not w10592;
w10594 <= not w10088 and w10593;
w10595 <= not w10270 and w10594;
w10596 <= not w10590 and not w10595;
w10597 <= not b(2) and not w10596;
w10598 <= b(0) and not b(38);
w10599 <= w153 and w10598;
w10600 <= w164 and w10599;
w10601 <= w340 and w10600;
w10602 <= w338 and w10601;
w10603 <= not w10270 and w10602;
w10604 <= a(26) and not w10603;
w10605 <= w36 and w10087;
w10606 <= w34 and w10605;
w10607 <= w45 and w10606;
w10608 <= w31 and w10607;
w10609 <= not w10270 and w10608;
w10610 <= not w10604 and not w10609;
w10611 <= b(1) and not w10610;
w10612 <= not b(1) and not w10609;
w10613 <= not w10604 and w10612;
w10614 <= not w10611 and not w10613;
w10615 <= not a(25) and b(0);
w10616 <= not w10614 and not w10615;
w10617 <= not b(1) and not w10610;
w10618 <= not w10616 and not w10617;
w10619 <= b(2) and not w10595;
w10620 <= not w10590 and w10619;
w10621 <= not w10597 and not w10620;
w10622 <= not w10618 and w10621;
w10623 <= not w10597 and not w10622;
w10624 <= b(3) and not w10587;
w10625 <= not w10581 and w10624;
w10626 <= not w10589 and not w10625;
w10627 <= not w10623 and w10626;
w10628 <= not w10589 and not w10627;
w10629 <= b(4) and not w10578;
w10630 <= not w10572 and w10629;
w10631 <= not w10580 and not w10630;
w10632 <= not w10628 and w10631;
w10633 <= not w10580 and not w10632;
w10634 <= b(5) and not w10569;
w10635 <= not w10563 and w10634;
w10636 <= not w10571 and not w10635;
w10637 <= not w10633 and w10636;
w10638 <= not w10571 and not w10637;
w10639 <= b(6) and not w10560;
w10640 <= not w10554 and w10639;
w10641 <= not w10562 and not w10640;
w10642 <= not w10638 and w10641;
w10643 <= not w10562 and not w10642;
w10644 <= b(7) and not w10551;
w10645 <= not w10545 and w10644;
w10646 <= not w10553 and not w10645;
w10647 <= not w10643 and w10646;
w10648 <= not w10553 and not w10647;
w10649 <= b(8) and not w10542;
w10650 <= not w10536 and w10649;
w10651 <= not w10544 and not w10650;
w10652 <= not w10648 and w10651;
w10653 <= not w10544 and not w10652;
w10654 <= b(9) and not w10533;
w10655 <= not w10527 and w10654;
w10656 <= not w10535 and not w10655;
w10657 <= not w10653 and w10656;
w10658 <= not w10535 and not w10657;
w10659 <= b(10) and not w10524;
w10660 <= not w10518 and w10659;
w10661 <= not w10526 and not w10660;
w10662 <= not w10658 and w10661;
w10663 <= not w10526 and not w10662;
w10664 <= b(11) and not w10515;
w10665 <= not w10509 and w10664;
w10666 <= not w10517 and not w10665;
w10667 <= not w10663 and w10666;
w10668 <= not w10517 and not w10667;
w10669 <= b(12) and not w10506;
w10670 <= not w10500 and w10669;
w10671 <= not w10508 and not w10670;
w10672 <= not w10668 and w10671;
w10673 <= not w10508 and not w10672;
w10674 <= b(13) and not w10497;
w10675 <= not w10491 and w10674;
w10676 <= not w10499 and not w10675;
w10677 <= not w10673 and w10676;
w10678 <= not w10499 and not w10677;
w10679 <= b(14) and not w10488;
w10680 <= not w10482 and w10679;
w10681 <= not w10490 and not w10680;
w10682 <= not w10678 and w10681;
w10683 <= not w10490 and not w10682;
w10684 <= b(15) and not w10479;
w10685 <= not w10473 and w10684;
w10686 <= not w10481 and not w10685;
w10687 <= not w10683 and w10686;
w10688 <= not w10481 and not w10687;
w10689 <= b(16) and not w10470;
w10690 <= not w10464 and w10689;
w10691 <= not w10472 and not w10690;
w10692 <= not w10688 and w10691;
w10693 <= not w10472 and not w10692;
w10694 <= b(17) and not w10461;
w10695 <= not w10455 and w10694;
w10696 <= not w10463 and not w10695;
w10697 <= not w10693 and w10696;
w10698 <= not w10463 and not w10697;
w10699 <= b(18) and not w10452;
w10700 <= not w10446 and w10699;
w10701 <= not w10454 and not w10700;
w10702 <= not w10698 and w10701;
w10703 <= not w10454 and not w10702;
w10704 <= b(19) and not w10443;
w10705 <= not w10437 and w10704;
w10706 <= not w10445 and not w10705;
w10707 <= not w10703 and w10706;
w10708 <= not w10445 and not w10707;
w10709 <= b(20) and not w10434;
w10710 <= not w10428 and w10709;
w10711 <= not w10436 and not w10710;
w10712 <= not w10708 and w10711;
w10713 <= not w10436 and not w10712;
w10714 <= b(21) and not w10425;
w10715 <= not w10419 and w10714;
w10716 <= not w10427 and not w10715;
w10717 <= not w10713 and w10716;
w10718 <= not w10427 and not w10717;
w10719 <= b(22) and not w10416;
w10720 <= not w10410 and w10719;
w10721 <= not w10418 and not w10720;
w10722 <= not w10718 and w10721;
w10723 <= not w10418 and not w10722;
w10724 <= b(23) and not w10407;
w10725 <= not w10401 and w10724;
w10726 <= not w10409 and not w10725;
w10727 <= not w10723 and w10726;
w10728 <= not w10409 and not w10727;
w10729 <= b(24) and not w10398;
w10730 <= not w10392 and w10729;
w10731 <= not w10400 and not w10730;
w10732 <= not w10728 and w10731;
w10733 <= not w10400 and not w10732;
w10734 <= b(25) and not w10389;
w10735 <= not w10383 and w10734;
w10736 <= not w10391 and not w10735;
w10737 <= not w10733 and w10736;
w10738 <= not w10391 and not w10737;
w10739 <= b(26) and not w10380;
w10740 <= not w10374 and w10739;
w10741 <= not w10382 and not w10740;
w10742 <= not w10738 and w10741;
w10743 <= not w10382 and not w10742;
w10744 <= b(27) and not w10371;
w10745 <= not w10365 and w10744;
w10746 <= not w10373 and not w10745;
w10747 <= not w10743 and w10746;
w10748 <= not w10373 and not w10747;
w10749 <= b(28) and not w10362;
w10750 <= not w10356 and w10749;
w10751 <= not w10364 and not w10750;
w10752 <= not w10748 and w10751;
w10753 <= not w10364 and not w10752;
w10754 <= b(29) and not w10353;
w10755 <= not w10347 and w10754;
w10756 <= not w10355 and not w10755;
w10757 <= not w10753 and w10756;
w10758 <= not w10355 and not w10757;
w10759 <= b(30) and not w10344;
w10760 <= not w10338 and w10759;
w10761 <= not w10346 and not w10760;
w10762 <= not w10758 and w10761;
w10763 <= not w10346 and not w10762;
w10764 <= b(31) and not w10335;
w10765 <= not w10329 and w10764;
w10766 <= not w10337 and not w10765;
w10767 <= not w10763 and w10766;
w10768 <= not w10337 and not w10767;
w10769 <= b(32) and not w10326;
w10770 <= not w10320 and w10769;
w10771 <= not w10328 and not w10770;
w10772 <= not w10768 and w10771;
w10773 <= not w10328 and not w10772;
w10774 <= b(33) and not w10317;
w10775 <= not w10311 and w10774;
w10776 <= not w10319 and not w10775;
w10777 <= not w10773 and w10776;
w10778 <= not w10319 and not w10777;
w10779 <= b(34) and not w10308;
w10780 <= not w10302 and w10779;
w10781 <= not w10310 and not w10780;
w10782 <= not w10778 and w10781;
w10783 <= not w10310 and not w10782;
w10784 <= b(35) and not w10299;
w10785 <= not w10293 and w10784;
w10786 <= not w10301 and not w10785;
w10787 <= not w10783 and w10786;
w10788 <= not w10301 and not w10787;
w10789 <= b(36) and not w10290;
w10790 <= not w10284 and w10789;
w10791 <= not w10292 and not w10790;
w10792 <= not w10788 and w10791;
w10793 <= not w10292 and not w10792;
w10794 <= b(37) and not w10281;
w10795 <= not w10275 and w10794;
w10796 <= not w10283 and not w10795;
w10797 <= not w10793 and w10796;
w10798 <= not w10283 and not w10797;
w10799 <= not w9763 and not w10274;
w10800 <= not w9765 and w10268;
w10801 <= not w10264 and w10800;
w10802 <= not w10265 and not w10268;
w10803 <= not w10801 and not w10802;
w10804 <= w10274 and not w10803;
w10805 <= not w10799 and not w10804;
w10806 <= not b(38) and not w10805;
w10807 <= b(38) and not w10799;
w10808 <= not w10804 and w10807;
w10809 <= w153 and w164;
w10810 <= w340 and w10809;
w10811 <= w338 and w10810;
w10812 <= not w10808 and w10811;
w10813 <= not w10806 and w10812;
w10814 <= not w10798 and w10813;
w10815 <= w10273 and not w10805;
w10816 <= not w10814 and not w10815;
w10817 <= not w10292 and w10796;
w10818 <= not w10792 and w10817;
w10819 <= not w10793 and not w10796;
w10820 <= not w10818 and not w10819;
w10821 <= not w10816 and not w10820;
w10822 <= not w10282 and not w10815;
w10823 <= not w10814 and w10822;
w10824 <= not w10821 and not w10823;
w10825 <= not w10283 and not w10808;
w10826 <= not w10806 and w10825;
w10827 <= not w10797 and w10826;
w10828 <= not w10806 and not w10808;
w10829 <= not w10798 and not w10828;
w10830 <= not w10827 and not w10829;
w10831 <= not w10816 and not w10830;
w10832 <= not w10805 and not w10815;
w10833 <= not w10814 and w10832;
w10834 <= not w10831 and not w10833;
w10835 <= not b(39) and not w10834;
w10836 <= not b(38) and not w10824;
w10837 <= not w10301 and w10791;
w10838 <= not w10787 and w10837;
w10839 <= not w10788 and not w10791;
w10840 <= not w10838 and not w10839;
w10841 <= not w10816 and not w10840;
w10842 <= not w10291 and not w10815;
w10843 <= not w10814 and w10842;
w10844 <= not w10841 and not w10843;
w10845 <= not b(37) and not w10844;
w10846 <= not w10310 and w10786;
w10847 <= not w10782 and w10846;
w10848 <= not w10783 and not w10786;
w10849 <= not w10847 and not w10848;
w10850 <= not w10816 and not w10849;
w10851 <= not w10300 and not w10815;
w10852 <= not w10814 and w10851;
w10853 <= not w10850 and not w10852;
w10854 <= not b(36) and not w10853;
w10855 <= not w10319 and w10781;
w10856 <= not w10777 and w10855;
w10857 <= not w10778 and not w10781;
w10858 <= not w10856 and not w10857;
w10859 <= not w10816 and not w10858;
w10860 <= not w10309 and not w10815;
w10861 <= not w10814 and w10860;
w10862 <= not w10859 and not w10861;
w10863 <= not b(35) and not w10862;
w10864 <= not w10328 and w10776;
w10865 <= not w10772 and w10864;
w10866 <= not w10773 and not w10776;
w10867 <= not w10865 and not w10866;
w10868 <= not w10816 and not w10867;
w10869 <= not w10318 and not w10815;
w10870 <= not w10814 and w10869;
w10871 <= not w10868 and not w10870;
w10872 <= not b(34) and not w10871;
w10873 <= not w10337 and w10771;
w10874 <= not w10767 and w10873;
w10875 <= not w10768 and not w10771;
w10876 <= not w10874 and not w10875;
w10877 <= not w10816 and not w10876;
w10878 <= not w10327 and not w10815;
w10879 <= not w10814 and w10878;
w10880 <= not w10877 and not w10879;
w10881 <= not b(33) and not w10880;
w10882 <= not w10346 and w10766;
w10883 <= not w10762 and w10882;
w10884 <= not w10763 and not w10766;
w10885 <= not w10883 and not w10884;
w10886 <= not w10816 and not w10885;
w10887 <= not w10336 and not w10815;
w10888 <= not w10814 and w10887;
w10889 <= not w10886 and not w10888;
w10890 <= not b(32) and not w10889;
w10891 <= not w10355 and w10761;
w10892 <= not w10757 and w10891;
w10893 <= not w10758 and not w10761;
w10894 <= not w10892 and not w10893;
w10895 <= not w10816 and not w10894;
w10896 <= not w10345 and not w10815;
w10897 <= not w10814 and w10896;
w10898 <= not w10895 and not w10897;
w10899 <= not b(31) and not w10898;
w10900 <= not w10364 and w10756;
w10901 <= not w10752 and w10900;
w10902 <= not w10753 and not w10756;
w10903 <= not w10901 and not w10902;
w10904 <= not w10816 and not w10903;
w10905 <= not w10354 and not w10815;
w10906 <= not w10814 and w10905;
w10907 <= not w10904 and not w10906;
w10908 <= not b(30) and not w10907;
w10909 <= not w10373 and w10751;
w10910 <= not w10747 and w10909;
w10911 <= not w10748 and not w10751;
w10912 <= not w10910 and not w10911;
w10913 <= not w10816 and not w10912;
w10914 <= not w10363 and not w10815;
w10915 <= not w10814 and w10914;
w10916 <= not w10913 and not w10915;
w10917 <= not b(29) and not w10916;
w10918 <= not w10382 and w10746;
w10919 <= not w10742 and w10918;
w10920 <= not w10743 and not w10746;
w10921 <= not w10919 and not w10920;
w10922 <= not w10816 and not w10921;
w10923 <= not w10372 and not w10815;
w10924 <= not w10814 and w10923;
w10925 <= not w10922 and not w10924;
w10926 <= not b(28) and not w10925;
w10927 <= not w10391 and w10741;
w10928 <= not w10737 and w10927;
w10929 <= not w10738 and not w10741;
w10930 <= not w10928 and not w10929;
w10931 <= not w10816 and not w10930;
w10932 <= not w10381 and not w10815;
w10933 <= not w10814 and w10932;
w10934 <= not w10931 and not w10933;
w10935 <= not b(27) and not w10934;
w10936 <= not w10400 and w10736;
w10937 <= not w10732 and w10936;
w10938 <= not w10733 and not w10736;
w10939 <= not w10937 and not w10938;
w10940 <= not w10816 and not w10939;
w10941 <= not w10390 and not w10815;
w10942 <= not w10814 and w10941;
w10943 <= not w10940 and not w10942;
w10944 <= not b(26) and not w10943;
w10945 <= not w10409 and w10731;
w10946 <= not w10727 and w10945;
w10947 <= not w10728 and not w10731;
w10948 <= not w10946 and not w10947;
w10949 <= not w10816 and not w10948;
w10950 <= not w10399 and not w10815;
w10951 <= not w10814 and w10950;
w10952 <= not w10949 and not w10951;
w10953 <= not b(25) and not w10952;
w10954 <= not w10418 and w10726;
w10955 <= not w10722 and w10954;
w10956 <= not w10723 and not w10726;
w10957 <= not w10955 and not w10956;
w10958 <= not w10816 and not w10957;
w10959 <= not w10408 and not w10815;
w10960 <= not w10814 and w10959;
w10961 <= not w10958 and not w10960;
w10962 <= not b(24) and not w10961;
w10963 <= not w10427 and w10721;
w10964 <= not w10717 and w10963;
w10965 <= not w10718 and not w10721;
w10966 <= not w10964 and not w10965;
w10967 <= not w10816 and not w10966;
w10968 <= not w10417 and not w10815;
w10969 <= not w10814 and w10968;
w10970 <= not w10967 and not w10969;
w10971 <= not b(23) and not w10970;
w10972 <= not w10436 and w10716;
w10973 <= not w10712 and w10972;
w10974 <= not w10713 and not w10716;
w10975 <= not w10973 and not w10974;
w10976 <= not w10816 and not w10975;
w10977 <= not w10426 and not w10815;
w10978 <= not w10814 and w10977;
w10979 <= not w10976 and not w10978;
w10980 <= not b(22) and not w10979;
w10981 <= not w10445 and w10711;
w10982 <= not w10707 and w10981;
w10983 <= not w10708 and not w10711;
w10984 <= not w10982 and not w10983;
w10985 <= not w10816 and not w10984;
w10986 <= not w10435 and not w10815;
w10987 <= not w10814 and w10986;
w10988 <= not w10985 and not w10987;
w10989 <= not b(21) and not w10988;
w10990 <= not w10454 and w10706;
w10991 <= not w10702 and w10990;
w10992 <= not w10703 and not w10706;
w10993 <= not w10991 and not w10992;
w10994 <= not w10816 and not w10993;
w10995 <= not w10444 and not w10815;
w10996 <= not w10814 and w10995;
w10997 <= not w10994 and not w10996;
w10998 <= not b(20) and not w10997;
w10999 <= not w10463 and w10701;
w11000 <= not w10697 and w10999;
w11001 <= not w10698 and not w10701;
w11002 <= not w11000 and not w11001;
w11003 <= not w10816 and not w11002;
w11004 <= not w10453 and not w10815;
w11005 <= not w10814 and w11004;
w11006 <= not w11003 and not w11005;
w11007 <= not b(19) and not w11006;
w11008 <= not w10472 and w10696;
w11009 <= not w10692 and w11008;
w11010 <= not w10693 and not w10696;
w11011 <= not w11009 and not w11010;
w11012 <= not w10816 and not w11011;
w11013 <= not w10462 and not w10815;
w11014 <= not w10814 and w11013;
w11015 <= not w11012 and not w11014;
w11016 <= not b(18) and not w11015;
w11017 <= not w10481 and w10691;
w11018 <= not w10687 and w11017;
w11019 <= not w10688 and not w10691;
w11020 <= not w11018 and not w11019;
w11021 <= not w10816 and not w11020;
w11022 <= not w10471 and not w10815;
w11023 <= not w10814 and w11022;
w11024 <= not w11021 and not w11023;
w11025 <= not b(17) and not w11024;
w11026 <= not w10490 and w10686;
w11027 <= not w10682 and w11026;
w11028 <= not w10683 and not w10686;
w11029 <= not w11027 and not w11028;
w11030 <= not w10816 and not w11029;
w11031 <= not w10480 and not w10815;
w11032 <= not w10814 and w11031;
w11033 <= not w11030 and not w11032;
w11034 <= not b(16) and not w11033;
w11035 <= not w10499 and w10681;
w11036 <= not w10677 and w11035;
w11037 <= not w10678 and not w10681;
w11038 <= not w11036 and not w11037;
w11039 <= not w10816 and not w11038;
w11040 <= not w10489 and not w10815;
w11041 <= not w10814 and w11040;
w11042 <= not w11039 and not w11041;
w11043 <= not b(15) and not w11042;
w11044 <= not w10508 and w10676;
w11045 <= not w10672 and w11044;
w11046 <= not w10673 and not w10676;
w11047 <= not w11045 and not w11046;
w11048 <= not w10816 and not w11047;
w11049 <= not w10498 and not w10815;
w11050 <= not w10814 and w11049;
w11051 <= not w11048 and not w11050;
w11052 <= not b(14) and not w11051;
w11053 <= not w10517 and w10671;
w11054 <= not w10667 and w11053;
w11055 <= not w10668 and not w10671;
w11056 <= not w11054 and not w11055;
w11057 <= not w10816 and not w11056;
w11058 <= not w10507 and not w10815;
w11059 <= not w10814 and w11058;
w11060 <= not w11057 and not w11059;
w11061 <= not b(13) and not w11060;
w11062 <= not w10526 and w10666;
w11063 <= not w10662 and w11062;
w11064 <= not w10663 and not w10666;
w11065 <= not w11063 and not w11064;
w11066 <= not w10816 and not w11065;
w11067 <= not w10516 and not w10815;
w11068 <= not w10814 and w11067;
w11069 <= not w11066 and not w11068;
w11070 <= not b(12) and not w11069;
w11071 <= not w10535 and w10661;
w11072 <= not w10657 and w11071;
w11073 <= not w10658 and not w10661;
w11074 <= not w11072 and not w11073;
w11075 <= not w10816 and not w11074;
w11076 <= not w10525 and not w10815;
w11077 <= not w10814 and w11076;
w11078 <= not w11075 and not w11077;
w11079 <= not b(11) and not w11078;
w11080 <= not w10544 and w10656;
w11081 <= not w10652 and w11080;
w11082 <= not w10653 and not w10656;
w11083 <= not w11081 and not w11082;
w11084 <= not w10816 and not w11083;
w11085 <= not w10534 and not w10815;
w11086 <= not w10814 and w11085;
w11087 <= not w11084 and not w11086;
w11088 <= not b(10) and not w11087;
w11089 <= not w10553 and w10651;
w11090 <= not w10647 and w11089;
w11091 <= not w10648 and not w10651;
w11092 <= not w11090 and not w11091;
w11093 <= not w10816 and not w11092;
w11094 <= not w10543 and not w10815;
w11095 <= not w10814 and w11094;
w11096 <= not w11093 and not w11095;
w11097 <= not b(9) and not w11096;
w11098 <= not w10562 and w10646;
w11099 <= not w10642 and w11098;
w11100 <= not w10643 and not w10646;
w11101 <= not w11099 and not w11100;
w11102 <= not w10816 and not w11101;
w11103 <= not w10552 and not w10815;
w11104 <= not w10814 and w11103;
w11105 <= not w11102 and not w11104;
w11106 <= not b(8) and not w11105;
w11107 <= not w10571 and w10641;
w11108 <= not w10637 and w11107;
w11109 <= not w10638 and not w10641;
w11110 <= not w11108 and not w11109;
w11111 <= not w10816 and not w11110;
w11112 <= not w10561 and not w10815;
w11113 <= not w10814 and w11112;
w11114 <= not w11111 and not w11113;
w11115 <= not b(7) and not w11114;
w11116 <= not w10580 and w10636;
w11117 <= not w10632 and w11116;
w11118 <= not w10633 and not w10636;
w11119 <= not w11117 and not w11118;
w11120 <= not w10816 and not w11119;
w11121 <= not w10570 and not w10815;
w11122 <= not w10814 and w11121;
w11123 <= not w11120 and not w11122;
w11124 <= not b(6) and not w11123;
w11125 <= not w10589 and w10631;
w11126 <= not w10627 and w11125;
w11127 <= not w10628 and not w10631;
w11128 <= not w11126 and not w11127;
w11129 <= not w10816 and not w11128;
w11130 <= not w10579 and not w10815;
w11131 <= not w10814 and w11130;
w11132 <= not w11129 and not w11131;
w11133 <= not b(5) and not w11132;
w11134 <= not w10597 and w10626;
w11135 <= not w10622 and w11134;
w11136 <= not w10623 and not w10626;
w11137 <= not w11135 and not w11136;
w11138 <= not w10816 and not w11137;
w11139 <= not w10588 and not w10815;
w11140 <= not w10814 and w11139;
w11141 <= not w11138 and not w11140;
w11142 <= not b(4) and not w11141;
w11143 <= not w10617 and w10621;
w11144 <= not w10616 and w11143;
w11145 <= not w10618 and not w10621;
w11146 <= not w11144 and not w11145;
w11147 <= not w10816 and not w11146;
w11148 <= not w10596 and not w10815;
w11149 <= not w10814 and w11148;
w11150 <= not w11147 and not w11149;
w11151 <= not b(3) and not w11150;
w11152 <= not w10613 and w10615;
w11153 <= not w10611 and w11152;
w11154 <= not w10616 and not w11153;
w11155 <= not w10816 and w11154;
w11156 <= not w10610 and not w10815;
w11157 <= not w10814 and w11156;
w11158 <= not w11155 and not w11157;
w11159 <= not b(2) and not w11158;
w11160 <= b(0) and not w10816;
w11161 <= a(25) and not w11160;
w11162 <= w10615 and not w10816;
w11163 <= not w11161 and not w11162;
w11164 <= b(1) and not w11163;
w11165 <= not b(1) and not w11162;
w11166 <= not w11161 and w11165;
w11167 <= not w11164 and not w11166;
w11168 <= not a(24) and b(0);
w11169 <= not w11167 and not w11168;
w11170 <= not b(1) and not w11163;
w11171 <= not w11169 and not w11170;
w11172 <= b(2) and not w11157;
w11173 <= not w11155 and w11172;
w11174 <= not w11159 and not w11173;
w11175 <= not w11171 and w11174;
w11176 <= not w11159 and not w11175;
w11177 <= b(3) and not w11149;
w11178 <= not w11147 and w11177;
w11179 <= not w11151 and not w11178;
w11180 <= not w11176 and w11179;
w11181 <= not w11151 and not w11180;
w11182 <= b(4) and not w11140;
w11183 <= not w11138 and w11182;
w11184 <= not w11142 and not w11183;
w11185 <= not w11181 and w11184;
w11186 <= not w11142 and not w11185;
w11187 <= b(5) and not w11131;
w11188 <= not w11129 and w11187;
w11189 <= not w11133 and not w11188;
w11190 <= not w11186 and w11189;
w11191 <= not w11133 and not w11190;
w11192 <= b(6) and not w11122;
w11193 <= not w11120 and w11192;
w11194 <= not w11124 and not w11193;
w11195 <= not w11191 and w11194;
w11196 <= not w11124 and not w11195;
w11197 <= b(7) and not w11113;
w11198 <= not w11111 and w11197;
w11199 <= not w11115 and not w11198;
w11200 <= not w11196 and w11199;
w11201 <= not w11115 and not w11200;
w11202 <= b(8) and not w11104;
w11203 <= not w11102 and w11202;
w11204 <= not w11106 and not w11203;
w11205 <= not w11201 and w11204;
w11206 <= not w11106 and not w11205;
w11207 <= b(9) and not w11095;
w11208 <= not w11093 and w11207;
w11209 <= not w11097 and not w11208;
w11210 <= not w11206 and w11209;
w11211 <= not w11097 and not w11210;
w11212 <= b(10) and not w11086;
w11213 <= not w11084 and w11212;
w11214 <= not w11088 and not w11213;
w11215 <= not w11211 and w11214;
w11216 <= not w11088 and not w11215;
w11217 <= b(11) and not w11077;
w11218 <= not w11075 and w11217;
w11219 <= not w11079 and not w11218;
w11220 <= not w11216 and w11219;
w11221 <= not w11079 and not w11220;
w11222 <= b(12) and not w11068;
w11223 <= not w11066 and w11222;
w11224 <= not w11070 and not w11223;
w11225 <= not w11221 and w11224;
w11226 <= not w11070 and not w11225;
w11227 <= b(13) and not w11059;
w11228 <= not w11057 and w11227;
w11229 <= not w11061 and not w11228;
w11230 <= not w11226 and w11229;
w11231 <= not w11061 and not w11230;
w11232 <= b(14) and not w11050;
w11233 <= not w11048 and w11232;
w11234 <= not w11052 and not w11233;
w11235 <= not w11231 and w11234;
w11236 <= not w11052 and not w11235;
w11237 <= b(15) and not w11041;
w11238 <= not w11039 and w11237;
w11239 <= not w11043 and not w11238;
w11240 <= not w11236 and w11239;
w11241 <= not w11043 and not w11240;
w11242 <= b(16) and not w11032;
w11243 <= not w11030 and w11242;
w11244 <= not w11034 and not w11243;
w11245 <= not w11241 and w11244;
w11246 <= not w11034 and not w11245;
w11247 <= b(17) and not w11023;
w11248 <= not w11021 and w11247;
w11249 <= not w11025 and not w11248;
w11250 <= not w11246 and w11249;
w11251 <= not w11025 and not w11250;
w11252 <= b(18) and not w11014;
w11253 <= not w11012 and w11252;
w11254 <= not w11016 and not w11253;
w11255 <= not w11251 and w11254;
w11256 <= not w11016 and not w11255;
w11257 <= b(19) and not w11005;
w11258 <= not w11003 and w11257;
w11259 <= not w11007 and not w11258;
w11260 <= not w11256 and w11259;
w11261 <= not w11007 and not w11260;
w11262 <= b(20) and not w10996;
w11263 <= not w10994 and w11262;
w11264 <= not w10998 and not w11263;
w11265 <= not w11261 and w11264;
w11266 <= not w10998 and not w11265;
w11267 <= b(21) and not w10987;
w11268 <= not w10985 and w11267;
w11269 <= not w10989 and not w11268;
w11270 <= not w11266 and w11269;
w11271 <= not w10989 and not w11270;
w11272 <= b(22) and not w10978;
w11273 <= not w10976 and w11272;
w11274 <= not w10980 and not w11273;
w11275 <= not w11271 and w11274;
w11276 <= not w10980 and not w11275;
w11277 <= b(23) and not w10969;
w11278 <= not w10967 and w11277;
w11279 <= not w10971 and not w11278;
w11280 <= not w11276 and w11279;
w11281 <= not w10971 and not w11280;
w11282 <= b(24) and not w10960;
w11283 <= not w10958 and w11282;
w11284 <= not w10962 and not w11283;
w11285 <= not w11281 and w11284;
w11286 <= not w10962 and not w11285;
w11287 <= b(25) and not w10951;
w11288 <= not w10949 and w11287;
w11289 <= not w10953 and not w11288;
w11290 <= not w11286 and w11289;
w11291 <= not w10953 and not w11290;
w11292 <= b(26) and not w10942;
w11293 <= not w10940 and w11292;
w11294 <= not w10944 and not w11293;
w11295 <= not w11291 and w11294;
w11296 <= not w10944 and not w11295;
w11297 <= b(27) and not w10933;
w11298 <= not w10931 and w11297;
w11299 <= not w10935 and not w11298;
w11300 <= not w11296 and w11299;
w11301 <= not w10935 and not w11300;
w11302 <= b(28) and not w10924;
w11303 <= not w10922 and w11302;
w11304 <= not w10926 and not w11303;
w11305 <= not w11301 and w11304;
w11306 <= not w10926 and not w11305;
w11307 <= b(29) and not w10915;
w11308 <= not w10913 and w11307;
w11309 <= not w10917 and not w11308;
w11310 <= not w11306 and w11309;
w11311 <= not w10917 and not w11310;
w11312 <= b(30) and not w10906;
w11313 <= not w10904 and w11312;
w11314 <= not w10908 and not w11313;
w11315 <= not w11311 and w11314;
w11316 <= not w10908 and not w11315;
w11317 <= b(31) and not w10897;
w11318 <= not w10895 and w11317;
w11319 <= not w10899 and not w11318;
w11320 <= not w11316 and w11319;
w11321 <= not w10899 and not w11320;
w11322 <= b(32) and not w10888;
w11323 <= not w10886 and w11322;
w11324 <= not w10890 and not w11323;
w11325 <= not w11321 and w11324;
w11326 <= not w10890 and not w11325;
w11327 <= b(33) and not w10879;
w11328 <= not w10877 and w11327;
w11329 <= not w10881 and not w11328;
w11330 <= not w11326 and w11329;
w11331 <= not w10881 and not w11330;
w11332 <= b(34) and not w10870;
w11333 <= not w10868 and w11332;
w11334 <= not w10872 and not w11333;
w11335 <= not w11331 and w11334;
w11336 <= not w10872 and not w11335;
w11337 <= b(35) and not w10861;
w11338 <= not w10859 and w11337;
w11339 <= not w10863 and not w11338;
w11340 <= not w11336 and w11339;
w11341 <= not w10863 and not w11340;
w11342 <= b(36) and not w10852;
w11343 <= not w10850 and w11342;
w11344 <= not w10854 and not w11343;
w11345 <= not w11341 and w11344;
w11346 <= not w10854 and not w11345;
w11347 <= b(37) and not w10843;
w11348 <= not w10841 and w11347;
w11349 <= not w10845 and not w11348;
w11350 <= not w11346 and w11349;
w11351 <= not w10845 and not w11350;
w11352 <= b(38) and not w10823;
w11353 <= not w10821 and w11352;
w11354 <= not w10836 and not w11353;
w11355 <= not w11351 and w11354;
w11356 <= not w10836 and not w11355;
w11357 <= b(39) and not w10833;
w11358 <= not w10831 and w11357;
w11359 <= not w10835 and not w11358;
w11360 <= not w11356 and w11359;
w11361 <= not w10835 and not w11360;
w11362 <= w81 and w83;
w11363 <= not w11361 and w11362;
w11364 <= not w10824 and not w11363;
w11365 <= not w10845 and w11354;
w11366 <= not w11350 and w11365;
w11367 <= not w11351 and not w11354;
w11368 <= not w11366 and not w11367;
w11369 <= w11362 and not w11368;
w11370 <= not w11361 and w11369;
w11371 <= not w11364 and not w11370;
w11372 <= not w10834 and not w11363;
w11373 <= not w10836 and w11359;
w11374 <= not w11355 and w11373;
w11375 <= not w11356 and not w11359;
w11376 <= not w11374 and not w11375;
w11377 <= w11363 and not w11376;
w11378 <= not w11372 and not w11377;
w11379 <= not b(40) and not w11378;
w11380 <= not b(39) and not w11371;
w11381 <= not w10844 and not w11363;
w11382 <= not w10854 and w11349;
w11383 <= not w11345 and w11382;
w11384 <= not w11346 and not w11349;
w11385 <= not w11383 and not w11384;
w11386 <= w11362 and not w11385;
w11387 <= not w11361 and w11386;
w11388 <= not w11381 and not w11387;
w11389 <= not b(38) and not w11388;
w11390 <= not w10853 and not w11363;
w11391 <= not w10863 and w11344;
w11392 <= not w11340 and w11391;
w11393 <= not w11341 and not w11344;
w11394 <= not w11392 and not w11393;
w11395 <= w11362 and not w11394;
w11396 <= not w11361 and w11395;
w11397 <= not w11390 and not w11396;
w11398 <= not b(37) and not w11397;
w11399 <= not w10862 and not w11363;
w11400 <= not w10872 and w11339;
w11401 <= not w11335 and w11400;
w11402 <= not w11336 and not w11339;
w11403 <= not w11401 and not w11402;
w11404 <= w11362 and not w11403;
w11405 <= not w11361 and w11404;
w11406 <= not w11399 and not w11405;
w11407 <= not b(36) and not w11406;
w11408 <= not w10871 and not w11363;
w11409 <= not w10881 and w11334;
w11410 <= not w11330 and w11409;
w11411 <= not w11331 and not w11334;
w11412 <= not w11410 and not w11411;
w11413 <= w11362 and not w11412;
w11414 <= not w11361 and w11413;
w11415 <= not w11408 and not w11414;
w11416 <= not b(35) and not w11415;
w11417 <= not w10880 and not w11363;
w11418 <= not w10890 and w11329;
w11419 <= not w11325 and w11418;
w11420 <= not w11326 and not w11329;
w11421 <= not w11419 and not w11420;
w11422 <= w11362 and not w11421;
w11423 <= not w11361 and w11422;
w11424 <= not w11417 and not w11423;
w11425 <= not b(34) and not w11424;
w11426 <= not w10889 and not w11363;
w11427 <= not w10899 and w11324;
w11428 <= not w11320 and w11427;
w11429 <= not w11321 and not w11324;
w11430 <= not w11428 and not w11429;
w11431 <= w11362 and not w11430;
w11432 <= not w11361 and w11431;
w11433 <= not w11426 and not w11432;
w11434 <= not b(33) and not w11433;
w11435 <= not w10898 and not w11363;
w11436 <= not w10908 and w11319;
w11437 <= not w11315 and w11436;
w11438 <= not w11316 and not w11319;
w11439 <= not w11437 and not w11438;
w11440 <= w11362 and not w11439;
w11441 <= not w11361 and w11440;
w11442 <= not w11435 and not w11441;
w11443 <= not b(32) and not w11442;
w11444 <= not w10907 and not w11363;
w11445 <= not w10917 and w11314;
w11446 <= not w11310 and w11445;
w11447 <= not w11311 and not w11314;
w11448 <= not w11446 and not w11447;
w11449 <= w11362 and not w11448;
w11450 <= not w11361 and w11449;
w11451 <= not w11444 and not w11450;
w11452 <= not b(31) and not w11451;
w11453 <= not w10916 and not w11363;
w11454 <= not w10926 and w11309;
w11455 <= not w11305 and w11454;
w11456 <= not w11306 and not w11309;
w11457 <= not w11455 and not w11456;
w11458 <= w11362 and not w11457;
w11459 <= not w11361 and w11458;
w11460 <= not w11453 and not w11459;
w11461 <= not b(30) and not w11460;
w11462 <= not w10925 and not w11363;
w11463 <= not w10935 and w11304;
w11464 <= not w11300 and w11463;
w11465 <= not w11301 and not w11304;
w11466 <= not w11464 and not w11465;
w11467 <= w11362 and not w11466;
w11468 <= not w11361 and w11467;
w11469 <= not w11462 and not w11468;
w11470 <= not b(29) and not w11469;
w11471 <= not w10934 and not w11363;
w11472 <= not w10944 and w11299;
w11473 <= not w11295 and w11472;
w11474 <= not w11296 and not w11299;
w11475 <= not w11473 and not w11474;
w11476 <= w11362 and not w11475;
w11477 <= not w11361 and w11476;
w11478 <= not w11471 and not w11477;
w11479 <= not b(28) and not w11478;
w11480 <= not w10943 and not w11363;
w11481 <= not w10953 and w11294;
w11482 <= not w11290 and w11481;
w11483 <= not w11291 and not w11294;
w11484 <= not w11482 and not w11483;
w11485 <= w11362 and not w11484;
w11486 <= not w11361 and w11485;
w11487 <= not w11480 and not w11486;
w11488 <= not b(27) and not w11487;
w11489 <= not w10952 and not w11363;
w11490 <= not w10962 and w11289;
w11491 <= not w11285 and w11490;
w11492 <= not w11286 and not w11289;
w11493 <= not w11491 and not w11492;
w11494 <= w11362 and not w11493;
w11495 <= not w11361 and w11494;
w11496 <= not w11489 and not w11495;
w11497 <= not b(26) and not w11496;
w11498 <= not w10961 and not w11363;
w11499 <= not w10971 and w11284;
w11500 <= not w11280 and w11499;
w11501 <= not w11281 and not w11284;
w11502 <= not w11500 and not w11501;
w11503 <= w11362 and not w11502;
w11504 <= not w11361 and w11503;
w11505 <= not w11498 and not w11504;
w11506 <= not b(25) and not w11505;
w11507 <= not w10970 and not w11363;
w11508 <= not w10980 and w11279;
w11509 <= not w11275 and w11508;
w11510 <= not w11276 and not w11279;
w11511 <= not w11509 and not w11510;
w11512 <= w11362 and not w11511;
w11513 <= not w11361 and w11512;
w11514 <= not w11507 and not w11513;
w11515 <= not b(24) and not w11514;
w11516 <= not w10979 and not w11363;
w11517 <= not w10989 and w11274;
w11518 <= not w11270 and w11517;
w11519 <= not w11271 and not w11274;
w11520 <= not w11518 and not w11519;
w11521 <= w11362 and not w11520;
w11522 <= not w11361 and w11521;
w11523 <= not w11516 and not w11522;
w11524 <= not b(23) and not w11523;
w11525 <= not w10988 and not w11363;
w11526 <= not w10998 and w11269;
w11527 <= not w11265 and w11526;
w11528 <= not w11266 and not w11269;
w11529 <= not w11527 and not w11528;
w11530 <= w11362 and not w11529;
w11531 <= not w11361 and w11530;
w11532 <= not w11525 and not w11531;
w11533 <= not b(22) and not w11532;
w11534 <= not w10997 and not w11363;
w11535 <= not w11007 and w11264;
w11536 <= not w11260 and w11535;
w11537 <= not w11261 and not w11264;
w11538 <= not w11536 and not w11537;
w11539 <= w11362 and not w11538;
w11540 <= not w11361 and w11539;
w11541 <= not w11534 and not w11540;
w11542 <= not b(21) and not w11541;
w11543 <= not w11006 and not w11363;
w11544 <= not w11016 and w11259;
w11545 <= not w11255 and w11544;
w11546 <= not w11256 and not w11259;
w11547 <= not w11545 and not w11546;
w11548 <= w11362 and not w11547;
w11549 <= not w11361 and w11548;
w11550 <= not w11543 and not w11549;
w11551 <= not b(20) and not w11550;
w11552 <= not w11015 and not w11363;
w11553 <= not w11025 and w11254;
w11554 <= not w11250 and w11553;
w11555 <= not w11251 and not w11254;
w11556 <= not w11554 and not w11555;
w11557 <= w11362 and not w11556;
w11558 <= not w11361 and w11557;
w11559 <= not w11552 and not w11558;
w11560 <= not b(19) and not w11559;
w11561 <= not w11024 and not w11363;
w11562 <= not w11034 and w11249;
w11563 <= not w11245 and w11562;
w11564 <= not w11246 and not w11249;
w11565 <= not w11563 and not w11564;
w11566 <= w11362 and not w11565;
w11567 <= not w11361 and w11566;
w11568 <= not w11561 and not w11567;
w11569 <= not b(18) and not w11568;
w11570 <= not w11033 and not w11363;
w11571 <= not w11043 and w11244;
w11572 <= not w11240 and w11571;
w11573 <= not w11241 and not w11244;
w11574 <= not w11572 and not w11573;
w11575 <= w11362 and not w11574;
w11576 <= not w11361 and w11575;
w11577 <= not w11570 and not w11576;
w11578 <= not b(17) and not w11577;
w11579 <= not w11042 and not w11363;
w11580 <= not w11052 and w11239;
w11581 <= not w11235 and w11580;
w11582 <= not w11236 and not w11239;
w11583 <= not w11581 and not w11582;
w11584 <= w11362 and not w11583;
w11585 <= not w11361 and w11584;
w11586 <= not w11579 and not w11585;
w11587 <= not b(16) and not w11586;
w11588 <= not w11051 and not w11363;
w11589 <= not w11061 and w11234;
w11590 <= not w11230 and w11589;
w11591 <= not w11231 and not w11234;
w11592 <= not w11590 and not w11591;
w11593 <= w11362 and not w11592;
w11594 <= not w11361 and w11593;
w11595 <= not w11588 and not w11594;
w11596 <= not b(15) and not w11595;
w11597 <= not w11060 and not w11363;
w11598 <= not w11070 and w11229;
w11599 <= not w11225 and w11598;
w11600 <= not w11226 and not w11229;
w11601 <= not w11599 and not w11600;
w11602 <= w11362 and not w11601;
w11603 <= not w11361 and w11602;
w11604 <= not w11597 and not w11603;
w11605 <= not b(14) and not w11604;
w11606 <= not w11069 and not w11363;
w11607 <= not w11079 and w11224;
w11608 <= not w11220 and w11607;
w11609 <= not w11221 and not w11224;
w11610 <= not w11608 and not w11609;
w11611 <= w11362 and not w11610;
w11612 <= not w11361 and w11611;
w11613 <= not w11606 and not w11612;
w11614 <= not b(13) and not w11613;
w11615 <= not w11078 and not w11363;
w11616 <= not w11088 and w11219;
w11617 <= not w11215 and w11616;
w11618 <= not w11216 and not w11219;
w11619 <= not w11617 and not w11618;
w11620 <= w11362 and not w11619;
w11621 <= not w11361 and w11620;
w11622 <= not w11615 and not w11621;
w11623 <= not b(12) and not w11622;
w11624 <= not w11087 and not w11363;
w11625 <= not w11097 and w11214;
w11626 <= not w11210 and w11625;
w11627 <= not w11211 and not w11214;
w11628 <= not w11626 and not w11627;
w11629 <= w11362 and not w11628;
w11630 <= not w11361 and w11629;
w11631 <= not w11624 and not w11630;
w11632 <= not b(11) and not w11631;
w11633 <= not w11096 and not w11363;
w11634 <= not w11106 and w11209;
w11635 <= not w11205 and w11634;
w11636 <= not w11206 and not w11209;
w11637 <= not w11635 and not w11636;
w11638 <= w11362 and not w11637;
w11639 <= not w11361 and w11638;
w11640 <= not w11633 and not w11639;
w11641 <= not b(10) and not w11640;
w11642 <= not w11105 and not w11363;
w11643 <= not w11115 and w11204;
w11644 <= not w11200 and w11643;
w11645 <= not w11201 and not w11204;
w11646 <= not w11644 and not w11645;
w11647 <= w11362 and not w11646;
w11648 <= not w11361 and w11647;
w11649 <= not w11642 and not w11648;
w11650 <= not b(9) and not w11649;
w11651 <= not w11114 and not w11363;
w11652 <= not w11124 and w11199;
w11653 <= not w11195 and w11652;
w11654 <= not w11196 and not w11199;
w11655 <= not w11653 and not w11654;
w11656 <= w11362 and not w11655;
w11657 <= not w11361 and w11656;
w11658 <= not w11651 and not w11657;
w11659 <= not b(8) and not w11658;
w11660 <= not w11123 and not w11363;
w11661 <= not w11133 and w11194;
w11662 <= not w11190 and w11661;
w11663 <= not w11191 and not w11194;
w11664 <= not w11662 and not w11663;
w11665 <= w11362 and not w11664;
w11666 <= not w11361 and w11665;
w11667 <= not w11660 and not w11666;
w11668 <= not b(7) and not w11667;
w11669 <= not w11132 and not w11363;
w11670 <= not w11142 and w11189;
w11671 <= not w11185 and w11670;
w11672 <= not w11186 and not w11189;
w11673 <= not w11671 and not w11672;
w11674 <= w11362 and not w11673;
w11675 <= not w11361 and w11674;
w11676 <= not w11669 and not w11675;
w11677 <= not b(6) and not w11676;
w11678 <= not w11141 and not w11363;
w11679 <= not w11151 and w11184;
w11680 <= not w11180 and w11679;
w11681 <= not w11181 and not w11184;
w11682 <= not w11680 and not w11681;
w11683 <= w11362 and not w11682;
w11684 <= not w11361 and w11683;
w11685 <= not w11678 and not w11684;
w11686 <= not b(5) and not w11685;
w11687 <= not w11150 and not w11363;
w11688 <= not w11159 and w11179;
w11689 <= not w11175 and w11688;
w11690 <= not w11176 and not w11179;
w11691 <= not w11689 and not w11690;
w11692 <= w11362 and not w11691;
w11693 <= not w11361 and w11692;
w11694 <= not w11687 and not w11693;
w11695 <= not b(4) and not w11694;
w11696 <= not w11158 and not w11363;
w11697 <= not w11170 and w11174;
w11698 <= not w11169 and w11697;
w11699 <= not w11171 and not w11174;
w11700 <= not w11698 and not w11699;
w11701 <= w11362 and not w11700;
w11702 <= not w11361 and w11701;
w11703 <= not w11696 and not w11702;
w11704 <= not b(3) and not w11703;
w11705 <= not w11163 and not w11363;
w11706 <= not w11166 and w11168;
w11707 <= not w11164 and w11706;
w11708 <= w11362 and not w11707;
w11709 <= not w11169 and w11708;
w11710 <= not w11361 and w11709;
w11711 <= not w11705 and not w11710;
w11712 <= not b(2) and not w11711;
w11713 <= b(0) and not b(40);
w11714 <= w164 and w11713;
w11715 <= w340 and w11714;
w11716 <= w338 and w11715;
w11717 <= not w11361 and w11716;
w11718 <= a(24) and not w11717;
w11719 <= w34 and w11168;
w11720 <= w45 and w11719;
w11721 <= w31 and w11720;
w11722 <= not w11361 and w11721;
w11723 <= not w11718 and not w11722;
w11724 <= b(1) and not w11723;
w11725 <= not b(1) and not w11722;
w11726 <= not w11718 and w11725;
w11727 <= not w11724 and not w11726;
w11728 <= not a(23) and b(0);
w11729 <= not w11727 and not w11728;
w11730 <= not b(1) and not w11723;
w11731 <= not w11729 and not w11730;
w11732 <= b(2) and not w11710;
w11733 <= not w11705 and w11732;
w11734 <= not w11712 and not w11733;
w11735 <= not w11731 and w11734;
w11736 <= not w11712 and not w11735;
w11737 <= b(3) and not w11702;
w11738 <= not w11696 and w11737;
w11739 <= not w11704 and not w11738;
w11740 <= not w11736 and w11739;
w11741 <= not w11704 and not w11740;
w11742 <= b(4) and not w11693;
w11743 <= not w11687 and w11742;
w11744 <= not w11695 and not w11743;
w11745 <= not w11741 and w11744;
w11746 <= not w11695 and not w11745;
w11747 <= b(5) and not w11684;
w11748 <= not w11678 and w11747;
w11749 <= not w11686 and not w11748;
w11750 <= not w11746 and w11749;
w11751 <= not w11686 and not w11750;
w11752 <= b(6) and not w11675;
w11753 <= not w11669 and w11752;
w11754 <= not w11677 and not w11753;
w11755 <= not w11751 and w11754;
w11756 <= not w11677 and not w11755;
w11757 <= b(7) and not w11666;
w11758 <= not w11660 and w11757;
w11759 <= not w11668 and not w11758;
w11760 <= not w11756 and w11759;
w11761 <= not w11668 and not w11760;
w11762 <= b(8) and not w11657;
w11763 <= not w11651 and w11762;
w11764 <= not w11659 and not w11763;
w11765 <= not w11761 and w11764;
w11766 <= not w11659 and not w11765;
w11767 <= b(9) and not w11648;
w11768 <= not w11642 and w11767;
w11769 <= not w11650 and not w11768;
w11770 <= not w11766 and w11769;
w11771 <= not w11650 and not w11770;
w11772 <= b(10) and not w11639;
w11773 <= not w11633 and w11772;
w11774 <= not w11641 and not w11773;
w11775 <= not w11771 and w11774;
w11776 <= not w11641 and not w11775;
w11777 <= b(11) and not w11630;
w11778 <= not w11624 and w11777;
w11779 <= not w11632 and not w11778;
w11780 <= not w11776 and w11779;
w11781 <= not w11632 and not w11780;
w11782 <= b(12) and not w11621;
w11783 <= not w11615 and w11782;
w11784 <= not w11623 and not w11783;
w11785 <= not w11781 and w11784;
w11786 <= not w11623 and not w11785;
w11787 <= b(13) and not w11612;
w11788 <= not w11606 and w11787;
w11789 <= not w11614 and not w11788;
w11790 <= not w11786 and w11789;
w11791 <= not w11614 and not w11790;
w11792 <= b(14) and not w11603;
w11793 <= not w11597 and w11792;
w11794 <= not w11605 and not w11793;
w11795 <= not w11791 and w11794;
w11796 <= not w11605 and not w11795;
w11797 <= b(15) and not w11594;
w11798 <= not w11588 and w11797;
w11799 <= not w11596 and not w11798;
w11800 <= not w11796 and w11799;
w11801 <= not w11596 and not w11800;
w11802 <= b(16) and not w11585;
w11803 <= not w11579 and w11802;
w11804 <= not w11587 and not w11803;
w11805 <= not w11801 and w11804;
w11806 <= not w11587 and not w11805;
w11807 <= b(17) and not w11576;
w11808 <= not w11570 and w11807;
w11809 <= not w11578 and not w11808;
w11810 <= not w11806 and w11809;
w11811 <= not w11578 and not w11810;
w11812 <= b(18) and not w11567;
w11813 <= not w11561 and w11812;
w11814 <= not w11569 and not w11813;
w11815 <= not w11811 and w11814;
w11816 <= not w11569 and not w11815;
w11817 <= b(19) and not w11558;
w11818 <= not w11552 and w11817;
w11819 <= not w11560 and not w11818;
w11820 <= not w11816 and w11819;
w11821 <= not w11560 and not w11820;
w11822 <= b(20) and not w11549;
w11823 <= not w11543 and w11822;
w11824 <= not w11551 and not w11823;
w11825 <= not w11821 and w11824;
w11826 <= not w11551 and not w11825;
w11827 <= b(21) and not w11540;
w11828 <= not w11534 and w11827;
w11829 <= not w11542 and not w11828;
w11830 <= not w11826 and w11829;
w11831 <= not w11542 and not w11830;
w11832 <= b(22) and not w11531;
w11833 <= not w11525 and w11832;
w11834 <= not w11533 and not w11833;
w11835 <= not w11831 and w11834;
w11836 <= not w11533 and not w11835;
w11837 <= b(23) and not w11522;
w11838 <= not w11516 and w11837;
w11839 <= not w11524 and not w11838;
w11840 <= not w11836 and w11839;
w11841 <= not w11524 and not w11840;
w11842 <= b(24) and not w11513;
w11843 <= not w11507 and w11842;
w11844 <= not w11515 and not w11843;
w11845 <= not w11841 and w11844;
w11846 <= not w11515 and not w11845;
w11847 <= b(25) and not w11504;
w11848 <= not w11498 and w11847;
w11849 <= not w11506 and not w11848;
w11850 <= not w11846 and w11849;
w11851 <= not w11506 and not w11850;
w11852 <= b(26) and not w11495;
w11853 <= not w11489 and w11852;
w11854 <= not w11497 and not w11853;
w11855 <= not w11851 and w11854;
w11856 <= not w11497 and not w11855;
w11857 <= b(27) and not w11486;
w11858 <= not w11480 and w11857;
w11859 <= not w11488 and not w11858;
w11860 <= not w11856 and w11859;
w11861 <= not w11488 and not w11860;
w11862 <= b(28) and not w11477;
w11863 <= not w11471 and w11862;
w11864 <= not w11479 and not w11863;
w11865 <= not w11861 and w11864;
w11866 <= not w11479 and not w11865;
w11867 <= b(29) and not w11468;
w11868 <= not w11462 and w11867;
w11869 <= not w11470 and not w11868;
w11870 <= not w11866 and w11869;
w11871 <= not w11470 and not w11870;
w11872 <= b(30) and not w11459;
w11873 <= not w11453 and w11872;
w11874 <= not w11461 and not w11873;
w11875 <= not w11871 and w11874;
w11876 <= not w11461 and not w11875;
w11877 <= b(31) and not w11450;
w11878 <= not w11444 and w11877;
w11879 <= not w11452 and not w11878;
w11880 <= not w11876 and w11879;
w11881 <= not w11452 and not w11880;
w11882 <= b(32) and not w11441;
w11883 <= not w11435 and w11882;
w11884 <= not w11443 and not w11883;
w11885 <= not w11881 and w11884;
w11886 <= not w11443 and not w11885;
w11887 <= b(33) and not w11432;
w11888 <= not w11426 and w11887;
w11889 <= not w11434 and not w11888;
w11890 <= not w11886 and w11889;
w11891 <= not w11434 and not w11890;
w11892 <= b(34) and not w11423;
w11893 <= not w11417 and w11892;
w11894 <= not w11425 and not w11893;
w11895 <= not w11891 and w11894;
w11896 <= not w11425 and not w11895;
w11897 <= b(35) and not w11414;
w11898 <= not w11408 and w11897;
w11899 <= not w11416 and not w11898;
w11900 <= not w11896 and w11899;
w11901 <= not w11416 and not w11900;
w11902 <= b(36) and not w11405;
w11903 <= not w11399 and w11902;
w11904 <= not w11407 and not w11903;
w11905 <= not w11901 and w11904;
w11906 <= not w11407 and not w11905;
w11907 <= b(37) and not w11396;
w11908 <= not w11390 and w11907;
w11909 <= not w11398 and not w11908;
w11910 <= not w11906 and w11909;
w11911 <= not w11398 and not w11910;
w11912 <= b(38) and not w11387;
w11913 <= not w11381 and w11912;
w11914 <= not w11389 and not w11913;
w11915 <= not w11911 and w11914;
w11916 <= not w11389 and not w11915;
w11917 <= b(39) and not w11370;
w11918 <= not w11364 and w11917;
w11919 <= not w11380 and not w11918;
w11920 <= not w11916 and w11919;
w11921 <= not w11380 and not w11920;
w11922 <= b(40) and not w11372;
w11923 <= not w11377 and w11922;
w11924 <= not w11379 and not w11923;
w11925 <= not w11921 and w11924;
w11926 <= not w11379 and not w11925;
w11927 <= w151 and w165;
w11928 <= not w11926 and w11927;
w11929 <= not w11371 and not w11928;
w11930 <= not w11389 and w11919;
w11931 <= not w11915 and w11930;
w11932 <= not w11916 and not w11919;
w11933 <= not w11931 and not w11932;
w11934 <= w11927 and not w11933;
w11935 <= not w11926 and w11934;
w11936 <= not w11929 and not w11935;
w11937 <= not b(40) and not w11936;
w11938 <= not w11388 and not w11928;
w11939 <= not w11398 and w11914;
w11940 <= not w11910 and w11939;
w11941 <= not w11911 and not w11914;
w11942 <= not w11940 and not w11941;
w11943 <= w11927 and not w11942;
w11944 <= not w11926 and w11943;
w11945 <= not w11938 and not w11944;
w11946 <= not b(39) and not w11945;
w11947 <= not w11397 and not w11928;
w11948 <= not w11407 and w11909;
w11949 <= not w11905 and w11948;
w11950 <= not w11906 and not w11909;
w11951 <= not w11949 and not w11950;
w11952 <= w11927 and not w11951;
w11953 <= not w11926 and w11952;
w11954 <= not w11947 and not w11953;
w11955 <= not b(38) and not w11954;
w11956 <= not w11406 and not w11928;
w11957 <= not w11416 and w11904;
w11958 <= not w11900 and w11957;
w11959 <= not w11901 and not w11904;
w11960 <= not w11958 and not w11959;
w11961 <= w11927 and not w11960;
w11962 <= not w11926 and w11961;
w11963 <= not w11956 and not w11962;
w11964 <= not b(37) and not w11963;
w11965 <= not w11415 and not w11928;
w11966 <= not w11425 and w11899;
w11967 <= not w11895 and w11966;
w11968 <= not w11896 and not w11899;
w11969 <= not w11967 and not w11968;
w11970 <= w11927 and not w11969;
w11971 <= not w11926 and w11970;
w11972 <= not w11965 and not w11971;
w11973 <= not b(36) and not w11972;
w11974 <= not w11424 and not w11928;
w11975 <= not w11434 and w11894;
w11976 <= not w11890 and w11975;
w11977 <= not w11891 and not w11894;
w11978 <= not w11976 and not w11977;
w11979 <= w11927 and not w11978;
w11980 <= not w11926 and w11979;
w11981 <= not w11974 and not w11980;
w11982 <= not b(35) and not w11981;
w11983 <= not w11433 and not w11928;
w11984 <= not w11443 and w11889;
w11985 <= not w11885 and w11984;
w11986 <= not w11886 and not w11889;
w11987 <= not w11985 and not w11986;
w11988 <= w11927 and not w11987;
w11989 <= not w11926 and w11988;
w11990 <= not w11983 and not w11989;
w11991 <= not b(34) and not w11990;
w11992 <= not w11442 and not w11928;
w11993 <= not w11452 and w11884;
w11994 <= not w11880 and w11993;
w11995 <= not w11881 and not w11884;
w11996 <= not w11994 and not w11995;
w11997 <= w11927 and not w11996;
w11998 <= not w11926 and w11997;
w11999 <= not w11992 and not w11998;
w12000 <= not b(33) and not w11999;
w12001 <= not w11451 and not w11928;
w12002 <= not w11461 and w11879;
w12003 <= not w11875 and w12002;
w12004 <= not w11876 and not w11879;
w12005 <= not w12003 and not w12004;
w12006 <= w11927 and not w12005;
w12007 <= not w11926 and w12006;
w12008 <= not w12001 and not w12007;
w12009 <= not b(32) and not w12008;
w12010 <= not w11460 and not w11928;
w12011 <= not w11470 and w11874;
w12012 <= not w11870 and w12011;
w12013 <= not w11871 and not w11874;
w12014 <= not w12012 and not w12013;
w12015 <= w11927 and not w12014;
w12016 <= not w11926 and w12015;
w12017 <= not w12010 and not w12016;
w12018 <= not b(31) and not w12017;
w12019 <= not w11469 and not w11928;
w12020 <= not w11479 and w11869;
w12021 <= not w11865 and w12020;
w12022 <= not w11866 and not w11869;
w12023 <= not w12021 and not w12022;
w12024 <= w11927 and not w12023;
w12025 <= not w11926 and w12024;
w12026 <= not w12019 and not w12025;
w12027 <= not b(30) and not w12026;
w12028 <= not w11478 and not w11928;
w12029 <= not w11488 and w11864;
w12030 <= not w11860 and w12029;
w12031 <= not w11861 and not w11864;
w12032 <= not w12030 and not w12031;
w12033 <= w11927 and not w12032;
w12034 <= not w11926 and w12033;
w12035 <= not w12028 and not w12034;
w12036 <= not b(29) and not w12035;
w12037 <= not w11487 and not w11928;
w12038 <= not w11497 and w11859;
w12039 <= not w11855 and w12038;
w12040 <= not w11856 and not w11859;
w12041 <= not w12039 and not w12040;
w12042 <= w11927 and not w12041;
w12043 <= not w11926 and w12042;
w12044 <= not w12037 and not w12043;
w12045 <= not b(28) and not w12044;
w12046 <= not w11496 and not w11928;
w12047 <= not w11506 and w11854;
w12048 <= not w11850 and w12047;
w12049 <= not w11851 and not w11854;
w12050 <= not w12048 and not w12049;
w12051 <= w11927 and not w12050;
w12052 <= not w11926 and w12051;
w12053 <= not w12046 and not w12052;
w12054 <= not b(27) and not w12053;
w12055 <= not w11505 and not w11928;
w12056 <= not w11515 and w11849;
w12057 <= not w11845 and w12056;
w12058 <= not w11846 and not w11849;
w12059 <= not w12057 and not w12058;
w12060 <= w11927 and not w12059;
w12061 <= not w11926 and w12060;
w12062 <= not w12055 and not w12061;
w12063 <= not b(26) and not w12062;
w12064 <= not w11514 and not w11928;
w12065 <= not w11524 and w11844;
w12066 <= not w11840 and w12065;
w12067 <= not w11841 and not w11844;
w12068 <= not w12066 and not w12067;
w12069 <= w11927 and not w12068;
w12070 <= not w11926 and w12069;
w12071 <= not w12064 and not w12070;
w12072 <= not b(25) and not w12071;
w12073 <= not w11523 and not w11928;
w12074 <= not w11533 and w11839;
w12075 <= not w11835 and w12074;
w12076 <= not w11836 and not w11839;
w12077 <= not w12075 and not w12076;
w12078 <= w11927 and not w12077;
w12079 <= not w11926 and w12078;
w12080 <= not w12073 and not w12079;
w12081 <= not b(24) and not w12080;
w12082 <= not w11532 and not w11928;
w12083 <= not w11542 and w11834;
w12084 <= not w11830 and w12083;
w12085 <= not w11831 and not w11834;
w12086 <= not w12084 and not w12085;
w12087 <= w11927 and not w12086;
w12088 <= not w11926 and w12087;
w12089 <= not w12082 and not w12088;
w12090 <= not b(23) and not w12089;
w12091 <= not w11541 and not w11928;
w12092 <= not w11551 and w11829;
w12093 <= not w11825 and w12092;
w12094 <= not w11826 and not w11829;
w12095 <= not w12093 and not w12094;
w12096 <= w11927 and not w12095;
w12097 <= not w11926 and w12096;
w12098 <= not w12091 and not w12097;
w12099 <= not b(22) and not w12098;
w12100 <= not w11550 and not w11928;
w12101 <= not w11560 and w11824;
w12102 <= not w11820 and w12101;
w12103 <= not w11821 and not w11824;
w12104 <= not w12102 and not w12103;
w12105 <= w11927 and not w12104;
w12106 <= not w11926 and w12105;
w12107 <= not w12100 and not w12106;
w12108 <= not b(21) and not w12107;
w12109 <= not w11559 and not w11928;
w12110 <= not w11569 and w11819;
w12111 <= not w11815 and w12110;
w12112 <= not w11816 and not w11819;
w12113 <= not w12111 and not w12112;
w12114 <= w11927 and not w12113;
w12115 <= not w11926 and w12114;
w12116 <= not w12109 and not w12115;
w12117 <= not b(20) and not w12116;
w12118 <= not w11568 and not w11928;
w12119 <= not w11578 and w11814;
w12120 <= not w11810 and w12119;
w12121 <= not w11811 and not w11814;
w12122 <= not w12120 and not w12121;
w12123 <= w11927 and not w12122;
w12124 <= not w11926 and w12123;
w12125 <= not w12118 and not w12124;
w12126 <= not b(19) and not w12125;
w12127 <= not w11577 and not w11928;
w12128 <= not w11587 and w11809;
w12129 <= not w11805 and w12128;
w12130 <= not w11806 and not w11809;
w12131 <= not w12129 and not w12130;
w12132 <= w11927 and not w12131;
w12133 <= not w11926 and w12132;
w12134 <= not w12127 and not w12133;
w12135 <= not b(18) and not w12134;
w12136 <= not w11586 and not w11928;
w12137 <= not w11596 and w11804;
w12138 <= not w11800 and w12137;
w12139 <= not w11801 and not w11804;
w12140 <= not w12138 and not w12139;
w12141 <= w11927 and not w12140;
w12142 <= not w11926 and w12141;
w12143 <= not w12136 and not w12142;
w12144 <= not b(17) and not w12143;
w12145 <= not w11595 and not w11928;
w12146 <= not w11605 and w11799;
w12147 <= not w11795 and w12146;
w12148 <= not w11796 and not w11799;
w12149 <= not w12147 and not w12148;
w12150 <= w11927 and not w12149;
w12151 <= not w11926 and w12150;
w12152 <= not w12145 and not w12151;
w12153 <= not b(16) and not w12152;
w12154 <= not w11604 and not w11928;
w12155 <= not w11614 and w11794;
w12156 <= not w11790 and w12155;
w12157 <= not w11791 and not w11794;
w12158 <= not w12156 and not w12157;
w12159 <= w11927 and not w12158;
w12160 <= not w11926 and w12159;
w12161 <= not w12154 and not w12160;
w12162 <= not b(15) and not w12161;
w12163 <= not w11613 and not w11928;
w12164 <= not w11623 and w11789;
w12165 <= not w11785 and w12164;
w12166 <= not w11786 and not w11789;
w12167 <= not w12165 and not w12166;
w12168 <= w11927 and not w12167;
w12169 <= not w11926 and w12168;
w12170 <= not w12163 and not w12169;
w12171 <= not b(14) and not w12170;
w12172 <= not w11622 and not w11928;
w12173 <= not w11632 and w11784;
w12174 <= not w11780 and w12173;
w12175 <= not w11781 and not w11784;
w12176 <= not w12174 and not w12175;
w12177 <= w11927 and not w12176;
w12178 <= not w11926 and w12177;
w12179 <= not w12172 and not w12178;
w12180 <= not b(13) and not w12179;
w12181 <= not w11631 and not w11928;
w12182 <= not w11641 and w11779;
w12183 <= not w11775 and w12182;
w12184 <= not w11776 and not w11779;
w12185 <= not w12183 and not w12184;
w12186 <= w11927 and not w12185;
w12187 <= not w11926 and w12186;
w12188 <= not w12181 and not w12187;
w12189 <= not b(12) and not w12188;
w12190 <= not w11640 and not w11928;
w12191 <= not w11650 and w11774;
w12192 <= not w11770 and w12191;
w12193 <= not w11771 and not w11774;
w12194 <= not w12192 and not w12193;
w12195 <= w11927 and not w12194;
w12196 <= not w11926 and w12195;
w12197 <= not w12190 and not w12196;
w12198 <= not b(11) and not w12197;
w12199 <= not w11649 and not w11928;
w12200 <= not w11659 and w11769;
w12201 <= not w11765 and w12200;
w12202 <= not w11766 and not w11769;
w12203 <= not w12201 and not w12202;
w12204 <= w11927 and not w12203;
w12205 <= not w11926 and w12204;
w12206 <= not w12199 and not w12205;
w12207 <= not b(10) and not w12206;
w12208 <= not w11658 and not w11928;
w12209 <= not w11668 and w11764;
w12210 <= not w11760 and w12209;
w12211 <= not w11761 and not w11764;
w12212 <= not w12210 and not w12211;
w12213 <= w11927 and not w12212;
w12214 <= not w11926 and w12213;
w12215 <= not w12208 and not w12214;
w12216 <= not b(9) and not w12215;
w12217 <= not w11667 and not w11928;
w12218 <= not w11677 and w11759;
w12219 <= not w11755 and w12218;
w12220 <= not w11756 and not w11759;
w12221 <= not w12219 and not w12220;
w12222 <= w11927 and not w12221;
w12223 <= not w11926 and w12222;
w12224 <= not w12217 and not w12223;
w12225 <= not b(8) and not w12224;
w12226 <= not w11676 and not w11928;
w12227 <= not w11686 and w11754;
w12228 <= not w11750 and w12227;
w12229 <= not w11751 and not w11754;
w12230 <= not w12228 and not w12229;
w12231 <= w11927 and not w12230;
w12232 <= not w11926 and w12231;
w12233 <= not w12226 and not w12232;
w12234 <= not b(7) and not w12233;
w12235 <= not w11685 and not w11928;
w12236 <= not w11695 and w11749;
w12237 <= not w11745 and w12236;
w12238 <= not w11746 and not w11749;
w12239 <= not w12237 and not w12238;
w12240 <= w11927 and not w12239;
w12241 <= not w11926 and w12240;
w12242 <= not w12235 and not w12241;
w12243 <= not b(6) and not w12242;
w12244 <= not w11694 and not w11928;
w12245 <= not w11704 and w11744;
w12246 <= not w11740 and w12245;
w12247 <= not w11741 and not w11744;
w12248 <= not w12246 and not w12247;
w12249 <= w11927 and not w12248;
w12250 <= not w11926 and w12249;
w12251 <= not w12244 and not w12250;
w12252 <= not b(5) and not w12251;
w12253 <= not w11703 and not w11928;
w12254 <= not w11712 and w11739;
w12255 <= not w11735 and w12254;
w12256 <= not w11736 and not w11739;
w12257 <= not w12255 and not w12256;
w12258 <= w11927 and not w12257;
w12259 <= not w11926 and w12258;
w12260 <= not w12253 and not w12259;
w12261 <= not b(4) and not w12260;
w12262 <= not w11711 and not w11928;
w12263 <= not w11730 and w11734;
w12264 <= not w11729 and w12263;
w12265 <= not w11731 and not w11734;
w12266 <= not w12264 and not w12265;
w12267 <= w11927 and not w12266;
w12268 <= not w11926 and w12267;
w12269 <= not w12262 and not w12268;
w12270 <= not b(3) and not w12269;
w12271 <= not w11723 and not w11928;
w12272 <= not w11726 and w11728;
w12273 <= not w11724 and w12272;
w12274 <= w11927 and not w12273;
w12275 <= not w11729 and w12274;
w12276 <= not w11926 and w12275;
w12277 <= not w12271 and not w12276;
w12278 <= not b(2) and not w12277;
w12279 <= b(0) and not b(41);
w12280 <= w33 and w12279;
w12281 <= w44 and w12280;
w12282 <= w81 and w12281;
w12283 <= not w11926 and w12282;
w12284 <= a(23) and not w12283;
w12285 <= w164 and w11728;
w12286 <= w340 and w12285;
w12287 <= w338 and w12286;
w12288 <= not w11926 and w12287;
w12289 <= not w12284 and not w12288;
w12290 <= b(1) and not w12289;
w12291 <= not b(1) and not w12288;
w12292 <= not w12284 and w12291;
w12293 <= not w12290 and not w12292;
w12294 <= not a(22) and b(0);
w12295 <= not w12293 and not w12294;
w12296 <= not b(1) and not w12289;
w12297 <= not w12295 and not w12296;
w12298 <= b(2) and not w12276;
w12299 <= not w12271 and w12298;
w12300 <= not w12278 and not w12299;
w12301 <= not w12297 and w12300;
w12302 <= not w12278 and not w12301;
w12303 <= b(3) and not w12268;
w12304 <= not w12262 and w12303;
w12305 <= not w12270 and not w12304;
w12306 <= not w12302 and w12305;
w12307 <= not w12270 and not w12306;
w12308 <= b(4) and not w12259;
w12309 <= not w12253 and w12308;
w12310 <= not w12261 and not w12309;
w12311 <= not w12307 and w12310;
w12312 <= not w12261 and not w12311;
w12313 <= b(5) and not w12250;
w12314 <= not w12244 and w12313;
w12315 <= not w12252 and not w12314;
w12316 <= not w12312 and w12315;
w12317 <= not w12252 and not w12316;
w12318 <= b(6) and not w12241;
w12319 <= not w12235 and w12318;
w12320 <= not w12243 and not w12319;
w12321 <= not w12317 and w12320;
w12322 <= not w12243 and not w12321;
w12323 <= b(7) and not w12232;
w12324 <= not w12226 and w12323;
w12325 <= not w12234 and not w12324;
w12326 <= not w12322 and w12325;
w12327 <= not w12234 and not w12326;
w12328 <= b(8) and not w12223;
w12329 <= not w12217 and w12328;
w12330 <= not w12225 and not w12329;
w12331 <= not w12327 and w12330;
w12332 <= not w12225 and not w12331;
w12333 <= b(9) and not w12214;
w12334 <= not w12208 and w12333;
w12335 <= not w12216 and not w12334;
w12336 <= not w12332 and w12335;
w12337 <= not w12216 and not w12336;
w12338 <= b(10) and not w12205;
w12339 <= not w12199 and w12338;
w12340 <= not w12207 and not w12339;
w12341 <= not w12337 and w12340;
w12342 <= not w12207 and not w12341;
w12343 <= b(11) and not w12196;
w12344 <= not w12190 and w12343;
w12345 <= not w12198 and not w12344;
w12346 <= not w12342 and w12345;
w12347 <= not w12198 and not w12346;
w12348 <= b(12) and not w12187;
w12349 <= not w12181 and w12348;
w12350 <= not w12189 and not w12349;
w12351 <= not w12347 and w12350;
w12352 <= not w12189 and not w12351;
w12353 <= b(13) and not w12178;
w12354 <= not w12172 and w12353;
w12355 <= not w12180 and not w12354;
w12356 <= not w12352 and w12355;
w12357 <= not w12180 and not w12356;
w12358 <= b(14) and not w12169;
w12359 <= not w12163 and w12358;
w12360 <= not w12171 and not w12359;
w12361 <= not w12357 and w12360;
w12362 <= not w12171 and not w12361;
w12363 <= b(15) and not w12160;
w12364 <= not w12154 and w12363;
w12365 <= not w12162 and not w12364;
w12366 <= not w12362 and w12365;
w12367 <= not w12162 and not w12366;
w12368 <= b(16) and not w12151;
w12369 <= not w12145 and w12368;
w12370 <= not w12153 and not w12369;
w12371 <= not w12367 and w12370;
w12372 <= not w12153 and not w12371;
w12373 <= b(17) and not w12142;
w12374 <= not w12136 and w12373;
w12375 <= not w12144 and not w12374;
w12376 <= not w12372 and w12375;
w12377 <= not w12144 and not w12376;
w12378 <= b(18) and not w12133;
w12379 <= not w12127 and w12378;
w12380 <= not w12135 and not w12379;
w12381 <= not w12377 and w12380;
w12382 <= not w12135 and not w12381;
w12383 <= b(19) and not w12124;
w12384 <= not w12118 and w12383;
w12385 <= not w12126 and not w12384;
w12386 <= not w12382 and w12385;
w12387 <= not w12126 and not w12386;
w12388 <= b(20) and not w12115;
w12389 <= not w12109 and w12388;
w12390 <= not w12117 and not w12389;
w12391 <= not w12387 and w12390;
w12392 <= not w12117 and not w12391;
w12393 <= b(21) and not w12106;
w12394 <= not w12100 and w12393;
w12395 <= not w12108 and not w12394;
w12396 <= not w12392 and w12395;
w12397 <= not w12108 and not w12396;
w12398 <= b(22) and not w12097;
w12399 <= not w12091 and w12398;
w12400 <= not w12099 and not w12399;
w12401 <= not w12397 and w12400;
w12402 <= not w12099 and not w12401;
w12403 <= b(23) and not w12088;
w12404 <= not w12082 and w12403;
w12405 <= not w12090 and not w12404;
w12406 <= not w12402 and w12405;
w12407 <= not w12090 and not w12406;
w12408 <= b(24) and not w12079;
w12409 <= not w12073 and w12408;
w12410 <= not w12081 and not w12409;
w12411 <= not w12407 and w12410;
w12412 <= not w12081 and not w12411;
w12413 <= b(25) and not w12070;
w12414 <= not w12064 and w12413;
w12415 <= not w12072 and not w12414;
w12416 <= not w12412 and w12415;
w12417 <= not w12072 and not w12416;
w12418 <= b(26) and not w12061;
w12419 <= not w12055 and w12418;
w12420 <= not w12063 and not w12419;
w12421 <= not w12417 and w12420;
w12422 <= not w12063 and not w12421;
w12423 <= b(27) and not w12052;
w12424 <= not w12046 and w12423;
w12425 <= not w12054 and not w12424;
w12426 <= not w12422 and w12425;
w12427 <= not w12054 and not w12426;
w12428 <= b(28) and not w12043;
w12429 <= not w12037 and w12428;
w12430 <= not w12045 and not w12429;
w12431 <= not w12427 and w12430;
w12432 <= not w12045 and not w12431;
w12433 <= b(29) and not w12034;
w12434 <= not w12028 and w12433;
w12435 <= not w12036 and not w12434;
w12436 <= not w12432 and w12435;
w12437 <= not w12036 and not w12436;
w12438 <= b(30) and not w12025;
w12439 <= not w12019 and w12438;
w12440 <= not w12027 and not w12439;
w12441 <= not w12437 and w12440;
w12442 <= not w12027 and not w12441;
w12443 <= b(31) and not w12016;
w12444 <= not w12010 and w12443;
w12445 <= not w12018 and not w12444;
w12446 <= not w12442 and w12445;
w12447 <= not w12018 and not w12446;
w12448 <= b(32) and not w12007;
w12449 <= not w12001 and w12448;
w12450 <= not w12009 and not w12449;
w12451 <= not w12447 and w12450;
w12452 <= not w12009 and not w12451;
w12453 <= b(33) and not w11998;
w12454 <= not w11992 and w12453;
w12455 <= not w12000 and not w12454;
w12456 <= not w12452 and w12455;
w12457 <= not w12000 and not w12456;
w12458 <= b(34) and not w11989;
w12459 <= not w11983 and w12458;
w12460 <= not w11991 and not w12459;
w12461 <= not w12457 and w12460;
w12462 <= not w11991 and not w12461;
w12463 <= b(35) and not w11980;
w12464 <= not w11974 and w12463;
w12465 <= not w11982 and not w12464;
w12466 <= not w12462 and w12465;
w12467 <= not w11982 and not w12466;
w12468 <= b(36) and not w11971;
w12469 <= not w11965 and w12468;
w12470 <= not w11973 and not w12469;
w12471 <= not w12467 and w12470;
w12472 <= not w11973 and not w12471;
w12473 <= b(37) and not w11962;
w12474 <= not w11956 and w12473;
w12475 <= not w11964 and not w12474;
w12476 <= not w12472 and w12475;
w12477 <= not w11964 and not w12476;
w12478 <= b(38) and not w11953;
w12479 <= not w11947 and w12478;
w12480 <= not w11955 and not w12479;
w12481 <= not w12477 and w12480;
w12482 <= not w11955 and not w12481;
w12483 <= b(39) and not w11944;
w12484 <= not w11938 and w12483;
w12485 <= not w11946 and not w12484;
w12486 <= not w12482 and w12485;
w12487 <= not w11946 and not w12486;
w12488 <= b(40) and not w11935;
w12489 <= not w11929 and w12488;
w12490 <= not w11937 and not w12489;
w12491 <= not w12487 and w12490;
w12492 <= not w11937 and not w12491;
w12493 <= not w11378 and not w11928;
w12494 <= not w11380 and w11924;
w12495 <= not w11920 and w12494;
w12496 <= not w11921 and not w11924;
w12497 <= not w12495 and not w12496;
w12498 <= w11928 and not w12497;
w12499 <= not w12493 and not w12498;
w12500 <= not b(41) and not w12499;
w12501 <= b(41) and not w12493;
w12502 <= not w12498 and w12501;
w12503 <= w33 and w44;
w12504 <= w81 and w12503;
w12505 <= not w12502 and w12504;
w12506 <= not w12500 and w12505;
w12507 <= not w12492 and w12506;
w12508 <= w11927 and not w12499;
w12509 <= not w12507 and not w12508;
w12510 <= not w11946 and w12490;
w12511 <= not w12486 and w12510;
w12512 <= not w12487 and not w12490;
w12513 <= not w12511 and not w12512;
w12514 <= not w12509 and not w12513;
w12515 <= not w11936 and not w12508;
w12516 <= not w12507 and w12515;
w12517 <= not w12514 and not w12516;
w12518 <= not w11937 and not w12502;
w12519 <= not w12500 and w12518;
w12520 <= not w12491 and w12519;
w12521 <= not w12500 and not w12502;
w12522 <= not w12492 and not w12521;
w12523 <= not w12520 and not w12522;
w12524 <= not w12509 and not w12523;
w12525 <= not w12499 and not w12508;
w12526 <= not w12507 and w12525;
w12527 <= not w12524 and not w12526;
w12528 <= not b(42) and not w12527;
w12529 <= not b(41) and not w12517;
w12530 <= not w11955 and w12485;
w12531 <= not w12481 and w12530;
w12532 <= not w12482 and not w12485;
w12533 <= not w12531 and not w12532;
w12534 <= not w12509 and not w12533;
w12535 <= not w11945 and not w12508;
w12536 <= not w12507 and w12535;
w12537 <= not w12534 and not w12536;
w12538 <= not b(40) and not w12537;
w12539 <= not w11964 and w12480;
w12540 <= not w12476 and w12539;
w12541 <= not w12477 and not w12480;
w12542 <= not w12540 and not w12541;
w12543 <= not w12509 and not w12542;
w12544 <= not w11954 and not w12508;
w12545 <= not w12507 and w12544;
w12546 <= not w12543 and not w12545;
w12547 <= not b(39) and not w12546;
w12548 <= not w11973 and w12475;
w12549 <= not w12471 and w12548;
w12550 <= not w12472 and not w12475;
w12551 <= not w12549 and not w12550;
w12552 <= not w12509 and not w12551;
w12553 <= not w11963 and not w12508;
w12554 <= not w12507 and w12553;
w12555 <= not w12552 and not w12554;
w12556 <= not b(38) and not w12555;
w12557 <= not w11982 and w12470;
w12558 <= not w12466 and w12557;
w12559 <= not w12467 and not w12470;
w12560 <= not w12558 and not w12559;
w12561 <= not w12509 and not w12560;
w12562 <= not w11972 and not w12508;
w12563 <= not w12507 and w12562;
w12564 <= not w12561 and not w12563;
w12565 <= not b(37) and not w12564;
w12566 <= not w11991 and w12465;
w12567 <= not w12461 and w12566;
w12568 <= not w12462 and not w12465;
w12569 <= not w12567 and not w12568;
w12570 <= not w12509 and not w12569;
w12571 <= not w11981 and not w12508;
w12572 <= not w12507 and w12571;
w12573 <= not w12570 and not w12572;
w12574 <= not b(36) and not w12573;
w12575 <= not w12000 and w12460;
w12576 <= not w12456 and w12575;
w12577 <= not w12457 and not w12460;
w12578 <= not w12576 and not w12577;
w12579 <= not w12509 and not w12578;
w12580 <= not w11990 and not w12508;
w12581 <= not w12507 and w12580;
w12582 <= not w12579 and not w12581;
w12583 <= not b(35) and not w12582;
w12584 <= not w12009 and w12455;
w12585 <= not w12451 and w12584;
w12586 <= not w12452 and not w12455;
w12587 <= not w12585 and not w12586;
w12588 <= not w12509 and not w12587;
w12589 <= not w11999 and not w12508;
w12590 <= not w12507 and w12589;
w12591 <= not w12588 and not w12590;
w12592 <= not b(34) and not w12591;
w12593 <= not w12018 and w12450;
w12594 <= not w12446 and w12593;
w12595 <= not w12447 and not w12450;
w12596 <= not w12594 and not w12595;
w12597 <= not w12509 and not w12596;
w12598 <= not w12008 and not w12508;
w12599 <= not w12507 and w12598;
w12600 <= not w12597 and not w12599;
w12601 <= not b(33) and not w12600;
w12602 <= not w12027 and w12445;
w12603 <= not w12441 and w12602;
w12604 <= not w12442 and not w12445;
w12605 <= not w12603 and not w12604;
w12606 <= not w12509 and not w12605;
w12607 <= not w12017 and not w12508;
w12608 <= not w12507 and w12607;
w12609 <= not w12606 and not w12608;
w12610 <= not b(32) and not w12609;
w12611 <= not w12036 and w12440;
w12612 <= not w12436 and w12611;
w12613 <= not w12437 and not w12440;
w12614 <= not w12612 and not w12613;
w12615 <= not w12509 and not w12614;
w12616 <= not w12026 and not w12508;
w12617 <= not w12507 and w12616;
w12618 <= not w12615 and not w12617;
w12619 <= not b(31) and not w12618;
w12620 <= not w12045 and w12435;
w12621 <= not w12431 and w12620;
w12622 <= not w12432 and not w12435;
w12623 <= not w12621 and not w12622;
w12624 <= not w12509 and not w12623;
w12625 <= not w12035 and not w12508;
w12626 <= not w12507 and w12625;
w12627 <= not w12624 and not w12626;
w12628 <= not b(30) and not w12627;
w12629 <= not w12054 and w12430;
w12630 <= not w12426 and w12629;
w12631 <= not w12427 and not w12430;
w12632 <= not w12630 and not w12631;
w12633 <= not w12509 and not w12632;
w12634 <= not w12044 and not w12508;
w12635 <= not w12507 and w12634;
w12636 <= not w12633 and not w12635;
w12637 <= not b(29) and not w12636;
w12638 <= not w12063 and w12425;
w12639 <= not w12421 and w12638;
w12640 <= not w12422 and not w12425;
w12641 <= not w12639 and not w12640;
w12642 <= not w12509 and not w12641;
w12643 <= not w12053 and not w12508;
w12644 <= not w12507 and w12643;
w12645 <= not w12642 and not w12644;
w12646 <= not b(28) and not w12645;
w12647 <= not w12072 and w12420;
w12648 <= not w12416 and w12647;
w12649 <= not w12417 and not w12420;
w12650 <= not w12648 and not w12649;
w12651 <= not w12509 and not w12650;
w12652 <= not w12062 and not w12508;
w12653 <= not w12507 and w12652;
w12654 <= not w12651 and not w12653;
w12655 <= not b(27) and not w12654;
w12656 <= not w12081 and w12415;
w12657 <= not w12411 and w12656;
w12658 <= not w12412 and not w12415;
w12659 <= not w12657 and not w12658;
w12660 <= not w12509 and not w12659;
w12661 <= not w12071 and not w12508;
w12662 <= not w12507 and w12661;
w12663 <= not w12660 and not w12662;
w12664 <= not b(26) and not w12663;
w12665 <= not w12090 and w12410;
w12666 <= not w12406 and w12665;
w12667 <= not w12407 and not w12410;
w12668 <= not w12666 and not w12667;
w12669 <= not w12509 and not w12668;
w12670 <= not w12080 and not w12508;
w12671 <= not w12507 and w12670;
w12672 <= not w12669 and not w12671;
w12673 <= not b(25) and not w12672;
w12674 <= not w12099 and w12405;
w12675 <= not w12401 and w12674;
w12676 <= not w12402 and not w12405;
w12677 <= not w12675 and not w12676;
w12678 <= not w12509 and not w12677;
w12679 <= not w12089 and not w12508;
w12680 <= not w12507 and w12679;
w12681 <= not w12678 and not w12680;
w12682 <= not b(24) and not w12681;
w12683 <= not w12108 and w12400;
w12684 <= not w12396 and w12683;
w12685 <= not w12397 and not w12400;
w12686 <= not w12684 and not w12685;
w12687 <= not w12509 and not w12686;
w12688 <= not w12098 and not w12508;
w12689 <= not w12507 and w12688;
w12690 <= not w12687 and not w12689;
w12691 <= not b(23) and not w12690;
w12692 <= not w12117 and w12395;
w12693 <= not w12391 and w12692;
w12694 <= not w12392 and not w12395;
w12695 <= not w12693 and not w12694;
w12696 <= not w12509 and not w12695;
w12697 <= not w12107 and not w12508;
w12698 <= not w12507 and w12697;
w12699 <= not w12696 and not w12698;
w12700 <= not b(22) and not w12699;
w12701 <= not w12126 and w12390;
w12702 <= not w12386 and w12701;
w12703 <= not w12387 and not w12390;
w12704 <= not w12702 and not w12703;
w12705 <= not w12509 and not w12704;
w12706 <= not w12116 and not w12508;
w12707 <= not w12507 and w12706;
w12708 <= not w12705 and not w12707;
w12709 <= not b(21) and not w12708;
w12710 <= not w12135 and w12385;
w12711 <= not w12381 and w12710;
w12712 <= not w12382 and not w12385;
w12713 <= not w12711 and not w12712;
w12714 <= not w12509 and not w12713;
w12715 <= not w12125 and not w12508;
w12716 <= not w12507 and w12715;
w12717 <= not w12714 and not w12716;
w12718 <= not b(20) and not w12717;
w12719 <= not w12144 and w12380;
w12720 <= not w12376 and w12719;
w12721 <= not w12377 and not w12380;
w12722 <= not w12720 and not w12721;
w12723 <= not w12509 and not w12722;
w12724 <= not w12134 and not w12508;
w12725 <= not w12507 and w12724;
w12726 <= not w12723 and not w12725;
w12727 <= not b(19) and not w12726;
w12728 <= not w12153 and w12375;
w12729 <= not w12371 and w12728;
w12730 <= not w12372 and not w12375;
w12731 <= not w12729 and not w12730;
w12732 <= not w12509 and not w12731;
w12733 <= not w12143 and not w12508;
w12734 <= not w12507 and w12733;
w12735 <= not w12732 and not w12734;
w12736 <= not b(18) and not w12735;
w12737 <= not w12162 and w12370;
w12738 <= not w12366 and w12737;
w12739 <= not w12367 and not w12370;
w12740 <= not w12738 and not w12739;
w12741 <= not w12509 and not w12740;
w12742 <= not w12152 and not w12508;
w12743 <= not w12507 and w12742;
w12744 <= not w12741 and not w12743;
w12745 <= not b(17) and not w12744;
w12746 <= not w12171 and w12365;
w12747 <= not w12361 and w12746;
w12748 <= not w12362 and not w12365;
w12749 <= not w12747 and not w12748;
w12750 <= not w12509 and not w12749;
w12751 <= not w12161 and not w12508;
w12752 <= not w12507 and w12751;
w12753 <= not w12750 and not w12752;
w12754 <= not b(16) and not w12753;
w12755 <= not w12180 and w12360;
w12756 <= not w12356 and w12755;
w12757 <= not w12357 and not w12360;
w12758 <= not w12756 and not w12757;
w12759 <= not w12509 and not w12758;
w12760 <= not w12170 and not w12508;
w12761 <= not w12507 and w12760;
w12762 <= not w12759 and not w12761;
w12763 <= not b(15) and not w12762;
w12764 <= not w12189 and w12355;
w12765 <= not w12351 and w12764;
w12766 <= not w12352 and not w12355;
w12767 <= not w12765 and not w12766;
w12768 <= not w12509 and not w12767;
w12769 <= not w12179 and not w12508;
w12770 <= not w12507 and w12769;
w12771 <= not w12768 and not w12770;
w12772 <= not b(14) and not w12771;
w12773 <= not w12198 and w12350;
w12774 <= not w12346 and w12773;
w12775 <= not w12347 and not w12350;
w12776 <= not w12774 and not w12775;
w12777 <= not w12509 and not w12776;
w12778 <= not w12188 and not w12508;
w12779 <= not w12507 and w12778;
w12780 <= not w12777 and not w12779;
w12781 <= not b(13) and not w12780;
w12782 <= not w12207 and w12345;
w12783 <= not w12341 and w12782;
w12784 <= not w12342 and not w12345;
w12785 <= not w12783 and not w12784;
w12786 <= not w12509 and not w12785;
w12787 <= not w12197 and not w12508;
w12788 <= not w12507 and w12787;
w12789 <= not w12786 and not w12788;
w12790 <= not b(12) and not w12789;
w12791 <= not w12216 and w12340;
w12792 <= not w12336 and w12791;
w12793 <= not w12337 and not w12340;
w12794 <= not w12792 and not w12793;
w12795 <= not w12509 and not w12794;
w12796 <= not w12206 and not w12508;
w12797 <= not w12507 and w12796;
w12798 <= not w12795 and not w12797;
w12799 <= not b(11) and not w12798;
w12800 <= not w12225 and w12335;
w12801 <= not w12331 and w12800;
w12802 <= not w12332 and not w12335;
w12803 <= not w12801 and not w12802;
w12804 <= not w12509 and not w12803;
w12805 <= not w12215 and not w12508;
w12806 <= not w12507 and w12805;
w12807 <= not w12804 and not w12806;
w12808 <= not b(10) and not w12807;
w12809 <= not w12234 and w12330;
w12810 <= not w12326 and w12809;
w12811 <= not w12327 and not w12330;
w12812 <= not w12810 and not w12811;
w12813 <= not w12509 and not w12812;
w12814 <= not w12224 and not w12508;
w12815 <= not w12507 and w12814;
w12816 <= not w12813 and not w12815;
w12817 <= not b(9) and not w12816;
w12818 <= not w12243 and w12325;
w12819 <= not w12321 and w12818;
w12820 <= not w12322 and not w12325;
w12821 <= not w12819 and not w12820;
w12822 <= not w12509 and not w12821;
w12823 <= not w12233 and not w12508;
w12824 <= not w12507 and w12823;
w12825 <= not w12822 and not w12824;
w12826 <= not b(8) and not w12825;
w12827 <= not w12252 and w12320;
w12828 <= not w12316 and w12827;
w12829 <= not w12317 and not w12320;
w12830 <= not w12828 and not w12829;
w12831 <= not w12509 and not w12830;
w12832 <= not w12242 and not w12508;
w12833 <= not w12507 and w12832;
w12834 <= not w12831 and not w12833;
w12835 <= not b(7) and not w12834;
w12836 <= not w12261 and w12315;
w12837 <= not w12311 and w12836;
w12838 <= not w12312 and not w12315;
w12839 <= not w12837 and not w12838;
w12840 <= not w12509 and not w12839;
w12841 <= not w12251 and not w12508;
w12842 <= not w12507 and w12841;
w12843 <= not w12840 and not w12842;
w12844 <= not b(6) and not w12843;
w12845 <= not w12270 and w12310;
w12846 <= not w12306 and w12845;
w12847 <= not w12307 and not w12310;
w12848 <= not w12846 and not w12847;
w12849 <= not w12509 and not w12848;
w12850 <= not w12260 and not w12508;
w12851 <= not w12507 and w12850;
w12852 <= not w12849 and not w12851;
w12853 <= not b(5) and not w12852;
w12854 <= not w12278 and w12305;
w12855 <= not w12301 and w12854;
w12856 <= not w12302 and not w12305;
w12857 <= not w12855 and not w12856;
w12858 <= not w12509 and not w12857;
w12859 <= not w12269 and not w12508;
w12860 <= not w12507 and w12859;
w12861 <= not w12858 and not w12860;
w12862 <= not b(4) and not w12861;
w12863 <= not w12296 and w12300;
w12864 <= not w12295 and w12863;
w12865 <= not w12297 and not w12300;
w12866 <= not w12864 and not w12865;
w12867 <= not w12509 and not w12866;
w12868 <= not w12277 and not w12508;
w12869 <= not w12507 and w12868;
w12870 <= not w12867 and not w12869;
w12871 <= not b(3) and not w12870;
w12872 <= not w12292 and w12294;
w12873 <= not w12290 and w12872;
w12874 <= not w12295 and not w12873;
w12875 <= not w12509 and w12874;
w12876 <= not w12289 and not w12508;
w12877 <= not w12507 and w12876;
w12878 <= not w12875 and not w12877;
w12879 <= not b(2) and not w12878;
w12880 <= b(0) and not w12509;
w12881 <= a(22) and not w12880;
w12882 <= w12294 and not w12509;
w12883 <= not w12881 and not w12882;
w12884 <= b(1) and not w12883;
w12885 <= not b(1) and not w12882;
w12886 <= not w12881 and w12885;
w12887 <= not w12884 and not w12886;
w12888 <= not a(21) and b(0);
w12889 <= not w12887 and not w12888;
w12890 <= not b(1) and not w12883;
w12891 <= not w12889 and not w12890;
w12892 <= b(2) and not w12877;
w12893 <= not w12875 and w12892;
w12894 <= not w12879 and not w12893;
w12895 <= not w12891 and w12894;
w12896 <= not w12879 and not w12895;
w12897 <= b(3) and not w12869;
w12898 <= not w12867 and w12897;
w12899 <= not w12871 and not w12898;
w12900 <= not w12896 and w12899;
w12901 <= not w12871 and not w12900;
w12902 <= b(4) and not w12860;
w12903 <= not w12858 and w12902;
w12904 <= not w12862 and not w12903;
w12905 <= not w12901 and w12904;
w12906 <= not w12862 and not w12905;
w12907 <= b(5) and not w12851;
w12908 <= not w12849 and w12907;
w12909 <= not w12853 and not w12908;
w12910 <= not w12906 and w12909;
w12911 <= not w12853 and not w12910;
w12912 <= b(6) and not w12842;
w12913 <= not w12840 and w12912;
w12914 <= not w12844 and not w12913;
w12915 <= not w12911 and w12914;
w12916 <= not w12844 and not w12915;
w12917 <= b(7) and not w12833;
w12918 <= not w12831 and w12917;
w12919 <= not w12835 and not w12918;
w12920 <= not w12916 and w12919;
w12921 <= not w12835 and not w12920;
w12922 <= b(8) and not w12824;
w12923 <= not w12822 and w12922;
w12924 <= not w12826 and not w12923;
w12925 <= not w12921 and w12924;
w12926 <= not w12826 and not w12925;
w12927 <= b(9) and not w12815;
w12928 <= not w12813 and w12927;
w12929 <= not w12817 and not w12928;
w12930 <= not w12926 and w12929;
w12931 <= not w12817 and not w12930;
w12932 <= b(10) and not w12806;
w12933 <= not w12804 and w12932;
w12934 <= not w12808 and not w12933;
w12935 <= not w12931 and w12934;
w12936 <= not w12808 and not w12935;
w12937 <= b(11) and not w12797;
w12938 <= not w12795 and w12937;
w12939 <= not w12799 and not w12938;
w12940 <= not w12936 and w12939;
w12941 <= not w12799 and not w12940;
w12942 <= b(12) and not w12788;
w12943 <= not w12786 and w12942;
w12944 <= not w12790 and not w12943;
w12945 <= not w12941 and w12944;
w12946 <= not w12790 and not w12945;
w12947 <= b(13) and not w12779;
w12948 <= not w12777 and w12947;
w12949 <= not w12781 and not w12948;
w12950 <= not w12946 and w12949;
w12951 <= not w12781 and not w12950;
w12952 <= b(14) and not w12770;
w12953 <= not w12768 and w12952;
w12954 <= not w12772 and not w12953;
w12955 <= not w12951 and w12954;
w12956 <= not w12772 and not w12955;
w12957 <= b(15) and not w12761;
w12958 <= not w12759 and w12957;
w12959 <= not w12763 and not w12958;
w12960 <= not w12956 and w12959;
w12961 <= not w12763 and not w12960;
w12962 <= b(16) and not w12752;
w12963 <= not w12750 and w12962;
w12964 <= not w12754 and not w12963;
w12965 <= not w12961 and w12964;
w12966 <= not w12754 and not w12965;
w12967 <= b(17) and not w12743;
w12968 <= not w12741 and w12967;
w12969 <= not w12745 and not w12968;
w12970 <= not w12966 and w12969;
w12971 <= not w12745 and not w12970;
w12972 <= b(18) and not w12734;
w12973 <= not w12732 and w12972;
w12974 <= not w12736 and not w12973;
w12975 <= not w12971 and w12974;
w12976 <= not w12736 and not w12975;
w12977 <= b(19) and not w12725;
w12978 <= not w12723 and w12977;
w12979 <= not w12727 and not w12978;
w12980 <= not w12976 and w12979;
w12981 <= not w12727 and not w12980;
w12982 <= b(20) and not w12716;
w12983 <= not w12714 and w12982;
w12984 <= not w12718 and not w12983;
w12985 <= not w12981 and w12984;
w12986 <= not w12718 and not w12985;
w12987 <= b(21) and not w12707;
w12988 <= not w12705 and w12987;
w12989 <= not w12709 and not w12988;
w12990 <= not w12986 and w12989;
w12991 <= not w12709 and not w12990;
w12992 <= b(22) and not w12698;
w12993 <= not w12696 and w12992;
w12994 <= not w12700 and not w12993;
w12995 <= not w12991 and w12994;
w12996 <= not w12700 and not w12995;
w12997 <= b(23) and not w12689;
w12998 <= not w12687 and w12997;
w12999 <= not w12691 and not w12998;
w13000 <= not w12996 and w12999;
w13001 <= not w12691 and not w13000;
w13002 <= b(24) and not w12680;
w13003 <= not w12678 and w13002;
w13004 <= not w12682 and not w13003;
w13005 <= not w13001 and w13004;
w13006 <= not w12682 and not w13005;
w13007 <= b(25) and not w12671;
w13008 <= not w12669 and w13007;
w13009 <= not w12673 and not w13008;
w13010 <= not w13006 and w13009;
w13011 <= not w12673 and not w13010;
w13012 <= b(26) and not w12662;
w13013 <= not w12660 and w13012;
w13014 <= not w12664 and not w13013;
w13015 <= not w13011 and w13014;
w13016 <= not w12664 and not w13015;
w13017 <= b(27) and not w12653;
w13018 <= not w12651 and w13017;
w13019 <= not w12655 and not w13018;
w13020 <= not w13016 and w13019;
w13021 <= not w12655 and not w13020;
w13022 <= b(28) and not w12644;
w13023 <= not w12642 and w13022;
w13024 <= not w12646 and not w13023;
w13025 <= not w13021 and w13024;
w13026 <= not w12646 and not w13025;
w13027 <= b(29) and not w12635;
w13028 <= not w12633 and w13027;
w13029 <= not w12637 and not w13028;
w13030 <= not w13026 and w13029;
w13031 <= not w12637 and not w13030;
w13032 <= b(30) and not w12626;
w13033 <= not w12624 and w13032;
w13034 <= not w12628 and not w13033;
w13035 <= not w13031 and w13034;
w13036 <= not w12628 and not w13035;
w13037 <= b(31) and not w12617;
w13038 <= not w12615 and w13037;
w13039 <= not w12619 and not w13038;
w13040 <= not w13036 and w13039;
w13041 <= not w12619 and not w13040;
w13042 <= b(32) and not w12608;
w13043 <= not w12606 and w13042;
w13044 <= not w12610 and not w13043;
w13045 <= not w13041 and w13044;
w13046 <= not w12610 and not w13045;
w13047 <= b(33) and not w12599;
w13048 <= not w12597 and w13047;
w13049 <= not w12601 and not w13048;
w13050 <= not w13046 and w13049;
w13051 <= not w12601 and not w13050;
w13052 <= b(34) and not w12590;
w13053 <= not w12588 and w13052;
w13054 <= not w12592 and not w13053;
w13055 <= not w13051 and w13054;
w13056 <= not w12592 and not w13055;
w13057 <= b(35) and not w12581;
w13058 <= not w12579 and w13057;
w13059 <= not w12583 and not w13058;
w13060 <= not w13056 and w13059;
w13061 <= not w12583 and not w13060;
w13062 <= b(36) and not w12572;
w13063 <= not w12570 and w13062;
w13064 <= not w12574 and not w13063;
w13065 <= not w13061 and w13064;
w13066 <= not w12574 and not w13065;
w13067 <= b(37) and not w12563;
w13068 <= not w12561 and w13067;
w13069 <= not w12565 and not w13068;
w13070 <= not w13066 and w13069;
w13071 <= not w12565 and not w13070;
w13072 <= b(38) and not w12554;
w13073 <= not w12552 and w13072;
w13074 <= not w12556 and not w13073;
w13075 <= not w13071 and w13074;
w13076 <= not w12556 and not w13075;
w13077 <= b(39) and not w12545;
w13078 <= not w12543 and w13077;
w13079 <= not w12547 and not w13078;
w13080 <= not w13076 and w13079;
w13081 <= not w12547 and not w13080;
w13082 <= b(40) and not w12536;
w13083 <= not w12534 and w13082;
w13084 <= not w12538 and not w13083;
w13085 <= not w13081 and w13084;
w13086 <= not w12538 and not w13085;
w13087 <= b(41) and not w12516;
w13088 <= not w12514 and w13087;
w13089 <= not w12529 and not w13088;
w13090 <= not w13086 and w13089;
w13091 <= not w12529 and not w13090;
w13092 <= b(42) and not w12526;
w13093 <= not w12524 and w13092;
w13094 <= not w12528 and not w13093;
w13095 <= not w13091 and w13094;
w13096 <= not w12528 and not w13095;
w13097 <= w161 and w163;
w13098 <= w151 and w13097;
w13099 <= not w13096 and w13098;
w13100 <= not w12517 and not w13099;
w13101 <= not w12538 and w13089;
w13102 <= not w13085 and w13101;
w13103 <= not w13086 and not w13089;
w13104 <= not w13102 and not w13103;
w13105 <= w13098 and not w13104;
w13106 <= not w13096 and w13105;
w13107 <= not w13100 and not w13106;
w13108 <= not b(42) and not w13107;
w13109 <= not w12537 and not w13099;
w13110 <= not w12547 and w13084;
w13111 <= not w13080 and w13110;
w13112 <= not w13081 and not w13084;
w13113 <= not w13111 and not w13112;
w13114 <= w13098 and not w13113;
w13115 <= not w13096 and w13114;
w13116 <= not w13109 and not w13115;
w13117 <= not b(41) and not w13116;
w13118 <= not w12546 and not w13099;
w13119 <= not w12556 and w13079;
w13120 <= not w13075 and w13119;
w13121 <= not w13076 and not w13079;
w13122 <= not w13120 and not w13121;
w13123 <= w13098 and not w13122;
w13124 <= not w13096 and w13123;
w13125 <= not w13118 and not w13124;
w13126 <= not b(40) and not w13125;
w13127 <= not w12555 and not w13099;
w13128 <= not w12565 and w13074;
w13129 <= not w13070 and w13128;
w13130 <= not w13071 and not w13074;
w13131 <= not w13129 and not w13130;
w13132 <= w13098 and not w13131;
w13133 <= not w13096 and w13132;
w13134 <= not w13127 and not w13133;
w13135 <= not b(39) and not w13134;
w13136 <= not w12564 and not w13099;
w13137 <= not w12574 and w13069;
w13138 <= not w13065 and w13137;
w13139 <= not w13066 and not w13069;
w13140 <= not w13138 and not w13139;
w13141 <= w13098 and not w13140;
w13142 <= not w13096 and w13141;
w13143 <= not w13136 and not w13142;
w13144 <= not b(38) and not w13143;
w13145 <= not w12573 and not w13099;
w13146 <= not w12583 and w13064;
w13147 <= not w13060 and w13146;
w13148 <= not w13061 and not w13064;
w13149 <= not w13147 and not w13148;
w13150 <= w13098 and not w13149;
w13151 <= not w13096 and w13150;
w13152 <= not w13145 and not w13151;
w13153 <= not b(37) and not w13152;
w13154 <= not w12582 and not w13099;
w13155 <= not w12592 and w13059;
w13156 <= not w13055 and w13155;
w13157 <= not w13056 and not w13059;
w13158 <= not w13156 and not w13157;
w13159 <= w13098 and not w13158;
w13160 <= not w13096 and w13159;
w13161 <= not w13154 and not w13160;
w13162 <= not b(36) and not w13161;
w13163 <= not w12591 and not w13099;
w13164 <= not w12601 and w13054;
w13165 <= not w13050 and w13164;
w13166 <= not w13051 and not w13054;
w13167 <= not w13165 and not w13166;
w13168 <= w13098 and not w13167;
w13169 <= not w13096 and w13168;
w13170 <= not w13163 and not w13169;
w13171 <= not b(35) and not w13170;
w13172 <= not w12600 and not w13099;
w13173 <= not w12610 and w13049;
w13174 <= not w13045 and w13173;
w13175 <= not w13046 and not w13049;
w13176 <= not w13174 and not w13175;
w13177 <= w13098 and not w13176;
w13178 <= not w13096 and w13177;
w13179 <= not w13172 and not w13178;
w13180 <= not b(34) and not w13179;
w13181 <= not w12609 and not w13099;
w13182 <= not w12619 and w13044;
w13183 <= not w13040 and w13182;
w13184 <= not w13041 and not w13044;
w13185 <= not w13183 and not w13184;
w13186 <= w13098 and not w13185;
w13187 <= not w13096 and w13186;
w13188 <= not w13181 and not w13187;
w13189 <= not b(33) and not w13188;
w13190 <= not w12618 and not w13099;
w13191 <= not w12628 and w13039;
w13192 <= not w13035 and w13191;
w13193 <= not w13036 and not w13039;
w13194 <= not w13192 and not w13193;
w13195 <= w13098 and not w13194;
w13196 <= not w13096 and w13195;
w13197 <= not w13190 and not w13196;
w13198 <= not b(32) and not w13197;
w13199 <= not w12627 and not w13099;
w13200 <= not w12637 and w13034;
w13201 <= not w13030 and w13200;
w13202 <= not w13031 and not w13034;
w13203 <= not w13201 and not w13202;
w13204 <= w13098 and not w13203;
w13205 <= not w13096 and w13204;
w13206 <= not w13199 and not w13205;
w13207 <= not b(31) and not w13206;
w13208 <= not w12636 and not w13099;
w13209 <= not w12646 and w13029;
w13210 <= not w13025 and w13209;
w13211 <= not w13026 and not w13029;
w13212 <= not w13210 and not w13211;
w13213 <= w13098 and not w13212;
w13214 <= not w13096 and w13213;
w13215 <= not w13208 and not w13214;
w13216 <= not b(30) and not w13215;
w13217 <= not w12645 and not w13099;
w13218 <= not w12655 and w13024;
w13219 <= not w13020 and w13218;
w13220 <= not w13021 and not w13024;
w13221 <= not w13219 and not w13220;
w13222 <= w13098 and not w13221;
w13223 <= not w13096 and w13222;
w13224 <= not w13217 and not w13223;
w13225 <= not b(29) and not w13224;
w13226 <= not w12654 and not w13099;
w13227 <= not w12664 and w13019;
w13228 <= not w13015 and w13227;
w13229 <= not w13016 and not w13019;
w13230 <= not w13228 and not w13229;
w13231 <= w13098 and not w13230;
w13232 <= not w13096 and w13231;
w13233 <= not w13226 and not w13232;
w13234 <= not b(28) and not w13233;
w13235 <= not w12663 and not w13099;
w13236 <= not w12673 and w13014;
w13237 <= not w13010 and w13236;
w13238 <= not w13011 and not w13014;
w13239 <= not w13237 and not w13238;
w13240 <= w13098 and not w13239;
w13241 <= not w13096 and w13240;
w13242 <= not w13235 and not w13241;
w13243 <= not b(27) and not w13242;
w13244 <= not w12672 and not w13099;
w13245 <= not w12682 and w13009;
w13246 <= not w13005 and w13245;
w13247 <= not w13006 and not w13009;
w13248 <= not w13246 and not w13247;
w13249 <= w13098 and not w13248;
w13250 <= not w13096 and w13249;
w13251 <= not w13244 and not w13250;
w13252 <= not b(26) and not w13251;
w13253 <= not w12681 and not w13099;
w13254 <= not w12691 and w13004;
w13255 <= not w13000 and w13254;
w13256 <= not w13001 and not w13004;
w13257 <= not w13255 and not w13256;
w13258 <= w13098 and not w13257;
w13259 <= not w13096 and w13258;
w13260 <= not w13253 and not w13259;
w13261 <= not b(25) and not w13260;
w13262 <= not w12690 and not w13099;
w13263 <= not w12700 and w12999;
w13264 <= not w12995 and w13263;
w13265 <= not w12996 and not w12999;
w13266 <= not w13264 and not w13265;
w13267 <= w13098 and not w13266;
w13268 <= not w13096 and w13267;
w13269 <= not w13262 and not w13268;
w13270 <= not b(24) and not w13269;
w13271 <= not w12699 and not w13099;
w13272 <= not w12709 and w12994;
w13273 <= not w12990 and w13272;
w13274 <= not w12991 and not w12994;
w13275 <= not w13273 and not w13274;
w13276 <= w13098 and not w13275;
w13277 <= not w13096 and w13276;
w13278 <= not w13271 and not w13277;
w13279 <= not b(23) and not w13278;
w13280 <= not w12708 and not w13099;
w13281 <= not w12718 and w12989;
w13282 <= not w12985 and w13281;
w13283 <= not w12986 and not w12989;
w13284 <= not w13282 and not w13283;
w13285 <= w13098 and not w13284;
w13286 <= not w13096 and w13285;
w13287 <= not w13280 and not w13286;
w13288 <= not b(22) and not w13287;
w13289 <= not w12717 and not w13099;
w13290 <= not w12727 and w12984;
w13291 <= not w12980 and w13290;
w13292 <= not w12981 and not w12984;
w13293 <= not w13291 and not w13292;
w13294 <= w13098 and not w13293;
w13295 <= not w13096 and w13294;
w13296 <= not w13289 and not w13295;
w13297 <= not b(21) and not w13296;
w13298 <= not w12726 and not w13099;
w13299 <= not w12736 and w12979;
w13300 <= not w12975 and w13299;
w13301 <= not w12976 and not w12979;
w13302 <= not w13300 and not w13301;
w13303 <= w13098 and not w13302;
w13304 <= not w13096 and w13303;
w13305 <= not w13298 and not w13304;
w13306 <= not b(20) and not w13305;
w13307 <= not w12735 and not w13099;
w13308 <= not w12745 and w12974;
w13309 <= not w12970 and w13308;
w13310 <= not w12971 and not w12974;
w13311 <= not w13309 and not w13310;
w13312 <= w13098 and not w13311;
w13313 <= not w13096 and w13312;
w13314 <= not w13307 and not w13313;
w13315 <= not b(19) and not w13314;
w13316 <= not w12744 and not w13099;
w13317 <= not w12754 and w12969;
w13318 <= not w12965 and w13317;
w13319 <= not w12966 and not w12969;
w13320 <= not w13318 and not w13319;
w13321 <= w13098 and not w13320;
w13322 <= not w13096 and w13321;
w13323 <= not w13316 and not w13322;
w13324 <= not b(18) and not w13323;
w13325 <= not w12753 and not w13099;
w13326 <= not w12763 and w12964;
w13327 <= not w12960 and w13326;
w13328 <= not w12961 and not w12964;
w13329 <= not w13327 and not w13328;
w13330 <= w13098 and not w13329;
w13331 <= not w13096 and w13330;
w13332 <= not w13325 and not w13331;
w13333 <= not b(17) and not w13332;
w13334 <= not w12762 and not w13099;
w13335 <= not w12772 and w12959;
w13336 <= not w12955 and w13335;
w13337 <= not w12956 and not w12959;
w13338 <= not w13336 and not w13337;
w13339 <= w13098 and not w13338;
w13340 <= not w13096 and w13339;
w13341 <= not w13334 and not w13340;
w13342 <= not b(16) and not w13341;
w13343 <= not w12771 and not w13099;
w13344 <= not w12781 and w12954;
w13345 <= not w12950 and w13344;
w13346 <= not w12951 and not w12954;
w13347 <= not w13345 and not w13346;
w13348 <= w13098 and not w13347;
w13349 <= not w13096 and w13348;
w13350 <= not w13343 and not w13349;
w13351 <= not b(15) and not w13350;
w13352 <= not w12780 and not w13099;
w13353 <= not w12790 and w12949;
w13354 <= not w12945 and w13353;
w13355 <= not w12946 and not w12949;
w13356 <= not w13354 and not w13355;
w13357 <= w13098 and not w13356;
w13358 <= not w13096 and w13357;
w13359 <= not w13352 and not w13358;
w13360 <= not b(14) and not w13359;
w13361 <= not w12789 and not w13099;
w13362 <= not w12799 and w12944;
w13363 <= not w12940 and w13362;
w13364 <= not w12941 and not w12944;
w13365 <= not w13363 and not w13364;
w13366 <= w13098 and not w13365;
w13367 <= not w13096 and w13366;
w13368 <= not w13361 and not w13367;
w13369 <= not b(13) and not w13368;
w13370 <= not w12798 and not w13099;
w13371 <= not w12808 and w12939;
w13372 <= not w12935 and w13371;
w13373 <= not w12936 and not w12939;
w13374 <= not w13372 and not w13373;
w13375 <= w13098 and not w13374;
w13376 <= not w13096 and w13375;
w13377 <= not w13370 and not w13376;
w13378 <= not b(12) and not w13377;
w13379 <= not w12807 and not w13099;
w13380 <= not w12817 and w12934;
w13381 <= not w12930 and w13380;
w13382 <= not w12931 and not w12934;
w13383 <= not w13381 and not w13382;
w13384 <= w13098 and not w13383;
w13385 <= not w13096 and w13384;
w13386 <= not w13379 and not w13385;
w13387 <= not b(11) and not w13386;
w13388 <= not w12816 and not w13099;
w13389 <= not w12826 and w12929;
w13390 <= not w12925 and w13389;
w13391 <= not w12926 and not w12929;
w13392 <= not w13390 and not w13391;
w13393 <= w13098 and not w13392;
w13394 <= not w13096 and w13393;
w13395 <= not w13388 and not w13394;
w13396 <= not b(10) and not w13395;
w13397 <= not w12825 and not w13099;
w13398 <= not w12835 and w12924;
w13399 <= not w12920 and w13398;
w13400 <= not w12921 and not w12924;
w13401 <= not w13399 and not w13400;
w13402 <= w13098 and not w13401;
w13403 <= not w13096 and w13402;
w13404 <= not w13397 and not w13403;
w13405 <= not b(9) and not w13404;
w13406 <= not w12834 and not w13099;
w13407 <= not w12844 and w12919;
w13408 <= not w12915 and w13407;
w13409 <= not w12916 and not w12919;
w13410 <= not w13408 and not w13409;
w13411 <= w13098 and not w13410;
w13412 <= not w13096 and w13411;
w13413 <= not w13406 and not w13412;
w13414 <= not b(8) and not w13413;
w13415 <= not w12843 and not w13099;
w13416 <= not w12853 and w12914;
w13417 <= not w12910 and w13416;
w13418 <= not w12911 and not w12914;
w13419 <= not w13417 and not w13418;
w13420 <= w13098 and not w13419;
w13421 <= not w13096 and w13420;
w13422 <= not w13415 and not w13421;
w13423 <= not b(7) and not w13422;
w13424 <= not w12852 and not w13099;
w13425 <= not w12862 and w12909;
w13426 <= not w12905 and w13425;
w13427 <= not w12906 and not w12909;
w13428 <= not w13426 and not w13427;
w13429 <= w13098 and not w13428;
w13430 <= not w13096 and w13429;
w13431 <= not w13424 and not w13430;
w13432 <= not b(6) and not w13431;
w13433 <= not w12861 and not w13099;
w13434 <= not w12871 and w12904;
w13435 <= not w12900 and w13434;
w13436 <= not w12901 and not w12904;
w13437 <= not w13435 and not w13436;
w13438 <= w13098 and not w13437;
w13439 <= not w13096 and w13438;
w13440 <= not w13433 and not w13439;
w13441 <= not b(5) and not w13440;
w13442 <= not w12870 and not w13099;
w13443 <= not w12879 and w12899;
w13444 <= not w12895 and w13443;
w13445 <= not w12896 and not w12899;
w13446 <= not w13444 and not w13445;
w13447 <= w13098 and not w13446;
w13448 <= not w13096 and w13447;
w13449 <= not w13442 and not w13448;
w13450 <= not b(4) and not w13449;
w13451 <= not w12878 and not w13099;
w13452 <= not w12890 and w12894;
w13453 <= not w12889 and w13452;
w13454 <= not w12891 and not w12894;
w13455 <= not w13453 and not w13454;
w13456 <= w13098 and not w13455;
w13457 <= not w13096 and w13456;
w13458 <= not w13451 and not w13457;
w13459 <= not b(3) and not w13458;
w13460 <= not w12883 and not w13099;
w13461 <= not w12886 and w12888;
w13462 <= not w12884 and w13461;
w13463 <= w13098 and not w13462;
w13464 <= not w12889 and w13463;
w13465 <= not w13096 and w13464;
w13466 <= not w13460 and not w13465;
w13467 <= not b(2) and not w13466;
w13468 <= b(0) and not b(43);
w13469 <= w44 and w13468;
w13470 <= w81 and w13469;
w13471 <= not w13096 and w13470;
w13472 <= a(21) and not w13471;
w13473 <= w163 and w12888;
w13474 <= w161 and w13473;
w13475 <= w151 and w13474;
w13476 <= not w13096 and w13475;
w13477 <= not w13472 and not w13476;
w13478 <= b(1) and not w13477;
w13479 <= not b(1) and not w13476;
w13480 <= not w13472 and w13479;
w13481 <= not w13478 and not w13480;
w13482 <= not a(20) and b(0);
w13483 <= not w13481 and not w13482;
w13484 <= not b(1) and not w13477;
w13485 <= not w13483 and not w13484;
w13486 <= b(2) and not w13465;
w13487 <= not w13460 and w13486;
w13488 <= not w13467 and not w13487;
w13489 <= not w13485 and w13488;
w13490 <= not w13467 and not w13489;
w13491 <= b(3) and not w13457;
w13492 <= not w13451 and w13491;
w13493 <= not w13459 and not w13492;
w13494 <= not w13490 and w13493;
w13495 <= not w13459 and not w13494;
w13496 <= b(4) and not w13448;
w13497 <= not w13442 and w13496;
w13498 <= not w13450 and not w13497;
w13499 <= not w13495 and w13498;
w13500 <= not w13450 and not w13499;
w13501 <= b(5) and not w13439;
w13502 <= not w13433 and w13501;
w13503 <= not w13441 and not w13502;
w13504 <= not w13500 and w13503;
w13505 <= not w13441 and not w13504;
w13506 <= b(6) and not w13430;
w13507 <= not w13424 and w13506;
w13508 <= not w13432 and not w13507;
w13509 <= not w13505 and w13508;
w13510 <= not w13432 and not w13509;
w13511 <= b(7) and not w13421;
w13512 <= not w13415 and w13511;
w13513 <= not w13423 and not w13512;
w13514 <= not w13510 and w13513;
w13515 <= not w13423 and not w13514;
w13516 <= b(8) and not w13412;
w13517 <= not w13406 and w13516;
w13518 <= not w13414 and not w13517;
w13519 <= not w13515 and w13518;
w13520 <= not w13414 and not w13519;
w13521 <= b(9) and not w13403;
w13522 <= not w13397 and w13521;
w13523 <= not w13405 and not w13522;
w13524 <= not w13520 and w13523;
w13525 <= not w13405 and not w13524;
w13526 <= b(10) and not w13394;
w13527 <= not w13388 and w13526;
w13528 <= not w13396 and not w13527;
w13529 <= not w13525 and w13528;
w13530 <= not w13396 and not w13529;
w13531 <= b(11) and not w13385;
w13532 <= not w13379 and w13531;
w13533 <= not w13387 and not w13532;
w13534 <= not w13530 and w13533;
w13535 <= not w13387 and not w13534;
w13536 <= b(12) and not w13376;
w13537 <= not w13370 and w13536;
w13538 <= not w13378 and not w13537;
w13539 <= not w13535 and w13538;
w13540 <= not w13378 and not w13539;
w13541 <= b(13) and not w13367;
w13542 <= not w13361 and w13541;
w13543 <= not w13369 and not w13542;
w13544 <= not w13540 and w13543;
w13545 <= not w13369 and not w13544;
w13546 <= b(14) and not w13358;
w13547 <= not w13352 and w13546;
w13548 <= not w13360 and not w13547;
w13549 <= not w13545 and w13548;
w13550 <= not w13360 and not w13549;
w13551 <= b(15) and not w13349;
w13552 <= not w13343 and w13551;
w13553 <= not w13351 and not w13552;
w13554 <= not w13550 and w13553;
w13555 <= not w13351 and not w13554;
w13556 <= b(16) and not w13340;
w13557 <= not w13334 and w13556;
w13558 <= not w13342 and not w13557;
w13559 <= not w13555 and w13558;
w13560 <= not w13342 and not w13559;
w13561 <= b(17) and not w13331;
w13562 <= not w13325 and w13561;
w13563 <= not w13333 and not w13562;
w13564 <= not w13560 and w13563;
w13565 <= not w13333 and not w13564;
w13566 <= b(18) and not w13322;
w13567 <= not w13316 and w13566;
w13568 <= not w13324 and not w13567;
w13569 <= not w13565 and w13568;
w13570 <= not w13324 and not w13569;
w13571 <= b(19) and not w13313;
w13572 <= not w13307 and w13571;
w13573 <= not w13315 and not w13572;
w13574 <= not w13570 and w13573;
w13575 <= not w13315 and not w13574;
w13576 <= b(20) and not w13304;
w13577 <= not w13298 and w13576;
w13578 <= not w13306 and not w13577;
w13579 <= not w13575 and w13578;
w13580 <= not w13306 and not w13579;
w13581 <= b(21) and not w13295;
w13582 <= not w13289 and w13581;
w13583 <= not w13297 and not w13582;
w13584 <= not w13580 and w13583;
w13585 <= not w13297 and not w13584;
w13586 <= b(22) and not w13286;
w13587 <= not w13280 and w13586;
w13588 <= not w13288 and not w13587;
w13589 <= not w13585 and w13588;
w13590 <= not w13288 and not w13589;
w13591 <= b(23) and not w13277;
w13592 <= not w13271 and w13591;
w13593 <= not w13279 and not w13592;
w13594 <= not w13590 and w13593;
w13595 <= not w13279 and not w13594;
w13596 <= b(24) and not w13268;
w13597 <= not w13262 and w13596;
w13598 <= not w13270 and not w13597;
w13599 <= not w13595 and w13598;
w13600 <= not w13270 and not w13599;
w13601 <= b(25) and not w13259;
w13602 <= not w13253 and w13601;
w13603 <= not w13261 and not w13602;
w13604 <= not w13600 and w13603;
w13605 <= not w13261 and not w13604;
w13606 <= b(26) and not w13250;
w13607 <= not w13244 and w13606;
w13608 <= not w13252 and not w13607;
w13609 <= not w13605 and w13608;
w13610 <= not w13252 and not w13609;
w13611 <= b(27) and not w13241;
w13612 <= not w13235 and w13611;
w13613 <= not w13243 and not w13612;
w13614 <= not w13610 and w13613;
w13615 <= not w13243 and not w13614;
w13616 <= b(28) and not w13232;
w13617 <= not w13226 and w13616;
w13618 <= not w13234 and not w13617;
w13619 <= not w13615 and w13618;
w13620 <= not w13234 and not w13619;
w13621 <= b(29) and not w13223;
w13622 <= not w13217 and w13621;
w13623 <= not w13225 and not w13622;
w13624 <= not w13620 and w13623;
w13625 <= not w13225 and not w13624;
w13626 <= b(30) and not w13214;
w13627 <= not w13208 and w13626;
w13628 <= not w13216 and not w13627;
w13629 <= not w13625 and w13628;
w13630 <= not w13216 and not w13629;
w13631 <= b(31) and not w13205;
w13632 <= not w13199 and w13631;
w13633 <= not w13207 and not w13632;
w13634 <= not w13630 and w13633;
w13635 <= not w13207 and not w13634;
w13636 <= b(32) and not w13196;
w13637 <= not w13190 and w13636;
w13638 <= not w13198 and not w13637;
w13639 <= not w13635 and w13638;
w13640 <= not w13198 and not w13639;
w13641 <= b(33) and not w13187;
w13642 <= not w13181 and w13641;
w13643 <= not w13189 and not w13642;
w13644 <= not w13640 and w13643;
w13645 <= not w13189 and not w13644;
w13646 <= b(34) and not w13178;
w13647 <= not w13172 and w13646;
w13648 <= not w13180 and not w13647;
w13649 <= not w13645 and w13648;
w13650 <= not w13180 and not w13649;
w13651 <= b(35) and not w13169;
w13652 <= not w13163 and w13651;
w13653 <= not w13171 and not w13652;
w13654 <= not w13650 and w13653;
w13655 <= not w13171 and not w13654;
w13656 <= b(36) and not w13160;
w13657 <= not w13154 and w13656;
w13658 <= not w13162 and not w13657;
w13659 <= not w13655 and w13658;
w13660 <= not w13162 and not w13659;
w13661 <= b(37) and not w13151;
w13662 <= not w13145 and w13661;
w13663 <= not w13153 and not w13662;
w13664 <= not w13660 and w13663;
w13665 <= not w13153 and not w13664;
w13666 <= b(38) and not w13142;
w13667 <= not w13136 and w13666;
w13668 <= not w13144 and not w13667;
w13669 <= not w13665 and w13668;
w13670 <= not w13144 and not w13669;
w13671 <= b(39) and not w13133;
w13672 <= not w13127 and w13671;
w13673 <= not w13135 and not w13672;
w13674 <= not w13670 and w13673;
w13675 <= not w13135 and not w13674;
w13676 <= b(40) and not w13124;
w13677 <= not w13118 and w13676;
w13678 <= not w13126 and not w13677;
w13679 <= not w13675 and w13678;
w13680 <= not w13126 and not w13679;
w13681 <= b(41) and not w13115;
w13682 <= not w13109 and w13681;
w13683 <= not w13117 and not w13682;
w13684 <= not w13680 and w13683;
w13685 <= not w13117 and not w13684;
w13686 <= b(42) and not w13106;
w13687 <= not w13100 and w13686;
w13688 <= not w13108 and not w13687;
w13689 <= not w13685 and w13688;
w13690 <= not w13108 and not w13689;
w13691 <= not w12527 and not w13099;
w13692 <= not w12529 and w13094;
w13693 <= not w13090 and w13692;
w13694 <= not w13091 and not w13094;
w13695 <= not w13693 and not w13694;
w13696 <= w13099 and not w13695;
w13697 <= not w13691 and not w13696;
w13698 <= not b(43) and not w13697;
w13699 <= b(43) and not w13691;
w13700 <= not w13696 and w13699;
w13701 <= w31 and w45;
w13702 <= not w13700 and w13701;
w13703 <= not w13698 and w13702;
w13704 <= not w13690 and w13703;
w13705 <= w13098 and not w13697;
w13706 <= not w13704 and not w13705;
w13707 <= not w13117 and w13688;
w13708 <= not w13684 and w13707;
w13709 <= not w13685 and not w13688;
w13710 <= not w13708 and not w13709;
w13711 <= not w13706 and not w13710;
w13712 <= not w13107 and not w13705;
w13713 <= not w13704 and w13712;
w13714 <= not w13711 and not w13713;
w13715 <= not b(43) and not w13714;
w13716 <= not w13126 and w13683;
w13717 <= not w13679 and w13716;
w13718 <= not w13680 and not w13683;
w13719 <= not w13717 and not w13718;
w13720 <= not w13706 and not w13719;
w13721 <= not w13116 and not w13705;
w13722 <= not w13704 and w13721;
w13723 <= not w13720 and not w13722;
w13724 <= not b(42) and not w13723;
w13725 <= not w13135 and w13678;
w13726 <= not w13674 and w13725;
w13727 <= not w13675 and not w13678;
w13728 <= not w13726 and not w13727;
w13729 <= not w13706 and not w13728;
w13730 <= not w13125 and not w13705;
w13731 <= not w13704 and w13730;
w13732 <= not w13729 and not w13731;
w13733 <= not b(41) and not w13732;
w13734 <= not w13144 and w13673;
w13735 <= not w13669 and w13734;
w13736 <= not w13670 and not w13673;
w13737 <= not w13735 and not w13736;
w13738 <= not w13706 and not w13737;
w13739 <= not w13134 and not w13705;
w13740 <= not w13704 and w13739;
w13741 <= not w13738 and not w13740;
w13742 <= not b(40) and not w13741;
w13743 <= not w13153 and w13668;
w13744 <= not w13664 and w13743;
w13745 <= not w13665 and not w13668;
w13746 <= not w13744 and not w13745;
w13747 <= not w13706 and not w13746;
w13748 <= not w13143 and not w13705;
w13749 <= not w13704 and w13748;
w13750 <= not w13747 and not w13749;
w13751 <= not b(39) and not w13750;
w13752 <= not w13162 and w13663;
w13753 <= not w13659 and w13752;
w13754 <= not w13660 and not w13663;
w13755 <= not w13753 and not w13754;
w13756 <= not w13706 and not w13755;
w13757 <= not w13152 and not w13705;
w13758 <= not w13704 and w13757;
w13759 <= not w13756 and not w13758;
w13760 <= not b(38) and not w13759;
w13761 <= not w13171 and w13658;
w13762 <= not w13654 and w13761;
w13763 <= not w13655 and not w13658;
w13764 <= not w13762 and not w13763;
w13765 <= not w13706 and not w13764;
w13766 <= not w13161 and not w13705;
w13767 <= not w13704 and w13766;
w13768 <= not w13765 and not w13767;
w13769 <= not b(37) and not w13768;
w13770 <= not w13180 and w13653;
w13771 <= not w13649 and w13770;
w13772 <= not w13650 and not w13653;
w13773 <= not w13771 and not w13772;
w13774 <= not w13706 and not w13773;
w13775 <= not w13170 and not w13705;
w13776 <= not w13704 and w13775;
w13777 <= not w13774 and not w13776;
w13778 <= not b(36) and not w13777;
w13779 <= not w13189 and w13648;
w13780 <= not w13644 and w13779;
w13781 <= not w13645 and not w13648;
w13782 <= not w13780 and not w13781;
w13783 <= not w13706 and not w13782;
w13784 <= not w13179 and not w13705;
w13785 <= not w13704 and w13784;
w13786 <= not w13783 and not w13785;
w13787 <= not b(35) and not w13786;
w13788 <= not w13198 and w13643;
w13789 <= not w13639 and w13788;
w13790 <= not w13640 and not w13643;
w13791 <= not w13789 and not w13790;
w13792 <= not w13706 and not w13791;
w13793 <= not w13188 and not w13705;
w13794 <= not w13704 and w13793;
w13795 <= not w13792 and not w13794;
w13796 <= not b(34) and not w13795;
w13797 <= not w13207 and w13638;
w13798 <= not w13634 and w13797;
w13799 <= not w13635 and not w13638;
w13800 <= not w13798 and not w13799;
w13801 <= not w13706 and not w13800;
w13802 <= not w13197 and not w13705;
w13803 <= not w13704 and w13802;
w13804 <= not w13801 and not w13803;
w13805 <= not b(33) and not w13804;
w13806 <= not w13216 and w13633;
w13807 <= not w13629 and w13806;
w13808 <= not w13630 and not w13633;
w13809 <= not w13807 and not w13808;
w13810 <= not w13706 and not w13809;
w13811 <= not w13206 and not w13705;
w13812 <= not w13704 and w13811;
w13813 <= not w13810 and not w13812;
w13814 <= not b(32) and not w13813;
w13815 <= not w13225 and w13628;
w13816 <= not w13624 and w13815;
w13817 <= not w13625 and not w13628;
w13818 <= not w13816 and not w13817;
w13819 <= not w13706 and not w13818;
w13820 <= not w13215 and not w13705;
w13821 <= not w13704 and w13820;
w13822 <= not w13819 and not w13821;
w13823 <= not b(31) and not w13822;
w13824 <= not w13234 and w13623;
w13825 <= not w13619 and w13824;
w13826 <= not w13620 and not w13623;
w13827 <= not w13825 and not w13826;
w13828 <= not w13706 and not w13827;
w13829 <= not w13224 and not w13705;
w13830 <= not w13704 and w13829;
w13831 <= not w13828 and not w13830;
w13832 <= not b(30) and not w13831;
w13833 <= not w13243 and w13618;
w13834 <= not w13614 and w13833;
w13835 <= not w13615 and not w13618;
w13836 <= not w13834 and not w13835;
w13837 <= not w13706 and not w13836;
w13838 <= not w13233 and not w13705;
w13839 <= not w13704 and w13838;
w13840 <= not w13837 and not w13839;
w13841 <= not b(29) and not w13840;
w13842 <= not w13252 and w13613;
w13843 <= not w13609 and w13842;
w13844 <= not w13610 and not w13613;
w13845 <= not w13843 and not w13844;
w13846 <= not w13706 and not w13845;
w13847 <= not w13242 and not w13705;
w13848 <= not w13704 and w13847;
w13849 <= not w13846 and not w13848;
w13850 <= not b(28) and not w13849;
w13851 <= not w13261 and w13608;
w13852 <= not w13604 and w13851;
w13853 <= not w13605 and not w13608;
w13854 <= not w13852 and not w13853;
w13855 <= not w13706 and not w13854;
w13856 <= not w13251 and not w13705;
w13857 <= not w13704 and w13856;
w13858 <= not w13855 and not w13857;
w13859 <= not b(27) and not w13858;
w13860 <= not w13270 and w13603;
w13861 <= not w13599 and w13860;
w13862 <= not w13600 and not w13603;
w13863 <= not w13861 and not w13862;
w13864 <= not w13706 and not w13863;
w13865 <= not w13260 and not w13705;
w13866 <= not w13704 and w13865;
w13867 <= not w13864 and not w13866;
w13868 <= not b(26) and not w13867;
w13869 <= not w13279 and w13598;
w13870 <= not w13594 and w13869;
w13871 <= not w13595 and not w13598;
w13872 <= not w13870 and not w13871;
w13873 <= not w13706 and not w13872;
w13874 <= not w13269 and not w13705;
w13875 <= not w13704 and w13874;
w13876 <= not w13873 and not w13875;
w13877 <= not b(25) and not w13876;
w13878 <= not w13288 and w13593;
w13879 <= not w13589 and w13878;
w13880 <= not w13590 and not w13593;
w13881 <= not w13879 and not w13880;
w13882 <= not w13706 and not w13881;
w13883 <= not w13278 and not w13705;
w13884 <= not w13704 and w13883;
w13885 <= not w13882 and not w13884;
w13886 <= not b(24) and not w13885;
w13887 <= not w13297 and w13588;
w13888 <= not w13584 and w13887;
w13889 <= not w13585 and not w13588;
w13890 <= not w13888 and not w13889;
w13891 <= not w13706 and not w13890;
w13892 <= not w13287 and not w13705;
w13893 <= not w13704 and w13892;
w13894 <= not w13891 and not w13893;
w13895 <= not b(23) and not w13894;
w13896 <= not w13306 and w13583;
w13897 <= not w13579 and w13896;
w13898 <= not w13580 and not w13583;
w13899 <= not w13897 and not w13898;
w13900 <= not w13706 and not w13899;
w13901 <= not w13296 and not w13705;
w13902 <= not w13704 and w13901;
w13903 <= not w13900 and not w13902;
w13904 <= not b(22) and not w13903;
w13905 <= not w13315 and w13578;
w13906 <= not w13574 and w13905;
w13907 <= not w13575 and not w13578;
w13908 <= not w13906 and not w13907;
w13909 <= not w13706 and not w13908;
w13910 <= not w13305 and not w13705;
w13911 <= not w13704 and w13910;
w13912 <= not w13909 and not w13911;
w13913 <= not b(21) and not w13912;
w13914 <= not w13324 and w13573;
w13915 <= not w13569 and w13914;
w13916 <= not w13570 and not w13573;
w13917 <= not w13915 and not w13916;
w13918 <= not w13706 and not w13917;
w13919 <= not w13314 and not w13705;
w13920 <= not w13704 and w13919;
w13921 <= not w13918 and not w13920;
w13922 <= not b(20) and not w13921;
w13923 <= not w13333 and w13568;
w13924 <= not w13564 and w13923;
w13925 <= not w13565 and not w13568;
w13926 <= not w13924 and not w13925;
w13927 <= not w13706 and not w13926;
w13928 <= not w13323 and not w13705;
w13929 <= not w13704 and w13928;
w13930 <= not w13927 and not w13929;
w13931 <= not b(19) and not w13930;
w13932 <= not w13342 and w13563;
w13933 <= not w13559 and w13932;
w13934 <= not w13560 and not w13563;
w13935 <= not w13933 and not w13934;
w13936 <= not w13706 and not w13935;
w13937 <= not w13332 and not w13705;
w13938 <= not w13704 and w13937;
w13939 <= not w13936 and not w13938;
w13940 <= not b(18) and not w13939;
w13941 <= not w13351 and w13558;
w13942 <= not w13554 and w13941;
w13943 <= not w13555 and not w13558;
w13944 <= not w13942 and not w13943;
w13945 <= not w13706 and not w13944;
w13946 <= not w13341 and not w13705;
w13947 <= not w13704 and w13946;
w13948 <= not w13945 and not w13947;
w13949 <= not b(17) and not w13948;
w13950 <= not w13360 and w13553;
w13951 <= not w13549 and w13950;
w13952 <= not w13550 and not w13553;
w13953 <= not w13951 and not w13952;
w13954 <= not w13706 and not w13953;
w13955 <= not w13350 and not w13705;
w13956 <= not w13704 and w13955;
w13957 <= not w13954 and not w13956;
w13958 <= not b(16) and not w13957;
w13959 <= not w13369 and w13548;
w13960 <= not w13544 and w13959;
w13961 <= not w13545 and not w13548;
w13962 <= not w13960 and not w13961;
w13963 <= not w13706 and not w13962;
w13964 <= not w13359 and not w13705;
w13965 <= not w13704 and w13964;
w13966 <= not w13963 and not w13965;
w13967 <= not b(15) and not w13966;
w13968 <= not w13378 and w13543;
w13969 <= not w13539 and w13968;
w13970 <= not w13540 and not w13543;
w13971 <= not w13969 and not w13970;
w13972 <= not w13706 and not w13971;
w13973 <= not w13368 and not w13705;
w13974 <= not w13704 and w13973;
w13975 <= not w13972 and not w13974;
w13976 <= not b(14) and not w13975;
w13977 <= not w13387 and w13538;
w13978 <= not w13534 and w13977;
w13979 <= not w13535 and not w13538;
w13980 <= not w13978 and not w13979;
w13981 <= not w13706 and not w13980;
w13982 <= not w13377 and not w13705;
w13983 <= not w13704 and w13982;
w13984 <= not w13981 and not w13983;
w13985 <= not b(13) and not w13984;
w13986 <= not w13396 and w13533;
w13987 <= not w13529 and w13986;
w13988 <= not w13530 and not w13533;
w13989 <= not w13987 and not w13988;
w13990 <= not w13706 and not w13989;
w13991 <= not w13386 and not w13705;
w13992 <= not w13704 and w13991;
w13993 <= not w13990 and not w13992;
w13994 <= not b(12) and not w13993;
w13995 <= not w13405 and w13528;
w13996 <= not w13524 and w13995;
w13997 <= not w13525 and not w13528;
w13998 <= not w13996 and not w13997;
w13999 <= not w13706 and not w13998;
w14000 <= not w13395 and not w13705;
w14001 <= not w13704 and w14000;
w14002 <= not w13999 and not w14001;
w14003 <= not b(11) and not w14002;
w14004 <= not w13414 and w13523;
w14005 <= not w13519 and w14004;
w14006 <= not w13520 and not w13523;
w14007 <= not w14005 and not w14006;
w14008 <= not w13706 and not w14007;
w14009 <= not w13404 and not w13705;
w14010 <= not w13704 and w14009;
w14011 <= not w14008 and not w14010;
w14012 <= not b(10) and not w14011;
w14013 <= not w13423 and w13518;
w14014 <= not w13514 and w14013;
w14015 <= not w13515 and not w13518;
w14016 <= not w14014 and not w14015;
w14017 <= not w13706 and not w14016;
w14018 <= not w13413 and not w13705;
w14019 <= not w13704 and w14018;
w14020 <= not w14017 and not w14019;
w14021 <= not b(9) and not w14020;
w14022 <= not w13432 and w13513;
w14023 <= not w13509 and w14022;
w14024 <= not w13510 and not w13513;
w14025 <= not w14023 and not w14024;
w14026 <= not w13706 and not w14025;
w14027 <= not w13422 and not w13705;
w14028 <= not w13704 and w14027;
w14029 <= not w14026 and not w14028;
w14030 <= not b(8) and not w14029;
w14031 <= not w13441 and w13508;
w14032 <= not w13504 and w14031;
w14033 <= not w13505 and not w13508;
w14034 <= not w14032 and not w14033;
w14035 <= not w13706 and not w14034;
w14036 <= not w13431 and not w13705;
w14037 <= not w13704 and w14036;
w14038 <= not w14035 and not w14037;
w14039 <= not b(7) and not w14038;
w14040 <= not w13450 and w13503;
w14041 <= not w13499 and w14040;
w14042 <= not w13500 and not w13503;
w14043 <= not w14041 and not w14042;
w14044 <= not w13706 and not w14043;
w14045 <= not w13440 and not w13705;
w14046 <= not w13704 and w14045;
w14047 <= not w14044 and not w14046;
w14048 <= not b(6) and not w14047;
w14049 <= not w13459 and w13498;
w14050 <= not w13494 and w14049;
w14051 <= not w13495 and not w13498;
w14052 <= not w14050 and not w14051;
w14053 <= not w13706 and not w14052;
w14054 <= not w13449 and not w13705;
w14055 <= not w13704 and w14054;
w14056 <= not w14053 and not w14055;
w14057 <= not b(5) and not w14056;
w14058 <= not w13467 and w13493;
w14059 <= not w13489 and w14058;
w14060 <= not w13490 and not w13493;
w14061 <= not w14059 and not w14060;
w14062 <= not w13706 and not w14061;
w14063 <= not w13458 and not w13705;
w14064 <= not w13704 and w14063;
w14065 <= not w14062 and not w14064;
w14066 <= not b(4) and not w14065;
w14067 <= not w13484 and w13488;
w14068 <= not w13483 and w14067;
w14069 <= not w13485 and not w13488;
w14070 <= not w14068 and not w14069;
w14071 <= not w13706 and not w14070;
w14072 <= not w13466 and not w13705;
w14073 <= not w13704 and w14072;
w14074 <= not w14071 and not w14073;
w14075 <= not b(3) and not w14074;
w14076 <= not w13480 and w13482;
w14077 <= not w13478 and w14076;
w14078 <= not w13483 and not w14077;
w14079 <= not w13706 and w14078;
w14080 <= not w13477 and not w13705;
w14081 <= not w13704 and w14080;
w14082 <= not w14079 and not w14081;
w14083 <= not b(2) and not w14082;
w14084 <= b(0) and not w13706;
w14085 <= a(20) and not w14084;
w14086 <= w13482 and not w13706;
w14087 <= not w14085 and not w14086;
w14088 <= b(1) and not w14087;
w14089 <= not b(1) and not w14086;
w14090 <= not w14085 and w14089;
w14091 <= not w14088 and not w14090;
w14092 <= not a(19) and b(0);
w14093 <= not w14091 and not w14092;
w14094 <= not b(1) and not w14087;
w14095 <= not w14093 and not w14094;
w14096 <= b(2) and not w14081;
w14097 <= not w14079 and w14096;
w14098 <= not w14083 and not w14097;
w14099 <= not w14095 and w14098;
w14100 <= not w14083 and not w14099;
w14101 <= b(3) and not w14073;
w14102 <= not w14071 and w14101;
w14103 <= not w14075 and not w14102;
w14104 <= not w14100 and w14103;
w14105 <= not w14075 and not w14104;
w14106 <= b(4) and not w14064;
w14107 <= not w14062 and w14106;
w14108 <= not w14066 and not w14107;
w14109 <= not w14105 and w14108;
w14110 <= not w14066 and not w14109;
w14111 <= b(5) and not w14055;
w14112 <= not w14053 and w14111;
w14113 <= not w14057 and not w14112;
w14114 <= not w14110 and w14113;
w14115 <= not w14057 and not w14114;
w14116 <= b(6) and not w14046;
w14117 <= not w14044 and w14116;
w14118 <= not w14048 and not w14117;
w14119 <= not w14115 and w14118;
w14120 <= not w14048 and not w14119;
w14121 <= b(7) and not w14037;
w14122 <= not w14035 and w14121;
w14123 <= not w14039 and not w14122;
w14124 <= not w14120 and w14123;
w14125 <= not w14039 and not w14124;
w14126 <= b(8) and not w14028;
w14127 <= not w14026 and w14126;
w14128 <= not w14030 and not w14127;
w14129 <= not w14125 and w14128;
w14130 <= not w14030 and not w14129;
w14131 <= b(9) and not w14019;
w14132 <= not w14017 and w14131;
w14133 <= not w14021 and not w14132;
w14134 <= not w14130 and w14133;
w14135 <= not w14021 and not w14134;
w14136 <= b(10) and not w14010;
w14137 <= not w14008 and w14136;
w14138 <= not w14012 and not w14137;
w14139 <= not w14135 and w14138;
w14140 <= not w14012 and not w14139;
w14141 <= b(11) and not w14001;
w14142 <= not w13999 and w14141;
w14143 <= not w14003 and not w14142;
w14144 <= not w14140 and w14143;
w14145 <= not w14003 and not w14144;
w14146 <= b(12) and not w13992;
w14147 <= not w13990 and w14146;
w14148 <= not w13994 and not w14147;
w14149 <= not w14145 and w14148;
w14150 <= not w13994 and not w14149;
w14151 <= b(13) and not w13983;
w14152 <= not w13981 and w14151;
w14153 <= not w13985 and not w14152;
w14154 <= not w14150 and w14153;
w14155 <= not w13985 and not w14154;
w14156 <= b(14) and not w13974;
w14157 <= not w13972 and w14156;
w14158 <= not w13976 and not w14157;
w14159 <= not w14155 and w14158;
w14160 <= not w13976 and not w14159;
w14161 <= b(15) and not w13965;
w14162 <= not w13963 and w14161;
w14163 <= not w13967 and not w14162;
w14164 <= not w14160 and w14163;
w14165 <= not w13967 and not w14164;
w14166 <= b(16) and not w13956;
w14167 <= not w13954 and w14166;
w14168 <= not w13958 and not w14167;
w14169 <= not w14165 and w14168;
w14170 <= not w13958 and not w14169;
w14171 <= b(17) and not w13947;
w14172 <= not w13945 and w14171;
w14173 <= not w13949 and not w14172;
w14174 <= not w14170 and w14173;
w14175 <= not w13949 and not w14174;
w14176 <= b(18) and not w13938;
w14177 <= not w13936 and w14176;
w14178 <= not w13940 and not w14177;
w14179 <= not w14175 and w14178;
w14180 <= not w13940 and not w14179;
w14181 <= b(19) and not w13929;
w14182 <= not w13927 and w14181;
w14183 <= not w13931 and not w14182;
w14184 <= not w14180 and w14183;
w14185 <= not w13931 and not w14184;
w14186 <= b(20) and not w13920;
w14187 <= not w13918 and w14186;
w14188 <= not w13922 and not w14187;
w14189 <= not w14185 and w14188;
w14190 <= not w13922 and not w14189;
w14191 <= b(21) and not w13911;
w14192 <= not w13909 and w14191;
w14193 <= not w13913 and not w14192;
w14194 <= not w14190 and w14193;
w14195 <= not w13913 and not w14194;
w14196 <= b(22) and not w13902;
w14197 <= not w13900 and w14196;
w14198 <= not w13904 and not w14197;
w14199 <= not w14195 and w14198;
w14200 <= not w13904 and not w14199;
w14201 <= b(23) and not w13893;
w14202 <= not w13891 and w14201;
w14203 <= not w13895 and not w14202;
w14204 <= not w14200 and w14203;
w14205 <= not w13895 and not w14204;
w14206 <= b(24) and not w13884;
w14207 <= not w13882 and w14206;
w14208 <= not w13886 and not w14207;
w14209 <= not w14205 and w14208;
w14210 <= not w13886 and not w14209;
w14211 <= b(25) and not w13875;
w14212 <= not w13873 and w14211;
w14213 <= not w13877 and not w14212;
w14214 <= not w14210 and w14213;
w14215 <= not w13877 and not w14214;
w14216 <= b(26) and not w13866;
w14217 <= not w13864 and w14216;
w14218 <= not w13868 and not w14217;
w14219 <= not w14215 and w14218;
w14220 <= not w13868 and not w14219;
w14221 <= b(27) and not w13857;
w14222 <= not w13855 and w14221;
w14223 <= not w13859 and not w14222;
w14224 <= not w14220 and w14223;
w14225 <= not w13859 and not w14224;
w14226 <= b(28) and not w13848;
w14227 <= not w13846 and w14226;
w14228 <= not w13850 and not w14227;
w14229 <= not w14225 and w14228;
w14230 <= not w13850 and not w14229;
w14231 <= b(29) and not w13839;
w14232 <= not w13837 and w14231;
w14233 <= not w13841 and not w14232;
w14234 <= not w14230 and w14233;
w14235 <= not w13841 and not w14234;
w14236 <= b(30) and not w13830;
w14237 <= not w13828 and w14236;
w14238 <= not w13832 and not w14237;
w14239 <= not w14235 and w14238;
w14240 <= not w13832 and not w14239;
w14241 <= b(31) and not w13821;
w14242 <= not w13819 and w14241;
w14243 <= not w13823 and not w14242;
w14244 <= not w14240 and w14243;
w14245 <= not w13823 and not w14244;
w14246 <= b(32) and not w13812;
w14247 <= not w13810 and w14246;
w14248 <= not w13814 and not w14247;
w14249 <= not w14245 and w14248;
w14250 <= not w13814 and not w14249;
w14251 <= b(33) and not w13803;
w14252 <= not w13801 and w14251;
w14253 <= not w13805 and not w14252;
w14254 <= not w14250 and w14253;
w14255 <= not w13805 and not w14254;
w14256 <= b(34) and not w13794;
w14257 <= not w13792 and w14256;
w14258 <= not w13796 and not w14257;
w14259 <= not w14255 and w14258;
w14260 <= not w13796 and not w14259;
w14261 <= b(35) and not w13785;
w14262 <= not w13783 and w14261;
w14263 <= not w13787 and not w14262;
w14264 <= not w14260 and w14263;
w14265 <= not w13787 and not w14264;
w14266 <= b(36) and not w13776;
w14267 <= not w13774 and w14266;
w14268 <= not w13778 and not w14267;
w14269 <= not w14265 and w14268;
w14270 <= not w13778 and not w14269;
w14271 <= b(37) and not w13767;
w14272 <= not w13765 and w14271;
w14273 <= not w13769 and not w14272;
w14274 <= not w14270 and w14273;
w14275 <= not w13769 and not w14274;
w14276 <= b(38) and not w13758;
w14277 <= not w13756 and w14276;
w14278 <= not w13760 and not w14277;
w14279 <= not w14275 and w14278;
w14280 <= not w13760 and not w14279;
w14281 <= b(39) and not w13749;
w14282 <= not w13747 and w14281;
w14283 <= not w13751 and not w14282;
w14284 <= not w14280 and w14283;
w14285 <= not w13751 and not w14284;
w14286 <= b(40) and not w13740;
w14287 <= not w13738 and w14286;
w14288 <= not w13742 and not w14287;
w14289 <= not w14285 and w14288;
w14290 <= not w13742 and not w14289;
w14291 <= b(41) and not w13731;
w14292 <= not w13729 and w14291;
w14293 <= not w13733 and not w14292;
w14294 <= not w14290 and w14293;
w14295 <= not w13733 and not w14294;
w14296 <= b(42) and not w13722;
w14297 <= not w13720 and w14296;
w14298 <= not w13724 and not w14297;
w14299 <= not w14295 and w14298;
w14300 <= not w13724 and not w14299;
w14301 <= b(43) and not w13713;
w14302 <= not w13711 and w14301;
w14303 <= not w13715 and not w14302;
w14304 <= not w14300 and w14303;
w14305 <= not w13715 and not w14304;
w14306 <= not w13108 and not w13700;
w14307 <= not w13698 and w14306;
w14308 <= not w13689 and w14307;
w14309 <= not w13698 and not w13700;
w14310 <= not w13690 and not w14309;
w14311 <= not w14308 and not w14310;
w14312 <= not w13706 and not w14311;
w14313 <= not w13697 and not w13705;
w14314 <= not w13704 and w14313;
w14315 <= not w14312 and not w14314;
w14316 <= not b(44) and not w14315;
w14317 <= b(44) and not w14314;
w14318 <= not w14312 and w14317;
w14319 <= w338 and w340;
w14320 <= not w14318 and w14319;
w14321 <= not w14316 and w14320;
w14322 <= not w14305 and w14321;
w14323 <= w13701 and not w14315;
w14324 <= not w14322 and not w14323;
w14325 <= not w13724 and w14303;
w14326 <= not w14299 and w14325;
w14327 <= not w14300 and not w14303;
w14328 <= not w14326 and not w14327;
w14329 <= not w14324 and not w14328;
w14330 <= not w13714 and not w14323;
w14331 <= not w14322 and w14330;
w14332 <= not w14329 and not w14331;
w14333 <= not w13715 and not w14318;
w14334 <= not w14316 and w14333;
w14335 <= not w14304 and w14334;
w14336 <= not w14316 and not w14318;
w14337 <= not w14305 and not w14336;
w14338 <= not w14335 and not w14337;
w14339 <= not w14324 and not w14338;
w14340 <= not w14315 and not w14323;
w14341 <= not w14322 and w14340;
w14342 <= not w14339 and not w14341;
w14343 <= not b(45) and not w14342;
w14344 <= not b(44) and not w14332;
w14345 <= not w13733 and w14298;
w14346 <= not w14294 and w14345;
w14347 <= not w14295 and not w14298;
w14348 <= not w14346 and not w14347;
w14349 <= not w14324 and not w14348;
w14350 <= not w13723 and not w14323;
w14351 <= not w14322 and w14350;
w14352 <= not w14349 and not w14351;
w14353 <= not b(43) and not w14352;
w14354 <= not w13742 and w14293;
w14355 <= not w14289 and w14354;
w14356 <= not w14290 and not w14293;
w14357 <= not w14355 and not w14356;
w14358 <= not w14324 and not w14357;
w14359 <= not w13732 and not w14323;
w14360 <= not w14322 and w14359;
w14361 <= not w14358 and not w14360;
w14362 <= not b(42) and not w14361;
w14363 <= not w13751 and w14288;
w14364 <= not w14284 and w14363;
w14365 <= not w14285 and not w14288;
w14366 <= not w14364 and not w14365;
w14367 <= not w14324 and not w14366;
w14368 <= not w13741 and not w14323;
w14369 <= not w14322 and w14368;
w14370 <= not w14367 and not w14369;
w14371 <= not b(41) and not w14370;
w14372 <= not w13760 and w14283;
w14373 <= not w14279 and w14372;
w14374 <= not w14280 and not w14283;
w14375 <= not w14373 and not w14374;
w14376 <= not w14324 and not w14375;
w14377 <= not w13750 and not w14323;
w14378 <= not w14322 and w14377;
w14379 <= not w14376 and not w14378;
w14380 <= not b(40) and not w14379;
w14381 <= not w13769 and w14278;
w14382 <= not w14274 and w14381;
w14383 <= not w14275 and not w14278;
w14384 <= not w14382 and not w14383;
w14385 <= not w14324 and not w14384;
w14386 <= not w13759 and not w14323;
w14387 <= not w14322 and w14386;
w14388 <= not w14385 and not w14387;
w14389 <= not b(39) and not w14388;
w14390 <= not w13778 and w14273;
w14391 <= not w14269 and w14390;
w14392 <= not w14270 and not w14273;
w14393 <= not w14391 and not w14392;
w14394 <= not w14324 and not w14393;
w14395 <= not w13768 and not w14323;
w14396 <= not w14322 and w14395;
w14397 <= not w14394 and not w14396;
w14398 <= not b(38) and not w14397;
w14399 <= not w13787 and w14268;
w14400 <= not w14264 and w14399;
w14401 <= not w14265 and not w14268;
w14402 <= not w14400 and not w14401;
w14403 <= not w14324 and not w14402;
w14404 <= not w13777 and not w14323;
w14405 <= not w14322 and w14404;
w14406 <= not w14403 and not w14405;
w14407 <= not b(37) and not w14406;
w14408 <= not w13796 and w14263;
w14409 <= not w14259 and w14408;
w14410 <= not w14260 and not w14263;
w14411 <= not w14409 and not w14410;
w14412 <= not w14324 and not w14411;
w14413 <= not w13786 and not w14323;
w14414 <= not w14322 and w14413;
w14415 <= not w14412 and not w14414;
w14416 <= not b(36) and not w14415;
w14417 <= not w13805 and w14258;
w14418 <= not w14254 and w14417;
w14419 <= not w14255 and not w14258;
w14420 <= not w14418 and not w14419;
w14421 <= not w14324 and not w14420;
w14422 <= not w13795 and not w14323;
w14423 <= not w14322 and w14422;
w14424 <= not w14421 and not w14423;
w14425 <= not b(35) and not w14424;
w14426 <= not w13814 and w14253;
w14427 <= not w14249 and w14426;
w14428 <= not w14250 and not w14253;
w14429 <= not w14427 and not w14428;
w14430 <= not w14324 and not w14429;
w14431 <= not w13804 and not w14323;
w14432 <= not w14322 and w14431;
w14433 <= not w14430 and not w14432;
w14434 <= not b(34) and not w14433;
w14435 <= not w13823 and w14248;
w14436 <= not w14244 and w14435;
w14437 <= not w14245 and not w14248;
w14438 <= not w14436 and not w14437;
w14439 <= not w14324 and not w14438;
w14440 <= not w13813 and not w14323;
w14441 <= not w14322 and w14440;
w14442 <= not w14439 and not w14441;
w14443 <= not b(33) and not w14442;
w14444 <= not w13832 and w14243;
w14445 <= not w14239 and w14444;
w14446 <= not w14240 and not w14243;
w14447 <= not w14445 and not w14446;
w14448 <= not w14324 and not w14447;
w14449 <= not w13822 and not w14323;
w14450 <= not w14322 and w14449;
w14451 <= not w14448 and not w14450;
w14452 <= not b(32) and not w14451;
w14453 <= not w13841 and w14238;
w14454 <= not w14234 and w14453;
w14455 <= not w14235 and not w14238;
w14456 <= not w14454 and not w14455;
w14457 <= not w14324 and not w14456;
w14458 <= not w13831 and not w14323;
w14459 <= not w14322 and w14458;
w14460 <= not w14457 and not w14459;
w14461 <= not b(31) and not w14460;
w14462 <= not w13850 and w14233;
w14463 <= not w14229 and w14462;
w14464 <= not w14230 and not w14233;
w14465 <= not w14463 and not w14464;
w14466 <= not w14324 and not w14465;
w14467 <= not w13840 and not w14323;
w14468 <= not w14322 and w14467;
w14469 <= not w14466 and not w14468;
w14470 <= not b(30) and not w14469;
w14471 <= not w13859 and w14228;
w14472 <= not w14224 and w14471;
w14473 <= not w14225 and not w14228;
w14474 <= not w14472 and not w14473;
w14475 <= not w14324 and not w14474;
w14476 <= not w13849 and not w14323;
w14477 <= not w14322 and w14476;
w14478 <= not w14475 and not w14477;
w14479 <= not b(29) and not w14478;
w14480 <= not w13868 and w14223;
w14481 <= not w14219 and w14480;
w14482 <= not w14220 and not w14223;
w14483 <= not w14481 and not w14482;
w14484 <= not w14324 and not w14483;
w14485 <= not w13858 and not w14323;
w14486 <= not w14322 and w14485;
w14487 <= not w14484 and not w14486;
w14488 <= not b(28) and not w14487;
w14489 <= not w13877 and w14218;
w14490 <= not w14214 and w14489;
w14491 <= not w14215 and not w14218;
w14492 <= not w14490 and not w14491;
w14493 <= not w14324 and not w14492;
w14494 <= not w13867 and not w14323;
w14495 <= not w14322 and w14494;
w14496 <= not w14493 and not w14495;
w14497 <= not b(27) and not w14496;
w14498 <= not w13886 and w14213;
w14499 <= not w14209 and w14498;
w14500 <= not w14210 and not w14213;
w14501 <= not w14499 and not w14500;
w14502 <= not w14324 and not w14501;
w14503 <= not w13876 and not w14323;
w14504 <= not w14322 and w14503;
w14505 <= not w14502 and not w14504;
w14506 <= not b(26) and not w14505;
w14507 <= not w13895 and w14208;
w14508 <= not w14204 and w14507;
w14509 <= not w14205 and not w14208;
w14510 <= not w14508 and not w14509;
w14511 <= not w14324 and not w14510;
w14512 <= not w13885 and not w14323;
w14513 <= not w14322 and w14512;
w14514 <= not w14511 and not w14513;
w14515 <= not b(25) and not w14514;
w14516 <= not w13904 and w14203;
w14517 <= not w14199 and w14516;
w14518 <= not w14200 and not w14203;
w14519 <= not w14517 and not w14518;
w14520 <= not w14324 and not w14519;
w14521 <= not w13894 and not w14323;
w14522 <= not w14322 and w14521;
w14523 <= not w14520 and not w14522;
w14524 <= not b(24) and not w14523;
w14525 <= not w13913 and w14198;
w14526 <= not w14194 and w14525;
w14527 <= not w14195 and not w14198;
w14528 <= not w14526 and not w14527;
w14529 <= not w14324 and not w14528;
w14530 <= not w13903 and not w14323;
w14531 <= not w14322 and w14530;
w14532 <= not w14529 and not w14531;
w14533 <= not b(23) and not w14532;
w14534 <= not w13922 and w14193;
w14535 <= not w14189 and w14534;
w14536 <= not w14190 and not w14193;
w14537 <= not w14535 and not w14536;
w14538 <= not w14324 and not w14537;
w14539 <= not w13912 and not w14323;
w14540 <= not w14322 and w14539;
w14541 <= not w14538 and not w14540;
w14542 <= not b(22) and not w14541;
w14543 <= not w13931 and w14188;
w14544 <= not w14184 and w14543;
w14545 <= not w14185 and not w14188;
w14546 <= not w14544 and not w14545;
w14547 <= not w14324 and not w14546;
w14548 <= not w13921 and not w14323;
w14549 <= not w14322 and w14548;
w14550 <= not w14547 and not w14549;
w14551 <= not b(21) and not w14550;
w14552 <= not w13940 and w14183;
w14553 <= not w14179 and w14552;
w14554 <= not w14180 and not w14183;
w14555 <= not w14553 and not w14554;
w14556 <= not w14324 and not w14555;
w14557 <= not w13930 and not w14323;
w14558 <= not w14322 and w14557;
w14559 <= not w14556 and not w14558;
w14560 <= not b(20) and not w14559;
w14561 <= not w13949 and w14178;
w14562 <= not w14174 and w14561;
w14563 <= not w14175 and not w14178;
w14564 <= not w14562 and not w14563;
w14565 <= not w14324 and not w14564;
w14566 <= not w13939 and not w14323;
w14567 <= not w14322 and w14566;
w14568 <= not w14565 and not w14567;
w14569 <= not b(19) and not w14568;
w14570 <= not w13958 and w14173;
w14571 <= not w14169 and w14570;
w14572 <= not w14170 and not w14173;
w14573 <= not w14571 and not w14572;
w14574 <= not w14324 and not w14573;
w14575 <= not w13948 and not w14323;
w14576 <= not w14322 and w14575;
w14577 <= not w14574 and not w14576;
w14578 <= not b(18) and not w14577;
w14579 <= not w13967 and w14168;
w14580 <= not w14164 and w14579;
w14581 <= not w14165 and not w14168;
w14582 <= not w14580 and not w14581;
w14583 <= not w14324 and not w14582;
w14584 <= not w13957 and not w14323;
w14585 <= not w14322 and w14584;
w14586 <= not w14583 and not w14585;
w14587 <= not b(17) and not w14586;
w14588 <= not w13976 and w14163;
w14589 <= not w14159 and w14588;
w14590 <= not w14160 and not w14163;
w14591 <= not w14589 and not w14590;
w14592 <= not w14324 and not w14591;
w14593 <= not w13966 and not w14323;
w14594 <= not w14322 and w14593;
w14595 <= not w14592 and not w14594;
w14596 <= not b(16) and not w14595;
w14597 <= not w13985 and w14158;
w14598 <= not w14154 and w14597;
w14599 <= not w14155 and not w14158;
w14600 <= not w14598 and not w14599;
w14601 <= not w14324 and not w14600;
w14602 <= not w13975 and not w14323;
w14603 <= not w14322 and w14602;
w14604 <= not w14601 and not w14603;
w14605 <= not b(15) and not w14604;
w14606 <= not w13994 and w14153;
w14607 <= not w14149 and w14606;
w14608 <= not w14150 and not w14153;
w14609 <= not w14607 and not w14608;
w14610 <= not w14324 and not w14609;
w14611 <= not w13984 and not w14323;
w14612 <= not w14322 and w14611;
w14613 <= not w14610 and not w14612;
w14614 <= not b(14) and not w14613;
w14615 <= not w14003 and w14148;
w14616 <= not w14144 and w14615;
w14617 <= not w14145 and not w14148;
w14618 <= not w14616 and not w14617;
w14619 <= not w14324 and not w14618;
w14620 <= not w13993 and not w14323;
w14621 <= not w14322 and w14620;
w14622 <= not w14619 and not w14621;
w14623 <= not b(13) and not w14622;
w14624 <= not w14012 and w14143;
w14625 <= not w14139 and w14624;
w14626 <= not w14140 and not w14143;
w14627 <= not w14625 and not w14626;
w14628 <= not w14324 and not w14627;
w14629 <= not w14002 and not w14323;
w14630 <= not w14322 and w14629;
w14631 <= not w14628 and not w14630;
w14632 <= not b(12) and not w14631;
w14633 <= not w14021 and w14138;
w14634 <= not w14134 and w14633;
w14635 <= not w14135 and not w14138;
w14636 <= not w14634 and not w14635;
w14637 <= not w14324 and not w14636;
w14638 <= not w14011 and not w14323;
w14639 <= not w14322 and w14638;
w14640 <= not w14637 and not w14639;
w14641 <= not b(11) and not w14640;
w14642 <= not w14030 and w14133;
w14643 <= not w14129 and w14642;
w14644 <= not w14130 and not w14133;
w14645 <= not w14643 and not w14644;
w14646 <= not w14324 and not w14645;
w14647 <= not w14020 and not w14323;
w14648 <= not w14322 and w14647;
w14649 <= not w14646 and not w14648;
w14650 <= not b(10) and not w14649;
w14651 <= not w14039 and w14128;
w14652 <= not w14124 and w14651;
w14653 <= not w14125 and not w14128;
w14654 <= not w14652 and not w14653;
w14655 <= not w14324 and not w14654;
w14656 <= not w14029 and not w14323;
w14657 <= not w14322 and w14656;
w14658 <= not w14655 and not w14657;
w14659 <= not b(9) and not w14658;
w14660 <= not w14048 and w14123;
w14661 <= not w14119 and w14660;
w14662 <= not w14120 and not w14123;
w14663 <= not w14661 and not w14662;
w14664 <= not w14324 and not w14663;
w14665 <= not w14038 and not w14323;
w14666 <= not w14322 and w14665;
w14667 <= not w14664 and not w14666;
w14668 <= not b(8) and not w14667;
w14669 <= not w14057 and w14118;
w14670 <= not w14114 and w14669;
w14671 <= not w14115 and not w14118;
w14672 <= not w14670 and not w14671;
w14673 <= not w14324 and not w14672;
w14674 <= not w14047 and not w14323;
w14675 <= not w14322 and w14674;
w14676 <= not w14673 and not w14675;
w14677 <= not b(7) and not w14676;
w14678 <= not w14066 and w14113;
w14679 <= not w14109 and w14678;
w14680 <= not w14110 and not w14113;
w14681 <= not w14679 and not w14680;
w14682 <= not w14324 and not w14681;
w14683 <= not w14056 and not w14323;
w14684 <= not w14322 and w14683;
w14685 <= not w14682 and not w14684;
w14686 <= not b(6) and not w14685;
w14687 <= not w14075 and w14108;
w14688 <= not w14104 and w14687;
w14689 <= not w14105 and not w14108;
w14690 <= not w14688 and not w14689;
w14691 <= not w14324 and not w14690;
w14692 <= not w14065 and not w14323;
w14693 <= not w14322 and w14692;
w14694 <= not w14691 and not w14693;
w14695 <= not b(5) and not w14694;
w14696 <= not w14083 and w14103;
w14697 <= not w14099 and w14696;
w14698 <= not w14100 and not w14103;
w14699 <= not w14697 and not w14698;
w14700 <= not w14324 and not w14699;
w14701 <= not w14074 and not w14323;
w14702 <= not w14322 and w14701;
w14703 <= not w14700 and not w14702;
w14704 <= not b(4) and not w14703;
w14705 <= not w14094 and w14098;
w14706 <= not w14093 and w14705;
w14707 <= not w14095 and not w14098;
w14708 <= not w14706 and not w14707;
w14709 <= not w14324 and not w14708;
w14710 <= not w14082 and not w14323;
w14711 <= not w14322 and w14710;
w14712 <= not w14709 and not w14711;
w14713 <= not b(3) and not w14712;
w14714 <= not w14090 and w14092;
w14715 <= not w14088 and w14714;
w14716 <= not w14093 and not w14715;
w14717 <= not w14324 and w14716;
w14718 <= not w14087 and not w14323;
w14719 <= not w14322 and w14718;
w14720 <= not w14717 and not w14719;
w14721 <= not b(2) and not w14720;
w14722 <= b(0) and not w14324;
w14723 <= a(19) and not w14722;
w14724 <= w14092 and not w14324;
w14725 <= not w14723 and not w14724;
w14726 <= b(1) and not w14725;
w14727 <= not b(1) and not w14724;
w14728 <= not w14723 and w14727;
w14729 <= not w14726 and not w14728;
w14730 <= not a(18) and b(0);
w14731 <= not w14729 and not w14730;
w14732 <= not b(1) and not w14725;
w14733 <= not w14731 and not w14732;
w14734 <= b(2) and not w14719;
w14735 <= not w14717 and w14734;
w14736 <= not w14721 and not w14735;
w14737 <= not w14733 and w14736;
w14738 <= not w14721 and not w14737;
w14739 <= b(3) and not w14711;
w14740 <= not w14709 and w14739;
w14741 <= not w14713 and not w14740;
w14742 <= not w14738 and w14741;
w14743 <= not w14713 and not w14742;
w14744 <= b(4) and not w14702;
w14745 <= not w14700 and w14744;
w14746 <= not w14704 and not w14745;
w14747 <= not w14743 and w14746;
w14748 <= not w14704 and not w14747;
w14749 <= b(5) and not w14693;
w14750 <= not w14691 and w14749;
w14751 <= not w14695 and not w14750;
w14752 <= not w14748 and w14751;
w14753 <= not w14695 and not w14752;
w14754 <= b(6) and not w14684;
w14755 <= not w14682 and w14754;
w14756 <= not w14686 and not w14755;
w14757 <= not w14753 and w14756;
w14758 <= not w14686 and not w14757;
w14759 <= b(7) and not w14675;
w14760 <= not w14673 and w14759;
w14761 <= not w14677 and not w14760;
w14762 <= not w14758 and w14761;
w14763 <= not w14677 and not w14762;
w14764 <= b(8) and not w14666;
w14765 <= not w14664 and w14764;
w14766 <= not w14668 and not w14765;
w14767 <= not w14763 and w14766;
w14768 <= not w14668 and not w14767;
w14769 <= b(9) and not w14657;
w14770 <= not w14655 and w14769;
w14771 <= not w14659 and not w14770;
w14772 <= not w14768 and w14771;
w14773 <= not w14659 and not w14772;
w14774 <= b(10) and not w14648;
w14775 <= not w14646 and w14774;
w14776 <= not w14650 and not w14775;
w14777 <= not w14773 and w14776;
w14778 <= not w14650 and not w14777;
w14779 <= b(11) and not w14639;
w14780 <= not w14637 and w14779;
w14781 <= not w14641 and not w14780;
w14782 <= not w14778 and w14781;
w14783 <= not w14641 and not w14782;
w14784 <= b(12) and not w14630;
w14785 <= not w14628 and w14784;
w14786 <= not w14632 and not w14785;
w14787 <= not w14783 and w14786;
w14788 <= not w14632 and not w14787;
w14789 <= b(13) and not w14621;
w14790 <= not w14619 and w14789;
w14791 <= not w14623 and not w14790;
w14792 <= not w14788 and w14791;
w14793 <= not w14623 and not w14792;
w14794 <= b(14) and not w14612;
w14795 <= not w14610 and w14794;
w14796 <= not w14614 and not w14795;
w14797 <= not w14793 and w14796;
w14798 <= not w14614 and not w14797;
w14799 <= b(15) and not w14603;
w14800 <= not w14601 and w14799;
w14801 <= not w14605 and not w14800;
w14802 <= not w14798 and w14801;
w14803 <= not w14605 and not w14802;
w14804 <= b(16) and not w14594;
w14805 <= not w14592 and w14804;
w14806 <= not w14596 and not w14805;
w14807 <= not w14803 and w14806;
w14808 <= not w14596 and not w14807;
w14809 <= b(17) and not w14585;
w14810 <= not w14583 and w14809;
w14811 <= not w14587 and not w14810;
w14812 <= not w14808 and w14811;
w14813 <= not w14587 and not w14812;
w14814 <= b(18) and not w14576;
w14815 <= not w14574 and w14814;
w14816 <= not w14578 and not w14815;
w14817 <= not w14813 and w14816;
w14818 <= not w14578 and not w14817;
w14819 <= b(19) and not w14567;
w14820 <= not w14565 and w14819;
w14821 <= not w14569 and not w14820;
w14822 <= not w14818 and w14821;
w14823 <= not w14569 and not w14822;
w14824 <= b(20) and not w14558;
w14825 <= not w14556 and w14824;
w14826 <= not w14560 and not w14825;
w14827 <= not w14823 and w14826;
w14828 <= not w14560 and not w14827;
w14829 <= b(21) and not w14549;
w14830 <= not w14547 and w14829;
w14831 <= not w14551 and not w14830;
w14832 <= not w14828 and w14831;
w14833 <= not w14551 and not w14832;
w14834 <= b(22) and not w14540;
w14835 <= not w14538 and w14834;
w14836 <= not w14542 and not w14835;
w14837 <= not w14833 and w14836;
w14838 <= not w14542 and not w14837;
w14839 <= b(23) and not w14531;
w14840 <= not w14529 and w14839;
w14841 <= not w14533 and not w14840;
w14842 <= not w14838 and w14841;
w14843 <= not w14533 and not w14842;
w14844 <= b(24) and not w14522;
w14845 <= not w14520 and w14844;
w14846 <= not w14524 and not w14845;
w14847 <= not w14843 and w14846;
w14848 <= not w14524 and not w14847;
w14849 <= b(25) and not w14513;
w14850 <= not w14511 and w14849;
w14851 <= not w14515 and not w14850;
w14852 <= not w14848 and w14851;
w14853 <= not w14515 and not w14852;
w14854 <= b(26) and not w14504;
w14855 <= not w14502 and w14854;
w14856 <= not w14506 and not w14855;
w14857 <= not w14853 and w14856;
w14858 <= not w14506 and not w14857;
w14859 <= b(27) and not w14495;
w14860 <= not w14493 and w14859;
w14861 <= not w14497 and not w14860;
w14862 <= not w14858 and w14861;
w14863 <= not w14497 and not w14862;
w14864 <= b(28) and not w14486;
w14865 <= not w14484 and w14864;
w14866 <= not w14488 and not w14865;
w14867 <= not w14863 and w14866;
w14868 <= not w14488 and not w14867;
w14869 <= b(29) and not w14477;
w14870 <= not w14475 and w14869;
w14871 <= not w14479 and not w14870;
w14872 <= not w14868 and w14871;
w14873 <= not w14479 and not w14872;
w14874 <= b(30) and not w14468;
w14875 <= not w14466 and w14874;
w14876 <= not w14470 and not w14875;
w14877 <= not w14873 and w14876;
w14878 <= not w14470 and not w14877;
w14879 <= b(31) and not w14459;
w14880 <= not w14457 and w14879;
w14881 <= not w14461 and not w14880;
w14882 <= not w14878 and w14881;
w14883 <= not w14461 and not w14882;
w14884 <= b(32) and not w14450;
w14885 <= not w14448 and w14884;
w14886 <= not w14452 and not w14885;
w14887 <= not w14883 and w14886;
w14888 <= not w14452 and not w14887;
w14889 <= b(33) and not w14441;
w14890 <= not w14439 and w14889;
w14891 <= not w14443 and not w14890;
w14892 <= not w14888 and w14891;
w14893 <= not w14443 and not w14892;
w14894 <= b(34) and not w14432;
w14895 <= not w14430 and w14894;
w14896 <= not w14434 and not w14895;
w14897 <= not w14893 and w14896;
w14898 <= not w14434 and not w14897;
w14899 <= b(35) and not w14423;
w14900 <= not w14421 and w14899;
w14901 <= not w14425 and not w14900;
w14902 <= not w14898 and w14901;
w14903 <= not w14425 and not w14902;
w14904 <= b(36) and not w14414;
w14905 <= not w14412 and w14904;
w14906 <= not w14416 and not w14905;
w14907 <= not w14903 and w14906;
w14908 <= not w14416 and not w14907;
w14909 <= b(37) and not w14405;
w14910 <= not w14403 and w14909;
w14911 <= not w14407 and not w14910;
w14912 <= not w14908 and w14911;
w14913 <= not w14407 and not w14912;
w14914 <= b(38) and not w14396;
w14915 <= not w14394 and w14914;
w14916 <= not w14398 and not w14915;
w14917 <= not w14913 and w14916;
w14918 <= not w14398 and not w14917;
w14919 <= b(39) and not w14387;
w14920 <= not w14385 and w14919;
w14921 <= not w14389 and not w14920;
w14922 <= not w14918 and w14921;
w14923 <= not w14389 and not w14922;
w14924 <= b(40) and not w14378;
w14925 <= not w14376 and w14924;
w14926 <= not w14380 and not w14925;
w14927 <= not w14923 and w14926;
w14928 <= not w14380 and not w14927;
w14929 <= b(41) and not w14369;
w14930 <= not w14367 and w14929;
w14931 <= not w14371 and not w14930;
w14932 <= not w14928 and w14931;
w14933 <= not w14371 and not w14932;
w14934 <= b(42) and not w14360;
w14935 <= not w14358 and w14934;
w14936 <= not w14362 and not w14935;
w14937 <= not w14933 and w14936;
w14938 <= not w14362 and not w14937;
w14939 <= b(43) and not w14351;
w14940 <= not w14349 and w14939;
w14941 <= not w14353 and not w14940;
w14942 <= not w14938 and w14941;
w14943 <= not w14353 and not w14942;
w14944 <= b(44) and not w14331;
w14945 <= not w14329 and w14944;
w14946 <= not w14344 and not w14945;
w14947 <= not w14943 and w14946;
w14948 <= not w14344 and not w14947;
w14949 <= b(45) and not w14341;
w14950 <= not w14339 and w14949;
w14951 <= not w14343 and not w14950;
w14952 <= not w14948 and w14951;
w14953 <= not w14343 and not w14952;
w14954 <= w41 and w43;
w14955 <= w31 and w14954;
w14956 <= not w14953 and w14955;
w14957 <= not w14332 and not w14956;
w14958 <= not w14353 and w14946;
w14959 <= not w14942 and w14958;
w14960 <= not w14943 and not w14946;
w14961 <= not w14959 and not w14960;
w14962 <= w14955 and not w14961;
w14963 <= not w14953 and w14962;
w14964 <= not w14957 and not w14963;
w14965 <= not b(45) and not w14964;
w14966 <= not w14352 and not w14956;
w14967 <= not w14362 and w14941;
w14968 <= not w14937 and w14967;
w14969 <= not w14938 and not w14941;
w14970 <= not w14968 and not w14969;
w14971 <= w14955 and not w14970;
w14972 <= not w14953 and w14971;
w14973 <= not w14966 and not w14972;
w14974 <= not b(44) and not w14973;
w14975 <= not w14361 and not w14956;
w14976 <= not w14371 and w14936;
w14977 <= not w14932 and w14976;
w14978 <= not w14933 and not w14936;
w14979 <= not w14977 and not w14978;
w14980 <= w14955 and not w14979;
w14981 <= not w14953 and w14980;
w14982 <= not w14975 and not w14981;
w14983 <= not b(43) and not w14982;
w14984 <= not w14370 and not w14956;
w14985 <= not w14380 and w14931;
w14986 <= not w14927 and w14985;
w14987 <= not w14928 and not w14931;
w14988 <= not w14986 and not w14987;
w14989 <= w14955 and not w14988;
w14990 <= not w14953 and w14989;
w14991 <= not w14984 and not w14990;
w14992 <= not b(42) and not w14991;
w14993 <= not w14379 and not w14956;
w14994 <= not w14389 and w14926;
w14995 <= not w14922 and w14994;
w14996 <= not w14923 and not w14926;
w14997 <= not w14995 and not w14996;
w14998 <= w14955 and not w14997;
w14999 <= not w14953 and w14998;
w15000 <= not w14993 and not w14999;
w15001 <= not b(41) and not w15000;
w15002 <= not w14388 and not w14956;
w15003 <= not w14398 and w14921;
w15004 <= not w14917 and w15003;
w15005 <= not w14918 and not w14921;
w15006 <= not w15004 and not w15005;
w15007 <= w14955 and not w15006;
w15008 <= not w14953 and w15007;
w15009 <= not w15002 and not w15008;
w15010 <= not b(40) and not w15009;
w15011 <= not w14397 and not w14956;
w15012 <= not w14407 and w14916;
w15013 <= not w14912 and w15012;
w15014 <= not w14913 and not w14916;
w15015 <= not w15013 and not w15014;
w15016 <= w14955 and not w15015;
w15017 <= not w14953 and w15016;
w15018 <= not w15011 and not w15017;
w15019 <= not b(39) and not w15018;
w15020 <= not w14406 and not w14956;
w15021 <= not w14416 and w14911;
w15022 <= not w14907 and w15021;
w15023 <= not w14908 and not w14911;
w15024 <= not w15022 and not w15023;
w15025 <= w14955 and not w15024;
w15026 <= not w14953 and w15025;
w15027 <= not w15020 and not w15026;
w15028 <= not b(38) and not w15027;
w15029 <= not w14415 and not w14956;
w15030 <= not w14425 and w14906;
w15031 <= not w14902 and w15030;
w15032 <= not w14903 and not w14906;
w15033 <= not w15031 and not w15032;
w15034 <= w14955 and not w15033;
w15035 <= not w14953 and w15034;
w15036 <= not w15029 and not w15035;
w15037 <= not b(37) and not w15036;
w15038 <= not w14424 and not w14956;
w15039 <= not w14434 and w14901;
w15040 <= not w14897 and w15039;
w15041 <= not w14898 and not w14901;
w15042 <= not w15040 and not w15041;
w15043 <= w14955 and not w15042;
w15044 <= not w14953 and w15043;
w15045 <= not w15038 and not w15044;
w15046 <= not b(36) and not w15045;
w15047 <= not w14433 and not w14956;
w15048 <= not w14443 and w14896;
w15049 <= not w14892 and w15048;
w15050 <= not w14893 and not w14896;
w15051 <= not w15049 and not w15050;
w15052 <= w14955 and not w15051;
w15053 <= not w14953 and w15052;
w15054 <= not w15047 and not w15053;
w15055 <= not b(35) and not w15054;
w15056 <= not w14442 and not w14956;
w15057 <= not w14452 and w14891;
w15058 <= not w14887 and w15057;
w15059 <= not w14888 and not w14891;
w15060 <= not w15058 and not w15059;
w15061 <= w14955 and not w15060;
w15062 <= not w14953 and w15061;
w15063 <= not w15056 and not w15062;
w15064 <= not b(34) and not w15063;
w15065 <= not w14451 and not w14956;
w15066 <= not w14461 and w14886;
w15067 <= not w14882 and w15066;
w15068 <= not w14883 and not w14886;
w15069 <= not w15067 and not w15068;
w15070 <= w14955 and not w15069;
w15071 <= not w14953 and w15070;
w15072 <= not w15065 and not w15071;
w15073 <= not b(33) and not w15072;
w15074 <= not w14460 and not w14956;
w15075 <= not w14470 and w14881;
w15076 <= not w14877 and w15075;
w15077 <= not w14878 and not w14881;
w15078 <= not w15076 and not w15077;
w15079 <= w14955 and not w15078;
w15080 <= not w14953 and w15079;
w15081 <= not w15074 and not w15080;
w15082 <= not b(32) and not w15081;
w15083 <= not w14469 and not w14956;
w15084 <= not w14479 and w14876;
w15085 <= not w14872 and w15084;
w15086 <= not w14873 and not w14876;
w15087 <= not w15085 and not w15086;
w15088 <= w14955 and not w15087;
w15089 <= not w14953 and w15088;
w15090 <= not w15083 and not w15089;
w15091 <= not b(31) and not w15090;
w15092 <= not w14478 and not w14956;
w15093 <= not w14488 and w14871;
w15094 <= not w14867 and w15093;
w15095 <= not w14868 and not w14871;
w15096 <= not w15094 and not w15095;
w15097 <= w14955 and not w15096;
w15098 <= not w14953 and w15097;
w15099 <= not w15092 and not w15098;
w15100 <= not b(30) and not w15099;
w15101 <= not w14487 and not w14956;
w15102 <= not w14497 and w14866;
w15103 <= not w14862 and w15102;
w15104 <= not w14863 and not w14866;
w15105 <= not w15103 and not w15104;
w15106 <= w14955 and not w15105;
w15107 <= not w14953 and w15106;
w15108 <= not w15101 and not w15107;
w15109 <= not b(29) and not w15108;
w15110 <= not w14496 and not w14956;
w15111 <= not w14506 and w14861;
w15112 <= not w14857 and w15111;
w15113 <= not w14858 and not w14861;
w15114 <= not w15112 and not w15113;
w15115 <= w14955 and not w15114;
w15116 <= not w14953 and w15115;
w15117 <= not w15110 and not w15116;
w15118 <= not b(28) and not w15117;
w15119 <= not w14505 and not w14956;
w15120 <= not w14515 and w14856;
w15121 <= not w14852 and w15120;
w15122 <= not w14853 and not w14856;
w15123 <= not w15121 and not w15122;
w15124 <= w14955 and not w15123;
w15125 <= not w14953 and w15124;
w15126 <= not w15119 and not w15125;
w15127 <= not b(27) and not w15126;
w15128 <= not w14514 and not w14956;
w15129 <= not w14524 and w14851;
w15130 <= not w14847 and w15129;
w15131 <= not w14848 and not w14851;
w15132 <= not w15130 and not w15131;
w15133 <= w14955 and not w15132;
w15134 <= not w14953 and w15133;
w15135 <= not w15128 and not w15134;
w15136 <= not b(26) and not w15135;
w15137 <= not w14523 and not w14956;
w15138 <= not w14533 and w14846;
w15139 <= not w14842 and w15138;
w15140 <= not w14843 and not w14846;
w15141 <= not w15139 and not w15140;
w15142 <= w14955 and not w15141;
w15143 <= not w14953 and w15142;
w15144 <= not w15137 and not w15143;
w15145 <= not b(25) and not w15144;
w15146 <= not w14532 and not w14956;
w15147 <= not w14542 and w14841;
w15148 <= not w14837 and w15147;
w15149 <= not w14838 and not w14841;
w15150 <= not w15148 and not w15149;
w15151 <= w14955 and not w15150;
w15152 <= not w14953 and w15151;
w15153 <= not w15146 and not w15152;
w15154 <= not b(24) and not w15153;
w15155 <= not w14541 and not w14956;
w15156 <= not w14551 and w14836;
w15157 <= not w14832 and w15156;
w15158 <= not w14833 and not w14836;
w15159 <= not w15157 and not w15158;
w15160 <= w14955 and not w15159;
w15161 <= not w14953 and w15160;
w15162 <= not w15155 and not w15161;
w15163 <= not b(23) and not w15162;
w15164 <= not w14550 and not w14956;
w15165 <= not w14560 and w14831;
w15166 <= not w14827 and w15165;
w15167 <= not w14828 and not w14831;
w15168 <= not w15166 and not w15167;
w15169 <= w14955 and not w15168;
w15170 <= not w14953 and w15169;
w15171 <= not w15164 and not w15170;
w15172 <= not b(22) and not w15171;
w15173 <= not w14559 and not w14956;
w15174 <= not w14569 and w14826;
w15175 <= not w14822 and w15174;
w15176 <= not w14823 and not w14826;
w15177 <= not w15175 and not w15176;
w15178 <= w14955 and not w15177;
w15179 <= not w14953 and w15178;
w15180 <= not w15173 and not w15179;
w15181 <= not b(21) and not w15180;
w15182 <= not w14568 and not w14956;
w15183 <= not w14578 and w14821;
w15184 <= not w14817 and w15183;
w15185 <= not w14818 and not w14821;
w15186 <= not w15184 and not w15185;
w15187 <= w14955 and not w15186;
w15188 <= not w14953 and w15187;
w15189 <= not w15182 and not w15188;
w15190 <= not b(20) and not w15189;
w15191 <= not w14577 and not w14956;
w15192 <= not w14587 and w14816;
w15193 <= not w14812 and w15192;
w15194 <= not w14813 and not w14816;
w15195 <= not w15193 and not w15194;
w15196 <= w14955 and not w15195;
w15197 <= not w14953 and w15196;
w15198 <= not w15191 and not w15197;
w15199 <= not b(19) and not w15198;
w15200 <= not w14586 and not w14956;
w15201 <= not w14596 and w14811;
w15202 <= not w14807 and w15201;
w15203 <= not w14808 and not w14811;
w15204 <= not w15202 and not w15203;
w15205 <= w14955 and not w15204;
w15206 <= not w14953 and w15205;
w15207 <= not w15200 and not w15206;
w15208 <= not b(18) and not w15207;
w15209 <= not w14595 and not w14956;
w15210 <= not w14605 and w14806;
w15211 <= not w14802 and w15210;
w15212 <= not w14803 and not w14806;
w15213 <= not w15211 and not w15212;
w15214 <= w14955 and not w15213;
w15215 <= not w14953 and w15214;
w15216 <= not w15209 and not w15215;
w15217 <= not b(17) and not w15216;
w15218 <= not w14604 and not w14956;
w15219 <= not w14614 and w14801;
w15220 <= not w14797 and w15219;
w15221 <= not w14798 and not w14801;
w15222 <= not w15220 and not w15221;
w15223 <= w14955 and not w15222;
w15224 <= not w14953 and w15223;
w15225 <= not w15218 and not w15224;
w15226 <= not b(16) and not w15225;
w15227 <= not w14613 and not w14956;
w15228 <= not w14623 and w14796;
w15229 <= not w14792 and w15228;
w15230 <= not w14793 and not w14796;
w15231 <= not w15229 and not w15230;
w15232 <= w14955 and not w15231;
w15233 <= not w14953 and w15232;
w15234 <= not w15227 and not w15233;
w15235 <= not b(15) and not w15234;
w15236 <= not w14622 and not w14956;
w15237 <= not w14632 and w14791;
w15238 <= not w14787 and w15237;
w15239 <= not w14788 and not w14791;
w15240 <= not w15238 and not w15239;
w15241 <= w14955 and not w15240;
w15242 <= not w14953 and w15241;
w15243 <= not w15236 and not w15242;
w15244 <= not b(14) and not w15243;
w15245 <= not w14631 and not w14956;
w15246 <= not w14641 and w14786;
w15247 <= not w14782 and w15246;
w15248 <= not w14783 and not w14786;
w15249 <= not w15247 and not w15248;
w15250 <= w14955 and not w15249;
w15251 <= not w14953 and w15250;
w15252 <= not w15245 and not w15251;
w15253 <= not b(13) and not w15252;
w15254 <= not w14640 and not w14956;
w15255 <= not w14650 and w14781;
w15256 <= not w14777 and w15255;
w15257 <= not w14778 and not w14781;
w15258 <= not w15256 and not w15257;
w15259 <= w14955 and not w15258;
w15260 <= not w14953 and w15259;
w15261 <= not w15254 and not w15260;
w15262 <= not b(12) and not w15261;
w15263 <= not w14649 and not w14956;
w15264 <= not w14659 and w14776;
w15265 <= not w14772 and w15264;
w15266 <= not w14773 and not w14776;
w15267 <= not w15265 and not w15266;
w15268 <= w14955 and not w15267;
w15269 <= not w14953 and w15268;
w15270 <= not w15263 and not w15269;
w15271 <= not b(11) and not w15270;
w15272 <= not w14658 and not w14956;
w15273 <= not w14668 and w14771;
w15274 <= not w14767 and w15273;
w15275 <= not w14768 and not w14771;
w15276 <= not w15274 and not w15275;
w15277 <= w14955 and not w15276;
w15278 <= not w14953 and w15277;
w15279 <= not w15272 and not w15278;
w15280 <= not b(10) and not w15279;
w15281 <= not w14667 and not w14956;
w15282 <= not w14677 and w14766;
w15283 <= not w14762 and w15282;
w15284 <= not w14763 and not w14766;
w15285 <= not w15283 and not w15284;
w15286 <= w14955 and not w15285;
w15287 <= not w14953 and w15286;
w15288 <= not w15281 and not w15287;
w15289 <= not b(9) and not w15288;
w15290 <= not w14676 and not w14956;
w15291 <= not w14686 and w14761;
w15292 <= not w14757 and w15291;
w15293 <= not w14758 and not w14761;
w15294 <= not w15292 and not w15293;
w15295 <= w14955 and not w15294;
w15296 <= not w14953 and w15295;
w15297 <= not w15290 and not w15296;
w15298 <= not b(8) and not w15297;
w15299 <= not w14685 and not w14956;
w15300 <= not w14695 and w14756;
w15301 <= not w14752 and w15300;
w15302 <= not w14753 and not w14756;
w15303 <= not w15301 and not w15302;
w15304 <= w14955 and not w15303;
w15305 <= not w14953 and w15304;
w15306 <= not w15299 and not w15305;
w15307 <= not b(7) and not w15306;
w15308 <= not w14694 and not w14956;
w15309 <= not w14704 and w14751;
w15310 <= not w14747 and w15309;
w15311 <= not w14748 and not w14751;
w15312 <= not w15310 and not w15311;
w15313 <= w14955 and not w15312;
w15314 <= not w14953 and w15313;
w15315 <= not w15308 and not w15314;
w15316 <= not b(6) and not w15315;
w15317 <= not w14703 and not w14956;
w15318 <= not w14713 and w14746;
w15319 <= not w14742 and w15318;
w15320 <= not w14743 and not w14746;
w15321 <= not w15319 and not w15320;
w15322 <= w14955 and not w15321;
w15323 <= not w14953 and w15322;
w15324 <= not w15317 and not w15323;
w15325 <= not b(5) and not w15324;
w15326 <= not w14712 and not w14956;
w15327 <= not w14721 and w14741;
w15328 <= not w14737 and w15327;
w15329 <= not w14738 and not w14741;
w15330 <= not w15328 and not w15329;
w15331 <= w14955 and not w15330;
w15332 <= not w14953 and w15331;
w15333 <= not w15326 and not w15332;
w15334 <= not b(4) and not w15333;
w15335 <= not w14720 and not w14956;
w15336 <= not w14732 and w14736;
w15337 <= not w14731 and w15336;
w15338 <= not w14733 and not w14736;
w15339 <= not w15337 and not w15338;
w15340 <= w14955 and not w15339;
w15341 <= not w14953 and w15340;
w15342 <= not w15335 and not w15341;
w15343 <= not b(3) and not w15342;
w15344 <= not w14725 and not w14956;
w15345 <= not w14728 and w14730;
w15346 <= not w14726 and w15345;
w15347 <= w14955 and not w15346;
w15348 <= not w14731 and w15347;
w15349 <= not w14953 and w15348;
w15350 <= not w15344 and not w15349;
w15351 <= not b(2) and not w15350;
w15352 <= b(0) and not b(46);
w15353 <= w160 and w15352;
w15354 <= w143 and w15353;
w15355 <= w338 and w15354;
w15356 <= not w14953 and w15355;
w15357 <= a(18) and not w15356;
w15358 <= w43 and w14730;
w15359 <= w41 and w15358;
w15360 <= w31 and w15359;
w15361 <= not w14953 and w15360;
w15362 <= not w15357 and not w15361;
w15363 <= b(1) and not w15362;
w15364 <= not b(1) and not w15361;
w15365 <= not w15357 and w15364;
w15366 <= not w15363 and not w15365;
w15367 <= not a(17) and b(0);
w15368 <= not w15366 and not w15367;
w15369 <= not b(1) and not w15362;
w15370 <= not w15368 and not w15369;
w15371 <= b(2) and not w15349;
w15372 <= not w15344 and w15371;
w15373 <= not w15351 and not w15372;
w15374 <= not w15370 and w15373;
w15375 <= not w15351 and not w15374;
w15376 <= b(3) and not w15341;
w15377 <= not w15335 and w15376;
w15378 <= not w15343 and not w15377;
w15379 <= not w15375 and w15378;
w15380 <= not w15343 and not w15379;
w15381 <= b(4) and not w15332;
w15382 <= not w15326 and w15381;
w15383 <= not w15334 and not w15382;
w15384 <= not w15380 and w15383;
w15385 <= not w15334 and not w15384;
w15386 <= b(5) and not w15323;
w15387 <= not w15317 and w15386;
w15388 <= not w15325 and not w15387;
w15389 <= not w15385 and w15388;
w15390 <= not w15325 and not w15389;
w15391 <= b(6) and not w15314;
w15392 <= not w15308 and w15391;
w15393 <= not w15316 and not w15392;
w15394 <= not w15390 and w15393;
w15395 <= not w15316 and not w15394;
w15396 <= b(7) and not w15305;
w15397 <= not w15299 and w15396;
w15398 <= not w15307 and not w15397;
w15399 <= not w15395 and w15398;
w15400 <= not w15307 and not w15399;
w15401 <= b(8) and not w15296;
w15402 <= not w15290 and w15401;
w15403 <= not w15298 and not w15402;
w15404 <= not w15400 and w15403;
w15405 <= not w15298 and not w15404;
w15406 <= b(9) and not w15287;
w15407 <= not w15281 and w15406;
w15408 <= not w15289 and not w15407;
w15409 <= not w15405 and w15408;
w15410 <= not w15289 and not w15409;
w15411 <= b(10) and not w15278;
w15412 <= not w15272 and w15411;
w15413 <= not w15280 and not w15412;
w15414 <= not w15410 and w15413;
w15415 <= not w15280 and not w15414;
w15416 <= b(11) and not w15269;
w15417 <= not w15263 and w15416;
w15418 <= not w15271 and not w15417;
w15419 <= not w15415 and w15418;
w15420 <= not w15271 and not w15419;
w15421 <= b(12) and not w15260;
w15422 <= not w15254 and w15421;
w15423 <= not w15262 and not w15422;
w15424 <= not w15420 and w15423;
w15425 <= not w15262 and not w15424;
w15426 <= b(13) and not w15251;
w15427 <= not w15245 and w15426;
w15428 <= not w15253 and not w15427;
w15429 <= not w15425 and w15428;
w15430 <= not w15253 and not w15429;
w15431 <= b(14) and not w15242;
w15432 <= not w15236 and w15431;
w15433 <= not w15244 and not w15432;
w15434 <= not w15430 and w15433;
w15435 <= not w15244 and not w15434;
w15436 <= b(15) and not w15233;
w15437 <= not w15227 and w15436;
w15438 <= not w15235 and not w15437;
w15439 <= not w15435 and w15438;
w15440 <= not w15235 and not w15439;
w15441 <= b(16) and not w15224;
w15442 <= not w15218 and w15441;
w15443 <= not w15226 and not w15442;
w15444 <= not w15440 and w15443;
w15445 <= not w15226 and not w15444;
w15446 <= b(17) and not w15215;
w15447 <= not w15209 and w15446;
w15448 <= not w15217 and not w15447;
w15449 <= not w15445 and w15448;
w15450 <= not w15217 and not w15449;
w15451 <= b(18) and not w15206;
w15452 <= not w15200 and w15451;
w15453 <= not w15208 and not w15452;
w15454 <= not w15450 and w15453;
w15455 <= not w15208 and not w15454;
w15456 <= b(19) and not w15197;
w15457 <= not w15191 and w15456;
w15458 <= not w15199 and not w15457;
w15459 <= not w15455 and w15458;
w15460 <= not w15199 and not w15459;
w15461 <= b(20) and not w15188;
w15462 <= not w15182 and w15461;
w15463 <= not w15190 and not w15462;
w15464 <= not w15460 and w15463;
w15465 <= not w15190 and not w15464;
w15466 <= b(21) and not w15179;
w15467 <= not w15173 and w15466;
w15468 <= not w15181 and not w15467;
w15469 <= not w15465 and w15468;
w15470 <= not w15181 and not w15469;
w15471 <= b(22) and not w15170;
w15472 <= not w15164 and w15471;
w15473 <= not w15172 and not w15472;
w15474 <= not w15470 and w15473;
w15475 <= not w15172 and not w15474;
w15476 <= b(23) and not w15161;
w15477 <= not w15155 and w15476;
w15478 <= not w15163 and not w15477;
w15479 <= not w15475 and w15478;
w15480 <= not w15163 and not w15479;
w15481 <= b(24) and not w15152;
w15482 <= not w15146 and w15481;
w15483 <= not w15154 and not w15482;
w15484 <= not w15480 and w15483;
w15485 <= not w15154 and not w15484;
w15486 <= b(25) and not w15143;
w15487 <= not w15137 and w15486;
w15488 <= not w15145 and not w15487;
w15489 <= not w15485 and w15488;
w15490 <= not w15145 and not w15489;
w15491 <= b(26) and not w15134;
w15492 <= not w15128 and w15491;
w15493 <= not w15136 and not w15492;
w15494 <= not w15490 and w15493;
w15495 <= not w15136 and not w15494;
w15496 <= b(27) and not w15125;
w15497 <= not w15119 and w15496;
w15498 <= not w15127 and not w15497;
w15499 <= not w15495 and w15498;
w15500 <= not w15127 and not w15499;
w15501 <= b(28) and not w15116;
w15502 <= not w15110 and w15501;
w15503 <= not w15118 and not w15502;
w15504 <= not w15500 and w15503;
w15505 <= not w15118 and not w15504;
w15506 <= b(29) and not w15107;
w15507 <= not w15101 and w15506;
w15508 <= not w15109 and not w15507;
w15509 <= not w15505 and w15508;
w15510 <= not w15109 and not w15509;
w15511 <= b(30) and not w15098;
w15512 <= not w15092 and w15511;
w15513 <= not w15100 and not w15512;
w15514 <= not w15510 and w15513;
w15515 <= not w15100 and not w15514;
w15516 <= b(31) and not w15089;
w15517 <= not w15083 and w15516;
w15518 <= not w15091 and not w15517;
w15519 <= not w15515 and w15518;
w15520 <= not w15091 and not w15519;
w15521 <= b(32) and not w15080;
w15522 <= not w15074 and w15521;
w15523 <= not w15082 and not w15522;
w15524 <= not w15520 and w15523;
w15525 <= not w15082 and not w15524;
w15526 <= b(33) and not w15071;
w15527 <= not w15065 and w15526;
w15528 <= not w15073 and not w15527;
w15529 <= not w15525 and w15528;
w15530 <= not w15073 and not w15529;
w15531 <= b(34) and not w15062;
w15532 <= not w15056 and w15531;
w15533 <= not w15064 and not w15532;
w15534 <= not w15530 and w15533;
w15535 <= not w15064 and not w15534;
w15536 <= b(35) and not w15053;
w15537 <= not w15047 and w15536;
w15538 <= not w15055 and not w15537;
w15539 <= not w15535 and w15538;
w15540 <= not w15055 and not w15539;
w15541 <= b(36) and not w15044;
w15542 <= not w15038 and w15541;
w15543 <= not w15046 and not w15542;
w15544 <= not w15540 and w15543;
w15545 <= not w15046 and not w15544;
w15546 <= b(37) and not w15035;
w15547 <= not w15029 and w15546;
w15548 <= not w15037 and not w15547;
w15549 <= not w15545 and w15548;
w15550 <= not w15037 and not w15549;
w15551 <= b(38) and not w15026;
w15552 <= not w15020 and w15551;
w15553 <= not w15028 and not w15552;
w15554 <= not w15550 and w15553;
w15555 <= not w15028 and not w15554;
w15556 <= b(39) and not w15017;
w15557 <= not w15011 and w15556;
w15558 <= not w15019 and not w15557;
w15559 <= not w15555 and w15558;
w15560 <= not w15019 and not w15559;
w15561 <= b(40) and not w15008;
w15562 <= not w15002 and w15561;
w15563 <= not w15010 and not w15562;
w15564 <= not w15560 and w15563;
w15565 <= not w15010 and not w15564;
w15566 <= b(41) and not w14999;
w15567 <= not w14993 and w15566;
w15568 <= not w15001 and not w15567;
w15569 <= not w15565 and w15568;
w15570 <= not w15001 and not w15569;
w15571 <= b(42) and not w14990;
w15572 <= not w14984 and w15571;
w15573 <= not w14992 and not w15572;
w15574 <= not w15570 and w15573;
w15575 <= not w14992 and not w15574;
w15576 <= b(43) and not w14981;
w15577 <= not w14975 and w15576;
w15578 <= not w14983 and not w15577;
w15579 <= not w15575 and w15578;
w15580 <= not w14983 and not w15579;
w15581 <= b(44) and not w14972;
w15582 <= not w14966 and w15581;
w15583 <= not w14974 and not w15582;
w15584 <= not w15580 and w15583;
w15585 <= not w14974 and not w15584;
w15586 <= b(45) and not w14963;
w15587 <= not w14957 and w15586;
w15588 <= not w14965 and not w15587;
w15589 <= not w15585 and w15588;
w15590 <= not w14965 and not w15589;
w15591 <= not w14342 and not w14956;
w15592 <= not w14344 and w14951;
w15593 <= not w14947 and w15592;
w15594 <= not w14948 and not w14951;
w15595 <= not w15593 and not w15594;
w15596 <= w14956 and not w15595;
w15597 <= not w15591 and not w15596;
w15598 <= not b(46) and not w15597;
w15599 <= b(46) and not w15591;
w15600 <= not w15596 and w15599;
w15601 <= w143 and w160;
w15602 <= w338 and w15601;
w15603 <= not w15600 and w15602;
w15604 <= not w15598 and w15603;
w15605 <= not w15590 and w15604;
w15606 <= w14955 and not w15597;
w15607 <= not w15605 and not w15606;
w15608 <= not w14974 and w15588;
w15609 <= not w15584 and w15608;
w15610 <= not w15585 and not w15588;
w15611 <= not w15609 and not w15610;
w15612 <= not w15607 and not w15611;
w15613 <= not w14964 and not w15606;
w15614 <= not w15605 and w15613;
w15615 <= not w15612 and not w15614;
w15616 <= not b(46) and not w15615;
w15617 <= not w14983 and w15583;
w15618 <= not w15579 and w15617;
w15619 <= not w15580 and not w15583;
w15620 <= not w15618 and not w15619;
w15621 <= not w15607 and not w15620;
w15622 <= not w14973 and not w15606;
w15623 <= not w15605 and w15622;
w15624 <= not w15621 and not w15623;
w15625 <= not b(45) and not w15624;
w15626 <= not w14992 and w15578;
w15627 <= not w15574 and w15626;
w15628 <= not w15575 and not w15578;
w15629 <= not w15627 and not w15628;
w15630 <= not w15607 and not w15629;
w15631 <= not w14982 and not w15606;
w15632 <= not w15605 and w15631;
w15633 <= not w15630 and not w15632;
w15634 <= not b(44) and not w15633;
w15635 <= not w15001 and w15573;
w15636 <= not w15569 and w15635;
w15637 <= not w15570 and not w15573;
w15638 <= not w15636 and not w15637;
w15639 <= not w15607 and not w15638;
w15640 <= not w14991 and not w15606;
w15641 <= not w15605 and w15640;
w15642 <= not w15639 and not w15641;
w15643 <= not b(43) and not w15642;
w15644 <= not w15010 and w15568;
w15645 <= not w15564 and w15644;
w15646 <= not w15565 and not w15568;
w15647 <= not w15645 and not w15646;
w15648 <= not w15607 and not w15647;
w15649 <= not w15000 and not w15606;
w15650 <= not w15605 and w15649;
w15651 <= not w15648 and not w15650;
w15652 <= not b(42) and not w15651;
w15653 <= not w15019 and w15563;
w15654 <= not w15559 and w15653;
w15655 <= not w15560 and not w15563;
w15656 <= not w15654 and not w15655;
w15657 <= not w15607 and not w15656;
w15658 <= not w15009 and not w15606;
w15659 <= not w15605 and w15658;
w15660 <= not w15657 and not w15659;
w15661 <= not b(41) and not w15660;
w15662 <= not w15028 and w15558;
w15663 <= not w15554 and w15662;
w15664 <= not w15555 and not w15558;
w15665 <= not w15663 and not w15664;
w15666 <= not w15607 and not w15665;
w15667 <= not w15018 and not w15606;
w15668 <= not w15605 and w15667;
w15669 <= not w15666 and not w15668;
w15670 <= not b(40) and not w15669;
w15671 <= not w15037 and w15553;
w15672 <= not w15549 and w15671;
w15673 <= not w15550 and not w15553;
w15674 <= not w15672 and not w15673;
w15675 <= not w15607 and not w15674;
w15676 <= not w15027 and not w15606;
w15677 <= not w15605 and w15676;
w15678 <= not w15675 and not w15677;
w15679 <= not b(39) and not w15678;
w15680 <= not w15046 and w15548;
w15681 <= not w15544 and w15680;
w15682 <= not w15545 and not w15548;
w15683 <= not w15681 and not w15682;
w15684 <= not w15607 and not w15683;
w15685 <= not w15036 and not w15606;
w15686 <= not w15605 and w15685;
w15687 <= not w15684 and not w15686;
w15688 <= not b(38) and not w15687;
w15689 <= not w15055 and w15543;
w15690 <= not w15539 and w15689;
w15691 <= not w15540 and not w15543;
w15692 <= not w15690 and not w15691;
w15693 <= not w15607 and not w15692;
w15694 <= not w15045 and not w15606;
w15695 <= not w15605 and w15694;
w15696 <= not w15693 and not w15695;
w15697 <= not b(37) and not w15696;
w15698 <= not w15064 and w15538;
w15699 <= not w15534 and w15698;
w15700 <= not w15535 and not w15538;
w15701 <= not w15699 and not w15700;
w15702 <= not w15607 and not w15701;
w15703 <= not w15054 and not w15606;
w15704 <= not w15605 and w15703;
w15705 <= not w15702 and not w15704;
w15706 <= not b(36) and not w15705;
w15707 <= not w15073 and w15533;
w15708 <= not w15529 and w15707;
w15709 <= not w15530 and not w15533;
w15710 <= not w15708 and not w15709;
w15711 <= not w15607 and not w15710;
w15712 <= not w15063 and not w15606;
w15713 <= not w15605 and w15712;
w15714 <= not w15711 and not w15713;
w15715 <= not b(35) and not w15714;
w15716 <= not w15082 and w15528;
w15717 <= not w15524 and w15716;
w15718 <= not w15525 and not w15528;
w15719 <= not w15717 and not w15718;
w15720 <= not w15607 and not w15719;
w15721 <= not w15072 and not w15606;
w15722 <= not w15605 and w15721;
w15723 <= not w15720 and not w15722;
w15724 <= not b(34) and not w15723;
w15725 <= not w15091 and w15523;
w15726 <= not w15519 and w15725;
w15727 <= not w15520 and not w15523;
w15728 <= not w15726 and not w15727;
w15729 <= not w15607 and not w15728;
w15730 <= not w15081 and not w15606;
w15731 <= not w15605 and w15730;
w15732 <= not w15729 and not w15731;
w15733 <= not b(33) and not w15732;
w15734 <= not w15100 and w15518;
w15735 <= not w15514 and w15734;
w15736 <= not w15515 and not w15518;
w15737 <= not w15735 and not w15736;
w15738 <= not w15607 and not w15737;
w15739 <= not w15090 and not w15606;
w15740 <= not w15605 and w15739;
w15741 <= not w15738 and not w15740;
w15742 <= not b(32) and not w15741;
w15743 <= not w15109 and w15513;
w15744 <= not w15509 and w15743;
w15745 <= not w15510 and not w15513;
w15746 <= not w15744 and not w15745;
w15747 <= not w15607 and not w15746;
w15748 <= not w15099 and not w15606;
w15749 <= not w15605 and w15748;
w15750 <= not w15747 and not w15749;
w15751 <= not b(31) and not w15750;
w15752 <= not w15118 and w15508;
w15753 <= not w15504 and w15752;
w15754 <= not w15505 and not w15508;
w15755 <= not w15753 and not w15754;
w15756 <= not w15607 and not w15755;
w15757 <= not w15108 and not w15606;
w15758 <= not w15605 and w15757;
w15759 <= not w15756 and not w15758;
w15760 <= not b(30) and not w15759;
w15761 <= not w15127 and w15503;
w15762 <= not w15499 and w15761;
w15763 <= not w15500 and not w15503;
w15764 <= not w15762 and not w15763;
w15765 <= not w15607 and not w15764;
w15766 <= not w15117 and not w15606;
w15767 <= not w15605 and w15766;
w15768 <= not w15765 and not w15767;
w15769 <= not b(29) and not w15768;
w15770 <= not w15136 and w15498;
w15771 <= not w15494 and w15770;
w15772 <= not w15495 and not w15498;
w15773 <= not w15771 and not w15772;
w15774 <= not w15607 and not w15773;
w15775 <= not w15126 and not w15606;
w15776 <= not w15605 and w15775;
w15777 <= not w15774 and not w15776;
w15778 <= not b(28) and not w15777;
w15779 <= not w15145 and w15493;
w15780 <= not w15489 and w15779;
w15781 <= not w15490 and not w15493;
w15782 <= not w15780 and not w15781;
w15783 <= not w15607 and not w15782;
w15784 <= not w15135 and not w15606;
w15785 <= not w15605 and w15784;
w15786 <= not w15783 and not w15785;
w15787 <= not b(27) and not w15786;
w15788 <= not w15154 and w15488;
w15789 <= not w15484 and w15788;
w15790 <= not w15485 and not w15488;
w15791 <= not w15789 and not w15790;
w15792 <= not w15607 and not w15791;
w15793 <= not w15144 and not w15606;
w15794 <= not w15605 and w15793;
w15795 <= not w15792 and not w15794;
w15796 <= not b(26) and not w15795;
w15797 <= not w15163 and w15483;
w15798 <= not w15479 and w15797;
w15799 <= not w15480 and not w15483;
w15800 <= not w15798 and not w15799;
w15801 <= not w15607 and not w15800;
w15802 <= not w15153 and not w15606;
w15803 <= not w15605 and w15802;
w15804 <= not w15801 and not w15803;
w15805 <= not b(25) and not w15804;
w15806 <= not w15172 and w15478;
w15807 <= not w15474 and w15806;
w15808 <= not w15475 and not w15478;
w15809 <= not w15807 and not w15808;
w15810 <= not w15607 and not w15809;
w15811 <= not w15162 and not w15606;
w15812 <= not w15605 and w15811;
w15813 <= not w15810 and not w15812;
w15814 <= not b(24) and not w15813;
w15815 <= not w15181 and w15473;
w15816 <= not w15469 and w15815;
w15817 <= not w15470 and not w15473;
w15818 <= not w15816 and not w15817;
w15819 <= not w15607 and not w15818;
w15820 <= not w15171 and not w15606;
w15821 <= not w15605 and w15820;
w15822 <= not w15819 and not w15821;
w15823 <= not b(23) and not w15822;
w15824 <= not w15190 and w15468;
w15825 <= not w15464 and w15824;
w15826 <= not w15465 and not w15468;
w15827 <= not w15825 and not w15826;
w15828 <= not w15607 and not w15827;
w15829 <= not w15180 and not w15606;
w15830 <= not w15605 and w15829;
w15831 <= not w15828 and not w15830;
w15832 <= not b(22) and not w15831;
w15833 <= not w15199 and w15463;
w15834 <= not w15459 and w15833;
w15835 <= not w15460 and not w15463;
w15836 <= not w15834 and not w15835;
w15837 <= not w15607 and not w15836;
w15838 <= not w15189 and not w15606;
w15839 <= not w15605 and w15838;
w15840 <= not w15837 and not w15839;
w15841 <= not b(21) and not w15840;
w15842 <= not w15208 and w15458;
w15843 <= not w15454 and w15842;
w15844 <= not w15455 and not w15458;
w15845 <= not w15843 and not w15844;
w15846 <= not w15607 and not w15845;
w15847 <= not w15198 and not w15606;
w15848 <= not w15605 and w15847;
w15849 <= not w15846 and not w15848;
w15850 <= not b(20) and not w15849;
w15851 <= not w15217 and w15453;
w15852 <= not w15449 and w15851;
w15853 <= not w15450 and not w15453;
w15854 <= not w15852 and not w15853;
w15855 <= not w15607 and not w15854;
w15856 <= not w15207 and not w15606;
w15857 <= not w15605 and w15856;
w15858 <= not w15855 and not w15857;
w15859 <= not b(19) and not w15858;
w15860 <= not w15226 and w15448;
w15861 <= not w15444 and w15860;
w15862 <= not w15445 and not w15448;
w15863 <= not w15861 and not w15862;
w15864 <= not w15607 and not w15863;
w15865 <= not w15216 and not w15606;
w15866 <= not w15605 and w15865;
w15867 <= not w15864 and not w15866;
w15868 <= not b(18) and not w15867;
w15869 <= not w15235 and w15443;
w15870 <= not w15439 and w15869;
w15871 <= not w15440 and not w15443;
w15872 <= not w15870 and not w15871;
w15873 <= not w15607 and not w15872;
w15874 <= not w15225 and not w15606;
w15875 <= not w15605 and w15874;
w15876 <= not w15873 and not w15875;
w15877 <= not b(17) and not w15876;
w15878 <= not w15244 and w15438;
w15879 <= not w15434 and w15878;
w15880 <= not w15435 and not w15438;
w15881 <= not w15879 and not w15880;
w15882 <= not w15607 and not w15881;
w15883 <= not w15234 and not w15606;
w15884 <= not w15605 and w15883;
w15885 <= not w15882 and not w15884;
w15886 <= not b(16) and not w15885;
w15887 <= not w15253 and w15433;
w15888 <= not w15429 and w15887;
w15889 <= not w15430 and not w15433;
w15890 <= not w15888 and not w15889;
w15891 <= not w15607 and not w15890;
w15892 <= not w15243 and not w15606;
w15893 <= not w15605 and w15892;
w15894 <= not w15891 and not w15893;
w15895 <= not b(15) and not w15894;
w15896 <= not w15262 and w15428;
w15897 <= not w15424 and w15896;
w15898 <= not w15425 and not w15428;
w15899 <= not w15897 and not w15898;
w15900 <= not w15607 and not w15899;
w15901 <= not w15252 and not w15606;
w15902 <= not w15605 and w15901;
w15903 <= not w15900 and not w15902;
w15904 <= not b(14) and not w15903;
w15905 <= not w15271 and w15423;
w15906 <= not w15419 and w15905;
w15907 <= not w15420 and not w15423;
w15908 <= not w15906 and not w15907;
w15909 <= not w15607 and not w15908;
w15910 <= not w15261 and not w15606;
w15911 <= not w15605 and w15910;
w15912 <= not w15909 and not w15911;
w15913 <= not b(13) and not w15912;
w15914 <= not w15280 and w15418;
w15915 <= not w15414 and w15914;
w15916 <= not w15415 and not w15418;
w15917 <= not w15915 and not w15916;
w15918 <= not w15607 and not w15917;
w15919 <= not w15270 and not w15606;
w15920 <= not w15605 and w15919;
w15921 <= not w15918 and not w15920;
w15922 <= not b(12) and not w15921;
w15923 <= not w15289 and w15413;
w15924 <= not w15409 and w15923;
w15925 <= not w15410 and not w15413;
w15926 <= not w15924 and not w15925;
w15927 <= not w15607 and not w15926;
w15928 <= not w15279 and not w15606;
w15929 <= not w15605 and w15928;
w15930 <= not w15927 and not w15929;
w15931 <= not b(11) and not w15930;
w15932 <= not w15298 and w15408;
w15933 <= not w15404 and w15932;
w15934 <= not w15405 and not w15408;
w15935 <= not w15933 and not w15934;
w15936 <= not w15607 and not w15935;
w15937 <= not w15288 and not w15606;
w15938 <= not w15605 and w15937;
w15939 <= not w15936 and not w15938;
w15940 <= not b(10) and not w15939;
w15941 <= not w15307 and w15403;
w15942 <= not w15399 and w15941;
w15943 <= not w15400 and not w15403;
w15944 <= not w15942 and not w15943;
w15945 <= not w15607 and not w15944;
w15946 <= not w15297 and not w15606;
w15947 <= not w15605 and w15946;
w15948 <= not w15945 and not w15947;
w15949 <= not b(9) and not w15948;
w15950 <= not w15316 and w15398;
w15951 <= not w15394 and w15950;
w15952 <= not w15395 and not w15398;
w15953 <= not w15951 and not w15952;
w15954 <= not w15607 and not w15953;
w15955 <= not w15306 and not w15606;
w15956 <= not w15605 and w15955;
w15957 <= not w15954 and not w15956;
w15958 <= not b(8) and not w15957;
w15959 <= not w15325 and w15393;
w15960 <= not w15389 and w15959;
w15961 <= not w15390 and not w15393;
w15962 <= not w15960 and not w15961;
w15963 <= not w15607 and not w15962;
w15964 <= not w15315 and not w15606;
w15965 <= not w15605 and w15964;
w15966 <= not w15963 and not w15965;
w15967 <= not b(7) and not w15966;
w15968 <= not w15334 and w15388;
w15969 <= not w15384 and w15968;
w15970 <= not w15385 and not w15388;
w15971 <= not w15969 and not w15970;
w15972 <= not w15607 and not w15971;
w15973 <= not w15324 and not w15606;
w15974 <= not w15605 and w15973;
w15975 <= not w15972 and not w15974;
w15976 <= not b(6) and not w15975;
w15977 <= not w15343 and w15383;
w15978 <= not w15379 and w15977;
w15979 <= not w15380 and not w15383;
w15980 <= not w15978 and not w15979;
w15981 <= not w15607 and not w15980;
w15982 <= not w15333 and not w15606;
w15983 <= not w15605 and w15982;
w15984 <= not w15981 and not w15983;
w15985 <= not b(5) and not w15984;
w15986 <= not w15351 and w15378;
w15987 <= not w15374 and w15986;
w15988 <= not w15375 and not w15378;
w15989 <= not w15987 and not w15988;
w15990 <= not w15607 and not w15989;
w15991 <= not w15342 and not w15606;
w15992 <= not w15605 and w15991;
w15993 <= not w15990 and not w15992;
w15994 <= not b(4) and not w15993;
w15995 <= not w15369 and w15373;
w15996 <= not w15368 and w15995;
w15997 <= not w15370 and not w15373;
w15998 <= not w15996 and not w15997;
w15999 <= not w15607 and not w15998;
w16000 <= not w15350 and not w15606;
w16001 <= not w15605 and w16000;
w16002 <= not w15999 and not w16001;
w16003 <= not b(3) and not w16002;
w16004 <= not w15365 and w15367;
w16005 <= not w15363 and w16004;
w16006 <= not w15368 and not w16005;
w16007 <= not w15607 and w16006;
w16008 <= not w15362 and not w15606;
w16009 <= not w15605 and w16008;
w16010 <= not w16007 and not w16009;
w16011 <= not b(2) and not w16010;
w16012 <= b(0) and not w15607;
w16013 <= a(17) and not w16012;
w16014 <= w15367 and not w15607;
w16015 <= not w16013 and not w16014;
w16016 <= b(1) and not w16015;
w16017 <= not b(1) and not w16014;
w16018 <= not w16013 and w16017;
w16019 <= not w16016 and not w16018;
w16020 <= not a(16) and b(0);
w16021 <= not w16019 and not w16020;
w16022 <= not b(1) and not w16015;
w16023 <= not w16021 and not w16022;
w16024 <= b(2) and not w16009;
w16025 <= not w16007 and w16024;
w16026 <= not w16011 and not w16025;
w16027 <= not w16023 and w16026;
w16028 <= not w16011 and not w16027;
w16029 <= b(3) and not w16001;
w16030 <= not w15999 and w16029;
w16031 <= not w16003 and not w16030;
w16032 <= not w16028 and w16031;
w16033 <= not w16003 and not w16032;
w16034 <= b(4) and not w15992;
w16035 <= not w15990 and w16034;
w16036 <= not w15994 and not w16035;
w16037 <= not w16033 and w16036;
w16038 <= not w15994 and not w16037;
w16039 <= b(5) and not w15983;
w16040 <= not w15981 and w16039;
w16041 <= not w15985 and not w16040;
w16042 <= not w16038 and w16041;
w16043 <= not w15985 and not w16042;
w16044 <= b(6) and not w15974;
w16045 <= not w15972 and w16044;
w16046 <= not w15976 and not w16045;
w16047 <= not w16043 and w16046;
w16048 <= not w15976 and not w16047;
w16049 <= b(7) and not w15965;
w16050 <= not w15963 and w16049;
w16051 <= not w15967 and not w16050;
w16052 <= not w16048 and w16051;
w16053 <= not w15967 and not w16052;
w16054 <= b(8) and not w15956;
w16055 <= not w15954 and w16054;
w16056 <= not w15958 and not w16055;
w16057 <= not w16053 and w16056;
w16058 <= not w15958 and not w16057;
w16059 <= b(9) and not w15947;
w16060 <= not w15945 and w16059;
w16061 <= not w15949 and not w16060;
w16062 <= not w16058 and w16061;
w16063 <= not w15949 and not w16062;
w16064 <= b(10) and not w15938;
w16065 <= not w15936 and w16064;
w16066 <= not w15940 and not w16065;
w16067 <= not w16063 and w16066;
w16068 <= not w15940 and not w16067;
w16069 <= b(11) and not w15929;
w16070 <= not w15927 and w16069;
w16071 <= not w15931 and not w16070;
w16072 <= not w16068 and w16071;
w16073 <= not w15931 and not w16072;
w16074 <= b(12) and not w15920;
w16075 <= not w15918 and w16074;
w16076 <= not w15922 and not w16075;
w16077 <= not w16073 and w16076;
w16078 <= not w15922 and not w16077;
w16079 <= b(13) and not w15911;
w16080 <= not w15909 and w16079;
w16081 <= not w15913 and not w16080;
w16082 <= not w16078 and w16081;
w16083 <= not w15913 and not w16082;
w16084 <= b(14) and not w15902;
w16085 <= not w15900 and w16084;
w16086 <= not w15904 and not w16085;
w16087 <= not w16083 and w16086;
w16088 <= not w15904 and not w16087;
w16089 <= b(15) and not w15893;
w16090 <= not w15891 and w16089;
w16091 <= not w15895 and not w16090;
w16092 <= not w16088 and w16091;
w16093 <= not w15895 and not w16092;
w16094 <= b(16) and not w15884;
w16095 <= not w15882 and w16094;
w16096 <= not w15886 and not w16095;
w16097 <= not w16093 and w16096;
w16098 <= not w15886 and not w16097;
w16099 <= b(17) and not w15875;
w16100 <= not w15873 and w16099;
w16101 <= not w15877 and not w16100;
w16102 <= not w16098 and w16101;
w16103 <= not w15877 and not w16102;
w16104 <= b(18) and not w15866;
w16105 <= not w15864 and w16104;
w16106 <= not w15868 and not w16105;
w16107 <= not w16103 and w16106;
w16108 <= not w15868 and not w16107;
w16109 <= b(19) and not w15857;
w16110 <= not w15855 and w16109;
w16111 <= not w15859 and not w16110;
w16112 <= not w16108 and w16111;
w16113 <= not w15859 and not w16112;
w16114 <= b(20) and not w15848;
w16115 <= not w15846 and w16114;
w16116 <= not w15850 and not w16115;
w16117 <= not w16113 and w16116;
w16118 <= not w15850 and not w16117;
w16119 <= b(21) and not w15839;
w16120 <= not w15837 and w16119;
w16121 <= not w15841 and not w16120;
w16122 <= not w16118 and w16121;
w16123 <= not w15841 and not w16122;
w16124 <= b(22) and not w15830;
w16125 <= not w15828 and w16124;
w16126 <= not w15832 and not w16125;
w16127 <= not w16123 and w16126;
w16128 <= not w15832 and not w16127;
w16129 <= b(23) and not w15821;
w16130 <= not w15819 and w16129;
w16131 <= not w15823 and not w16130;
w16132 <= not w16128 and w16131;
w16133 <= not w15823 and not w16132;
w16134 <= b(24) and not w15812;
w16135 <= not w15810 and w16134;
w16136 <= not w15814 and not w16135;
w16137 <= not w16133 and w16136;
w16138 <= not w15814 and not w16137;
w16139 <= b(25) and not w15803;
w16140 <= not w15801 and w16139;
w16141 <= not w15805 and not w16140;
w16142 <= not w16138 and w16141;
w16143 <= not w15805 and not w16142;
w16144 <= b(26) and not w15794;
w16145 <= not w15792 and w16144;
w16146 <= not w15796 and not w16145;
w16147 <= not w16143 and w16146;
w16148 <= not w15796 and not w16147;
w16149 <= b(27) and not w15785;
w16150 <= not w15783 and w16149;
w16151 <= not w15787 and not w16150;
w16152 <= not w16148 and w16151;
w16153 <= not w15787 and not w16152;
w16154 <= b(28) and not w15776;
w16155 <= not w15774 and w16154;
w16156 <= not w15778 and not w16155;
w16157 <= not w16153 and w16156;
w16158 <= not w15778 and not w16157;
w16159 <= b(29) and not w15767;
w16160 <= not w15765 and w16159;
w16161 <= not w15769 and not w16160;
w16162 <= not w16158 and w16161;
w16163 <= not w15769 and not w16162;
w16164 <= b(30) and not w15758;
w16165 <= not w15756 and w16164;
w16166 <= not w15760 and not w16165;
w16167 <= not w16163 and w16166;
w16168 <= not w15760 and not w16167;
w16169 <= b(31) and not w15749;
w16170 <= not w15747 and w16169;
w16171 <= not w15751 and not w16170;
w16172 <= not w16168 and w16171;
w16173 <= not w15751 and not w16172;
w16174 <= b(32) and not w15740;
w16175 <= not w15738 and w16174;
w16176 <= not w15742 and not w16175;
w16177 <= not w16173 and w16176;
w16178 <= not w15742 and not w16177;
w16179 <= b(33) and not w15731;
w16180 <= not w15729 and w16179;
w16181 <= not w15733 and not w16180;
w16182 <= not w16178 and w16181;
w16183 <= not w15733 and not w16182;
w16184 <= b(34) and not w15722;
w16185 <= not w15720 and w16184;
w16186 <= not w15724 and not w16185;
w16187 <= not w16183 and w16186;
w16188 <= not w15724 and not w16187;
w16189 <= b(35) and not w15713;
w16190 <= not w15711 and w16189;
w16191 <= not w15715 and not w16190;
w16192 <= not w16188 and w16191;
w16193 <= not w15715 and not w16192;
w16194 <= b(36) and not w15704;
w16195 <= not w15702 and w16194;
w16196 <= not w15706 and not w16195;
w16197 <= not w16193 and w16196;
w16198 <= not w15706 and not w16197;
w16199 <= b(37) and not w15695;
w16200 <= not w15693 and w16199;
w16201 <= not w15697 and not w16200;
w16202 <= not w16198 and w16201;
w16203 <= not w15697 and not w16202;
w16204 <= b(38) and not w15686;
w16205 <= not w15684 and w16204;
w16206 <= not w15688 and not w16205;
w16207 <= not w16203 and w16206;
w16208 <= not w15688 and not w16207;
w16209 <= b(39) and not w15677;
w16210 <= not w15675 and w16209;
w16211 <= not w15679 and not w16210;
w16212 <= not w16208 and w16211;
w16213 <= not w15679 and not w16212;
w16214 <= b(40) and not w15668;
w16215 <= not w15666 and w16214;
w16216 <= not w15670 and not w16215;
w16217 <= not w16213 and w16216;
w16218 <= not w15670 and not w16217;
w16219 <= b(41) and not w15659;
w16220 <= not w15657 and w16219;
w16221 <= not w15661 and not w16220;
w16222 <= not w16218 and w16221;
w16223 <= not w15661 and not w16222;
w16224 <= b(42) and not w15650;
w16225 <= not w15648 and w16224;
w16226 <= not w15652 and not w16225;
w16227 <= not w16223 and w16226;
w16228 <= not w15652 and not w16227;
w16229 <= b(43) and not w15641;
w16230 <= not w15639 and w16229;
w16231 <= not w15643 and not w16230;
w16232 <= not w16228 and w16231;
w16233 <= not w15643 and not w16232;
w16234 <= b(44) and not w15632;
w16235 <= not w15630 and w16234;
w16236 <= not w15634 and not w16235;
w16237 <= not w16233 and w16236;
w16238 <= not w15634 and not w16237;
w16239 <= b(45) and not w15623;
w16240 <= not w15621 and w16239;
w16241 <= not w15625 and not w16240;
w16242 <= not w16238 and w16241;
w16243 <= not w15625 and not w16242;
w16244 <= b(46) and not w15614;
w16245 <= not w15612 and w16244;
w16246 <= not w15616 and not w16245;
w16247 <= not w16243 and w16246;
w16248 <= not w15616 and not w16247;
w16249 <= not w14965 and not w15600;
w16250 <= not w15598 and w16249;
w16251 <= not w15589 and w16250;
w16252 <= not w15598 and not w15600;
w16253 <= not w15590 and not w16252;
w16254 <= not w16251 and not w16253;
w16255 <= not w15607 and not w16254;
w16256 <= not w15597 and not w15606;
w16257 <= not w15605 and w16256;
w16258 <= not w16255 and not w16257;
w16259 <= not b(47) and not w16258;
w16260 <= b(47) and not w16257;
w16261 <= not w16255 and w16260;
w16262 <= w81 and not w16261;
w16263 <= not w16259 and w16262;
w16264 <= not w16248 and w16263;
w16265 <= w15602 and not w16258;
w16266 <= not w16264 and not w16265;
w16267 <= not w15625 and w16246;
w16268 <= not w16242 and w16267;
w16269 <= not w16243 and not w16246;
w16270 <= not w16268 and not w16269;
w16271 <= not w16266 and not w16270;
w16272 <= not w15615 and not w16265;
w16273 <= not w16264 and w16272;
w16274 <= not w16271 and not w16273;
w16275 <= not w15616 and not w16261;
w16276 <= not w16259 and w16275;
w16277 <= not w16247 and w16276;
w16278 <= not w16259 and not w16261;
w16279 <= not w16248 and not w16278;
w16280 <= not w16277 and not w16279;
w16281 <= not w16266 and not w16280;
w16282 <= not w16258 and not w16265;
w16283 <= not w16264 and w16282;
w16284 <= not w16281 and not w16283;
w16285 <= not b(48) and not w16284;
w16286 <= not b(47) and not w16274;
w16287 <= not w15634 and w16241;
w16288 <= not w16237 and w16287;
w16289 <= not w16238 and not w16241;
w16290 <= not w16288 and not w16289;
w16291 <= not w16266 and not w16290;
w16292 <= not w15624 and not w16265;
w16293 <= not w16264 and w16292;
w16294 <= not w16291 and not w16293;
w16295 <= not b(46) and not w16294;
w16296 <= not w15643 and w16236;
w16297 <= not w16232 and w16296;
w16298 <= not w16233 and not w16236;
w16299 <= not w16297 and not w16298;
w16300 <= not w16266 and not w16299;
w16301 <= not w15633 and not w16265;
w16302 <= not w16264 and w16301;
w16303 <= not w16300 and not w16302;
w16304 <= not b(45) and not w16303;
w16305 <= not w15652 and w16231;
w16306 <= not w16227 and w16305;
w16307 <= not w16228 and not w16231;
w16308 <= not w16306 and not w16307;
w16309 <= not w16266 and not w16308;
w16310 <= not w15642 and not w16265;
w16311 <= not w16264 and w16310;
w16312 <= not w16309 and not w16311;
w16313 <= not b(44) and not w16312;
w16314 <= not w15661 and w16226;
w16315 <= not w16222 and w16314;
w16316 <= not w16223 and not w16226;
w16317 <= not w16315 and not w16316;
w16318 <= not w16266 and not w16317;
w16319 <= not w15651 and not w16265;
w16320 <= not w16264 and w16319;
w16321 <= not w16318 and not w16320;
w16322 <= not b(43) and not w16321;
w16323 <= not w15670 and w16221;
w16324 <= not w16217 and w16323;
w16325 <= not w16218 and not w16221;
w16326 <= not w16324 and not w16325;
w16327 <= not w16266 and not w16326;
w16328 <= not w15660 and not w16265;
w16329 <= not w16264 and w16328;
w16330 <= not w16327 and not w16329;
w16331 <= not b(42) and not w16330;
w16332 <= not w15679 and w16216;
w16333 <= not w16212 and w16332;
w16334 <= not w16213 and not w16216;
w16335 <= not w16333 and not w16334;
w16336 <= not w16266 and not w16335;
w16337 <= not w15669 and not w16265;
w16338 <= not w16264 and w16337;
w16339 <= not w16336 and not w16338;
w16340 <= not b(41) and not w16339;
w16341 <= not w15688 and w16211;
w16342 <= not w16207 and w16341;
w16343 <= not w16208 and not w16211;
w16344 <= not w16342 and not w16343;
w16345 <= not w16266 and not w16344;
w16346 <= not w15678 and not w16265;
w16347 <= not w16264 and w16346;
w16348 <= not w16345 and not w16347;
w16349 <= not b(40) and not w16348;
w16350 <= not w15697 and w16206;
w16351 <= not w16202 and w16350;
w16352 <= not w16203 and not w16206;
w16353 <= not w16351 and not w16352;
w16354 <= not w16266 and not w16353;
w16355 <= not w15687 and not w16265;
w16356 <= not w16264 and w16355;
w16357 <= not w16354 and not w16356;
w16358 <= not b(39) and not w16357;
w16359 <= not w15706 and w16201;
w16360 <= not w16197 and w16359;
w16361 <= not w16198 and not w16201;
w16362 <= not w16360 and not w16361;
w16363 <= not w16266 and not w16362;
w16364 <= not w15696 and not w16265;
w16365 <= not w16264 and w16364;
w16366 <= not w16363 and not w16365;
w16367 <= not b(38) and not w16366;
w16368 <= not w15715 and w16196;
w16369 <= not w16192 and w16368;
w16370 <= not w16193 and not w16196;
w16371 <= not w16369 and not w16370;
w16372 <= not w16266 and not w16371;
w16373 <= not w15705 and not w16265;
w16374 <= not w16264 and w16373;
w16375 <= not w16372 and not w16374;
w16376 <= not b(37) and not w16375;
w16377 <= not w15724 and w16191;
w16378 <= not w16187 and w16377;
w16379 <= not w16188 and not w16191;
w16380 <= not w16378 and not w16379;
w16381 <= not w16266 and not w16380;
w16382 <= not w15714 and not w16265;
w16383 <= not w16264 and w16382;
w16384 <= not w16381 and not w16383;
w16385 <= not b(36) and not w16384;
w16386 <= not w15733 and w16186;
w16387 <= not w16182 and w16386;
w16388 <= not w16183 and not w16186;
w16389 <= not w16387 and not w16388;
w16390 <= not w16266 and not w16389;
w16391 <= not w15723 and not w16265;
w16392 <= not w16264 and w16391;
w16393 <= not w16390 and not w16392;
w16394 <= not b(35) and not w16393;
w16395 <= not w15742 and w16181;
w16396 <= not w16177 and w16395;
w16397 <= not w16178 and not w16181;
w16398 <= not w16396 and not w16397;
w16399 <= not w16266 and not w16398;
w16400 <= not w15732 and not w16265;
w16401 <= not w16264 and w16400;
w16402 <= not w16399 and not w16401;
w16403 <= not b(34) and not w16402;
w16404 <= not w15751 and w16176;
w16405 <= not w16172 and w16404;
w16406 <= not w16173 and not w16176;
w16407 <= not w16405 and not w16406;
w16408 <= not w16266 and not w16407;
w16409 <= not w15741 and not w16265;
w16410 <= not w16264 and w16409;
w16411 <= not w16408 and not w16410;
w16412 <= not b(33) and not w16411;
w16413 <= not w15760 and w16171;
w16414 <= not w16167 and w16413;
w16415 <= not w16168 and not w16171;
w16416 <= not w16414 and not w16415;
w16417 <= not w16266 and not w16416;
w16418 <= not w15750 and not w16265;
w16419 <= not w16264 and w16418;
w16420 <= not w16417 and not w16419;
w16421 <= not b(32) and not w16420;
w16422 <= not w15769 and w16166;
w16423 <= not w16162 and w16422;
w16424 <= not w16163 and not w16166;
w16425 <= not w16423 and not w16424;
w16426 <= not w16266 and not w16425;
w16427 <= not w15759 and not w16265;
w16428 <= not w16264 and w16427;
w16429 <= not w16426 and not w16428;
w16430 <= not b(31) and not w16429;
w16431 <= not w15778 and w16161;
w16432 <= not w16157 and w16431;
w16433 <= not w16158 and not w16161;
w16434 <= not w16432 and not w16433;
w16435 <= not w16266 and not w16434;
w16436 <= not w15768 and not w16265;
w16437 <= not w16264 and w16436;
w16438 <= not w16435 and not w16437;
w16439 <= not b(30) and not w16438;
w16440 <= not w15787 and w16156;
w16441 <= not w16152 and w16440;
w16442 <= not w16153 and not w16156;
w16443 <= not w16441 and not w16442;
w16444 <= not w16266 and not w16443;
w16445 <= not w15777 and not w16265;
w16446 <= not w16264 and w16445;
w16447 <= not w16444 and not w16446;
w16448 <= not b(29) and not w16447;
w16449 <= not w15796 and w16151;
w16450 <= not w16147 and w16449;
w16451 <= not w16148 and not w16151;
w16452 <= not w16450 and not w16451;
w16453 <= not w16266 and not w16452;
w16454 <= not w15786 and not w16265;
w16455 <= not w16264 and w16454;
w16456 <= not w16453 and not w16455;
w16457 <= not b(28) and not w16456;
w16458 <= not w15805 and w16146;
w16459 <= not w16142 and w16458;
w16460 <= not w16143 and not w16146;
w16461 <= not w16459 and not w16460;
w16462 <= not w16266 and not w16461;
w16463 <= not w15795 and not w16265;
w16464 <= not w16264 and w16463;
w16465 <= not w16462 and not w16464;
w16466 <= not b(27) and not w16465;
w16467 <= not w15814 and w16141;
w16468 <= not w16137 and w16467;
w16469 <= not w16138 and not w16141;
w16470 <= not w16468 and not w16469;
w16471 <= not w16266 and not w16470;
w16472 <= not w15804 and not w16265;
w16473 <= not w16264 and w16472;
w16474 <= not w16471 and not w16473;
w16475 <= not b(26) and not w16474;
w16476 <= not w15823 and w16136;
w16477 <= not w16132 and w16476;
w16478 <= not w16133 and not w16136;
w16479 <= not w16477 and not w16478;
w16480 <= not w16266 and not w16479;
w16481 <= not w15813 and not w16265;
w16482 <= not w16264 and w16481;
w16483 <= not w16480 and not w16482;
w16484 <= not b(25) and not w16483;
w16485 <= not w15832 and w16131;
w16486 <= not w16127 and w16485;
w16487 <= not w16128 and not w16131;
w16488 <= not w16486 and not w16487;
w16489 <= not w16266 and not w16488;
w16490 <= not w15822 and not w16265;
w16491 <= not w16264 and w16490;
w16492 <= not w16489 and not w16491;
w16493 <= not b(24) and not w16492;
w16494 <= not w15841 and w16126;
w16495 <= not w16122 and w16494;
w16496 <= not w16123 and not w16126;
w16497 <= not w16495 and not w16496;
w16498 <= not w16266 and not w16497;
w16499 <= not w15831 and not w16265;
w16500 <= not w16264 and w16499;
w16501 <= not w16498 and not w16500;
w16502 <= not b(23) and not w16501;
w16503 <= not w15850 and w16121;
w16504 <= not w16117 and w16503;
w16505 <= not w16118 and not w16121;
w16506 <= not w16504 and not w16505;
w16507 <= not w16266 and not w16506;
w16508 <= not w15840 and not w16265;
w16509 <= not w16264 and w16508;
w16510 <= not w16507 and not w16509;
w16511 <= not b(22) and not w16510;
w16512 <= not w15859 and w16116;
w16513 <= not w16112 and w16512;
w16514 <= not w16113 and not w16116;
w16515 <= not w16513 and not w16514;
w16516 <= not w16266 and not w16515;
w16517 <= not w15849 and not w16265;
w16518 <= not w16264 and w16517;
w16519 <= not w16516 and not w16518;
w16520 <= not b(21) and not w16519;
w16521 <= not w15868 and w16111;
w16522 <= not w16107 and w16521;
w16523 <= not w16108 and not w16111;
w16524 <= not w16522 and not w16523;
w16525 <= not w16266 and not w16524;
w16526 <= not w15858 and not w16265;
w16527 <= not w16264 and w16526;
w16528 <= not w16525 and not w16527;
w16529 <= not b(20) and not w16528;
w16530 <= not w15877 and w16106;
w16531 <= not w16102 and w16530;
w16532 <= not w16103 and not w16106;
w16533 <= not w16531 and not w16532;
w16534 <= not w16266 and not w16533;
w16535 <= not w15867 and not w16265;
w16536 <= not w16264 and w16535;
w16537 <= not w16534 and not w16536;
w16538 <= not b(19) and not w16537;
w16539 <= not w15886 and w16101;
w16540 <= not w16097 and w16539;
w16541 <= not w16098 and not w16101;
w16542 <= not w16540 and not w16541;
w16543 <= not w16266 and not w16542;
w16544 <= not w15876 and not w16265;
w16545 <= not w16264 and w16544;
w16546 <= not w16543 and not w16545;
w16547 <= not b(18) and not w16546;
w16548 <= not w15895 and w16096;
w16549 <= not w16092 and w16548;
w16550 <= not w16093 and not w16096;
w16551 <= not w16549 and not w16550;
w16552 <= not w16266 and not w16551;
w16553 <= not w15885 and not w16265;
w16554 <= not w16264 and w16553;
w16555 <= not w16552 and not w16554;
w16556 <= not b(17) and not w16555;
w16557 <= not w15904 and w16091;
w16558 <= not w16087 and w16557;
w16559 <= not w16088 and not w16091;
w16560 <= not w16558 and not w16559;
w16561 <= not w16266 and not w16560;
w16562 <= not w15894 and not w16265;
w16563 <= not w16264 and w16562;
w16564 <= not w16561 and not w16563;
w16565 <= not b(16) and not w16564;
w16566 <= not w15913 and w16086;
w16567 <= not w16082 and w16566;
w16568 <= not w16083 and not w16086;
w16569 <= not w16567 and not w16568;
w16570 <= not w16266 and not w16569;
w16571 <= not w15903 and not w16265;
w16572 <= not w16264 and w16571;
w16573 <= not w16570 and not w16572;
w16574 <= not b(15) and not w16573;
w16575 <= not w15922 and w16081;
w16576 <= not w16077 and w16575;
w16577 <= not w16078 and not w16081;
w16578 <= not w16576 and not w16577;
w16579 <= not w16266 and not w16578;
w16580 <= not w15912 and not w16265;
w16581 <= not w16264 and w16580;
w16582 <= not w16579 and not w16581;
w16583 <= not b(14) and not w16582;
w16584 <= not w15931 and w16076;
w16585 <= not w16072 and w16584;
w16586 <= not w16073 and not w16076;
w16587 <= not w16585 and not w16586;
w16588 <= not w16266 and not w16587;
w16589 <= not w15921 and not w16265;
w16590 <= not w16264 and w16589;
w16591 <= not w16588 and not w16590;
w16592 <= not b(13) and not w16591;
w16593 <= not w15940 and w16071;
w16594 <= not w16067 and w16593;
w16595 <= not w16068 and not w16071;
w16596 <= not w16594 and not w16595;
w16597 <= not w16266 and not w16596;
w16598 <= not w15930 and not w16265;
w16599 <= not w16264 and w16598;
w16600 <= not w16597 and not w16599;
w16601 <= not b(12) and not w16600;
w16602 <= not w15949 and w16066;
w16603 <= not w16062 and w16602;
w16604 <= not w16063 and not w16066;
w16605 <= not w16603 and not w16604;
w16606 <= not w16266 and not w16605;
w16607 <= not w15939 and not w16265;
w16608 <= not w16264 and w16607;
w16609 <= not w16606 and not w16608;
w16610 <= not b(11) and not w16609;
w16611 <= not w15958 and w16061;
w16612 <= not w16057 and w16611;
w16613 <= not w16058 and not w16061;
w16614 <= not w16612 and not w16613;
w16615 <= not w16266 and not w16614;
w16616 <= not w15948 and not w16265;
w16617 <= not w16264 and w16616;
w16618 <= not w16615 and not w16617;
w16619 <= not b(10) and not w16618;
w16620 <= not w15967 and w16056;
w16621 <= not w16052 and w16620;
w16622 <= not w16053 and not w16056;
w16623 <= not w16621 and not w16622;
w16624 <= not w16266 and not w16623;
w16625 <= not w15957 and not w16265;
w16626 <= not w16264 and w16625;
w16627 <= not w16624 and not w16626;
w16628 <= not b(9) and not w16627;
w16629 <= not w15976 and w16051;
w16630 <= not w16047 and w16629;
w16631 <= not w16048 and not w16051;
w16632 <= not w16630 and not w16631;
w16633 <= not w16266 and not w16632;
w16634 <= not w15966 and not w16265;
w16635 <= not w16264 and w16634;
w16636 <= not w16633 and not w16635;
w16637 <= not b(8) and not w16636;
w16638 <= not w15985 and w16046;
w16639 <= not w16042 and w16638;
w16640 <= not w16043 and not w16046;
w16641 <= not w16639 and not w16640;
w16642 <= not w16266 and not w16641;
w16643 <= not w15975 and not w16265;
w16644 <= not w16264 and w16643;
w16645 <= not w16642 and not w16644;
w16646 <= not b(7) and not w16645;
w16647 <= not w15994 and w16041;
w16648 <= not w16037 and w16647;
w16649 <= not w16038 and not w16041;
w16650 <= not w16648 and not w16649;
w16651 <= not w16266 and not w16650;
w16652 <= not w15984 and not w16265;
w16653 <= not w16264 and w16652;
w16654 <= not w16651 and not w16653;
w16655 <= not b(6) and not w16654;
w16656 <= not w16003 and w16036;
w16657 <= not w16032 and w16656;
w16658 <= not w16033 and not w16036;
w16659 <= not w16657 and not w16658;
w16660 <= not w16266 and not w16659;
w16661 <= not w15993 and not w16265;
w16662 <= not w16264 and w16661;
w16663 <= not w16660 and not w16662;
w16664 <= not b(5) and not w16663;
w16665 <= not w16011 and w16031;
w16666 <= not w16027 and w16665;
w16667 <= not w16028 and not w16031;
w16668 <= not w16666 and not w16667;
w16669 <= not w16266 and not w16668;
w16670 <= not w16002 and not w16265;
w16671 <= not w16264 and w16670;
w16672 <= not w16669 and not w16671;
w16673 <= not b(4) and not w16672;
w16674 <= not w16022 and w16026;
w16675 <= not w16021 and w16674;
w16676 <= not w16023 and not w16026;
w16677 <= not w16675 and not w16676;
w16678 <= not w16266 and not w16677;
w16679 <= not w16010 and not w16265;
w16680 <= not w16264 and w16679;
w16681 <= not w16678 and not w16680;
w16682 <= not b(3) and not w16681;
w16683 <= not w16018 and w16020;
w16684 <= not w16016 and w16683;
w16685 <= not w16021 and not w16684;
w16686 <= not w16266 and w16685;
w16687 <= not w16015 and not w16265;
w16688 <= not w16264 and w16687;
w16689 <= not w16686 and not w16688;
w16690 <= not b(2) and not w16689;
w16691 <= b(0) and not w16266;
w16692 <= a(16) and not w16691;
w16693 <= w16020 and not w16266;
w16694 <= not w16692 and not w16693;
w16695 <= b(1) and not w16694;
w16696 <= not b(1) and not w16693;
w16697 <= not w16692 and w16696;
w16698 <= not w16695 and not w16697;
w16699 <= not a(15) and b(0);
w16700 <= not w16698 and not w16699;
w16701 <= not b(1) and not w16694;
w16702 <= not w16700 and not w16701;
w16703 <= b(2) and not w16688;
w16704 <= not w16686 and w16703;
w16705 <= not w16690 and not w16704;
w16706 <= not w16702 and w16705;
w16707 <= not w16690 and not w16706;
w16708 <= b(3) and not w16680;
w16709 <= not w16678 and w16708;
w16710 <= not w16682 and not w16709;
w16711 <= not w16707 and w16710;
w16712 <= not w16682 and not w16711;
w16713 <= b(4) and not w16671;
w16714 <= not w16669 and w16713;
w16715 <= not w16673 and not w16714;
w16716 <= not w16712 and w16715;
w16717 <= not w16673 and not w16716;
w16718 <= b(5) and not w16662;
w16719 <= not w16660 and w16718;
w16720 <= not w16664 and not w16719;
w16721 <= not w16717 and w16720;
w16722 <= not w16664 and not w16721;
w16723 <= b(6) and not w16653;
w16724 <= not w16651 and w16723;
w16725 <= not w16655 and not w16724;
w16726 <= not w16722 and w16725;
w16727 <= not w16655 and not w16726;
w16728 <= b(7) and not w16644;
w16729 <= not w16642 and w16728;
w16730 <= not w16646 and not w16729;
w16731 <= not w16727 and w16730;
w16732 <= not w16646 and not w16731;
w16733 <= b(8) and not w16635;
w16734 <= not w16633 and w16733;
w16735 <= not w16637 and not w16734;
w16736 <= not w16732 and w16735;
w16737 <= not w16637 and not w16736;
w16738 <= b(9) and not w16626;
w16739 <= not w16624 and w16738;
w16740 <= not w16628 and not w16739;
w16741 <= not w16737 and w16740;
w16742 <= not w16628 and not w16741;
w16743 <= b(10) and not w16617;
w16744 <= not w16615 and w16743;
w16745 <= not w16619 and not w16744;
w16746 <= not w16742 and w16745;
w16747 <= not w16619 and not w16746;
w16748 <= b(11) and not w16608;
w16749 <= not w16606 and w16748;
w16750 <= not w16610 and not w16749;
w16751 <= not w16747 and w16750;
w16752 <= not w16610 and not w16751;
w16753 <= b(12) and not w16599;
w16754 <= not w16597 and w16753;
w16755 <= not w16601 and not w16754;
w16756 <= not w16752 and w16755;
w16757 <= not w16601 and not w16756;
w16758 <= b(13) and not w16590;
w16759 <= not w16588 and w16758;
w16760 <= not w16592 and not w16759;
w16761 <= not w16757 and w16760;
w16762 <= not w16592 and not w16761;
w16763 <= b(14) and not w16581;
w16764 <= not w16579 and w16763;
w16765 <= not w16583 and not w16764;
w16766 <= not w16762 and w16765;
w16767 <= not w16583 and not w16766;
w16768 <= b(15) and not w16572;
w16769 <= not w16570 and w16768;
w16770 <= not w16574 and not w16769;
w16771 <= not w16767 and w16770;
w16772 <= not w16574 and not w16771;
w16773 <= b(16) and not w16563;
w16774 <= not w16561 and w16773;
w16775 <= not w16565 and not w16774;
w16776 <= not w16772 and w16775;
w16777 <= not w16565 and not w16776;
w16778 <= b(17) and not w16554;
w16779 <= not w16552 and w16778;
w16780 <= not w16556 and not w16779;
w16781 <= not w16777 and w16780;
w16782 <= not w16556 and not w16781;
w16783 <= b(18) and not w16545;
w16784 <= not w16543 and w16783;
w16785 <= not w16547 and not w16784;
w16786 <= not w16782 and w16785;
w16787 <= not w16547 and not w16786;
w16788 <= b(19) and not w16536;
w16789 <= not w16534 and w16788;
w16790 <= not w16538 and not w16789;
w16791 <= not w16787 and w16790;
w16792 <= not w16538 and not w16791;
w16793 <= b(20) and not w16527;
w16794 <= not w16525 and w16793;
w16795 <= not w16529 and not w16794;
w16796 <= not w16792 and w16795;
w16797 <= not w16529 and not w16796;
w16798 <= b(21) and not w16518;
w16799 <= not w16516 and w16798;
w16800 <= not w16520 and not w16799;
w16801 <= not w16797 and w16800;
w16802 <= not w16520 and not w16801;
w16803 <= b(22) and not w16509;
w16804 <= not w16507 and w16803;
w16805 <= not w16511 and not w16804;
w16806 <= not w16802 and w16805;
w16807 <= not w16511 and not w16806;
w16808 <= b(23) and not w16500;
w16809 <= not w16498 and w16808;
w16810 <= not w16502 and not w16809;
w16811 <= not w16807 and w16810;
w16812 <= not w16502 and not w16811;
w16813 <= b(24) and not w16491;
w16814 <= not w16489 and w16813;
w16815 <= not w16493 and not w16814;
w16816 <= not w16812 and w16815;
w16817 <= not w16493 and not w16816;
w16818 <= b(25) and not w16482;
w16819 <= not w16480 and w16818;
w16820 <= not w16484 and not w16819;
w16821 <= not w16817 and w16820;
w16822 <= not w16484 and not w16821;
w16823 <= b(26) and not w16473;
w16824 <= not w16471 and w16823;
w16825 <= not w16475 and not w16824;
w16826 <= not w16822 and w16825;
w16827 <= not w16475 and not w16826;
w16828 <= b(27) and not w16464;
w16829 <= not w16462 and w16828;
w16830 <= not w16466 and not w16829;
w16831 <= not w16827 and w16830;
w16832 <= not w16466 and not w16831;
w16833 <= b(28) and not w16455;
w16834 <= not w16453 and w16833;
w16835 <= not w16457 and not w16834;
w16836 <= not w16832 and w16835;
w16837 <= not w16457 and not w16836;
w16838 <= b(29) and not w16446;
w16839 <= not w16444 and w16838;
w16840 <= not w16448 and not w16839;
w16841 <= not w16837 and w16840;
w16842 <= not w16448 and not w16841;
w16843 <= b(30) and not w16437;
w16844 <= not w16435 and w16843;
w16845 <= not w16439 and not w16844;
w16846 <= not w16842 and w16845;
w16847 <= not w16439 and not w16846;
w16848 <= b(31) and not w16428;
w16849 <= not w16426 and w16848;
w16850 <= not w16430 and not w16849;
w16851 <= not w16847 and w16850;
w16852 <= not w16430 and not w16851;
w16853 <= b(32) and not w16419;
w16854 <= not w16417 and w16853;
w16855 <= not w16421 and not w16854;
w16856 <= not w16852 and w16855;
w16857 <= not w16421 and not w16856;
w16858 <= b(33) and not w16410;
w16859 <= not w16408 and w16858;
w16860 <= not w16412 and not w16859;
w16861 <= not w16857 and w16860;
w16862 <= not w16412 and not w16861;
w16863 <= b(34) and not w16401;
w16864 <= not w16399 and w16863;
w16865 <= not w16403 and not w16864;
w16866 <= not w16862 and w16865;
w16867 <= not w16403 and not w16866;
w16868 <= b(35) and not w16392;
w16869 <= not w16390 and w16868;
w16870 <= not w16394 and not w16869;
w16871 <= not w16867 and w16870;
w16872 <= not w16394 and not w16871;
w16873 <= b(36) and not w16383;
w16874 <= not w16381 and w16873;
w16875 <= not w16385 and not w16874;
w16876 <= not w16872 and w16875;
w16877 <= not w16385 and not w16876;
w16878 <= b(37) and not w16374;
w16879 <= not w16372 and w16878;
w16880 <= not w16376 and not w16879;
w16881 <= not w16877 and w16880;
w16882 <= not w16376 and not w16881;
w16883 <= b(38) and not w16365;
w16884 <= not w16363 and w16883;
w16885 <= not w16367 and not w16884;
w16886 <= not w16882 and w16885;
w16887 <= not w16367 and not w16886;
w16888 <= b(39) and not w16356;
w16889 <= not w16354 and w16888;
w16890 <= not w16358 and not w16889;
w16891 <= not w16887 and w16890;
w16892 <= not w16358 and not w16891;
w16893 <= b(40) and not w16347;
w16894 <= not w16345 and w16893;
w16895 <= not w16349 and not w16894;
w16896 <= not w16892 and w16895;
w16897 <= not w16349 and not w16896;
w16898 <= b(41) and not w16338;
w16899 <= not w16336 and w16898;
w16900 <= not w16340 and not w16899;
w16901 <= not w16897 and w16900;
w16902 <= not w16340 and not w16901;
w16903 <= b(42) and not w16329;
w16904 <= not w16327 and w16903;
w16905 <= not w16331 and not w16904;
w16906 <= not w16902 and w16905;
w16907 <= not w16331 and not w16906;
w16908 <= b(43) and not w16320;
w16909 <= not w16318 and w16908;
w16910 <= not w16322 and not w16909;
w16911 <= not w16907 and w16910;
w16912 <= not w16322 and not w16911;
w16913 <= b(44) and not w16311;
w16914 <= not w16309 and w16913;
w16915 <= not w16313 and not w16914;
w16916 <= not w16912 and w16915;
w16917 <= not w16313 and not w16916;
w16918 <= b(45) and not w16302;
w16919 <= not w16300 and w16918;
w16920 <= not w16304 and not w16919;
w16921 <= not w16917 and w16920;
w16922 <= not w16304 and not w16921;
w16923 <= b(46) and not w16293;
w16924 <= not w16291 and w16923;
w16925 <= not w16295 and not w16924;
w16926 <= not w16922 and w16925;
w16927 <= not w16295 and not w16926;
w16928 <= b(47) and not w16273;
w16929 <= not w16271 and w16928;
w16930 <= not w16286 and not w16929;
w16931 <= not w16927 and w16930;
w16932 <= not w16286 and not w16931;
w16933 <= b(48) and not w16283;
w16934 <= not w16281 and w16933;
w16935 <= not w16285 and not w16934;
w16936 <= not w16932 and w16935;
w16937 <= not w16285 and not w16936;
w16938 <= w151 and not w16937;
w16939 <= not w16274 and not w16938;
w16940 <= not w16295 and w16930;
w16941 <= not w16926 and w16940;
w16942 <= not w16927 and not w16930;
w16943 <= not w16941 and not w16942;
w16944 <= w151 and not w16943;
w16945 <= not w16937 and w16944;
w16946 <= not w16939 and not w16945;
w16947 <= not b(48) and not w16946;
w16948 <= not w16294 and not w16938;
w16949 <= not w16304 and w16925;
w16950 <= not w16921 and w16949;
w16951 <= not w16922 and not w16925;
w16952 <= not w16950 and not w16951;
w16953 <= w151 and not w16952;
w16954 <= not w16937 and w16953;
w16955 <= not w16948 and not w16954;
w16956 <= not b(47) and not w16955;
w16957 <= not w16303 and not w16938;
w16958 <= not w16313 and w16920;
w16959 <= not w16916 and w16958;
w16960 <= not w16917 and not w16920;
w16961 <= not w16959 and not w16960;
w16962 <= w151 and not w16961;
w16963 <= not w16937 and w16962;
w16964 <= not w16957 and not w16963;
w16965 <= not b(46) and not w16964;
w16966 <= not w16312 and not w16938;
w16967 <= not w16322 and w16915;
w16968 <= not w16911 and w16967;
w16969 <= not w16912 and not w16915;
w16970 <= not w16968 and not w16969;
w16971 <= w151 and not w16970;
w16972 <= not w16937 and w16971;
w16973 <= not w16966 and not w16972;
w16974 <= not b(45) and not w16973;
w16975 <= not w16321 and not w16938;
w16976 <= not w16331 and w16910;
w16977 <= not w16906 and w16976;
w16978 <= not w16907 and not w16910;
w16979 <= not w16977 and not w16978;
w16980 <= w151 and not w16979;
w16981 <= not w16937 and w16980;
w16982 <= not w16975 and not w16981;
w16983 <= not b(44) and not w16982;
w16984 <= not w16330 and not w16938;
w16985 <= not w16340 and w16905;
w16986 <= not w16901 and w16985;
w16987 <= not w16902 and not w16905;
w16988 <= not w16986 and not w16987;
w16989 <= w151 and not w16988;
w16990 <= not w16937 and w16989;
w16991 <= not w16984 and not w16990;
w16992 <= not b(43) and not w16991;
w16993 <= not w16339 and not w16938;
w16994 <= not w16349 and w16900;
w16995 <= not w16896 and w16994;
w16996 <= not w16897 and not w16900;
w16997 <= not w16995 and not w16996;
w16998 <= w151 and not w16997;
w16999 <= not w16937 and w16998;
w17000 <= not w16993 and not w16999;
w17001 <= not b(42) and not w17000;
w17002 <= not w16348 and not w16938;
w17003 <= not w16358 and w16895;
w17004 <= not w16891 and w17003;
w17005 <= not w16892 and not w16895;
w17006 <= not w17004 and not w17005;
w17007 <= w151 and not w17006;
w17008 <= not w16937 and w17007;
w17009 <= not w17002 and not w17008;
w17010 <= not b(41) and not w17009;
w17011 <= not w16357 and not w16938;
w17012 <= not w16367 and w16890;
w17013 <= not w16886 and w17012;
w17014 <= not w16887 and not w16890;
w17015 <= not w17013 and not w17014;
w17016 <= w151 and not w17015;
w17017 <= not w16937 and w17016;
w17018 <= not w17011 and not w17017;
w17019 <= not b(40) and not w17018;
w17020 <= not w16366 and not w16938;
w17021 <= not w16376 and w16885;
w17022 <= not w16881 and w17021;
w17023 <= not w16882 and not w16885;
w17024 <= not w17022 and not w17023;
w17025 <= w151 and not w17024;
w17026 <= not w16937 and w17025;
w17027 <= not w17020 and not w17026;
w17028 <= not b(39) and not w17027;
w17029 <= not w16375 and not w16938;
w17030 <= not w16385 and w16880;
w17031 <= not w16876 and w17030;
w17032 <= not w16877 and not w16880;
w17033 <= not w17031 and not w17032;
w17034 <= w151 and not w17033;
w17035 <= not w16937 and w17034;
w17036 <= not w17029 and not w17035;
w17037 <= not b(38) and not w17036;
w17038 <= not w16384 and not w16938;
w17039 <= not w16394 and w16875;
w17040 <= not w16871 and w17039;
w17041 <= not w16872 and not w16875;
w17042 <= not w17040 and not w17041;
w17043 <= w151 and not w17042;
w17044 <= not w16937 and w17043;
w17045 <= not w17038 and not w17044;
w17046 <= not b(37) and not w17045;
w17047 <= not w16393 and not w16938;
w17048 <= not w16403 and w16870;
w17049 <= not w16866 and w17048;
w17050 <= not w16867 and not w16870;
w17051 <= not w17049 and not w17050;
w17052 <= w151 and not w17051;
w17053 <= not w16937 and w17052;
w17054 <= not w17047 and not w17053;
w17055 <= not b(36) and not w17054;
w17056 <= not w16402 and not w16938;
w17057 <= not w16412 and w16865;
w17058 <= not w16861 and w17057;
w17059 <= not w16862 and not w16865;
w17060 <= not w17058 and not w17059;
w17061 <= w151 and not w17060;
w17062 <= not w16937 and w17061;
w17063 <= not w17056 and not w17062;
w17064 <= not b(35) and not w17063;
w17065 <= not w16411 and not w16938;
w17066 <= not w16421 and w16860;
w17067 <= not w16856 and w17066;
w17068 <= not w16857 and not w16860;
w17069 <= not w17067 and not w17068;
w17070 <= w151 and not w17069;
w17071 <= not w16937 and w17070;
w17072 <= not w17065 and not w17071;
w17073 <= not b(34) and not w17072;
w17074 <= not w16420 and not w16938;
w17075 <= not w16430 and w16855;
w17076 <= not w16851 and w17075;
w17077 <= not w16852 and not w16855;
w17078 <= not w17076 and not w17077;
w17079 <= w151 and not w17078;
w17080 <= not w16937 and w17079;
w17081 <= not w17074 and not w17080;
w17082 <= not b(33) and not w17081;
w17083 <= not w16429 and not w16938;
w17084 <= not w16439 and w16850;
w17085 <= not w16846 and w17084;
w17086 <= not w16847 and not w16850;
w17087 <= not w17085 and not w17086;
w17088 <= w151 and not w17087;
w17089 <= not w16937 and w17088;
w17090 <= not w17083 and not w17089;
w17091 <= not b(32) and not w17090;
w17092 <= not w16438 and not w16938;
w17093 <= not w16448 and w16845;
w17094 <= not w16841 and w17093;
w17095 <= not w16842 and not w16845;
w17096 <= not w17094 and not w17095;
w17097 <= w151 and not w17096;
w17098 <= not w16937 and w17097;
w17099 <= not w17092 and not w17098;
w17100 <= not b(31) and not w17099;
w17101 <= not w16447 and not w16938;
w17102 <= not w16457 and w16840;
w17103 <= not w16836 and w17102;
w17104 <= not w16837 and not w16840;
w17105 <= not w17103 and not w17104;
w17106 <= w151 and not w17105;
w17107 <= not w16937 and w17106;
w17108 <= not w17101 and not w17107;
w17109 <= not b(30) and not w17108;
w17110 <= not w16456 and not w16938;
w17111 <= not w16466 and w16835;
w17112 <= not w16831 and w17111;
w17113 <= not w16832 and not w16835;
w17114 <= not w17112 and not w17113;
w17115 <= w151 and not w17114;
w17116 <= not w16937 and w17115;
w17117 <= not w17110 and not w17116;
w17118 <= not b(29) and not w17117;
w17119 <= not w16465 and not w16938;
w17120 <= not w16475 and w16830;
w17121 <= not w16826 and w17120;
w17122 <= not w16827 and not w16830;
w17123 <= not w17121 and not w17122;
w17124 <= w151 and not w17123;
w17125 <= not w16937 and w17124;
w17126 <= not w17119 and not w17125;
w17127 <= not b(28) and not w17126;
w17128 <= not w16474 and not w16938;
w17129 <= not w16484 and w16825;
w17130 <= not w16821 and w17129;
w17131 <= not w16822 and not w16825;
w17132 <= not w17130 and not w17131;
w17133 <= w151 and not w17132;
w17134 <= not w16937 and w17133;
w17135 <= not w17128 and not w17134;
w17136 <= not b(27) and not w17135;
w17137 <= not w16483 and not w16938;
w17138 <= not w16493 and w16820;
w17139 <= not w16816 and w17138;
w17140 <= not w16817 and not w16820;
w17141 <= not w17139 and not w17140;
w17142 <= w151 and not w17141;
w17143 <= not w16937 and w17142;
w17144 <= not w17137 and not w17143;
w17145 <= not b(26) and not w17144;
w17146 <= not w16492 and not w16938;
w17147 <= not w16502 and w16815;
w17148 <= not w16811 and w17147;
w17149 <= not w16812 and not w16815;
w17150 <= not w17148 and not w17149;
w17151 <= w151 and not w17150;
w17152 <= not w16937 and w17151;
w17153 <= not w17146 and not w17152;
w17154 <= not b(25) and not w17153;
w17155 <= not w16501 and not w16938;
w17156 <= not w16511 and w16810;
w17157 <= not w16806 and w17156;
w17158 <= not w16807 and not w16810;
w17159 <= not w17157 and not w17158;
w17160 <= w151 and not w17159;
w17161 <= not w16937 and w17160;
w17162 <= not w17155 and not w17161;
w17163 <= not b(24) and not w17162;
w17164 <= not w16510 and not w16938;
w17165 <= not w16520 and w16805;
w17166 <= not w16801 and w17165;
w17167 <= not w16802 and not w16805;
w17168 <= not w17166 and not w17167;
w17169 <= w151 and not w17168;
w17170 <= not w16937 and w17169;
w17171 <= not w17164 and not w17170;
w17172 <= not b(23) and not w17171;
w17173 <= not w16519 and not w16938;
w17174 <= not w16529 and w16800;
w17175 <= not w16796 and w17174;
w17176 <= not w16797 and not w16800;
w17177 <= not w17175 and not w17176;
w17178 <= w151 and not w17177;
w17179 <= not w16937 and w17178;
w17180 <= not w17173 and not w17179;
w17181 <= not b(22) and not w17180;
w17182 <= not w16528 and not w16938;
w17183 <= not w16538 and w16795;
w17184 <= not w16791 and w17183;
w17185 <= not w16792 and not w16795;
w17186 <= not w17184 and not w17185;
w17187 <= w151 and not w17186;
w17188 <= not w16937 and w17187;
w17189 <= not w17182 and not w17188;
w17190 <= not b(21) and not w17189;
w17191 <= not w16537 and not w16938;
w17192 <= not w16547 and w16790;
w17193 <= not w16786 and w17192;
w17194 <= not w16787 and not w16790;
w17195 <= not w17193 and not w17194;
w17196 <= w151 and not w17195;
w17197 <= not w16937 and w17196;
w17198 <= not w17191 and not w17197;
w17199 <= not b(20) and not w17198;
w17200 <= not w16546 and not w16938;
w17201 <= not w16556 and w16785;
w17202 <= not w16781 and w17201;
w17203 <= not w16782 and not w16785;
w17204 <= not w17202 and not w17203;
w17205 <= w151 and not w17204;
w17206 <= not w16937 and w17205;
w17207 <= not w17200 and not w17206;
w17208 <= not b(19) and not w17207;
w17209 <= not w16555 and not w16938;
w17210 <= not w16565 and w16780;
w17211 <= not w16776 and w17210;
w17212 <= not w16777 and not w16780;
w17213 <= not w17211 and not w17212;
w17214 <= w151 and not w17213;
w17215 <= not w16937 and w17214;
w17216 <= not w17209 and not w17215;
w17217 <= not b(18) and not w17216;
w17218 <= not w16564 and not w16938;
w17219 <= not w16574 and w16775;
w17220 <= not w16771 and w17219;
w17221 <= not w16772 and not w16775;
w17222 <= not w17220 and not w17221;
w17223 <= w151 and not w17222;
w17224 <= not w16937 and w17223;
w17225 <= not w17218 and not w17224;
w17226 <= not b(17) and not w17225;
w17227 <= not w16573 and not w16938;
w17228 <= not w16583 and w16770;
w17229 <= not w16766 and w17228;
w17230 <= not w16767 and not w16770;
w17231 <= not w17229 and not w17230;
w17232 <= w151 and not w17231;
w17233 <= not w16937 and w17232;
w17234 <= not w17227 and not w17233;
w17235 <= not b(16) and not w17234;
w17236 <= not w16582 and not w16938;
w17237 <= not w16592 and w16765;
w17238 <= not w16761 and w17237;
w17239 <= not w16762 and not w16765;
w17240 <= not w17238 and not w17239;
w17241 <= w151 and not w17240;
w17242 <= not w16937 and w17241;
w17243 <= not w17236 and not w17242;
w17244 <= not b(15) and not w17243;
w17245 <= not w16591 and not w16938;
w17246 <= not w16601 and w16760;
w17247 <= not w16756 and w17246;
w17248 <= not w16757 and not w16760;
w17249 <= not w17247 and not w17248;
w17250 <= w151 and not w17249;
w17251 <= not w16937 and w17250;
w17252 <= not w17245 and not w17251;
w17253 <= not b(14) and not w17252;
w17254 <= not w16600 and not w16938;
w17255 <= not w16610 and w16755;
w17256 <= not w16751 and w17255;
w17257 <= not w16752 and not w16755;
w17258 <= not w17256 and not w17257;
w17259 <= w151 and not w17258;
w17260 <= not w16937 and w17259;
w17261 <= not w17254 and not w17260;
w17262 <= not b(13) and not w17261;
w17263 <= not w16609 and not w16938;
w17264 <= not w16619 and w16750;
w17265 <= not w16746 and w17264;
w17266 <= not w16747 and not w16750;
w17267 <= not w17265 and not w17266;
w17268 <= w151 and not w17267;
w17269 <= not w16937 and w17268;
w17270 <= not w17263 and not w17269;
w17271 <= not b(12) and not w17270;
w17272 <= not w16618 and not w16938;
w17273 <= not w16628 and w16745;
w17274 <= not w16741 and w17273;
w17275 <= not w16742 and not w16745;
w17276 <= not w17274 and not w17275;
w17277 <= w151 and not w17276;
w17278 <= not w16937 and w17277;
w17279 <= not w17272 and not w17278;
w17280 <= not b(11) and not w17279;
w17281 <= not w16627 and not w16938;
w17282 <= not w16637 and w16740;
w17283 <= not w16736 and w17282;
w17284 <= not w16737 and not w16740;
w17285 <= not w17283 and not w17284;
w17286 <= w151 and not w17285;
w17287 <= not w16937 and w17286;
w17288 <= not w17281 and not w17287;
w17289 <= not b(10) and not w17288;
w17290 <= not w16636 and not w16938;
w17291 <= not w16646 and w16735;
w17292 <= not w16731 and w17291;
w17293 <= not w16732 and not w16735;
w17294 <= not w17292 and not w17293;
w17295 <= w151 and not w17294;
w17296 <= not w16937 and w17295;
w17297 <= not w17290 and not w17296;
w17298 <= not b(9) and not w17297;
w17299 <= not w16645 and not w16938;
w17300 <= not w16655 and w16730;
w17301 <= not w16726 and w17300;
w17302 <= not w16727 and not w16730;
w17303 <= not w17301 and not w17302;
w17304 <= w151 and not w17303;
w17305 <= not w16937 and w17304;
w17306 <= not w17299 and not w17305;
w17307 <= not b(8) and not w17306;
w17308 <= not w16654 and not w16938;
w17309 <= not w16664 and w16725;
w17310 <= not w16721 and w17309;
w17311 <= not w16722 and not w16725;
w17312 <= not w17310 and not w17311;
w17313 <= w151 and not w17312;
w17314 <= not w16937 and w17313;
w17315 <= not w17308 and not w17314;
w17316 <= not b(7) and not w17315;
w17317 <= not w16663 and not w16938;
w17318 <= not w16673 and w16720;
w17319 <= not w16716 and w17318;
w17320 <= not w16717 and not w16720;
w17321 <= not w17319 and not w17320;
w17322 <= w151 and not w17321;
w17323 <= not w16937 and w17322;
w17324 <= not w17317 and not w17323;
w17325 <= not b(6) and not w17324;
w17326 <= not w16672 and not w16938;
w17327 <= not w16682 and w16715;
w17328 <= not w16711 and w17327;
w17329 <= not w16712 and not w16715;
w17330 <= not w17328 and not w17329;
w17331 <= w151 and not w17330;
w17332 <= not w16937 and w17331;
w17333 <= not w17326 and not w17332;
w17334 <= not b(5) and not w17333;
w17335 <= not w16681 and not w16938;
w17336 <= not w16690 and w16710;
w17337 <= not w16706 and w17336;
w17338 <= not w16707 and not w16710;
w17339 <= not w17337 and not w17338;
w17340 <= w151 and not w17339;
w17341 <= not w16937 and w17340;
w17342 <= not w17335 and not w17341;
w17343 <= not b(4) and not w17342;
w17344 <= not w16689 and not w16938;
w17345 <= not w16701 and w16705;
w17346 <= not w16700 and w17345;
w17347 <= not w16702 and not w16705;
w17348 <= not w17346 and not w17347;
w17349 <= w151 and not w17348;
w17350 <= not w16937 and w17349;
w17351 <= not w17344 and not w17350;
w17352 <= not b(3) and not w17351;
w17353 <= not w16694 and not w16938;
w17354 <= not w16697 and w16699;
w17355 <= not w16695 and w17354;
w17356 <= w151 and not w17355;
w17357 <= not w16700 and w17356;
w17358 <= not w16937 and w17357;
w17359 <= not w17353 and not w17358;
w17360 <= not b(2) and not w17359;
w17361 <= b(0) and not b(49);
w17362 <= w40 and w17361;
w17363 <= w29 and w17362;
w17364 <= w80 and w17363;
w17365 <= not w16937 and w17364;
w17366 <= a(15) and not w17365;
w17367 <= w143 and w16699;
w17368 <= w338 and w17367;
w17369 <= not w16937 and w17368;
w17370 <= not w17366 and not w17369;
w17371 <= b(1) and not w17370;
w17372 <= not b(1) and not w17369;
w17373 <= not w17366 and w17372;
w17374 <= not w17371 and not w17373;
w17375 <= not a(14) and b(0);
w17376 <= not w17374 and not w17375;
w17377 <= not b(1) and not w17370;
w17378 <= not w17376 and not w17377;
w17379 <= b(2) and not w17358;
w17380 <= not w17353 and w17379;
w17381 <= not w17360 and not w17380;
w17382 <= not w17378 and w17381;
w17383 <= not w17360 and not w17382;
w17384 <= b(3) and not w17350;
w17385 <= not w17344 and w17384;
w17386 <= not w17352 and not w17385;
w17387 <= not w17383 and w17386;
w17388 <= not w17352 and not w17387;
w17389 <= b(4) and not w17341;
w17390 <= not w17335 and w17389;
w17391 <= not w17343 and not w17390;
w17392 <= not w17388 and w17391;
w17393 <= not w17343 and not w17392;
w17394 <= b(5) and not w17332;
w17395 <= not w17326 and w17394;
w17396 <= not w17334 and not w17395;
w17397 <= not w17393 and w17396;
w17398 <= not w17334 and not w17397;
w17399 <= b(6) and not w17323;
w17400 <= not w17317 and w17399;
w17401 <= not w17325 and not w17400;
w17402 <= not w17398 and w17401;
w17403 <= not w17325 and not w17402;
w17404 <= b(7) and not w17314;
w17405 <= not w17308 and w17404;
w17406 <= not w17316 and not w17405;
w17407 <= not w17403 and w17406;
w17408 <= not w17316 and not w17407;
w17409 <= b(8) and not w17305;
w17410 <= not w17299 and w17409;
w17411 <= not w17307 and not w17410;
w17412 <= not w17408 and w17411;
w17413 <= not w17307 and not w17412;
w17414 <= b(9) and not w17296;
w17415 <= not w17290 and w17414;
w17416 <= not w17298 and not w17415;
w17417 <= not w17413 and w17416;
w17418 <= not w17298 and not w17417;
w17419 <= b(10) and not w17287;
w17420 <= not w17281 and w17419;
w17421 <= not w17289 and not w17420;
w17422 <= not w17418 and w17421;
w17423 <= not w17289 and not w17422;
w17424 <= b(11) and not w17278;
w17425 <= not w17272 and w17424;
w17426 <= not w17280 and not w17425;
w17427 <= not w17423 and w17426;
w17428 <= not w17280 and not w17427;
w17429 <= b(12) and not w17269;
w17430 <= not w17263 and w17429;
w17431 <= not w17271 and not w17430;
w17432 <= not w17428 and w17431;
w17433 <= not w17271 and not w17432;
w17434 <= b(13) and not w17260;
w17435 <= not w17254 and w17434;
w17436 <= not w17262 and not w17435;
w17437 <= not w17433 and w17436;
w17438 <= not w17262 and not w17437;
w17439 <= b(14) and not w17251;
w17440 <= not w17245 and w17439;
w17441 <= not w17253 and not w17440;
w17442 <= not w17438 and w17441;
w17443 <= not w17253 and not w17442;
w17444 <= b(15) and not w17242;
w17445 <= not w17236 and w17444;
w17446 <= not w17244 and not w17445;
w17447 <= not w17443 and w17446;
w17448 <= not w17244 and not w17447;
w17449 <= b(16) and not w17233;
w17450 <= not w17227 and w17449;
w17451 <= not w17235 and not w17450;
w17452 <= not w17448 and w17451;
w17453 <= not w17235 and not w17452;
w17454 <= b(17) and not w17224;
w17455 <= not w17218 and w17454;
w17456 <= not w17226 and not w17455;
w17457 <= not w17453 and w17456;
w17458 <= not w17226 and not w17457;
w17459 <= b(18) and not w17215;
w17460 <= not w17209 and w17459;
w17461 <= not w17217 and not w17460;
w17462 <= not w17458 and w17461;
w17463 <= not w17217 and not w17462;
w17464 <= b(19) and not w17206;
w17465 <= not w17200 and w17464;
w17466 <= not w17208 and not w17465;
w17467 <= not w17463 and w17466;
w17468 <= not w17208 and not w17467;
w17469 <= b(20) and not w17197;
w17470 <= not w17191 and w17469;
w17471 <= not w17199 and not w17470;
w17472 <= not w17468 and w17471;
w17473 <= not w17199 and not w17472;
w17474 <= b(21) and not w17188;
w17475 <= not w17182 and w17474;
w17476 <= not w17190 and not w17475;
w17477 <= not w17473 and w17476;
w17478 <= not w17190 and not w17477;
w17479 <= b(22) and not w17179;
w17480 <= not w17173 and w17479;
w17481 <= not w17181 and not w17480;
w17482 <= not w17478 and w17481;
w17483 <= not w17181 and not w17482;
w17484 <= b(23) and not w17170;
w17485 <= not w17164 and w17484;
w17486 <= not w17172 and not w17485;
w17487 <= not w17483 and w17486;
w17488 <= not w17172 and not w17487;
w17489 <= b(24) and not w17161;
w17490 <= not w17155 and w17489;
w17491 <= not w17163 and not w17490;
w17492 <= not w17488 and w17491;
w17493 <= not w17163 and not w17492;
w17494 <= b(25) and not w17152;
w17495 <= not w17146 and w17494;
w17496 <= not w17154 and not w17495;
w17497 <= not w17493 and w17496;
w17498 <= not w17154 and not w17497;
w17499 <= b(26) and not w17143;
w17500 <= not w17137 and w17499;
w17501 <= not w17145 and not w17500;
w17502 <= not w17498 and w17501;
w17503 <= not w17145 and not w17502;
w17504 <= b(27) and not w17134;
w17505 <= not w17128 and w17504;
w17506 <= not w17136 and not w17505;
w17507 <= not w17503 and w17506;
w17508 <= not w17136 and not w17507;
w17509 <= b(28) and not w17125;
w17510 <= not w17119 and w17509;
w17511 <= not w17127 and not w17510;
w17512 <= not w17508 and w17511;
w17513 <= not w17127 and not w17512;
w17514 <= b(29) and not w17116;
w17515 <= not w17110 and w17514;
w17516 <= not w17118 and not w17515;
w17517 <= not w17513 and w17516;
w17518 <= not w17118 and not w17517;
w17519 <= b(30) and not w17107;
w17520 <= not w17101 and w17519;
w17521 <= not w17109 and not w17520;
w17522 <= not w17518 and w17521;
w17523 <= not w17109 and not w17522;
w17524 <= b(31) and not w17098;
w17525 <= not w17092 and w17524;
w17526 <= not w17100 and not w17525;
w17527 <= not w17523 and w17526;
w17528 <= not w17100 and not w17527;
w17529 <= b(32) and not w17089;
w17530 <= not w17083 and w17529;
w17531 <= not w17091 and not w17530;
w17532 <= not w17528 and w17531;
w17533 <= not w17091 and not w17532;
w17534 <= b(33) and not w17080;
w17535 <= not w17074 and w17534;
w17536 <= not w17082 and not w17535;
w17537 <= not w17533 and w17536;
w17538 <= not w17082 and not w17537;
w17539 <= b(34) and not w17071;
w17540 <= not w17065 and w17539;
w17541 <= not w17073 and not w17540;
w17542 <= not w17538 and w17541;
w17543 <= not w17073 and not w17542;
w17544 <= b(35) and not w17062;
w17545 <= not w17056 and w17544;
w17546 <= not w17064 and not w17545;
w17547 <= not w17543 and w17546;
w17548 <= not w17064 and not w17547;
w17549 <= b(36) and not w17053;
w17550 <= not w17047 and w17549;
w17551 <= not w17055 and not w17550;
w17552 <= not w17548 and w17551;
w17553 <= not w17055 and not w17552;
w17554 <= b(37) and not w17044;
w17555 <= not w17038 and w17554;
w17556 <= not w17046 and not w17555;
w17557 <= not w17553 and w17556;
w17558 <= not w17046 and not w17557;
w17559 <= b(38) and not w17035;
w17560 <= not w17029 and w17559;
w17561 <= not w17037 and not w17560;
w17562 <= not w17558 and w17561;
w17563 <= not w17037 and not w17562;
w17564 <= b(39) and not w17026;
w17565 <= not w17020 and w17564;
w17566 <= not w17028 and not w17565;
w17567 <= not w17563 and w17566;
w17568 <= not w17028 and not w17567;
w17569 <= b(40) and not w17017;
w17570 <= not w17011 and w17569;
w17571 <= not w17019 and not w17570;
w17572 <= not w17568 and w17571;
w17573 <= not w17019 and not w17572;
w17574 <= b(41) and not w17008;
w17575 <= not w17002 and w17574;
w17576 <= not w17010 and not w17575;
w17577 <= not w17573 and w17576;
w17578 <= not w17010 and not w17577;
w17579 <= b(42) and not w16999;
w17580 <= not w16993 and w17579;
w17581 <= not w17001 and not w17580;
w17582 <= not w17578 and w17581;
w17583 <= not w17001 and not w17582;
w17584 <= b(43) and not w16990;
w17585 <= not w16984 and w17584;
w17586 <= not w16992 and not w17585;
w17587 <= not w17583 and w17586;
w17588 <= not w16992 and not w17587;
w17589 <= b(44) and not w16981;
w17590 <= not w16975 and w17589;
w17591 <= not w16983 and not w17590;
w17592 <= not w17588 and w17591;
w17593 <= not w16983 and not w17592;
w17594 <= b(45) and not w16972;
w17595 <= not w16966 and w17594;
w17596 <= not w16974 and not w17595;
w17597 <= not w17593 and w17596;
w17598 <= not w16974 and not w17597;
w17599 <= b(46) and not w16963;
w17600 <= not w16957 and w17599;
w17601 <= not w16965 and not w17600;
w17602 <= not w17598 and w17601;
w17603 <= not w16965 and not w17602;
w17604 <= b(47) and not w16954;
w17605 <= not w16948 and w17604;
w17606 <= not w16956 and not w17605;
w17607 <= not w17603 and w17606;
w17608 <= not w16956 and not w17607;
w17609 <= b(48) and not w16945;
w17610 <= not w16939 and w17609;
w17611 <= not w16947 and not w17610;
w17612 <= not w17608 and w17611;
w17613 <= not w16947 and not w17612;
w17614 <= not w16284 and not w16938;
w17615 <= not w16286 and w16935;
w17616 <= not w16931 and w17615;
w17617 <= not w16932 and not w16935;
w17618 <= not w17616 and not w17617;
w17619 <= w16938 and not w17618;
w17620 <= not w17614 and not w17619;
w17621 <= not b(49) and not w17620;
w17622 <= b(49) and not w17614;
w17623 <= not w17619 and w17622;
w17624 <= w29 and w40;
w17625 <= w80 and w17624;
w17626 <= not w17623 and w17625;
w17627 <= not w17621 and w17626;
w17628 <= not w17613 and w17627;
w17629 <= w151 and not w17620;
w17630 <= not w17628 and not w17629;
w17631 <= not w16956 and w17611;
w17632 <= not w17607 and w17631;
w17633 <= not w17608 and not w17611;
w17634 <= not w17632 and not w17633;
w17635 <= not w17630 and not w17634;
w17636 <= not w16946 and not w17629;
w17637 <= not w17628 and w17636;
w17638 <= not w17635 and not w17637;
w17639 <= not b(49) and not w17638;
w17640 <= not w16965 and w17606;
w17641 <= not w17602 and w17640;
w17642 <= not w17603 and not w17606;
w17643 <= not w17641 and not w17642;
w17644 <= not w17630 and not w17643;
w17645 <= not w16955 and not w17629;
w17646 <= not w17628 and w17645;
w17647 <= not w17644 and not w17646;
w17648 <= not b(48) and not w17647;
w17649 <= not w16974 and w17601;
w17650 <= not w17597 and w17649;
w17651 <= not w17598 and not w17601;
w17652 <= not w17650 and not w17651;
w17653 <= not w17630 and not w17652;
w17654 <= not w16964 and not w17629;
w17655 <= not w17628 and w17654;
w17656 <= not w17653 and not w17655;
w17657 <= not b(47) and not w17656;
w17658 <= not w16983 and w17596;
w17659 <= not w17592 and w17658;
w17660 <= not w17593 and not w17596;
w17661 <= not w17659 and not w17660;
w17662 <= not w17630 and not w17661;
w17663 <= not w16973 and not w17629;
w17664 <= not w17628 and w17663;
w17665 <= not w17662 and not w17664;
w17666 <= not b(46) and not w17665;
w17667 <= not w16992 and w17591;
w17668 <= not w17587 and w17667;
w17669 <= not w17588 and not w17591;
w17670 <= not w17668 and not w17669;
w17671 <= not w17630 and not w17670;
w17672 <= not w16982 and not w17629;
w17673 <= not w17628 and w17672;
w17674 <= not w17671 and not w17673;
w17675 <= not b(45) and not w17674;
w17676 <= not w17001 and w17586;
w17677 <= not w17582 and w17676;
w17678 <= not w17583 and not w17586;
w17679 <= not w17677 and not w17678;
w17680 <= not w17630 and not w17679;
w17681 <= not w16991 and not w17629;
w17682 <= not w17628 and w17681;
w17683 <= not w17680 and not w17682;
w17684 <= not b(44) and not w17683;
w17685 <= not w17010 and w17581;
w17686 <= not w17577 and w17685;
w17687 <= not w17578 and not w17581;
w17688 <= not w17686 and not w17687;
w17689 <= not w17630 and not w17688;
w17690 <= not w17000 and not w17629;
w17691 <= not w17628 and w17690;
w17692 <= not w17689 and not w17691;
w17693 <= not b(43) and not w17692;
w17694 <= not w17019 and w17576;
w17695 <= not w17572 and w17694;
w17696 <= not w17573 and not w17576;
w17697 <= not w17695 and not w17696;
w17698 <= not w17630 and not w17697;
w17699 <= not w17009 and not w17629;
w17700 <= not w17628 and w17699;
w17701 <= not w17698 and not w17700;
w17702 <= not b(42) and not w17701;
w17703 <= not w17028 and w17571;
w17704 <= not w17567 and w17703;
w17705 <= not w17568 and not w17571;
w17706 <= not w17704 and not w17705;
w17707 <= not w17630 and not w17706;
w17708 <= not w17018 and not w17629;
w17709 <= not w17628 and w17708;
w17710 <= not w17707 and not w17709;
w17711 <= not b(41) and not w17710;
w17712 <= not w17037 and w17566;
w17713 <= not w17562 and w17712;
w17714 <= not w17563 and not w17566;
w17715 <= not w17713 and not w17714;
w17716 <= not w17630 and not w17715;
w17717 <= not w17027 and not w17629;
w17718 <= not w17628 and w17717;
w17719 <= not w17716 and not w17718;
w17720 <= not b(40) and not w17719;
w17721 <= not w17046 and w17561;
w17722 <= not w17557 and w17721;
w17723 <= not w17558 and not w17561;
w17724 <= not w17722 and not w17723;
w17725 <= not w17630 and not w17724;
w17726 <= not w17036 and not w17629;
w17727 <= not w17628 and w17726;
w17728 <= not w17725 and not w17727;
w17729 <= not b(39) and not w17728;
w17730 <= not w17055 and w17556;
w17731 <= not w17552 and w17730;
w17732 <= not w17553 and not w17556;
w17733 <= not w17731 and not w17732;
w17734 <= not w17630 and not w17733;
w17735 <= not w17045 and not w17629;
w17736 <= not w17628 and w17735;
w17737 <= not w17734 and not w17736;
w17738 <= not b(38) and not w17737;
w17739 <= not w17064 and w17551;
w17740 <= not w17547 and w17739;
w17741 <= not w17548 and not w17551;
w17742 <= not w17740 and not w17741;
w17743 <= not w17630 and not w17742;
w17744 <= not w17054 and not w17629;
w17745 <= not w17628 and w17744;
w17746 <= not w17743 and not w17745;
w17747 <= not b(37) and not w17746;
w17748 <= not w17073 and w17546;
w17749 <= not w17542 and w17748;
w17750 <= not w17543 and not w17546;
w17751 <= not w17749 and not w17750;
w17752 <= not w17630 and not w17751;
w17753 <= not w17063 and not w17629;
w17754 <= not w17628 and w17753;
w17755 <= not w17752 and not w17754;
w17756 <= not b(36) and not w17755;
w17757 <= not w17082 and w17541;
w17758 <= not w17537 and w17757;
w17759 <= not w17538 and not w17541;
w17760 <= not w17758 and not w17759;
w17761 <= not w17630 and not w17760;
w17762 <= not w17072 and not w17629;
w17763 <= not w17628 and w17762;
w17764 <= not w17761 and not w17763;
w17765 <= not b(35) and not w17764;
w17766 <= not w17091 and w17536;
w17767 <= not w17532 and w17766;
w17768 <= not w17533 and not w17536;
w17769 <= not w17767 and not w17768;
w17770 <= not w17630 and not w17769;
w17771 <= not w17081 and not w17629;
w17772 <= not w17628 and w17771;
w17773 <= not w17770 and not w17772;
w17774 <= not b(34) and not w17773;
w17775 <= not w17100 and w17531;
w17776 <= not w17527 and w17775;
w17777 <= not w17528 and not w17531;
w17778 <= not w17776 and not w17777;
w17779 <= not w17630 and not w17778;
w17780 <= not w17090 and not w17629;
w17781 <= not w17628 and w17780;
w17782 <= not w17779 and not w17781;
w17783 <= not b(33) and not w17782;
w17784 <= not w17109 and w17526;
w17785 <= not w17522 and w17784;
w17786 <= not w17523 and not w17526;
w17787 <= not w17785 and not w17786;
w17788 <= not w17630 and not w17787;
w17789 <= not w17099 and not w17629;
w17790 <= not w17628 and w17789;
w17791 <= not w17788 and not w17790;
w17792 <= not b(32) and not w17791;
w17793 <= not w17118 and w17521;
w17794 <= not w17517 and w17793;
w17795 <= not w17518 and not w17521;
w17796 <= not w17794 and not w17795;
w17797 <= not w17630 and not w17796;
w17798 <= not w17108 and not w17629;
w17799 <= not w17628 and w17798;
w17800 <= not w17797 and not w17799;
w17801 <= not b(31) and not w17800;
w17802 <= not w17127 and w17516;
w17803 <= not w17512 and w17802;
w17804 <= not w17513 and not w17516;
w17805 <= not w17803 and not w17804;
w17806 <= not w17630 and not w17805;
w17807 <= not w17117 and not w17629;
w17808 <= not w17628 and w17807;
w17809 <= not w17806 and not w17808;
w17810 <= not b(30) and not w17809;
w17811 <= not w17136 and w17511;
w17812 <= not w17507 and w17811;
w17813 <= not w17508 and not w17511;
w17814 <= not w17812 and not w17813;
w17815 <= not w17630 and not w17814;
w17816 <= not w17126 and not w17629;
w17817 <= not w17628 and w17816;
w17818 <= not w17815 and not w17817;
w17819 <= not b(29) and not w17818;
w17820 <= not w17145 and w17506;
w17821 <= not w17502 and w17820;
w17822 <= not w17503 and not w17506;
w17823 <= not w17821 and not w17822;
w17824 <= not w17630 and not w17823;
w17825 <= not w17135 and not w17629;
w17826 <= not w17628 and w17825;
w17827 <= not w17824 and not w17826;
w17828 <= not b(28) and not w17827;
w17829 <= not w17154 and w17501;
w17830 <= not w17497 and w17829;
w17831 <= not w17498 and not w17501;
w17832 <= not w17830 and not w17831;
w17833 <= not w17630 and not w17832;
w17834 <= not w17144 and not w17629;
w17835 <= not w17628 and w17834;
w17836 <= not w17833 and not w17835;
w17837 <= not b(27) and not w17836;
w17838 <= not w17163 and w17496;
w17839 <= not w17492 and w17838;
w17840 <= not w17493 and not w17496;
w17841 <= not w17839 and not w17840;
w17842 <= not w17630 and not w17841;
w17843 <= not w17153 and not w17629;
w17844 <= not w17628 and w17843;
w17845 <= not w17842 and not w17844;
w17846 <= not b(26) and not w17845;
w17847 <= not w17172 and w17491;
w17848 <= not w17487 and w17847;
w17849 <= not w17488 and not w17491;
w17850 <= not w17848 and not w17849;
w17851 <= not w17630 and not w17850;
w17852 <= not w17162 and not w17629;
w17853 <= not w17628 and w17852;
w17854 <= not w17851 and not w17853;
w17855 <= not b(25) and not w17854;
w17856 <= not w17181 and w17486;
w17857 <= not w17482 and w17856;
w17858 <= not w17483 and not w17486;
w17859 <= not w17857 and not w17858;
w17860 <= not w17630 and not w17859;
w17861 <= not w17171 and not w17629;
w17862 <= not w17628 and w17861;
w17863 <= not w17860 and not w17862;
w17864 <= not b(24) and not w17863;
w17865 <= not w17190 and w17481;
w17866 <= not w17477 and w17865;
w17867 <= not w17478 and not w17481;
w17868 <= not w17866 and not w17867;
w17869 <= not w17630 and not w17868;
w17870 <= not w17180 and not w17629;
w17871 <= not w17628 and w17870;
w17872 <= not w17869 and not w17871;
w17873 <= not b(23) and not w17872;
w17874 <= not w17199 and w17476;
w17875 <= not w17472 and w17874;
w17876 <= not w17473 and not w17476;
w17877 <= not w17875 and not w17876;
w17878 <= not w17630 and not w17877;
w17879 <= not w17189 and not w17629;
w17880 <= not w17628 and w17879;
w17881 <= not w17878 and not w17880;
w17882 <= not b(22) and not w17881;
w17883 <= not w17208 and w17471;
w17884 <= not w17467 and w17883;
w17885 <= not w17468 and not w17471;
w17886 <= not w17884 and not w17885;
w17887 <= not w17630 and not w17886;
w17888 <= not w17198 and not w17629;
w17889 <= not w17628 and w17888;
w17890 <= not w17887 and not w17889;
w17891 <= not b(21) and not w17890;
w17892 <= not w17217 and w17466;
w17893 <= not w17462 and w17892;
w17894 <= not w17463 and not w17466;
w17895 <= not w17893 and not w17894;
w17896 <= not w17630 and not w17895;
w17897 <= not w17207 and not w17629;
w17898 <= not w17628 and w17897;
w17899 <= not w17896 and not w17898;
w17900 <= not b(20) and not w17899;
w17901 <= not w17226 and w17461;
w17902 <= not w17457 and w17901;
w17903 <= not w17458 and not w17461;
w17904 <= not w17902 and not w17903;
w17905 <= not w17630 and not w17904;
w17906 <= not w17216 and not w17629;
w17907 <= not w17628 and w17906;
w17908 <= not w17905 and not w17907;
w17909 <= not b(19) and not w17908;
w17910 <= not w17235 and w17456;
w17911 <= not w17452 and w17910;
w17912 <= not w17453 and not w17456;
w17913 <= not w17911 and not w17912;
w17914 <= not w17630 and not w17913;
w17915 <= not w17225 and not w17629;
w17916 <= not w17628 and w17915;
w17917 <= not w17914 and not w17916;
w17918 <= not b(18) and not w17917;
w17919 <= not w17244 and w17451;
w17920 <= not w17447 and w17919;
w17921 <= not w17448 and not w17451;
w17922 <= not w17920 and not w17921;
w17923 <= not w17630 and not w17922;
w17924 <= not w17234 and not w17629;
w17925 <= not w17628 and w17924;
w17926 <= not w17923 and not w17925;
w17927 <= not b(17) and not w17926;
w17928 <= not w17253 and w17446;
w17929 <= not w17442 and w17928;
w17930 <= not w17443 and not w17446;
w17931 <= not w17929 and not w17930;
w17932 <= not w17630 and not w17931;
w17933 <= not w17243 and not w17629;
w17934 <= not w17628 and w17933;
w17935 <= not w17932 and not w17934;
w17936 <= not b(16) and not w17935;
w17937 <= not w17262 and w17441;
w17938 <= not w17437 and w17937;
w17939 <= not w17438 and not w17441;
w17940 <= not w17938 and not w17939;
w17941 <= not w17630 and not w17940;
w17942 <= not w17252 and not w17629;
w17943 <= not w17628 and w17942;
w17944 <= not w17941 and not w17943;
w17945 <= not b(15) and not w17944;
w17946 <= not w17271 and w17436;
w17947 <= not w17432 and w17946;
w17948 <= not w17433 and not w17436;
w17949 <= not w17947 and not w17948;
w17950 <= not w17630 and not w17949;
w17951 <= not w17261 and not w17629;
w17952 <= not w17628 and w17951;
w17953 <= not w17950 and not w17952;
w17954 <= not b(14) and not w17953;
w17955 <= not w17280 and w17431;
w17956 <= not w17427 and w17955;
w17957 <= not w17428 and not w17431;
w17958 <= not w17956 and not w17957;
w17959 <= not w17630 and not w17958;
w17960 <= not w17270 and not w17629;
w17961 <= not w17628 and w17960;
w17962 <= not w17959 and not w17961;
w17963 <= not b(13) and not w17962;
w17964 <= not w17289 and w17426;
w17965 <= not w17422 and w17964;
w17966 <= not w17423 and not w17426;
w17967 <= not w17965 and not w17966;
w17968 <= not w17630 and not w17967;
w17969 <= not w17279 and not w17629;
w17970 <= not w17628 and w17969;
w17971 <= not w17968 and not w17970;
w17972 <= not b(12) and not w17971;
w17973 <= not w17298 and w17421;
w17974 <= not w17417 and w17973;
w17975 <= not w17418 and not w17421;
w17976 <= not w17974 and not w17975;
w17977 <= not w17630 and not w17976;
w17978 <= not w17288 and not w17629;
w17979 <= not w17628 and w17978;
w17980 <= not w17977 and not w17979;
w17981 <= not b(11) and not w17980;
w17982 <= not w17307 and w17416;
w17983 <= not w17412 and w17982;
w17984 <= not w17413 and not w17416;
w17985 <= not w17983 and not w17984;
w17986 <= not w17630 and not w17985;
w17987 <= not w17297 and not w17629;
w17988 <= not w17628 and w17987;
w17989 <= not w17986 and not w17988;
w17990 <= not b(10) and not w17989;
w17991 <= not w17316 and w17411;
w17992 <= not w17407 and w17991;
w17993 <= not w17408 and not w17411;
w17994 <= not w17992 and not w17993;
w17995 <= not w17630 and not w17994;
w17996 <= not w17306 and not w17629;
w17997 <= not w17628 and w17996;
w17998 <= not w17995 and not w17997;
w17999 <= not b(9) and not w17998;
w18000 <= not w17325 and w17406;
w18001 <= not w17402 and w18000;
w18002 <= not w17403 and not w17406;
w18003 <= not w18001 and not w18002;
w18004 <= not w17630 and not w18003;
w18005 <= not w17315 and not w17629;
w18006 <= not w17628 and w18005;
w18007 <= not w18004 and not w18006;
w18008 <= not b(8) and not w18007;
w18009 <= not w17334 and w17401;
w18010 <= not w17397 and w18009;
w18011 <= not w17398 and not w17401;
w18012 <= not w18010 and not w18011;
w18013 <= not w17630 and not w18012;
w18014 <= not w17324 and not w17629;
w18015 <= not w17628 and w18014;
w18016 <= not w18013 and not w18015;
w18017 <= not b(7) and not w18016;
w18018 <= not w17343 and w17396;
w18019 <= not w17392 and w18018;
w18020 <= not w17393 and not w17396;
w18021 <= not w18019 and not w18020;
w18022 <= not w17630 and not w18021;
w18023 <= not w17333 and not w17629;
w18024 <= not w17628 and w18023;
w18025 <= not w18022 and not w18024;
w18026 <= not b(6) and not w18025;
w18027 <= not w17352 and w17391;
w18028 <= not w17387 and w18027;
w18029 <= not w17388 and not w17391;
w18030 <= not w18028 and not w18029;
w18031 <= not w17630 and not w18030;
w18032 <= not w17342 and not w17629;
w18033 <= not w17628 and w18032;
w18034 <= not w18031 and not w18033;
w18035 <= not b(5) and not w18034;
w18036 <= not w17360 and w17386;
w18037 <= not w17382 and w18036;
w18038 <= not w17383 and not w17386;
w18039 <= not w18037 and not w18038;
w18040 <= not w17630 and not w18039;
w18041 <= not w17351 and not w17629;
w18042 <= not w17628 and w18041;
w18043 <= not w18040 and not w18042;
w18044 <= not b(4) and not w18043;
w18045 <= not w17377 and w17381;
w18046 <= not w17376 and w18045;
w18047 <= not w17378 and not w17381;
w18048 <= not w18046 and not w18047;
w18049 <= not w17630 and not w18048;
w18050 <= not w17359 and not w17629;
w18051 <= not w17628 and w18050;
w18052 <= not w18049 and not w18051;
w18053 <= not b(3) and not w18052;
w18054 <= not w17373 and w17375;
w18055 <= not w17371 and w18054;
w18056 <= not w17376 and not w18055;
w18057 <= not w17630 and w18056;
w18058 <= not w17370 and not w17629;
w18059 <= not w17628 and w18058;
w18060 <= not w18057 and not w18059;
w18061 <= not b(2) and not w18060;
w18062 <= b(0) and not w17630;
w18063 <= a(14) and not w18062;
w18064 <= w17375 and not w17630;
w18065 <= not w18063 and not w18064;
w18066 <= b(1) and not w18065;
w18067 <= not b(1) and not w18064;
w18068 <= not w18063 and w18067;
w18069 <= not w18066 and not w18068;
w18070 <= not a(13) and b(0);
w18071 <= not w18069 and not w18070;
w18072 <= not b(1) and not w18065;
w18073 <= not w18071 and not w18072;
w18074 <= b(2) and not w18059;
w18075 <= not w18057 and w18074;
w18076 <= not w18061 and not w18075;
w18077 <= not w18073 and w18076;
w18078 <= not w18061 and not w18077;
w18079 <= b(3) and not w18051;
w18080 <= not w18049 and w18079;
w18081 <= not w18053 and not w18080;
w18082 <= not w18078 and w18081;
w18083 <= not w18053 and not w18082;
w18084 <= b(4) and not w18042;
w18085 <= not w18040 and w18084;
w18086 <= not w18044 and not w18085;
w18087 <= not w18083 and w18086;
w18088 <= not w18044 and not w18087;
w18089 <= b(5) and not w18033;
w18090 <= not w18031 and w18089;
w18091 <= not w18035 and not w18090;
w18092 <= not w18088 and w18091;
w18093 <= not w18035 and not w18092;
w18094 <= b(6) and not w18024;
w18095 <= not w18022 and w18094;
w18096 <= not w18026 and not w18095;
w18097 <= not w18093 and w18096;
w18098 <= not w18026 and not w18097;
w18099 <= b(7) and not w18015;
w18100 <= not w18013 and w18099;
w18101 <= not w18017 and not w18100;
w18102 <= not w18098 and w18101;
w18103 <= not w18017 and not w18102;
w18104 <= b(8) and not w18006;
w18105 <= not w18004 and w18104;
w18106 <= not w18008 and not w18105;
w18107 <= not w18103 and w18106;
w18108 <= not w18008 and not w18107;
w18109 <= b(9) and not w17997;
w18110 <= not w17995 and w18109;
w18111 <= not w17999 and not w18110;
w18112 <= not w18108 and w18111;
w18113 <= not w17999 and not w18112;
w18114 <= b(10) and not w17988;
w18115 <= not w17986 and w18114;
w18116 <= not w17990 and not w18115;
w18117 <= not w18113 and w18116;
w18118 <= not w17990 and not w18117;
w18119 <= b(11) and not w17979;
w18120 <= not w17977 and w18119;
w18121 <= not w17981 and not w18120;
w18122 <= not w18118 and w18121;
w18123 <= not w17981 and not w18122;
w18124 <= b(12) and not w17970;
w18125 <= not w17968 and w18124;
w18126 <= not w17972 and not w18125;
w18127 <= not w18123 and w18126;
w18128 <= not w17972 and not w18127;
w18129 <= b(13) and not w17961;
w18130 <= not w17959 and w18129;
w18131 <= not w17963 and not w18130;
w18132 <= not w18128 and w18131;
w18133 <= not w17963 and not w18132;
w18134 <= b(14) and not w17952;
w18135 <= not w17950 and w18134;
w18136 <= not w17954 and not w18135;
w18137 <= not w18133 and w18136;
w18138 <= not w17954 and not w18137;
w18139 <= b(15) and not w17943;
w18140 <= not w17941 and w18139;
w18141 <= not w17945 and not w18140;
w18142 <= not w18138 and w18141;
w18143 <= not w17945 and not w18142;
w18144 <= b(16) and not w17934;
w18145 <= not w17932 and w18144;
w18146 <= not w17936 and not w18145;
w18147 <= not w18143 and w18146;
w18148 <= not w17936 and not w18147;
w18149 <= b(17) and not w17925;
w18150 <= not w17923 and w18149;
w18151 <= not w17927 and not w18150;
w18152 <= not w18148 and w18151;
w18153 <= not w17927 and not w18152;
w18154 <= b(18) and not w17916;
w18155 <= not w17914 and w18154;
w18156 <= not w17918 and not w18155;
w18157 <= not w18153 and w18156;
w18158 <= not w17918 and not w18157;
w18159 <= b(19) and not w17907;
w18160 <= not w17905 and w18159;
w18161 <= not w17909 and not w18160;
w18162 <= not w18158 and w18161;
w18163 <= not w17909 and not w18162;
w18164 <= b(20) and not w17898;
w18165 <= not w17896 and w18164;
w18166 <= not w17900 and not w18165;
w18167 <= not w18163 and w18166;
w18168 <= not w17900 and not w18167;
w18169 <= b(21) and not w17889;
w18170 <= not w17887 and w18169;
w18171 <= not w17891 and not w18170;
w18172 <= not w18168 and w18171;
w18173 <= not w17891 and not w18172;
w18174 <= b(22) and not w17880;
w18175 <= not w17878 and w18174;
w18176 <= not w17882 and not w18175;
w18177 <= not w18173 and w18176;
w18178 <= not w17882 and not w18177;
w18179 <= b(23) and not w17871;
w18180 <= not w17869 and w18179;
w18181 <= not w17873 and not w18180;
w18182 <= not w18178 and w18181;
w18183 <= not w17873 and not w18182;
w18184 <= b(24) and not w17862;
w18185 <= not w17860 and w18184;
w18186 <= not w17864 and not w18185;
w18187 <= not w18183 and w18186;
w18188 <= not w17864 and not w18187;
w18189 <= b(25) and not w17853;
w18190 <= not w17851 and w18189;
w18191 <= not w17855 and not w18190;
w18192 <= not w18188 and w18191;
w18193 <= not w17855 and not w18192;
w18194 <= b(26) and not w17844;
w18195 <= not w17842 and w18194;
w18196 <= not w17846 and not w18195;
w18197 <= not w18193 and w18196;
w18198 <= not w17846 and not w18197;
w18199 <= b(27) and not w17835;
w18200 <= not w17833 and w18199;
w18201 <= not w17837 and not w18200;
w18202 <= not w18198 and w18201;
w18203 <= not w17837 and not w18202;
w18204 <= b(28) and not w17826;
w18205 <= not w17824 and w18204;
w18206 <= not w17828 and not w18205;
w18207 <= not w18203 and w18206;
w18208 <= not w17828 and not w18207;
w18209 <= b(29) and not w17817;
w18210 <= not w17815 and w18209;
w18211 <= not w17819 and not w18210;
w18212 <= not w18208 and w18211;
w18213 <= not w17819 and not w18212;
w18214 <= b(30) and not w17808;
w18215 <= not w17806 and w18214;
w18216 <= not w17810 and not w18215;
w18217 <= not w18213 and w18216;
w18218 <= not w17810 and not w18217;
w18219 <= b(31) and not w17799;
w18220 <= not w17797 and w18219;
w18221 <= not w17801 and not w18220;
w18222 <= not w18218 and w18221;
w18223 <= not w17801 and not w18222;
w18224 <= b(32) and not w17790;
w18225 <= not w17788 and w18224;
w18226 <= not w17792 and not w18225;
w18227 <= not w18223 and w18226;
w18228 <= not w17792 and not w18227;
w18229 <= b(33) and not w17781;
w18230 <= not w17779 and w18229;
w18231 <= not w17783 and not w18230;
w18232 <= not w18228 and w18231;
w18233 <= not w17783 and not w18232;
w18234 <= b(34) and not w17772;
w18235 <= not w17770 and w18234;
w18236 <= not w17774 and not w18235;
w18237 <= not w18233 and w18236;
w18238 <= not w17774 and not w18237;
w18239 <= b(35) and not w17763;
w18240 <= not w17761 and w18239;
w18241 <= not w17765 and not w18240;
w18242 <= not w18238 and w18241;
w18243 <= not w17765 and not w18242;
w18244 <= b(36) and not w17754;
w18245 <= not w17752 and w18244;
w18246 <= not w17756 and not w18245;
w18247 <= not w18243 and w18246;
w18248 <= not w17756 and not w18247;
w18249 <= b(37) and not w17745;
w18250 <= not w17743 and w18249;
w18251 <= not w17747 and not w18250;
w18252 <= not w18248 and w18251;
w18253 <= not w17747 and not w18252;
w18254 <= b(38) and not w17736;
w18255 <= not w17734 and w18254;
w18256 <= not w17738 and not w18255;
w18257 <= not w18253 and w18256;
w18258 <= not w17738 and not w18257;
w18259 <= b(39) and not w17727;
w18260 <= not w17725 and w18259;
w18261 <= not w17729 and not w18260;
w18262 <= not w18258 and w18261;
w18263 <= not w17729 and not w18262;
w18264 <= b(40) and not w17718;
w18265 <= not w17716 and w18264;
w18266 <= not w17720 and not w18265;
w18267 <= not w18263 and w18266;
w18268 <= not w17720 and not w18267;
w18269 <= b(41) and not w17709;
w18270 <= not w17707 and w18269;
w18271 <= not w17711 and not w18270;
w18272 <= not w18268 and w18271;
w18273 <= not w17711 and not w18272;
w18274 <= b(42) and not w17700;
w18275 <= not w17698 and w18274;
w18276 <= not w17702 and not w18275;
w18277 <= not w18273 and w18276;
w18278 <= not w17702 and not w18277;
w18279 <= b(43) and not w17691;
w18280 <= not w17689 and w18279;
w18281 <= not w17693 and not w18280;
w18282 <= not w18278 and w18281;
w18283 <= not w17693 and not w18282;
w18284 <= b(44) and not w17682;
w18285 <= not w17680 and w18284;
w18286 <= not w17684 and not w18285;
w18287 <= not w18283 and w18286;
w18288 <= not w17684 and not w18287;
w18289 <= b(45) and not w17673;
w18290 <= not w17671 and w18289;
w18291 <= not w17675 and not w18290;
w18292 <= not w18288 and w18291;
w18293 <= not w17675 and not w18292;
w18294 <= b(46) and not w17664;
w18295 <= not w17662 and w18294;
w18296 <= not w17666 and not w18295;
w18297 <= not w18293 and w18296;
w18298 <= not w17666 and not w18297;
w18299 <= b(47) and not w17655;
w18300 <= not w17653 and w18299;
w18301 <= not w17657 and not w18300;
w18302 <= not w18298 and w18301;
w18303 <= not w17657 and not w18302;
w18304 <= b(48) and not w17646;
w18305 <= not w17644 and w18304;
w18306 <= not w17648 and not w18305;
w18307 <= not w18303 and w18306;
w18308 <= not w17648 and not w18307;
w18309 <= b(49) and not w17637;
w18310 <= not w17635 and w18309;
w18311 <= not w17639 and not w18310;
w18312 <= not w18308 and w18311;
w18313 <= not w17639 and not w18312;
w18314 <= not w16947 and not w17623;
w18315 <= not w17621 and w18314;
w18316 <= not w17612 and w18315;
w18317 <= not w17621 and not w17623;
w18318 <= not w17613 and not w18317;
w18319 <= not w18316 and not w18318;
w18320 <= not w17630 and not w18319;
w18321 <= not w17620 and not w17629;
w18322 <= not w17628 and w18321;
w18323 <= not w18320 and not w18322;
w18324 <= not b(50) and not w18323;
w18325 <= b(50) and not w18322;
w18326 <= not w18320 and w18325;
w18327 <= w140 and w142;
w18328 <= w150 and w18327;
w18329 <= not w18326 and w18328;
w18330 <= not w18324 and w18329;
w18331 <= not w18313 and w18330;
w18332 <= w17625 and not w18323;
w18333 <= not w18331 and not w18332;
w18334 <= not w17648 and w18311;
w18335 <= not w18307 and w18334;
w18336 <= not w18308 and not w18311;
w18337 <= not w18335 and not w18336;
w18338 <= not w18333 and not w18337;
w18339 <= not w17638 and not w18332;
w18340 <= not w18331 and w18339;
w18341 <= not w18338 and not w18340;
w18342 <= not w17639 and not w18326;
w18343 <= not w18324 and w18342;
w18344 <= not w18312 and w18343;
w18345 <= not w18324 and not w18326;
w18346 <= not w18313 and not w18345;
w18347 <= not w18344 and not w18346;
w18348 <= not w18333 and not w18347;
w18349 <= not w18323 and not w18332;
w18350 <= not w18331 and w18349;
w18351 <= not w18348 and not w18350;
w18352 <= not b(51) and not w18351;
w18353 <= not b(50) and not w18341;
w18354 <= not w17657 and w18306;
w18355 <= not w18302 and w18354;
w18356 <= not w18303 and not w18306;
w18357 <= not w18355 and not w18356;
w18358 <= not w18333 and not w18357;
w18359 <= not w17647 and not w18332;
w18360 <= not w18331 and w18359;
w18361 <= not w18358 and not w18360;
w18362 <= not b(49) and not w18361;
w18363 <= not w17666 and w18301;
w18364 <= not w18297 and w18363;
w18365 <= not w18298 and not w18301;
w18366 <= not w18364 and not w18365;
w18367 <= not w18333 and not w18366;
w18368 <= not w17656 and not w18332;
w18369 <= not w18331 and w18368;
w18370 <= not w18367 and not w18369;
w18371 <= not b(48) and not w18370;
w18372 <= not w17675 and w18296;
w18373 <= not w18292 and w18372;
w18374 <= not w18293 and not w18296;
w18375 <= not w18373 and not w18374;
w18376 <= not w18333 and not w18375;
w18377 <= not w17665 and not w18332;
w18378 <= not w18331 and w18377;
w18379 <= not w18376 and not w18378;
w18380 <= not b(47) and not w18379;
w18381 <= not w17684 and w18291;
w18382 <= not w18287 and w18381;
w18383 <= not w18288 and not w18291;
w18384 <= not w18382 and not w18383;
w18385 <= not w18333 and not w18384;
w18386 <= not w17674 and not w18332;
w18387 <= not w18331 and w18386;
w18388 <= not w18385 and not w18387;
w18389 <= not b(46) and not w18388;
w18390 <= not w17693 and w18286;
w18391 <= not w18282 and w18390;
w18392 <= not w18283 and not w18286;
w18393 <= not w18391 and not w18392;
w18394 <= not w18333 and not w18393;
w18395 <= not w17683 and not w18332;
w18396 <= not w18331 and w18395;
w18397 <= not w18394 and not w18396;
w18398 <= not b(45) and not w18397;
w18399 <= not w17702 and w18281;
w18400 <= not w18277 and w18399;
w18401 <= not w18278 and not w18281;
w18402 <= not w18400 and not w18401;
w18403 <= not w18333 and not w18402;
w18404 <= not w17692 and not w18332;
w18405 <= not w18331 and w18404;
w18406 <= not w18403 and not w18405;
w18407 <= not b(44) and not w18406;
w18408 <= not w17711 and w18276;
w18409 <= not w18272 and w18408;
w18410 <= not w18273 and not w18276;
w18411 <= not w18409 and not w18410;
w18412 <= not w18333 and not w18411;
w18413 <= not w17701 and not w18332;
w18414 <= not w18331 and w18413;
w18415 <= not w18412 and not w18414;
w18416 <= not b(43) and not w18415;
w18417 <= not w17720 and w18271;
w18418 <= not w18267 and w18417;
w18419 <= not w18268 and not w18271;
w18420 <= not w18418 and not w18419;
w18421 <= not w18333 and not w18420;
w18422 <= not w17710 and not w18332;
w18423 <= not w18331 and w18422;
w18424 <= not w18421 and not w18423;
w18425 <= not b(42) and not w18424;
w18426 <= not w17729 and w18266;
w18427 <= not w18262 and w18426;
w18428 <= not w18263 and not w18266;
w18429 <= not w18427 and not w18428;
w18430 <= not w18333 and not w18429;
w18431 <= not w17719 and not w18332;
w18432 <= not w18331 and w18431;
w18433 <= not w18430 and not w18432;
w18434 <= not b(41) and not w18433;
w18435 <= not w17738 and w18261;
w18436 <= not w18257 and w18435;
w18437 <= not w18258 and not w18261;
w18438 <= not w18436 and not w18437;
w18439 <= not w18333 and not w18438;
w18440 <= not w17728 and not w18332;
w18441 <= not w18331 and w18440;
w18442 <= not w18439 and not w18441;
w18443 <= not b(40) and not w18442;
w18444 <= not w17747 and w18256;
w18445 <= not w18252 and w18444;
w18446 <= not w18253 and not w18256;
w18447 <= not w18445 and not w18446;
w18448 <= not w18333 and not w18447;
w18449 <= not w17737 and not w18332;
w18450 <= not w18331 and w18449;
w18451 <= not w18448 and not w18450;
w18452 <= not b(39) and not w18451;
w18453 <= not w17756 and w18251;
w18454 <= not w18247 and w18453;
w18455 <= not w18248 and not w18251;
w18456 <= not w18454 and not w18455;
w18457 <= not w18333 and not w18456;
w18458 <= not w17746 and not w18332;
w18459 <= not w18331 and w18458;
w18460 <= not w18457 and not w18459;
w18461 <= not b(38) and not w18460;
w18462 <= not w17765 and w18246;
w18463 <= not w18242 and w18462;
w18464 <= not w18243 and not w18246;
w18465 <= not w18463 and not w18464;
w18466 <= not w18333 and not w18465;
w18467 <= not w17755 and not w18332;
w18468 <= not w18331 and w18467;
w18469 <= not w18466 and not w18468;
w18470 <= not b(37) and not w18469;
w18471 <= not w17774 and w18241;
w18472 <= not w18237 and w18471;
w18473 <= not w18238 and not w18241;
w18474 <= not w18472 and not w18473;
w18475 <= not w18333 and not w18474;
w18476 <= not w17764 and not w18332;
w18477 <= not w18331 and w18476;
w18478 <= not w18475 and not w18477;
w18479 <= not b(36) and not w18478;
w18480 <= not w17783 and w18236;
w18481 <= not w18232 and w18480;
w18482 <= not w18233 and not w18236;
w18483 <= not w18481 and not w18482;
w18484 <= not w18333 and not w18483;
w18485 <= not w17773 and not w18332;
w18486 <= not w18331 and w18485;
w18487 <= not w18484 and not w18486;
w18488 <= not b(35) and not w18487;
w18489 <= not w17792 and w18231;
w18490 <= not w18227 and w18489;
w18491 <= not w18228 and not w18231;
w18492 <= not w18490 and not w18491;
w18493 <= not w18333 and not w18492;
w18494 <= not w17782 and not w18332;
w18495 <= not w18331 and w18494;
w18496 <= not w18493 and not w18495;
w18497 <= not b(34) and not w18496;
w18498 <= not w17801 and w18226;
w18499 <= not w18222 and w18498;
w18500 <= not w18223 and not w18226;
w18501 <= not w18499 and not w18500;
w18502 <= not w18333 and not w18501;
w18503 <= not w17791 and not w18332;
w18504 <= not w18331 and w18503;
w18505 <= not w18502 and not w18504;
w18506 <= not b(33) and not w18505;
w18507 <= not w17810 and w18221;
w18508 <= not w18217 and w18507;
w18509 <= not w18218 and not w18221;
w18510 <= not w18508 and not w18509;
w18511 <= not w18333 and not w18510;
w18512 <= not w17800 and not w18332;
w18513 <= not w18331 and w18512;
w18514 <= not w18511 and not w18513;
w18515 <= not b(32) and not w18514;
w18516 <= not w17819 and w18216;
w18517 <= not w18212 and w18516;
w18518 <= not w18213 and not w18216;
w18519 <= not w18517 and not w18518;
w18520 <= not w18333 and not w18519;
w18521 <= not w17809 and not w18332;
w18522 <= not w18331 and w18521;
w18523 <= not w18520 and not w18522;
w18524 <= not b(31) and not w18523;
w18525 <= not w17828 and w18211;
w18526 <= not w18207 and w18525;
w18527 <= not w18208 and not w18211;
w18528 <= not w18526 and not w18527;
w18529 <= not w18333 and not w18528;
w18530 <= not w17818 and not w18332;
w18531 <= not w18331 and w18530;
w18532 <= not w18529 and not w18531;
w18533 <= not b(30) and not w18532;
w18534 <= not w17837 and w18206;
w18535 <= not w18202 and w18534;
w18536 <= not w18203 and not w18206;
w18537 <= not w18535 and not w18536;
w18538 <= not w18333 and not w18537;
w18539 <= not w17827 and not w18332;
w18540 <= not w18331 and w18539;
w18541 <= not w18538 and not w18540;
w18542 <= not b(29) and not w18541;
w18543 <= not w17846 and w18201;
w18544 <= not w18197 and w18543;
w18545 <= not w18198 and not w18201;
w18546 <= not w18544 and not w18545;
w18547 <= not w18333 and not w18546;
w18548 <= not w17836 and not w18332;
w18549 <= not w18331 and w18548;
w18550 <= not w18547 and not w18549;
w18551 <= not b(28) and not w18550;
w18552 <= not w17855 and w18196;
w18553 <= not w18192 and w18552;
w18554 <= not w18193 and not w18196;
w18555 <= not w18553 and not w18554;
w18556 <= not w18333 and not w18555;
w18557 <= not w17845 and not w18332;
w18558 <= not w18331 and w18557;
w18559 <= not w18556 and not w18558;
w18560 <= not b(27) and not w18559;
w18561 <= not w17864 and w18191;
w18562 <= not w18187 and w18561;
w18563 <= not w18188 and not w18191;
w18564 <= not w18562 and not w18563;
w18565 <= not w18333 and not w18564;
w18566 <= not w17854 and not w18332;
w18567 <= not w18331 and w18566;
w18568 <= not w18565 and not w18567;
w18569 <= not b(26) and not w18568;
w18570 <= not w17873 and w18186;
w18571 <= not w18182 and w18570;
w18572 <= not w18183 and not w18186;
w18573 <= not w18571 and not w18572;
w18574 <= not w18333 and not w18573;
w18575 <= not w17863 and not w18332;
w18576 <= not w18331 and w18575;
w18577 <= not w18574 and not w18576;
w18578 <= not b(25) and not w18577;
w18579 <= not w17882 and w18181;
w18580 <= not w18177 and w18579;
w18581 <= not w18178 and not w18181;
w18582 <= not w18580 and not w18581;
w18583 <= not w18333 and not w18582;
w18584 <= not w17872 and not w18332;
w18585 <= not w18331 and w18584;
w18586 <= not w18583 and not w18585;
w18587 <= not b(24) and not w18586;
w18588 <= not w17891 and w18176;
w18589 <= not w18172 and w18588;
w18590 <= not w18173 and not w18176;
w18591 <= not w18589 and not w18590;
w18592 <= not w18333 and not w18591;
w18593 <= not w17881 and not w18332;
w18594 <= not w18331 and w18593;
w18595 <= not w18592 and not w18594;
w18596 <= not b(23) and not w18595;
w18597 <= not w17900 and w18171;
w18598 <= not w18167 and w18597;
w18599 <= not w18168 and not w18171;
w18600 <= not w18598 and not w18599;
w18601 <= not w18333 and not w18600;
w18602 <= not w17890 and not w18332;
w18603 <= not w18331 and w18602;
w18604 <= not w18601 and not w18603;
w18605 <= not b(22) and not w18604;
w18606 <= not w17909 and w18166;
w18607 <= not w18162 and w18606;
w18608 <= not w18163 and not w18166;
w18609 <= not w18607 and not w18608;
w18610 <= not w18333 and not w18609;
w18611 <= not w17899 and not w18332;
w18612 <= not w18331 and w18611;
w18613 <= not w18610 and not w18612;
w18614 <= not b(21) and not w18613;
w18615 <= not w17918 and w18161;
w18616 <= not w18157 and w18615;
w18617 <= not w18158 and not w18161;
w18618 <= not w18616 and not w18617;
w18619 <= not w18333 and not w18618;
w18620 <= not w17908 and not w18332;
w18621 <= not w18331 and w18620;
w18622 <= not w18619 and not w18621;
w18623 <= not b(20) and not w18622;
w18624 <= not w17927 and w18156;
w18625 <= not w18152 and w18624;
w18626 <= not w18153 and not w18156;
w18627 <= not w18625 and not w18626;
w18628 <= not w18333 and not w18627;
w18629 <= not w17917 and not w18332;
w18630 <= not w18331 and w18629;
w18631 <= not w18628 and not w18630;
w18632 <= not b(19) and not w18631;
w18633 <= not w17936 and w18151;
w18634 <= not w18147 and w18633;
w18635 <= not w18148 and not w18151;
w18636 <= not w18634 and not w18635;
w18637 <= not w18333 and not w18636;
w18638 <= not w17926 and not w18332;
w18639 <= not w18331 and w18638;
w18640 <= not w18637 and not w18639;
w18641 <= not b(18) and not w18640;
w18642 <= not w17945 and w18146;
w18643 <= not w18142 and w18642;
w18644 <= not w18143 and not w18146;
w18645 <= not w18643 and not w18644;
w18646 <= not w18333 and not w18645;
w18647 <= not w17935 and not w18332;
w18648 <= not w18331 and w18647;
w18649 <= not w18646 and not w18648;
w18650 <= not b(17) and not w18649;
w18651 <= not w17954 and w18141;
w18652 <= not w18137 and w18651;
w18653 <= not w18138 and not w18141;
w18654 <= not w18652 and not w18653;
w18655 <= not w18333 and not w18654;
w18656 <= not w17944 and not w18332;
w18657 <= not w18331 and w18656;
w18658 <= not w18655 and not w18657;
w18659 <= not b(16) and not w18658;
w18660 <= not w17963 and w18136;
w18661 <= not w18132 and w18660;
w18662 <= not w18133 and not w18136;
w18663 <= not w18661 and not w18662;
w18664 <= not w18333 and not w18663;
w18665 <= not w17953 and not w18332;
w18666 <= not w18331 and w18665;
w18667 <= not w18664 and not w18666;
w18668 <= not b(15) and not w18667;
w18669 <= not w17972 and w18131;
w18670 <= not w18127 and w18669;
w18671 <= not w18128 and not w18131;
w18672 <= not w18670 and not w18671;
w18673 <= not w18333 and not w18672;
w18674 <= not w17962 and not w18332;
w18675 <= not w18331 and w18674;
w18676 <= not w18673 and not w18675;
w18677 <= not b(14) and not w18676;
w18678 <= not w17981 and w18126;
w18679 <= not w18122 and w18678;
w18680 <= not w18123 and not w18126;
w18681 <= not w18679 and not w18680;
w18682 <= not w18333 and not w18681;
w18683 <= not w17971 and not w18332;
w18684 <= not w18331 and w18683;
w18685 <= not w18682 and not w18684;
w18686 <= not b(13) and not w18685;
w18687 <= not w17990 and w18121;
w18688 <= not w18117 and w18687;
w18689 <= not w18118 and not w18121;
w18690 <= not w18688 and not w18689;
w18691 <= not w18333 and not w18690;
w18692 <= not w17980 and not w18332;
w18693 <= not w18331 and w18692;
w18694 <= not w18691 and not w18693;
w18695 <= not b(12) and not w18694;
w18696 <= not w17999 and w18116;
w18697 <= not w18112 and w18696;
w18698 <= not w18113 and not w18116;
w18699 <= not w18697 and not w18698;
w18700 <= not w18333 and not w18699;
w18701 <= not w17989 and not w18332;
w18702 <= not w18331 and w18701;
w18703 <= not w18700 and not w18702;
w18704 <= not b(11) and not w18703;
w18705 <= not w18008 and w18111;
w18706 <= not w18107 and w18705;
w18707 <= not w18108 and not w18111;
w18708 <= not w18706 and not w18707;
w18709 <= not w18333 and not w18708;
w18710 <= not w17998 and not w18332;
w18711 <= not w18331 and w18710;
w18712 <= not w18709 and not w18711;
w18713 <= not b(10) and not w18712;
w18714 <= not w18017 and w18106;
w18715 <= not w18102 and w18714;
w18716 <= not w18103 and not w18106;
w18717 <= not w18715 and not w18716;
w18718 <= not w18333 and not w18717;
w18719 <= not w18007 and not w18332;
w18720 <= not w18331 and w18719;
w18721 <= not w18718 and not w18720;
w18722 <= not b(9) and not w18721;
w18723 <= not w18026 and w18101;
w18724 <= not w18097 and w18723;
w18725 <= not w18098 and not w18101;
w18726 <= not w18724 and not w18725;
w18727 <= not w18333 and not w18726;
w18728 <= not w18016 and not w18332;
w18729 <= not w18331 and w18728;
w18730 <= not w18727 and not w18729;
w18731 <= not b(8) and not w18730;
w18732 <= not w18035 and w18096;
w18733 <= not w18092 and w18732;
w18734 <= not w18093 and not w18096;
w18735 <= not w18733 and not w18734;
w18736 <= not w18333 and not w18735;
w18737 <= not w18025 and not w18332;
w18738 <= not w18331 and w18737;
w18739 <= not w18736 and not w18738;
w18740 <= not b(7) and not w18739;
w18741 <= not w18044 and w18091;
w18742 <= not w18087 and w18741;
w18743 <= not w18088 and not w18091;
w18744 <= not w18742 and not w18743;
w18745 <= not w18333 and not w18744;
w18746 <= not w18034 and not w18332;
w18747 <= not w18331 and w18746;
w18748 <= not w18745 and not w18747;
w18749 <= not b(6) and not w18748;
w18750 <= not w18053 and w18086;
w18751 <= not w18082 and w18750;
w18752 <= not w18083 and not w18086;
w18753 <= not w18751 and not w18752;
w18754 <= not w18333 and not w18753;
w18755 <= not w18043 and not w18332;
w18756 <= not w18331 and w18755;
w18757 <= not w18754 and not w18756;
w18758 <= not b(5) and not w18757;
w18759 <= not w18061 and w18081;
w18760 <= not w18077 and w18759;
w18761 <= not w18078 and not w18081;
w18762 <= not w18760 and not w18761;
w18763 <= not w18333 and not w18762;
w18764 <= not w18052 and not w18332;
w18765 <= not w18331 and w18764;
w18766 <= not w18763 and not w18765;
w18767 <= not b(4) and not w18766;
w18768 <= not w18072 and w18076;
w18769 <= not w18071 and w18768;
w18770 <= not w18073 and not w18076;
w18771 <= not w18769 and not w18770;
w18772 <= not w18333 and not w18771;
w18773 <= not w18060 and not w18332;
w18774 <= not w18331 and w18773;
w18775 <= not w18772 and not w18774;
w18776 <= not b(3) and not w18775;
w18777 <= not w18068 and w18070;
w18778 <= not w18066 and w18777;
w18779 <= not w18071 and not w18778;
w18780 <= not w18333 and w18779;
w18781 <= not w18065 and not w18332;
w18782 <= not w18331 and w18781;
w18783 <= not w18780 and not w18782;
w18784 <= not b(2) and not w18783;
w18785 <= b(0) and not w18333;
w18786 <= a(13) and not w18785;
w18787 <= w18070 and not w18333;
w18788 <= not w18786 and not w18787;
w18789 <= b(1) and not w18788;
w18790 <= not b(1) and not w18787;
w18791 <= not w18786 and w18790;
w18792 <= not w18789 and not w18791;
w18793 <= not a(12) and b(0);
w18794 <= not w18792 and not w18793;
w18795 <= not b(1) and not w18788;
w18796 <= not w18794 and not w18795;
w18797 <= b(2) and not w18782;
w18798 <= not w18780 and w18797;
w18799 <= not w18784 and not w18798;
w18800 <= not w18796 and w18799;
w18801 <= not w18784 and not w18800;
w18802 <= b(3) and not w18774;
w18803 <= not w18772 and w18802;
w18804 <= not w18776 and not w18803;
w18805 <= not w18801 and w18804;
w18806 <= not w18776 and not w18805;
w18807 <= b(4) and not w18765;
w18808 <= not w18763 and w18807;
w18809 <= not w18767 and not w18808;
w18810 <= not w18806 and w18809;
w18811 <= not w18767 and not w18810;
w18812 <= b(5) and not w18756;
w18813 <= not w18754 and w18812;
w18814 <= not w18758 and not w18813;
w18815 <= not w18811 and w18814;
w18816 <= not w18758 and not w18815;
w18817 <= b(6) and not w18747;
w18818 <= not w18745 and w18817;
w18819 <= not w18749 and not w18818;
w18820 <= not w18816 and w18819;
w18821 <= not w18749 and not w18820;
w18822 <= b(7) and not w18738;
w18823 <= not w18736 and w18822;
w18824 <= not w18740 and not w18823;
w18825 <= not w18821 and w18824;
w18826 <= not w18740 and not w18825;
w18827 <= b(8) and not w18729;
w18828 <= not w18727 and w18827;
w18829 <= not w18731 and not w18828;
w18830 <= not w18826 and w18829;
w18831 <= not w18731 and not w18830;
w18832 <= b(9) and not w18720;
w18833 <= not w18718 and w18832;
w18834 <= not w18722 and not w18833;
w18835 <= not w18831 and w18834;
w18836 <= not w18722 and not w18835;
w18837 <= b(10) and not w18711;
w18838 <= not w18709 and w18837;
w18839 <= not w18713 and not w18838;
w18840 <= not w18836 and w18839;
w18841 <= not w18713 and not w18840;
w18842 <= b(11) and not w18702;
w18843 <= not w18700 and w18842;
w18844 <= not w18704 and not w18843;
w18845 <= not w18841 and w18844;
w18846 <= not w18704 and not w18845;
w18847 <= b(12) and not w18693;
w18848 <= not w18691 and w18847;
w18849 <= not w18695 and not w18848;
w18850 <= not w18846 and w18849;
w18851 <= not w18695 and not w18850;
w18852 <= b(13) and not w18684;
w18853 <= not w18682 and w18852;
w18854 <= not w18686 and not w18853;
w18855 <= not w18851 and w18854;
w18856 <= not w18686 and not w18855;
w18857 <= b(14) and not w18675;
w18858 <= not w18673 and w18857;
w18859 <= not w18677 and not w18858;
w18860 <= not w18856 and w18859;
w18861 <= not w18677 and not w18860;
w18862 <= b(15) and not w18666;
w18863 <= not w18664 and w18862;
w18864 <= not w18668 and not w18863;
w18865 <= not w18861 and w18864;
w18866 <= not w18668 and not w18865;
w18867 <= b(16) and not w18657;
w18868 <= not w18655 and w18867;
w18869 <= not w18659 and not w18868;
w18870 <= not w18866 and w18869;
w18871 <= not w18659 and not w18870;
w18872 <= b(17) and not w18648;
w18873 <= not w18646 and w18872;
w18874 <= not w18650 and not w18873;
w18875 <= not w18871 and w18874;
w18876 <= not w18650 and not w18875;
w18877 <= b(18) and not w18639;
w18878 <= not w18637 and w18877;
w18879 <= not w18641 and not w18878;
w18880 <= not w18876 and w18879;
w18881 <= not w18641 and not w18880;
w18882 <= b(19) and not w18630;
w18883 <= not w18628 and w18882;
w18884 <= not w18632 and not w18883;
w18885 <= not w18881 and w18884;
w18886 <= not w18632 and not w18885;
w18887 <= b(20) and not w18621;
w18888 <= not w18619 and w18887;
w18889 <= not w18623 and not w18888;
w18890 <= not w18886 and w18889;
w18891 <= not w18623 and not w18890;
w18892 <= b(21) and not w18612;
w18893 <= not w18610 and w18892;
w18894 <= not w18614 and not w18893;
w18895 <= not w18891 and w18894;
w18896 <= not w18614 and not w18895;
w18897 <= b(22) and not w18603;
w18898 <= not w18601 and w18897;
w18899 <= not w18605 and not w18898;
w18900 <= not w18896 and w18899;
w18901 <= not w18605 and not w18900;
w18902 <= b(23) and not w18594;
w18903 <= not w18592 and w18902;
w18904 <= not w18596 and not w18903;
w18905 <= not w18901 and w18904;
w18906 <= not w18596 and not w18905;
w18907 <= b(24) and not w18585;
w18908 <= not w18583 and w18907;
w18909 <= not w18587 and not w18908;
w18910 <= not w18906 and w18909;
w18911 <= not w18587 and not w18910;
w18912 <= b(25) and not w18576;
w18913 <= not w18574 and w18912;
w18914 <= not w18578 and not w18913;
w18915 <= not w18911 and w18914;
w18916 <= not w18578 and not w18915;
w18917 <= b(26) and not w18567;
w18918 <= not w18565 and w18917;
w18919 <= not w18569 and not w18918;
w18920 <= not w18916 and w18919;
w18921 <= not w18569 and not w18920;
w18922 <= b(27) and not w18558;
w18923 <= not w18556 and w18922;
w18924 <= not w18560 and not w18923;
w18925 <= not w18921 and w18924;
w18926 <= not w18560 and not w18925;
w18927 <= b(28) and not w18549;
w18928 <= not w18547 and w18927;
w18929 <= not w18551 and not w18928;
w18930 <= not w18926 and w18929;
w18931 <= not w18551 and not w18930;
w18932 <= b(29) and not w18540;
w18933 <= not w18538 and w18932;
w18934 <= not w18542 and not w18933;
w18935 <= not w18931 and w18934;
w18936 <= not w18542 and not w18935;
w18937 <= b(30) and not w18531;
w18938 <= not w18529 and w18937;
w18939 <= not w18533 and not w18938;
w18940 <= not w18936 and w18939;
w18941 <= not w18533 and not w18940;
w18942 <= b(31) and not w18522;
w18943 <= not w18520 and w18942;
w18944 <= not w18524 and not w18943;
w18945 <= not w18941 and w18944;
w18946 <= not w18524 and not w18945;
w18947 <= b(32) and not w18513;
w18948 <= not w18511 and w18947;
w18949 <= not w18515 and not w18948;
w18950 <= not w18946 and w18949;
w18951 <= not w18515 and not w18950;
w18952 <= b(33) and not w18504;
w18953 <= not w18502 and w18952;
w18954 <= not w18506 and not w18953;
w18955 <= not w18951 and w18954;
w18956 <= not w18506 and not w18955;
w18957 <= b(34) and not w18495;
w18958 <= not w18493 and w18957;
w18959 <= not w18497 and not w18958;
w18960 <= not w18956 and w18959;
w18961 <= not w18497 and not w18960;
w18962 <= b(35) and not w18486;
w18963 <= not w18484 and w18962;
w18964 <= not w18488 and not w18963;
w18965 <= not w18961 and w18964;
w18966 <= not w18488 and not w18965;
w18967 <= b(36) and not w18477;
w18968 <= not w18475 and w18967;
w18969 <= not w18479 and not w18968;
w18970 <= not w18966 and w18969;
w18971 <= not w18479 and not w18970;
w18972 <= b(37) and not w18468;
w18973 <= not w18466 and w18972;
w18974 <= not w18470 and not w18973;
w18975 <= not w18971 and w18974;
w18976 <= not w18470 and not w18975;
w18977 <= b(38) and not w18459;
w18978 <= not w18457 and w18977;
w18979 <= not w18461 and not w18978;
w18980 <= not w18976 and w18979;
w18981 <= not w18461 and not w18980;
w18982 <= b(39) and not w18450;
w18983 <= not w18448 and w18982;
w18984 <= not w18452 and not w18983;
w18985 <= not w18981 and w18984;
w18986 <= not w18452 and not w18985;
w18987 <= b(40) and not w18441;
w18988 <= not w18439 and w18987;
w18989 <= not w18443 and not w18988;
w18990 <= not w18986 and w18989;
w18991 <= not w18443 and not w18990;
w18992 <= b(41) and not w18432;
w18993 <= not w18430 and w18992;
w18994 <= not w18434 and not w18993;
w18995 <= not w18991 and w18994;
w18996 <= not w18434 and not w18995;
w18997 <= b(42) and not w18423;
w18998 <= not w18421 and w18997;
w18999 <= not w18425 and not w18998;
w19000 <= not w18996 and w18999;
w19001 <= not w18425 and not w19000;
w19002 <= b(43) and not w18414;
w19003 <= not w18412 and w19002;
w19004 <= not w18416 and not w19003;
w19005 <= not w19001 and w19004;
w19006 <= not w18416 and not w19005;
w19007 <= b(44) and not w18405;
w19008 <= not w18403 and w19007;
w19009 <= not w18407 and not w19008;
w19010 <= not w19006 and w19009;
w19011 <= not w18407 and not w19010;
w19012 <= b(45) and not w18396;
w19013 <= not w18394 and w19012;
w19014 <= not w18398 and not w19013;
w19015 <= not w19011 and w19014;
w19016 <= not w18398 and not w19015;
w19017 <= b(46) and not w18387;
w19018 <= not w18385 and w19017;
w19019 <= not w18389 and not w19018;
w19020 <= not w19016 and w19019;
w19021 <= not w18389 and not w19020;
w19022 <= b(47) and not w18378;
w19023 <= not w18376 and w19022;
w19024 <= not w18380 and not w19023;
w19025 <= not w19021 and w19024;
w19026 <= not w18380 and not w19025;
w19027 <= b(48) and not w18369;
w19028 <= not w18367 and w19027;
w19029 <= not w18371 and not w19028;
w19030 <= not w19026 and w19029;
w19031 <= not w18371 and not w19030;
w19032 <= b(49) and not w18360;
w19033 <= not w18358 and w19032;
w19034 <= not w18362 and not w19033;
w19035 <= not w19031 and w19034;
w19036 <= not w18362 and not w19035;
w19037 <= b(50) and not w18340;
w19038 <= not w18338 and w19037;
w19039 <= not w18353 and not w19038;
w19040 <= not w19036 and w19039;
w19041 <= not w18353 and not w19040;
w19042 <= b(51) and not w18350;
w19043 <= not w18348 and w19042;
w19044 <= not w18352 and not w19043;
w19045 <= not w19041 and w19044;
w19046 <= not w18352 and not w19045;
w19047 <= w31 and not w19046;
w19048 <= not w18341 and not w19047;
w19049 <= not w18362 and w19039;
w19050 <= not w19035 and w19049;
w19051 <= not w19036 and not w19039;
w19052 <= not w19050 and not w19051;
w19053 <= w31 and not w19052;
w19054 <= not w19046 and w19053;
w19055 <= not w19048 and not w19054;
w19056 <= not b(51) and not w19055;
w19057 <= not w18361 and not w19047;
w19058 <= not w18371 and w19034;
w19059 <= not w19030 and w19058;
w19060 <= not w19031 and not w19034;
w19061 <= not w19059 and not w19060;
w19062 <= w31 and not w19061;
w19063 <= not w19046 and w19062;
w19064 <= not w19057 and not w19063;
w19065 <= not b(50) and not w19064;
w19066 <= not w18370 and not w19047;
w19067 <= not w18380 and w19029;
w19068 <= not w19025 and w19067;
w19069 <= not w19026 and not w19029;
w19070 <= not w19068 and not w19069;
w19071 <= w31 and not w19070;
w19072 <= not w19046 and w19071;
w19073 <= not w19066 and not w19072;
w19074 <= not b(49) and not w19073;
w19075 <= not w18379 and not w19047;
w19076 <= not w18389 and w19024;
w19077 <= not w19020 and w19076;
w19078 <= not w19021 and not w19024;
w19079 <= not w19077 and not w19078;
w19080 <= w31 and not w19079;
w19081 <= not w19046 and w19080;
w19082 <= not w19075 and not w19081;
w19083 <= not b(48) and not w19082;
w19084 <= not w18388 and not w19047;
w19085 <= not w18398 and w19019;
w19086 <= not w19015 and w19085;
w19087 <= not w19016 and not w19019;
w19088 <= not w19086 and not w19087;
w19089 <= w31 and not w19088;
w19090 <= not w19046 and w19089;
w19091 <= not w19084 and not w19090;
w19092 <= not b(47) and not w19091;
w19093 <= not w18397 and not w19047;
w19094 <= not w18407 and w19014;
w19095 <= not w19010 and w19094;
w19096 <= not w19011 and not w19014;
w19097 <= not w19095 and not w19096;
w19098 <= w31 and not w19097;
w19099 <= not w19046 and w19098;
w19100 <= not w19093 and not w19099;
w19101 <= not b(46) and not w19100;
w19102 <= not w18406 and not w19047;
w19103 <= not w18416 and w19009;
w19104 <= not w19005 and w19103;
w19105 <= not w19006 and not w19009;
w19106 <= not w19104 and not w19105;
w19107 <= w31 and not w19106;
w19108 <= not w19046 and w19107;
w19109 <= not w19102 and not w19108;
w19110 <= not b(45) and not w19109;
w19111 <= not w18415 and not w19047;
w19112 <= not w18425 and w19004;
w19113 <= not w19000 and w19112;
w19114 <= not w19001 and not w19004;
w19115 <= not w19113 and not w19114;
w19116 <= w31 and not w19115;
w19117 <= not w19046 and w19116;
w19118 <= not w19111 and not w19117;
w19119 <= not b(44) and not w19118;
w19120 <= not w18424 and not w19047;
w19121 <= not w18434 and w18999;
w19122 <= not w18995 and w19121;
w19123 <= not w18996 and not w18999;
w19124 <= not w19122 and not w19123;
w19125 <= w31 and not w19124;
w19126 <= not w19046 and w19125;
w19127 <= not w19120 and not w19126;
w19128 <= not b(43) and not w19127;
w19129 <= not w18433 and not w19047;
w19130 <= not w18443 and w18994;
w19131 <= not w18990 and w19130;
w19132 <= not w18991 and not w18994;
w19133 <= not w19131 and not w19132;
w19134 <= w31 and not w19133;
w19135 <= not w19046 and w19134;
w19136 <= not w19129 and not w19135;
w19137 <= not b(42) and not w19136;
w19138 <= not w18442 and not w19047;
w19139 <= not w18452 and w18989;
w19140 <= not w18985 and w19139;
w19141 <= not w18986 and not w18989;
w19142 <= not w19140 and not w19141;
w19143 <= w31 and not w19142;
w19144 <= not w19046 and w19143;
w19145 <= not w19138 and not w19144;
w19146 <= not b(41) and not w19145;
w19147 <= not w18451 and not w19047;
w19148 <= not w18461 and w18984;
w19149 <= not w18980 and w19148;
w19150 <= not w18981 and not w18984;
w19151 <= not w19149 and not w19150;
w19152 <= w31 and not w19151;
w19153 <= not w19046 and w19152;
w19154 <= not w19147 and not w19153;
w19155 <= not b(40) and not w19154;
w19156 <= not w18460 and not w19047;
w19157 <= not w18470 and w18979;
w19158 <= not w18975 and w19157;
w19159 <= not w18976 and not w18979;
w19160 <= not w19158 and not w19159;
w19161 <= w31 and not w19160;
w19162 <= not w19046 and w19161;
w19163 <= not w19156 and not w19162;
w19164 <= not b(39) and not w19163;
w19165 <= not w18469 and not w19047;
w19166 <= not w18479 and w18974;
w19167 <= not w18970 and w19166;
w19168 <= not w18971 and not w18974;
w19169 <= not w19167 and not w19168;
w19170 <= w31 and not w19169;
w19171 <= not w19046 and w19170;
w19172 <= not w19165 and not w19171;
w19173 <= not b(38) and not w19172;
w19174 <= not w18478 and not w19047;
w19175 <= not w18488 and w18969;
w19176 <= not w18965 and w19175;
w19177 <= not w18966 and not w18969;
w19178 <= not w19176 and not w19177;
w19179 <= w31 and not w19178;
w19180 <= not w19046 and w19179;
w19181 <= not w19174 and not w19180;
w19182 <= not b(37) and not w19181;
w19183 <= not w18487 and not w19047;
w19184 <= not w18497 and w18964;
w19185 <= not w18960 and w19184;
w19186 <= not w18961 and not w18964;
w19187 <= not w19185 and not w19186;
w19188 <= w31 and not w19187;
w19189 <= not w19046 and w19188;
w19190 <= not w19183 and not w19189;
w19191 <= not b(36) and not w19190;
w19192 <= not w18496 and not w19047;
w19193 <= not w18506 and w18959;
w19194 <= not w18955 and w19193;
w19195 <= not w18956 and not w18959;
w19196 <= not w19194 and not w19195;
w19197 <= w31 and not w19196;
w19198 <= not w19046 and w19197;
w19199 <= not w19192 and not w19198;
w19200 <= not b(35) and not w19199;
w19201 <= not w18505 and not w19047;
w19202 <= not w18515 and w18954;
w19203 <= not w18950 and w19202;
w19204 <= not w18951 and not w18954;
w19205 <= not w19203 and not w19204;
w19206 <= w31 and not w19205;
w19207 <= not w19046 and w19206;
w19208 <= not w19201 and not w19207;
w19209 <= not b(34) and not w19208;
w19210 <= not w18514 and not w19047;
w19211 <= not w18524 and w18949;
w19212 <= not w18945 and w19211;
w19213 <= not w18946 and not w18949;
w19214 <= not w19212 and not w19213;
w19215 <= w31 and not w19214;
w19216 <= not w19046 and w19215;
w19217 <= not w19210 and not w19216;
w19218 <= not b(33) and not w19217;
w19219 <= not w18523 and not w19047;
w19220 <= not w18533 and w18944;
w19221 <= not w18940 and w19220;
w19222 <= not w18941 and not w18944;
w19223 <= not w19221 and not w19222;
w19224 <= w31 and not w19223;
w19225 <= not w19046 and w19224;
w19226 <= not w19219 and not w19225;
w19227 <= not b(32) and not w19226;
w19228 <= not w18532 and not w19047;
w19229 <= not w18542 and w18939;
w19230 <= not w18935 and w19229;
w19231 <= not w18936 and not w18939;
w19232 <= not w19230 and not w19231;
w19233 <= w31 and not w19232;
w19234 <= not w19046 and w19233;
w19235 <= not w19228 and not w19234;
w19236 <= not b(31) and not w19235;
w19237 <= not w18541 and not w19047;
w19238 <= not w18551 and w18934;
w19239 <= not w18930 and w19238;
w19240 <= not w18931 and not w18934;
w19241 <= not w19239 and not w19240;
w19242 <= w31 and not w19241;
w19243 <= not w19046 and w19242;
w19244 <= not w19237 and not w19243;
w19245 <= not b(30) and not w19244;
w19246 <= not w18550 and not w19047;
w19247 <= not w18560 and w18929;
w19248 <= not w18925 and w19247;
w19249 <= not w18926 and not w18929;
w19250 <= not w19248 and not w19249;
w19251 <= w31 and not w19250;
w19252 <= not w19046 and w19251;
w19253 <= not w19246 and not w19252;
w19254 <= not b(29) and not w19253;
w19255 <= not w18559 and not w19047;
w19256 <= not w18569 and w18924;
w19257 <= not w18920 and w19256;
w19258 <= not w18921 and not w18924;
w19259 <= not w19257 and not w19258;
w19260 <= w31 and not w19259;
w19261 <= not w19046 and w19260;
w19262 <= not w19255 and not w19261;
w19263 <= not b(28) and not w19262;
w19264 <= not w18568 and not w19047;
w19265 <= not w18578 and w18919;
w19266 <= not w18915 and w19265;
w19267 <= not w18916 and not w18919;
w19268 <= not w19266 and not w19267;
w19269 <= w31 and not w19268;
w19270 <= not w19046 and w19269;
w19271 <= not w19264 and not w19270;
w19272 <= not b(27) and not w19271;
w19273 <= not w18577 and not w19047;
w19274 <= not w18587 and w18914;
w19275 <= not w18910 and w19274;
w19276 <= not w18911 and not w18914;
w19277 <= not w19275 and not w19276;
w19278 <= w31 and not w19277;
w19279 <= not w19046 and w19278;
w19280 <= not w19273 and not w19279;
w19281 <= not b(26) and not w19280;
w19282 <= not w18586 and not w19047;
w19283 <= not w18596 and w18909;
w19284 <= not w18905 and w19283;
w19285 <= not w18906 and not w18909;
w19286 <= not w19284 and not w19285;
w19287 <= w31 and not w19286;
w19288 <= not w19046 and w19287;
w19289 <= not w19282 and not w19288;
w19290 <= not b(25) and not w19289;
w19291 <= not w18595 and not w19047;
w19292 <= not w18605 and w18904;
w19293 <= not w18900 and w19292;
w19294 <= not w18901 and not w18904;
w19295 <= not w19293 and not w19294;
w19296 <= w31 and not w19295;
w19297 <= not w19046 and w19296;
w19298 <= not w19291 and not w19297;
w19299 <= not b(24) and not w19298;
w19300 <= not w18604 and not w19047;
w19301 <= not w18614 and w18899;
w19302 <= not w18895 and w19301;
w19303 <= not w18896 and not w18899;
w19304 <= not w19302 and not w19303;
w19305 <= w31 and not w19304;
w19306 <= not w19046 and w19305;
w19307 <= not w19300 and not w19306;
w19308 <= not b(23) and not w19307;
w19309 <= not w18613 and not w19047;
w19310 <= not w18623 and w18894;
w19311 <= not w18890 and w19310;
w19312 <= not w18891 and not w18894;
w19313 <= not w19311 and not w19312;
w19314 <= w31 and not w19313;
w19315 <= not w19046 and w19314;
w19316 <= not w19309 and not w19315;
w19317 <= not b(22) and not w19316;
w19318 <= not w18622 and not w19047;
w19319 <= not w18632 and w18889;
w19320 <= not w18885 and w19319;
w19321 <= not w18886 and not w18889;
w19322 <= not w19320 and not w19321;
w19323 <= w31 and not w19322;
w19324 <= not w19046 and w19323;
w19325 <= not w19318 and not w19324;
w19326 <= not b(21) and not w19325;
w19327 <= not w18631 and not w19047;
w19328 <= not w18641 and w18884;
w19329 <= not w18880 and w19328;
w19330 <= not w18881 and not w18884;
w19331 <= not w19329 and not w19330;
w19332 <= w31 and not w19331;
w19333 <= not w19046 and w19332;
w19334 <= not w19327 and not w19333;
w19335 <= not b(20) and not w19334;
w19336 <= not w18640 and not w19047;
w19337 <= not w18650 and w18879;
w19338 <= not w18875 and w19337;
w19339 <= not w18876 and not w18879;
w19340 <= not w19338 and not w19339;
w19341 <= w31 and not w19340;
w19342 <= not w19046 and w19341;
w19343 <= not w19336 and not w19342;
w19344 <= not b(19) and not w19343;
w19345 <= not w18649 and not w19047;
w19346 <= not w18659 and w18874;
w19347 <= not w18870 and w19346;
w19348 <= not w18871 and not w18874;
w19349 <= not w19347 and not w19348;
w19350 <= w31 and not w19349;
w19351 <= not w19046 and w19350;
w19352 <= not w19345 and not w19351;
w19353 <= not b(18) and not w19352;
w19354 <= not w18658 and not w19047;
w19355 <= not w18668 and w18869;
w19356 <= not w18865 and w19355;
w19357 <= not w18866 and not w18869;
w19358 <= not w19356 and not w19357;
w19359 <= w31 and not w19358;
w19360 <= not w19046 and w19359;
w19361 <= not w19354 and not w19360;
w19362 <= not b(17) and not w19361;
w19363 <= not w18667 and not w19047;
w19364 <= not w18677 and w18864;
w19365 <= not w18860 and w19364;
w19366 <= not w18861 and not w18864;
w19367 <= not w19365 and not w19366;
w19368 <= w31 and not w19367;
w19369 <= not w19046 and w19368;
w19370 <= not w19363 and not w19369;
w19371 <= not b(16) and not w19370;
w19372 <= not w18676 and not w19047;
w19373 <= not w18686 and w18859;
w19374 <= not w18855 and w19373;
w19375 <= not w18856 and not w18859;
w19376 <= not w19374 and not w19375;
w19377 <= w31 and not w19376;
w19378 <= not w19046 and w19377;
w19379 <= not w19372 and not w19378;
w19380 <= not b(15) and not w19379;
w19381 <= not w18685 and not w19047;
w19382 <= not w18695 and w18854;
w19383 <= not w18850 and w19382;
w19384 <= not w18851 and not w18854;
w19385 <= not w19383 and not w19384;
w19386 <= w31 and not w19385;
w19387 <= not w19046 and w19386;
w19388 <= not w19381 and not w19387;
w19389 <= not b(14) and not w19388;
w19390 <= not w18694 and not w19047;
w19391 <= not w18704 and w18849;
w19392 <= not w18845 and w19391;
w19393 <= not w18846 and not w18849;
w19394 <= not w19392 and not w19393;
w19395 <= w31 and not w19394;
w19396 <= not w19046 and w19395;
w19397 <= not w19390 and not w19396;
w19398 <= not b(13) and not w19397;
w19399 <= not w18703 and not w19047;
w19400 <= not w18713 and w18844;
w19401 <= not w18840 and w19400;
w19402 <= not w18841 and not w18844;
w19403 <= not w19401 and not w19402;
w19404 <= w31 and not w19403;
w19405 <= not w19046 and w19404;
w19406 <= not w19399 and not w19405;
w19407 <= not b(12) and not w19406;
w19408 <= not w18712 and not w19047;
w19409 <= not w18722 and w18839;
w19410 <= not w18835 and w19409;
w19411 <= not w18836 and not w18839;
w19412 <= not w19410 and not w19411;
w19413 <= w31 and not w19412;
w19414 <= not w19046 and w19413;
w19415 <= not w19408 and not w19414;
w19416 <= not b(11) and not w19415;
w19417 <= not w18721 and not w19047;
w19418 <= not w18731 and w18834;
w19419 <= not w18830 and w19418;
w19420 <= not w18831 and not w18834;
w19421 <= not w19419 and not w19420;
w19422 <= w31 and not w19421;
w19423 <= not w19046 and w19422;
w19424 <= not w19417 and not w19423;
w19425 <= not b(10) and not w19424;
w19426 <= not w18730 and not w19047;
w19427 <= not w18740 and w18829;
w19428 <= not w18825 and w19427;
w19429 <= not w18826 and not w18829;
w19430 <= not w19428 and not w19429;
w19431 <= w31 and not w19430;
w19432 <= not w19046 and w19431;
w19433 <= not w19426 and not w19432;
w19434 <= not b(9) and not w19433;
w19435 <= not w18739 and not w19047;
w19436 <= not w18749 and w18824;
w19437 <= not w18820 and w19436;
w19438 <= not w18821 and not w18824;
w19439 <= not w19437 and not w19438;
w19440 <= w31 and not w19439;
w19441 <= not w19046 and w19440;
w19442 <= not w19435 and not w19441;
w19443 <= not b(8) and not w19442;
w19444 <= not w18748 and not w19047;
w19445 <= not w18758 and w18819;
w19446 <= not w18815 and w19445;
w19447 <= not w18816 and not w18819;
w19448 <= not w19446 and not w19447;
w19449 <= w31 and not w19448;
w19450 <= not w19046 and w19449;
w19451 <= not w19444 and not w19450;
w19452 <= not b(7) and not w19451;
w19453 <= not w18757 and not w19047;
w19454 <= not w18767 and w18814;
w19455 <= not w18810 and w19454;
w19456 <= not w18811 and not w18814;
w19457 <= not w19455 and not w19456;
w19458 <= w31 and not w19457;
w19459 <= not w19046 and w19458;
w19460 <= not w19453 and not w19459;
w19461 <= not b(6) and not w19460;
w19462 <= not w18766 and not w19047;
w19463 <= not w18776 and w18809;
w19464 <= not w18805 and w19463;
w19465 <= not w18806 and not w18809;
w19466 <= not w19464 and not w19465;
w19467 <= w31 and not w19466;
w19468 <= not w19046 and w19467;
w19469 <= not w19462 and not w19468;
w19470 <= not b(5) and not w19469;
w19471 <= not w18775 and not w19047;
w19472 <= not w18784 and w18804;
w19473 <= not w18800 and w19472;
w19474 <= not w18801 and not w18804;
w19475 <= not w19473 and not w19474;
w19476 <= w31 and not w19475;
w19477 <= not w19046 and w19476;
w19478 <= not w19471 and not w19477;
w19479 <= not b(4) and not w19478;
w19480 <= not w18783 and not w19047;
w19481 <= not w18795 and w18799;
w19482 <= not w18794 and w19481;
w19483 <= not w18796 and not w18799;
w19484 <= not w19482 and not w19483;
w19485 <= w31 and not w19484;
w19486 <= not w19046 and w19485;
w19487 <= not w19480 and not w19486;
w19488 <= not b(3) and not w19487;
w19489 <= not w18788 and not w19047;
w19490 <= not w18791 and w18793;
w19491 <= not w18789 and w19490;
w19492 <= w31 and not w19491;
w19493 <= not w18794 and w19492;
w19494 <= not w19046 and w19493;
w19495 <= not w19489 and not w19494;
w19496 <= not b(2) and not w19495;
w19497 <= b(0) and not b(52);
w19498 <= w140 and w19497;
w19499 <= w150 and w19498;
w19500 <= not w19046 and w19499;
w19501 <= a(12) and not w19500;
w19502 <= w29 and w18793;
w19503 <= w80 and w19502;
w19504 <= not w19046 and w19503;
w19505 <= not w19501 and not w19504;
w19506 <= b(1) and not w19505;
w19507 <= not b(1) and not w19504;
w19508 <= not w19501 and w19507;
w19509 <= not w19506 and not w19508;
w19510 <= not a(11) and b(0);
w19511 <= not w19509 and not w19510;
w19512 <= not b(1) and not w19505;
w19513 <= not w19511 and not w19512;
w19514 <= b(2) and not w19494;
w19515 <= not w19489 and w19514;
w19516 <= not w19496 and not w19515;
w19517 <= not w19513 and w19516;
w19518 <= not w19496 and not w19517;
w19519 <= b(3) and not w19486;
w19520 <= not w19480 and w19519;
w19521 <= not w19488 and not w19520;
w19522 <= not w19518 and w19521;
w19523 <= not w19488 and not w19522;
w19524 <= b(4) and not w19477;
w19525 <= not w19471 and w19524;
w19526 <= not w19479 and not w19525;
w19527 <= not w19523 and w19526;
w19528 <= not w19479 and not w19527;
w19529 <= b(5) and not w19468;
w19530 <= not w19462 and w19529;
w19531 <= not w19470 and not w19530;
w19532 <= not w19528 and w19531;
w19533 <= not w19470 and not w19532;
w19534 <= b(6) and not w19459;
w19535 <= not w19453 and w19534;
w19536 <= not w19461 and not w19535;
w19537 <= not w19533 and w19536;
w19538 <= not w19461 and not w19537;
w19539 <= b(7) and not w19450;
w19540 <= not w19444 and w19539;
w19541 <= not w19452 and not w19540;
w19542 <= not w19538 and w19541;
w19543 <= not w19452 and not w19542;
w19544 <= b(8) and not w19441;
w19545 <= not w19435 and w19544;
w19546 <= not w19443 and not w19545;
w19547 <= not w19543 and w19546;
w19548 <= not w19443 and not w19547;
w19549 <= b(9) and not w19432;
w19550 <= not w19426 and w19549;
w19551 <= not w19434 and not w19550;
w19552 <= not w19548 and w19551;
w19553 <= not w19434 and not w19552;
w19554 <= b(10) and not w19423;
w19555 <= not w19417 and w19554;
w19556 <= not w19425 and not w19555;
w19557 <= not w19553 and w19556;
w19558 <= not w19425 and not w19557;
w19559 <= b(11) and not w19414;
w19560 <= not w19408 and w19559;
w19561 <= not w19416 and not w19560;
w19562 <= not w19558 and w19561;
w19563 <= not w19416 and not w19562;
w19564 <= b(12) and not w19405;
w19565 <= not w19399 and w19564;
w19566 <= not w19407 and not w19565;
w19567 <= not w19563 and w19566;
w19568 <= not w19407 and not w19567;
w19569 <= b(13) and not w19396;
w19570 <= not w19390 and w19569;
w19571 <= not w19398 and not w19570;
w19572 <= not w19568 and w19571;
w19573 <= not w19398 and not w19572;
w19574 <= b(14) and not w19387;
w19575 <= not w19381 and w19574;
w19576 <= not w19389 and not w19575;
w19577 <= not w19573 and w19576;
w19578 <= not w19389 and not w19577;
w19579 <= b(15) and not w19378;
w19580 <= not w19372 and w19579;
w19581 <= not w19380 and not w19580;
w19582 <= not w19578 and w19581;
w19583 <= not w19380 and not w19582;
w19584 <= b(16) and not w19369;
w19585 <= not w19363 and w19584;
w19586 <= not w19371 and not w19585;
w19587 <= not w19583 and w19586;
w19588 <= not w19371 and not w19587;
w19589 <= b(17) and not w19360;
w19590 <= not w19354 and w19589;
w19591 <= not w19362 and not w19590;
w19592 <= not w19588 and w19591;
w19593 <= not w19362 and not w19592;
w19594 <= b(18) and not w19351;
w19595 <= not w19345 and w19594;
w19596 <= not w19353 and not w19595;
w19597 <= not w19593 and w19596;
w19598 <= not w19353 and not w19597;
w19599 <= b(19) and not w19342;
w19600 <= not w19336 and w19599;
w19601 <= not w19344 and not w19600;
w19602 <= not w19598 and w19601;
w19603 <= not w19344 and not w19602;
w19604 <= b(20) and not w19333;
w19605 <= not w19327 and w19604;
w19606 <= not w19335 and not w19605;
w19607 <= not w19603 and w19606;
w19608 <= not w19335 and not w19607;
w19609 <= b(21) and not w19324;
w19610 <= not w19318 and w19609;
w19611 <= not w19326 and not w19610;
w19612 <= not w19608 and w19611;
w19613 <= not w19326 and not w19612;
w19614 <= b(22) and not w19315;
w19615 <= not w19309 and w19614;
w19616 <= not w19317 and not w19615;
w19617 <= not w19613 and w19616;
w19618 <= not w19317 and not w19617;
w19619 <= b(23) and not w19306;
w19620 <= not w19300 and w19619;
w19621 <= not w19308 and not w19620;
w19622 <= not w19618 and w19621;
w19623 <= not w19308 and not w19622;
w19624 <= b(24) and not w19297;
w19625 <= not w19291 and w19624;
w19626 <= not w19299 and not w19625;
w19627 <= not w19623 and w19626;
w19628 <= not w19299 and not w19627;
w19629 <= b(25) and not w19288;
w19630 <= not w19282 and w19629;
w19631 <= not w19290 and not w19630;
w19632 <= not w19628 and w19631;
w19633 <= not w19290 and not w19632;
w19634 <= b(26) and not w19279;
w19635 <= not w19273 and w19634;
w19636 <= not w19281 and not w19635;
w19637 <= not w19633 and w19636;
w19638 <= not w19281 and not w19637;
w19639 <= b(27) and not w19270;
w19640 <= not w19264 and w19639;
w19641 <= not w19272 and not w19640;
w19642 <= not w19638 and w19641;
w19643 <= not w19272 and not w19642;
w19644 <= b(28) and not w19261;
w19645 <= not w19255 and w19644;
w19646 <= not w19263 and not w19645;
w19647 <= not w19643 and w19646;
w19648 <= not w19263 and not w19647;
w19649 <= b(29) and not w19252;
w19650 <= not w19246 and w19649;
w19651 <= not w19254 and not w19650;
w19652 <= not w19648 and w19651;
w19653 <= not w19254 and not w19652;
w19654 <= b(30) and not w19243;
w19655 <= not w19237 and w19654;
w19656 <= not w19245 and not w19655;
w19657 <= not w19653 and w19656;
w19658 <= not w19245 and not w19657;
w19659 <= b(31) and not w19234;
w19660 <= not w19228 and w19659;
w19661 <= not w19236 and not w19660;
w19662 <= not w19658 and w19661;
w19663 <= not w19236 and not w19662;
w19664 <= b(32) and not w19225;
w19665 <= not w19219 and w19664;
w19666 <= not w19227 and not w19665;
w19667 <= not w19663 and w19666;
w19668 <= not w19227 and not w19667;
w19669 <= b(33) and not w19216;
w19670 <= not w19210 and w19669;
w19671 <= not w19218 and not w19670;
w19672 <= not w19668 and w19671;
w19673 <= not w19218 and not w19672;
w19674 <= b(34) and not w19207;
w19675 <= not w19201 and w19674;
w19676 <= not w19209 and not w19675;
w19677 <= not w19673 and w19676;
w19678 <= not w19209 and not w19677;
w19679 <= b(35) and not w19198;
w19680 <= not w19192 and w19679;
w19681 <= not w19200 and not w19680;
w19682 <= not w19678 and w19681;
w19683 <= not w19200 and not w19682;
w19684 <= b(36) and not w19189;
w19685 <= not w19183 and w19684;
w19686 <= not w19191 and not w19685;
w19687 <= not w19683 and w19686;
w19688 <= not w19191 and not w19687;
w19689 <= b(37) and not w19180;
w19690 <= not w19174 and w19689;
w19691 <= not w19182 and not w19690;
w19692 <= not w19688 and w19691;
w19693 <= not w19182 and not w19692;
w19694 <= b(38) and not w19171;
w19695 <= not w19165 and w19694;
w19696 <= not w19173 and not w19695;
w19697 <= not w19693 and w19696;
w19698 <= not w19173 and not w19697;
w19699 <= b(39) and not w19162;
w19700 <= not w19156 and w19699;
w19701 <= not w19164 and not w19700;
w19702 <= not w19698 and w19701;
w19703 <= not w19164 and not w19702;
w19704 <= b(40) and not w19153;
w19705 <= not w19147 and w19704;
w19706 <= not w19155 and not w19705;
w19707 <= not w19703 and w19706;
w19708 <= not w19155 and not w19707;
w19709 <= b(41) and not w19144;
w19710 <= not w19138 and w19709;
w19711 <= not w19146 and not w19710;
w19712 <= not w19708 and w19711;
w19713 <= not w19146 and not w19712;
w19714 <= b(42) and not w19135;
w19715 <= not w19129 and w19714;
w19716 <= not w19137 and not w19715;
w19717 <= not w19713 and w19716;
w19718 <= not w19137 and not w19717;
w19719 <= b(43) and not w19126;
w19720 <= not w19120 and w19719;
w19721 <= not w19128 and not w19720;
w19722 <= not w19718 and w19721;
w19723 <= not w19128 and not w19722;
w19724 <= b(44) and not w19117;
w19725 <= not w19111 and w19724;
w19726 <= not w19119 and not w19725;
w19727 <= not w19723 and w19726;
w19728 <= not w19119 and not w19727;
w19729 <= b(45) and not w19108;
w19730 <= not w19102 and w19729;
w19731 <= not w19110 and not w19730;
w19732 <= not w19728 and w19731;
w19733 <= not w19110 and not w19732;
w19734 <= b(46) and not w19099;
w19735 <= not w19093 and w19734;
w19736 <= not w19101 and not w19735;
w19737 <= not w19733 and w19736;
w19738 <= not w19101 and not w19737;
w19739 <= b(47) and not w19090;
w19740 <= not w19084 and w19739;
w19741 <= not w19092 and not w19740;
w19742 <= not w19738 and w19741;
w19743 <= not w19092 and not w19742;
w19744 <= b(48) and not w19081;
w19745 <= not w19075 and w19744;
w19746 <= not w19083 and not w19745;
w19747 <= not w19743 and w19746;
w19748 <= not w19083 and not w19747;
w19749 <= b(49) and not w19072;
w19750 <= not w19066 and w19749;
w19751 <= not w19074 and not w19750;
w19752 <= not w19748 and w19751;
w19753 <= not w19074 and not w19752;
w19754 <= b(50) and not w19063;
w19755 <= not w19057 and w19754;
w19756 <= not w19065 and not w19755;
w19757 <= not w19753 and w19756;
w19758 <= not w19065 and not w19757;
w19759 <= b(51) and not w19054;
w19760 <= not w19048 and w19759;
w19761 <= not w19056 and not w19760;
w19762 <= not w19758 and w19761;
w19763 <= not w19056 and not w19762;
w19764 <= not w18351 and not w19047;
w19765 <= not w18353 and w19044;
w19766 <= not w19040 and w19765;
w19767 <= not w19041 and not w19044;
w19768 <= not w19766 and not w19767;
w19769 <= w19047 and not w19768;
w19770 <= not w19764 and not w19769;
w19771 <= not b(52) and not w19770;
w19772 <= b(52) and not w19764;
w19773 <= not w19769 and w19772;
w19774 <= w338 and not w19773;
w19775 <= not w19771 and w19774;
w19776 <= not w19763 and w19775;
w19777 <= w31 and not w19770;
w19778 <= not w19776 and not w19777;
w19779 <= not w19065 and w19761;
w19780 <= not w19757 and w19779;
w19781 <= not w19758 and not w19761;
w19782 <= not w19780 and not w19781;
w19783 <= not w19778 and not w19782;
w19784 <= not w19055 and not w19777;
w19785 <= not w19776 and w19784;
w19786 <= not w19783 and not w19785;
w19787 <= not b(52) and not w19786;
w19788 <= not w19074 and w19756;
w19789 <= not w19752 and w19788;
w19790 <= not w19753 and not w19756;
w19791 <= not w19789 and not w19790;
w19792 <= not w19778 and not w19791;
w19793 <= not w19064 and not w19777;
w19794 <= not w19776 and w19793;
w19795 <= not w19792 and not w19794;
w19796 <= not b(51) and not w19795;
w19797 <= not w19083 and w19751;
w19798 <= not w19747 and w19797;
w19799 <= not w19748 and not w19751;
w19800 <= not w19798 and not w19799;
w19801 <= not w19778 and not w19800;
w19802 <= not w19073 and not w19777;
w19803 <= not w19776 and w19802;
w19804 <= not w19801 and not w19803;
w19805 <= not b(50) and not w19804;
w19806 <= not w19092 and w19746;
w19807 <= not w19742 and w19806;
w19808 <= not w19743 and not w19746;
w19809 <= not w19807 and not w19808;
w19810 <= not w19778 and not w19809;
w19811 <= not w19082 and not w19777;
w19812 <= not w19776 and w19811;
w19813 <= not w19810 and not w19812;
w19814 <= not b(49) and not w19813;
w19815 <= not w19101 and w19741;
w19816 <= not w19737 and w19815;
w19817 <= not w19738 and not w19741;
w19818 <= not w19816 and not w19817;
w19819 <= not w19778 and not w19818;
w19820 <= not w19091 and not w19777;
w19821 <= not w19776 and w19820;
w19822 <= not w19819 and not w19821;
w19823 <= not b(48) and not w19822;
w19824 <= not w19110 and w19736;
w19825 <= not w19732 and w19824;
w19826 <= not w19733 and not w19736;
w19827 <= not w19825 and not w19826;
w19828 <= not w19778 and not w19827;
w19829 <= not w19100 and not w19777;
w19830 <= not w19776 and w19829;
w19831 <= not w19828 and not w19830;
w19832 <= not b(47) and not w19831;
w19833 <= not w19119 and w19731;
w19834 <= not w19727 and w19833;
w19835 <= not w19728 and not w19731;
w19836 <= not w19834 and not w19835;
w19837 <= not w19778 and not w19836;
w19838 <= not w19109 and not w19777;
w19839 <= not w19776 and w19838;
w19840 <= not w19837 and not w19839;
w19841 <= not b(46) and not w19840;
w19842 <= not w19128 and w19726;
w19843 <= not w19722 and w19842;
w19844 <= not w19723 and not w19726;
w19845 <= not w19843 and not w19844;
w19846 <= not w19778 and not w19845;
w19847 <= not w19118 and not w19777;
w19848 <= not w19776 and w19847;
w19849 <= not w19846 and not w19848;
w19850 <= not b(45) and not w19849;
w19851 <= not w19137 and w19721;
w19852 <= not w19717 and w19851;
w19853 <= not w19718 and not w19721;
w19854 <= not w19852 and not w19853;
w19855 <= not w19778 and not w19854;
w19856 <= not w19127 and not w19777;
w19857 <= not w19776 and w19856;
w19858 <= not w19855 and not w19857;
w19859 <= not b(44) and not w19858;
w19860 <= not w19146 and w19716;
w19861 <= not w19712 and w19860;
w19862 <= not w19713 and not w19716;
w19863 <= not w19861 and not w19862;
w19864 <= not w19778 and not w19863;
w19865 <= not w19136 and not w19777;
w19866 <= not w19776 and w19865;
w19867 <= not w19864 and not w19866;
w19868 <= not b(43) and not w19867;
w19869 <= not w19155 and w19711;
w19870 <= not w19707 and w19869;
w19871 <= not w19708 and not w19711;
w19872 <= not w19870 and not w19871;
w19873 <= not w19778 and not w19872;
w19874 <= not w19145 and not w19777;
w19875 <= not w19776 and w19874;
w19876 <= not w19873 and not w19875;
w19877 <= not b(42) and not w19876;
w19878 <= not w19164 and w19706;
w19879 <= not w19702 and w19878;
w19880 <= not w19703 and not w19706;
w19881 <= not w19879 and not w19880;
w19882 <= not w19778 and not w19881;
w19883 <= not w19154 and not w19777;
w19884 <= not w19776 and w19883;
w19885 <= not w19882 and not w19884;
w19886 <= not b(41) and not w19885;
w19887 <= not w19173 and w19701;
w19888 <= not w19697 and w19887;
w19889 <= not w19698 and not w19701;
w19890 <= not w19888 and not w19889;
w19891 <= not w19778 and not w19890;
w19892 <= not w19163 and not w19777;
w19893 <= not w19776 and w19892;
w19894 <= not w19891 and not w19893;
w19895 <= not b(40) and not w19894;
w19896 <= not w19182 and w19696;
w19897 <= not w19692 and w19896;
w19898 <= not w19693 and not w19696;
w19899 <= not w19897 and not w19898;
w19900 <= not w19778 and not w19899;
w19901 <= not w19172 and not w19777;
w19902 <= not w19776 and w19901;
w19903 <= not w19900 and not w19902;
w19904 <= not b(39) and not w19903;
w19905 <= not w19191 and w19691;
w19906 <= not w19687 and w19905;
w19907 <= not w19688 and not w19691;
w19908 <= not w19906 and not w19907;
w19909 <= not w19778 and not w19908;
w19910 <= not w19181 and not w19777;
w19911 <= not w19776 and w19910;
w19912 <= not w19909 and not w19911;
w19913 <= not b(38) and not w19912;
w19914 <= not w19200 and w19686;
w19915 <= not w19682 and w19914;
w19916 <= not w19683 and not w19686;
w19917 <= not w19915 and not w19916;
w19918 <= not w19778 and not w19917;
w19919 <= not w19190 and not w19777;
w19920 <= not w19776 and w19919;
w19921 <= not w19918 and not w19920;
w19922 <= not b(37) and not w19921;
w19923 <= not w19209 and w19681;
w19924 <= not w19677 and w19923;
w19925 <= not w19678 and not w19681;
w19926 <= not w19924 and not w19925;
w19927 <= not w19778 and not w19926;
w19928 <= not w19199 and not w19777;
w19929 <= not w19776 and w19928;
w19930 <= not w19927 and not w19929;
w19931 <= not b(36) and not w19930;
w19932 <= not w19218 and w19676;
w19933 <= not w19672 and w19932;
w19934 <= not w19673 and not w19676;
w19935 <= not w19933 and not w19934;
w19936 <= not w19778 and not w19935;
w19937 <= not w19208 and not w19777;
w19938 <= not w19776 and w19937;
w19939 <= not w19936 and not w19938;
w19940 <= not b(35) and not w19939;
w19941 <= not w19227 and w19671;
w19942 <= not w19667 and w19941;
w19943 <= not w19668 and not w19671;
w19944 <= not w19942 and not w19943;
w19945 <= not w19778 and not w19944;
w19946 <= not w19217 and not w19777;
w19947 <= not w19776 and w19946;
w19948 <= not w19945 and not w19947;
w19949 <= not b(34) and not w19948;
w19950 <= not w19236 and w19666;
w19951 <= not w19662 and w19950;
w19952 <= not w19663 and not w19666;
w19953 <= not w19951 and not w19952;
w19954 <= not w19778 and not w19953;
w19955 <= not w19226 and not w19777;
w19956 <= not w19776 and w19955;
w19957 <= not w19954 and not w19956;
w19958 <= not b(33) and not w19957;
w19959 <= not w19245 and w19661;
w19960 <= not w19657 and w19959;
w19961 <= not w19658 and not w19661;
w19962 <= not w19960 and not w19961;
w19963 <= not w19778 and not w19962;
w19964 <= not w19235 and not w19777;
w19965 <= not w19776 and w19964;
w19966 <= not w19963 and not w19965;
w19967 <= not b(32) and not w19966;
w19968 <= not w19254 and w19656;
w19969 <= not w19652 and w19968;
w19970 <= not w19653 and not w19656;
w19971 <= not w19969 and not w19970;
w19972 <= not w19778 and not w19971;
w19973 <= not w19244 and not w19777;
w19974 <= not w19776 and w19973;
w19975 <= not w19972 and not w19974;
w19976 <= not b(31) and not w19975;
w19977 <= not w19263 and w19651;
w19978 <= not w19647 and w19977;
w19979 <= not w19648 and not w19651;
w19980 <= not w19978 and not w19979;
w19981 <= not w19778 and not w19980;
w19982 <= not w19253 and not w19777;
w19983 <= not w19776 and w19982;
w19984 <= not w19981 and not w19983;
w19985 <= not b(30) and not w19984;
w19986 <= not w19272 and w19646;
w19987 <= not w19642 and w19986;
w19988 <= not w19643 and not w19646;
w19989 <= not w19987 and not w19988;
w19990 <= not w19778 and not w19989;
w19991 <= not w19262 and not w19777;
w19992 <= not w19776 and w19991;
w19993 <= not w19990 and not w19992;
w19994 <= not b(29) and not w19993;
w19995 <= not w19281 and w19641;
w19996 <= not w19637 and w19995;
w19997 <= not w19638 and not w19641;
w19998 <= not w19996 and not w19997;
w19999 <= not w19778 and not w19998;
w20000 <= not w19271 and not w19777;
w20001 <= not w19776 and w20000;
w20002 <= not w19999 and not w20001;
w20003 <= not b(28) and not w20002;
w20004 <= not w19290 and w19636;
w20005 <= not w19632 and w20004;
w20006 <= not w19633 and not w19636;
w20007 <= not w20005 and not w20006;
w20008 <= not w19778 and not w20007;
w20009 <= not w19280 and not w19777;
w20010 <= not w19776 and w20009;
w20011 <= not w20008 and not w20010;
w20012 <= not b(27) and not w20011;
w20013 <= not w19299 and w19631;
w20014 <= not w19627 and w20013;
w20015 <= not w19628 and not w19631;
w20016 <= not w20014 and not w20015;
w20017 <= not w19778 and not w20016;
w20018 <= not w19289 and not w19777;
w20019 <= not w19776 and w20018;
w20020 <= not w20017 and not w20019;
w20021 <= not b(26) and not w20020;
w20022 <= not w19308 and w19626;
w20023 <= not w19622 and w20022;
w20024 <= not w19623 and not w19626;
w20025 <= not w20023 and not w20024;
w20026 <= not w19778 and not w20025;
w20027 <= not w19298 and not w19777;
w20028 <= not w19776 and w20027;
w20029 <= not w20026 and not w20028;
w20030 <= not b(25) and not w20029;
w20031 <= not w19317 and w19621;
w20032 <= not w19617 and w20031;
w20033 <= not w19618 and not w19621;
w20034 <= not w20032 and not w20033;
w20035 <= not w19778 and not w20034;
w20036 <= not w19307 and not w19777;
w20037 <= not w19776 and w20036;
w20038 <= not w20035 and not w20037;
w20039 <= not b(24) and not w20038;
w20040 <= not w19326 and w19616;
w20041 <= not w19612 and w20040;
w20042 <= not w19613 and not w19616;
w20043 <= not w20041 and not w20042;
w20044 <= not w19778 and not w20043;
w20045 <= not w19316 and not w19777;
w20046 <= not w19776 and w20045;
w20047 <= not w20044 and not w20046;
w20048 <= not b(23) and not w20047;
w20049 <= not w19335 and w19611;
w20050 <= not w19607 and w20049;
w20051 <= not w19608 and not w19611;
w20052 <= not w20050 and not w20051;
w20053 <= not w19778 and not w20052;
w20054 <= not w19325 and not w19777;
w20055 <= not w19776 and w20054;
w20056 <= not w20053 and not w20055;
w20057 <= not b(22) and not w20056;
w20058 <= not w19344 and w19606;
w20059 <= not w19602 and w20058;
w20060 <= not w19603 and not w19606;
w20061 <= not w20059 and not w20060;
w20062 <= not w19778 and not w20061;
w20063 <= not w19334 and not w19777;
w20064 <= not w19776 and w20063;
w20065 <= not w20062 and not w20064;
w20066 <= not b(21) and not w20065;
w20067 <= not w19353 and w19601;
w20068 <= not w19597 and w20067;
w20069 <= not w19598 and not w19601;
w20070 <= not w20068 and not w20069;
w20071 <= not w19778 and not w20070;
w20072 <= not w19343 and not w19777;
w20073 <= not w19776 and w20072;
w20074 <= not w20071 and not w20073;
w20075 <= not b(20) and not w20074;
w20076 <= not w19362 and w19596;
w20077 <= not w19592 and w20076;
w20078 <= not w19593 and not w19596;
w20079 <= not w20077 and not w20078;
w20080 <= not w19778 and not w20079;
w20081 <= not w19352 and not w19777;
w20082 <= not w19776 and w20081;
w20083 <= not w20080 and not w20082;
w20084 <= not b(19) and not w20083;
w20085 <= not w19371 and w19591;
w20086 <= not w19587 and w20085;
w20087 <= not w19588 and not w19591;
w20088 <= not w20086 and not w20087;
w20089 <= not w19778 and not w20088;
w20090 <= not w19361 and not w19777;
w20091 <= not w19776 and w20090;
w20092 <= not w20089 and not w20091;
w20093 <= not b(18) and not w20092;
w20094 <= not w19380 and w19586;
w20095 <= not w19582 and w20094;
w20096 <= not w19583 and not w19586;
w20097 <= not w20095 and not w20096;
w20098 <= not w19778 and not w20097;
w20099 <= not w19370 and not w19777;
w20100 <= not w19776 and w20099;
w20101 <= not w20098 and not w20100;
w20102 <= not b(17) and not w20101;
w20103 <= not w19389 and w19581;
w20104 <= not w19577 and w20103;
w20105 <= not w19578 and not w19581;
w20106 <= not w20104 and not w20105;
w20107 <= not w19778 and not w20106;
w20108 <= not w19379 and not w19777;
w20109 <= not w19776 and w20108;
w20110 <= not w20107 and not w20109;
w20111 <= not b(16) and not w20110;
w20112 <= not w19398 and w19576;
w20113 <= not w19572 and w20112;
w20114 <= not w19573 and not w19576;
w20115 <= not w20113 and not w20114;
w20116 <= not w19778 and not w20115;
w20117 <= not w19388 and not w19777;
w20118 <= not w19776 and w20117;
w20119 <= not w20116 and not w20118;
w20120 <= not b(15) and not w20119;
w20121 <= not w19407 and w19571;
w20122 <= not w19567 and w20121;
w20123 <= not w19568 and not w19571;
w20124 <= not w20122 and not w20123;
w20125 <= not w19778 and not w20124;
w20126 <= not w19397 and not w19777;
w20127 <= not w19776 and w20126;
w20128 <= not w20125 and not w20127;
w20129 <= not b(14) and not w20128;
w20130 <= not w19416 and w19566;
w20131 <= not w19562 and w20130;
w20132 <= not w19563 and not w19566;
w20133 <= not w20131 and not w20132;
w20134 <= not w19778 and not w20133;
w20135 <= not w19406 and not w19777;
w20136 <= not w19776 and w20135;
w20137 <= not w20134 and not w20136;
w20138 <= not b(13) and not w20137;
w20139 <= not w19425 and w19561;
w20140 <= not w19557 and w20139;
w20141 <= not w19558 and not w19561;
w20142 <= not w20140 and not w20141;
w20143 <= not w19778 and not w20142;
w20144 <= not w19415 and not w19777;
w20145 <= not w19776 and w20144;
w20146 <= not w20143 and not w20145;
w20147 <= not b(12) and not w20146;
w20148 <= not w19434 and w19556;
w20149 <= not w19552 and w20148;
w20150 <= not w19553 and not w19556;
w20151 <= not w20149 and not w20150;
w20152 <= not w19778 and not w20151;
w20153 <= not w19424 and not w19777;
w20154 <= not w19776 and w20153;
w20155 <= not w20152 and not w20154;
w20156 <= not b(11) and not w20155;
w20157 <= not w19443 and w19551;
w20158 <= not w19547 and w20157;
w20159 <= not w19548 and not w19551;
w20160 <= not w20158 and not w20159;
w20161 <= not w19778 and not w20160;
w20162 <= not w19433 and not w19777;
w20163 <= not w19776 and w20162;
w20164 <= not w20161 and not w20163;
w20165 <= not b(10) and not w20164;
w20166 <= not w19452 and w19546;
w20167 <= not w19542 and w20166;
w20168 <= not w19543 and not w19546;
w20169 <= not w20167 and not w20168;
w20170 <= not w19778 and not w20169;
w20171 <= not w19442 and not w19777;
w20172 <= not w19776 and w20171;
w20173 <= not w20170 and not w20172;
w20174 <= not b(9) and not w20173;
w20175 <= not w19461 and w19541;
w20176 <= not w19537 and w20175;
w20177 <= not w19538 and not w19541;
w20178 <= not w20176 and not w20177;
w20179 <= not w19778 and not w20178;
w20180 <= not w19451 and not w19777;
w20181 <= not w19776 and w20180;
w20182 <= not w20179 and not w20181;
w20183 <= not b(8) and not w20182;
w20184 <= not w19470 and w19536;
w20185 <= not w19532 and w20184;
w20186 <= not w19533 and not w19536;
w20187 <= not w20185 and not w20186;
w20188 <= not w19778 and not w20187;
w20189 <= not w19460 and not w19777;
w20190 <= not w19776 and w20189;
w20191 <= not w20188 and not w20190;
w20192 <= not b(7) and not w20191;
w20193 <= not w19479 and w19531;
w20194 <= not w19527 and w20193;
w20195 <= not w19528 and not w19531;
w20196 <= not w20194 and not w20195;
w20197 <= not w19778 and not w20196;
w20198 <= not w19469 and not w19777;
w20199 <= not w19776 and w20198;
w20200 <= not w20197 and not w20199;
w20201 <= not b(6) and not w20200;
w20202 <= not w19488 and w19526;
w20203 <= not w19522 and w20202;
w20204 <= not w19523 and not w19526;
w20205 <= not w20203 and not w20204;
w20206 <= not w19778 and not w20205;
w20207 <= not w19478 and not w19777;
w20208 <= not w19776 and w20207;
w20209 <= not w20206 and not w20208;
w20210 <= not b(5) and not w20209;
w20211 <= not w19496 and w19521;
w20212 <= not w19517 and w20211;
w20213 <= not w19518 and not w19521;
w20214 <= not w20212 and not w20213;
w20215 <= not w19778 and not w20214;
w20216 <= not w19487 and not w19777;
w20217 <= not w19776 and w20216;
w20218 <= not w20215 and not w20217;
w20219 <= not b(4) and not w20218;
w20220 <= not w19512 and w19516;
w20221 <= not w19511 and w20220;
w20222 <= not w19513 and not w19516;
w20223 <= not w20221 and not w20222;
w20224 <= not w19778 and not w20223;
w20225 <= not w19495 and not w19777;
w20226 <= not w19776 and w20225;
w20227 <= not w20224 and not w20226;
w20228 <= not b(3) and not w20227;
w20229 <= not w19508 and w19510;
w20230 <= not w19506 and w20229;
w20231 <= not w19511 and not w20230;
w20232 <= not w19778 and w20231;
w20233 <= not w19505 and not w19777;
w20234 <= not w19776 and w20233;
w20235 <= not w20232 and not w20234;
w20236 <= not b(2) and not w20235;
w20237 <= b(0) and not w19778;
w20238 <= a(11) and not w20237;
w20239 <= w19510 and not w19778;
w20240 <= not w20238 and not w20239;
w20241 <= b(1) and not w20240;
w20242 <= not b(1) and not w20239;
w20243 <= not w20238 and w20242;
w20244 <= not w20241 and not w20243;
w20245 <= not a(10) and b(0);
w20246 <= not w20244 and not w20245;
w20247 <= not b(1) and not w20240;
w20248 <= not w20246 and not w20247;
w20249 <= b(2) and not w20234;
w20250 <= not w20232 and w20249;
w20251 <= not w20236 and not w20250;
w20252 <= not w20248 and w20251;
w20253 <= not w20236 and not w20252;
w20254 <= b(3) and not w20226;
w20255 <= not w20224 and w20254;
w20256 <= not w20228 and not w20255;
w20257 <= not w20253 and w20256;
w20258 <= not w20228 and not w20257;
w20259 <= b(4) and not w20217;
w20260 <= not w20215 and w20259;
w20261 <= not w20219 and not w20260;
w20262 <= not w20258 and w20261;
w20263 <= not w20219 and not w20262;
w20264 <= b(5) and not w20208;
w20265 <= not w20206 and w20264;
w20266 <= not w20210 and not w20265;
w20267 <= not w20263 and w20266;
w20268 <= not w20210 and not w20267;
w20269 <= b(6) and not w20199;
w20270 <= not w20197 and w20269;
w20271 <= not w20201 and not w20270;
w20272 <= not w20268 and w20271;
w20273 <= not w20201 and not w20272;
w20274 <= b(7) and not w20190;
w20275 <= not w20188 and w20274;
w20276 <= not w20192 and not w20275;
w20277 <= not w20273 and w20276;
w20278 <= not w20192 and not w20277;
w20279 <= b(8) and not w20181;
w20280 <= not w20179 and w20279;
w20281 <= not w20183 and not w20280;
w20282 <= not w20278 and w20281;
w20283 <= not w20183 and not w20282;
w20284 <= b(9) and not w20172;
w20285 <= not w20170 and w20284;
w20286 <= not w20174 and not w20285;
w20287 <= not w20283 and w20286;
w20288 <= not w20174 and not w20287;
w20289 <= b(10) and not w20163;
w20290 <= not w20161 and w20289;
w20291 <= not w20165 and not w20290;
w20292 <= not w20288 and w20291;
w20293 <= not w20165 and not w20292;
w20294 <= b(11) and not w20154;
w20295 <= not w20152 and w20294;
w20296 <= not w20156 and not w20295;
w20297 <= not w20293 and w20296;
w20298 <= not w20156 and not w20297;
w20299 <= b(12) and not w20145;
w20300 <= not w20143 and w20299;
w20301 <= not w20147 and not w20300;
w20302 <= not w20298 and w20301;
w20303 <= not w20147 and not w20302;
w20304 <= b(13) and not w20136;
w20305 <= not w20134 and w20304;
w20306 <= not w20138 and not w20305;
w20307 <= not w20303 and w20306;
w20308 <= not w20138 and not w20307;
w20309 <= b(14) and not w20127;
w20310 <= not w20125 and w20309;
w20311 <= not w20129 and not w20310;
w20312 <= not w20308 and w20311;
w20313 <= not w20129 and not w20312;
w20314 <= b(15) and not w20118;
w20315 <= not w20116 and w20314;
w20316 <= not w20120 and not w20315;
w20317 <= not w20313 and w20316;
w20318 <= not w20120 and not w20317;
w20319 <= b(16) and not w20109;
w20320 <= not w20107 and w20319;
w20321 <= not w20111 and not w20320;
w20322 <= not w20318 and w20321;
w20323 <= not w20111 and not w20322;
w20324 <= b(17) and not w20100;
w20325 <= not w20098 and w20324;
w20326 <= not w20102 and not w20325;
w20327 <= not w20323 and w20326;
w20328 <= not w20102 and not w20327;
w20329 <= b(18) and not w20091;
w20330 <= not w20089 and w20329;
w20331 <= not w20093 and not w20330;
w20332 <= not w20328 and w20331;
w20333 <= not w20093 and not w20332;
w20334 <= b(19) and not w20082;
w20335 <= not w20080 and w20334;
w20336 <= not w20084 and not w20335;
w20337 <= not w20333 and w20336;
w20338 <= not w20084 and not w20337;
w20339 <= b(20) and not w20073;
w20340 <= not w20071 and w20339;
w20341 <= not w20075 and not w20340;
w20342 <= not w20338 and w20341;
w20343 <= not w20075 and not w20342;
w20344 <= b(21) and not w20064;
w20345 <= not w20062 and w20344;
w20346 <= not w20066 and not w20345;
w20347 <= not w20343 and w20346;
w20348 <= not w20066 and not w20347;
w20349 <= b(22) and not w20055;
w20350 <= not w20053 and w20349;
w20351 <= not w20057 and not w20350;
w20352 <= not w20348 and w20351;
w20353 <= not w20057 and not w20352;
w20354 <= b(23) and not w20046;
w20355 <= not w20044 and w20354;
w20356 <= not w20048 and not w20355;
w20357 <= not w20353 and w20356;
w20358 <= not w20048 and not w20357;
w20359 <= b(24) and not w20037;
w20360 <= not w20035 and w20359;
w20361 <= not w20039 and not w20360;
w20362 <= not w20358 and w20361;
w20363 <= not w20039 and not w20362;
w20364 <= b(25) and not w20028;
w20365 <= not w20026 and w20364;
w20366 <= not w20030 and not w20365;
w20367 <= not w20363 and w20366;
w20368 <= not w20030 and not w20367;
w20369 <= b(26) and not w20019;
w20370 <= not w20017 and w20369;
w20371 <= not w20021 and not w20370;
w20372 <= not w20368 and w20371;
w20373 <= not w20021 and not w20372;
w20374 <= b(27) and not w20010;
w20375 <= not w20008 and w20374;
w20376 <= not w20012 and not w20375;
w20377 <= not w20373 and w20376;
w20378 <= not w20012 and not w20377;
w20379 <= b(28) and not w20001;
w20380 <= not w19999 and w20379;
w20381 <= not w20003 and not w20380;
w20382 <= not w20378 and w20381;
w20383 <= not w20003 and not w20382;
w20384 <= b(29) and not w19992;
w20385 <= not w19990 and w20384;
w20386 <= not w19994 and not w20385;
w20387 <= not w20383 and w20386;
w20388 <= not w19994 and not w20387;
w20389 <= b(30) and not w19983;
w20390 <= not w19981 and w20389;
w20391 <= not w19985 and not w20390;
w20392 <= not w20388 and w20391;
w20393 <= not w19985 and not w20392;
w20394 <= b(31) and not w19974;
w20395 <= not w19972 and w20394;
w20396 <= not w19976 and not w20395;
w20397 <= not w20393 and w20396;
w20398 <= not w19976 and not w20397;
w20399 <= b(32) and not w19965;
w20400 <= not w19963 and w20399;
w20401 <= not w19967 and not w20400;
w20402 <= not w20398 and w20401;
w20403 <= not w19967 and not w20402;
w20404 <= b(33) and not w19956;
w20405 <= not w19954 and w20404;
w20406 <= not w19958 and not w20405;
w20407 <= not w20403 and w20406;
w20408 <= not w19958 and not w20407;
w20409 <= b(34) and not w19947;
w20410 <= not w19945 and w20409;
w20411 <= not w19949 and not w20410;
w20412 <= not w20408 and w20411;
w20413 <= not w19949 and not w20412;
w20414 <= b(35) and not w19938;
w20415 <= not w19936 and w20414;
w20416 <= not w19940 and not w20415;
w20417 <= not w20413 and w20416;
w20418 <= not w19940 and not w20417;
w20419 <= b(36) and not w19929;
w20420 <= not w19927 and w20419;
w20421 <= not w19931 and not w20420;
w20422 <= not w20418 and w20421;
w20423 <= not w19931 and not w20422;
w20424 <= b(37) and not w19920;
w20425 <= not w19918 and w20424;
w20426 <= not w19922 and not w20425;
w20427 <= not w20423 and w20426;
w20428 <= not w19922 and not w20427;
w20429 <= b(38) and not w19911;
w20430 <= not w19909 and w20429;
w20431 <= not w19913 and not w20430;
w20432 <= not w20428 and w20431;
w20433 <= not w19913 and not w20432;
w20434 <= b(39) and not w19902;
w20435 <= not w19900 and w20434;
w20436 <= not w19904 and not w20435;
w20437 <= not w20433 and w20436;
w20438 <= not w19904 and not w20437;
w20439 <= b(40) and not w19893;
w20440 <= not w19891 and w20439;
w20441 <= not w19895 and not w20440;
w20442 <= not w20438 and w20441;
w20443 <= not w19895 and not w20442;
w20444 <= b(41) and not w19884;
w20445 <= not w19882 and w20444;
w20446 <= not w19886 and not w20445;
w20447 <= not w20443 and w20446;
w20448 <= not w19886 and not w20447;
w20449 <= b(42) and not w19875;
w20450 <= not w19873 and w20449;
w20451 <= not w19877 and not w20450;
w20452 <= not w20448 and w20451;
w20453 <= not w19877 and not w20452;
w20454 <= b(43) and not w19866;
w20455 <= not w19864 and w20454;
w20456 <= not w19868 and not w20455;
w20457 <= not w20453 and w20456;
w20458 <= not w19868 and not w20457;
w20459 <= b(44) and not w19857;
w20460 <= not w19855 and w20459;
w20461 <= not w19859 and not w20460;
w20462 <= not w20458 and w20461;
w20463 <= not w19859 and not w20462;
w20464 <= b(45) and not w19848;
w20465 <= not w19846 and w20464;
w20466 <= not w19850 and not w20465;
w20467 <= not w20463 and w20466;
w20468 <= not w19850 and not w20467;
w20469 <= b(46) and not w19839;
w20470 <= not w19837 and w20469;
w20471 <= not w19841 and not w20470;
w20472 <= not w20468 and w20471;
w20473 <= not w19841 and not w20472;
w20474 <= b(47) and not w19830;
w20475 <= not w19828 and w20474;
w20476 <= not w19832 and not w20475;
w20477 <= not w20473 and w20476;
w20478 <= not w19832 and not w20477;
w20479 <= b(48) and not w19821;
w20480 <= not w19819 and w20479;
w20481 <= not w19823 and not w20480;
w20482 <= not w20478 and w20481;
w20483 <= not w19823 and not w20482;
w20484 <= b(49) and not w19812;
w20485 <= not w19810 and w20484;
w20486 <= not w19814 and not w20485;
w20487 <= not w20483 and w20486;
w20488 <= not w19814 and not w20487;
w20489 <= b(50) and not w19803;
w20490 <= not w19801 and w20489;
w20491 <= not w19805 and not w20490;
w20492 <= not w20488 and w20491;
w20493 <= not w19805 and not w20492;
w20494 <= b(51) and not w19794;
w20495 <= not w19792 and w20494;
w20496 <= not w19796 and not w20495;
w20497 <= not w20493 and w20496;
w20498 <= not w19796 and not w20497;
w20499 <= b(52) and not w19785;
w20500 <= not w19783 and w20499;
w20501 <= not w19787 and not w20500;
w20502 <= not w20498 and w20501;
w20503 <= not w19787 and not w20502;
w20504 <= not w19056 and not w19773;
w20505 <= not w19771 and w20504;
w20506 <= not w19762 and w20505;
w20507 <= not w19771 and not w19773;
w20508 <= not w19763 and not w20507;
w20509 <= not w20506 and not w20508;
w20510 <= not w19778 and not w20509;
w20511 <= not w19770 and not w19777;
w20512 <= not w19776 and w20511;
w20513 <= not w20510 and not w20512;
w20514 <= not b(53) and not w20513;
w20515 <= b(53) and not w20512;
w20516 <= not w20510 and w20515;
w20517 <= w26 and w28;
w20518 <= w23 and w20517;
w20519 <= not w20516 and w20518;
w20520 <= not w20514 and w20519;
w20521 <= not w20503 and w20520;
w20522 <= w338 and not w20513;
w20523 <= not w20521 and not w20522;
w20524 <= not w19796 and w20501;
w20525 <= not w20497 and w20524;
w20526 <= not w20498 and not w20501;
w20527 <= not w20525 and not w20526;
w20528 <= not w20523 and not w20527;
w20529 <= not w19786 and not w20522;
w20530 <= not w20521 and w20529;
w20531 <= not w20528 and not w20530;
w20532 <= not w19787 and not w20516;
w20533 <= not w20514 and w20532;
w20534 <= not w20502 and w20533;
w20535 <= not w20514 and not w20516;
w20536 <= not w20503 and not w20535;
w20537 <= not w20534 and not w20536;
w20538 <= not w20523 and not w20537;
w20539 <= not w20513 and not w20522;
w20540 <= not w20521 and w20539;
w20541 <= not w20538 and not w20540;
w20542 <= not b(54) and not w20541;
w20543 <= not b(53) and not w20531;
w20544 <= not w19805 and w20496;
w20545 <= not w20492 and w20544;
w20546 <= not w20493 and not w20496;
w20547 <= not w20545 and not w20546;
w20548 <= not w20523 and not w20547;
w20549 <= not w19795 and not w20522;
w20550 <= not w20521 and w20549;
w20551 <= not w20548 and not w20550;
w20552 <= not b(52) and not w20551;
w20553 <= not w19814 and w20491;
w20554 <= not w20487 and w20553;
w20555 <= not w20488 and not w20491;
w20556 <= not w20554 and not w20555;
w20557 <= not w20523 and not w20556;
w20558 <= not w19804 and not w20522;
w20559 <= not w20521 and w20558;
w20560 <= not w20557 and not w20559;
w20561 <= not b(51) and not w20560;
w20562 <= not w19823 and w20486;
w20563 <= not w20482 and w20562;
w20564 <= not w20483 and not w20486;
w20565 <= not w20563 and not w20564;
w20566 <= not w20523 and not w20565;
w20567 <= not w19813 and not w20522;
w20568 <= not w20521 and w20567;
w20569 <= not w20566 and not w20568;
w20570 <= not b(50) and not w20569;
w20571 <= not w19832 and w20481;
w20572 <= not w20477 and w20571;
w20573 <= not w20478 and not w20481;
w20574 <= not w20572 and not w20573;
w20575 <= not w20523 and not w20574;
w20576 <= not w19822 and not w20522;
w20577 <= not w20521 and w20576;
w20578 <= not w20575 and not w20577;
w20579 <= not b(49) and not w20578;
w20580 <= not w19841 and w20476;
w20581 <= not w20472 and w20580;
w20582 <= not w20473 and not w20476;
w20583 <= not w20581 and not w20582;
w20584 <= not w20523 and not w20583;
w20585 <= not w19831 and not w20522;
w20586 <= not w20521 and w20585;
w20587 <= not w20584 and not w20586;
w20588 <= not b(48) and not w20587;
w20589 <= not w19850 and w20471;
w20590 <= not w20467 and w20589;
w20591 <= not w20468 and not w20471;
w20592 <= not w20590 and not w20591;
w20593 <= not w20523 and not w20592;
w20594 <= not w19840 and not w20522;
w20595 <= not w20521 and w20594;
w20596 <= not w20593 and not w20595;
w20597 <= not b(47) and not w20596;
w20598 <= not w19859 and w20466;
w20599 <= not w20462 and w20598;
w20600 <= not w20463 and not w20466;
w20601 <= not w20599 and not w20600;
w20602 <= not w20523 and not w20601;
w20603 <= not w19849 and not w20522;
w20604 <= not w20521 and w20603;
w20605 <= not w20602 and not w20604;
w20606 <= not b(46) and not w20605;
w20607 <= not w19868 and w20461;
w20608 <= not w20457 and w20607;
w20609 <= not w20458 and not w20461;
w20610 <= not w20608 and not w20609;
w20611 <= not w20523 and not w20610;
w20612 <= not w19858 and not w20522;
w20613 <= not w20521 and w20612;
w20614 <= not w20611 and not w20613;
w20615 <= not b(45) and not w20614;
w20616 <= not w19877 and w20456;
w20617 <= not w20452 and w20616;
w20618 <= not w20453 and not w20456;
w20619 <= not w20617 and not w20618;
w20620 <= not w20523 and not w20619;
w20621 <= not w19867 and not w20522;
w20622 <= not w20521 and w20621;
w20623 <= not w20620 and not w20622;
w20624 <= not b(44) and not w20623;
w20625 <= not w19886 and w20451;
w20626 <= not w20447 and w20625;
w20627 <= not w20448 and not w20451;
w20628 <= not w20626 and not w20627;
w20629 <= not w20523 and not w20628;
w20630 <= not w19876 and not w20522;
w20631 <= not w20521 and w20630;
w20632 <= not w20629 and not w20631;
w20633 <= not b(43) and not w20632;
w20634 <= not w19895 and w20446;
w20635 <= not w20442 and w20634;
w20636 <= not w20443 and not w20446;
w20637 <= not w20635 and not w20636;
w20638 <= not w20523 and not w20637;
w20639 <= not w19885 and not w20522;
w20640 <= not w20521 and w20639;
w20641 <= not w20638 and not w20640;
w20642 <= not b(42) and not w20641;
w20643 <= not w19904 and w20441;
w20644 <= not w20437 and w20643;
w20645 <= not w20438 and not w20441;
w20646 <= not w20644 and not w20645;
w20647 <= not w20523 and not w20646;
w20648 <= not w19894 and not w20522;
w20649 <= not w20521 and w20648;
w20650 <= not w20647 and not w20649;
w20651 <= not b(41) and not w20650;
w20652 <= not w19913 and w20436;
w20653 <= not w20432 and w20652;
w20654 <= not w20433 and not w20436;
w20655 <= not w20653 and not w20654;
w20656 <= not w20523 and not w20655;
w20657 <= not w19903 and not w20522;
w20658 <= not w20521 and w20657;
w20659 <= not w20656 and not w20658;
w20660 <= not b(40) and not w20659;
w20661 <= not w19922 and w20431;
w20662 <= not w20427 and w20661;
w20663 <= not w20428 and not w20431;
w20664 <= not w20662 and not w20663;
w20665 <= not w20523 and not w20664;
w20666 <= not w19912 and not w20522;
w20667 <= not w20521 and w20666;
w20668 <= not w20665 and not w20667;
w20669 <= not b(39) and not w20668;
w20670 <= not w19931 and w20426;
w20671 <= not w20422 and w20670;
w20672 <= not w20423 and not w20426;
w20673 <= not w20671 and not w20672;
w20674 <= not w20523 and not w20673;
w20675 <= not w19921 and not w20522;
w20676 <= not w20521 and w20675;
w20677 <= not w20674 and not w20676;
w20678 <= not b(38) and not w20677;
w20679 <= not w19940 and w20421;
w20680 <= not w20417 and w20679;
w20681 <= not w20418 and not w20421;
w20682 <= not w20680 and not w20681;
w20683 <= not w20523 and not w20682;
w20684 <= not w19930 and not w20522;
w20685 <= not w20521 and w20684;
w20686 <= not w20683 and not w20685;
w20687 <= not b(37) and not w20686;
w20688 <= not w19949 and w20416;
w20689 <= not w20412 and w20688;
w20690 <= not w20413 and not w20416;
w20691 <= not w20689 and not w20690;
w20692 <= not w20523 and not w20691;
w20693 <= not w19939 and not w20522;
w20694 <= not w20521 and w20693;
w20695 <= not w20692 and not w20694;
w20696 <= not b(36) and not w20695;
w20697 <= not w19958 and w20411;
w20698 <= not w20407 and w20697;
w20699 <= not w20408 and not w20411;
w20700 <= not w20698 and not w20699;
w20701 <= not w20523 and not w20700;
w20702 <= not w19948 and not w20522;
w20703 <= not w20521 and w20702;
w20704 <= not w20701 and not w20703;
w20705 <= not b(35) and not w20704;
w20706 <= not w19967 and w20406;
w20707 <= not w20402 and w20706;
w20708 <= not w20403 and not w20406;
w20709 <= not w20707 and not w20708;
w20710 <= not w20523 and not w20709;
w20711 <= not w19957 and not w20522;
w20712 <= not w20521 and w20711;
w20713 <= not w20710 and not w20712;
w20714 <= not b(34) and not w20713;
w20715 <= not w19976 and w20401;
w20716 <= not w20397 and w20715;
w20717 <= not w20398 and not w20401;
w20718 <= not w20716 and not w20717;
w20719 <= not w20523 and not w20718;
w20720 <= not w19966 and not w20522;
w20721 <= not w20521 and w20720;
w20722 <= not w20719 and not w20721;
w20723 <= not b(33) and not w20722;
w20724 <= not w19985 and w20396;
w20725 <= not w20392 and w20724;
w20726 <= not w20393 and not w20396;
w20727 <= not w20725 and not w20726;
w20728 <= not w20523 and not w20727;
w20729 <= not w19975 and not w20522;
w20730 <= not w20521 and w20729;
w20731 <= not w20728 and not w20730;
w20732 <= not b(32) and not w20731;
w20733 <= not w19994 and w20391;
w20734 <= not w20387 and w20733;
w20735 <= not w20388 and not w20391;
w20736 <= not w20734 and not w20735;
w20737 <= not w20523 and not w20736;
w20738 <= not w19984 and not w20522;
w20739 <= not w20521 and w20738;
w20740 <= not w20737 and not w20739;
w20741 <= not b(31) and not w20740;
w20742 <= not w20003 and w20386;
w20743 <= not w20382 and w20742;
w20744 <= not w20383 and not w20386;
w20745 <= not w20743 and not w20744;
w20746 <= not w20523 and not w20745;
w20747 <= not w19993 and not w20522;
w20748 <= not w20521 and w20747;
w20749 <= not w20746 and not w20748;
w20750 <= not b(30) and not w20749;
w20751 <= not w20012 and w20381;
w20752 <= not w20377 and w20751;
w20753 <= not w20378 and not w20381;
w20754 <= not w20752 and not w20753;
w20755 <= not w20523 and not w20754;
w20756 <= not w20002 and not w20522;
w20757 <= not w20521 and w20756;
w20758 <= not w20755 and not w20757;
w20759 <= not b(29) and not w20758;
w20760 <= not w20021 and w20376;
w20761 <= not w20372 and w20760;
w20762 <= not w20373 and not w20376;
w20763 <= not w20761 and not w20762;
w20764 <= not w20523 and not w20763;
w20765 <= not w20011 and not w20522;
w20766 <= not w20521 and w20765;
w20767 <= not w20764 and not w20766;
w20768 <= not b(28) and not w20767;
w20769 <= not w20030 and w20371;
w20770 <= not w20367 and w20769;
w20771 <= not w20368 and not w20371;
w20772 <= not w20770 and not w20771;
w20773 <= not w20523 and not w20772;
w20774 <= not w20020 and not w20522;
w20775 <= not w20521 and w20774;
w20776 <= not w20773 and not w20775;
w20777 <= not b(27) and not w20776;
w20778 <= not w20039 and w20366;
w20779 <= not w20362 and w20778;
w20780 <= not w20363 and not w20366;
w20781 <= not w20779 and not w20780;
w20782 <= not w20523 and not w20781;
w20783 <= not w20029 and not w20522;
w20784 <= not w20521 and w20783;
w20785 <= not w20782 and not w20784;
w20786 <= not b(26) and not w20785;
w20787 <= not w20048 and w20361;
w20788 <= not w20357 and w20787;
w20789 <= not w20358 and not w20361;
w20790 <= not w20788 and not w20789;
w20791 <= not w20523 and not w20790;
w20792 <= not w20038 and not w20522;
w20793 <= not w20521 and w20792;
w20794 <= not w20791 and not w20793;
w20795 <= not b(25) and not w20794;
w20796 <= not w20057 and w20356;
w20797 <= not w20352 and w20796;
w20798 <= not w20353 and not w20356;
w20799 <= not w20797 and not w20798;
w20800 <= not w20523 and not w20799;
w20801 <= not w20047 and not w20522;
w20802 <= not w20521 and w20801;
w20803 <= not w20800 and not w20802;
w20804 <= not b(24) and not w20803;
w20805 <= not w20066 and w20351;
w20806 <= not w20347 and w20805;
w20807 <= not w20348 and not w20351;
w20808 <= not w20806 and not w20807;
w20809 <= not w20523 and not w20808;
w20810 <= not w20056 and not w20522;
w20811 <= not w20521 and w20810;
w20812 <= not w20809 and not w20811;
w20813 <= not b(23) and not w20812;
w20814 <= not w20075 and w20346;
w20815 <= not w20342 and w20814;
w20816 <= not w20343 and not w20346;
w20817 <= not w20815 and not w20816;
w20818 <= not w20523 and not w20817;
w20819 <= not w20065 and not w20522;
w20820 <= not w20521 and w20819;
w20821 <= not w20818 and not w20820;
w20822 <= not b(22) and not w20821;
w20823 <= not w20084 and w20341;
w20824 <= not w20337 and w20823;
w20825 <= not w20338 and not w20341;
w20826 <= not w20824 and not w20825;
w20827 <= not w20523 and not w20826;
w20828 <= not w20074 and not w20522;
w20829 <= not w20521 and w20828;
w20830 <= not w20827 and not w20829;
w20831 <= not b(21) and not w20830;
w20832 <= not w20093 and w20336;
w20833 <= not w20332 and w20832;
w20834 <= not w20333 and not w20336;
w20835 <= not w20833 and not w20834;
w20836 <= not w20523 and not w20835;
w20837 <= not w20083 and not w20522;
w20838 <= not w20521 and w20837;
w20839 <= not w20836 and not w20838;
w20840 <= not b(20) and not w20839;
w20841 <= not w20102 and w20331;
w20842 <= not w20327 and w20841;
w20843 <= not w20328 and not w20331;
w20844 <= not w20842 and not w20843;
w20845 <= not w20523 and not w20844;
w20846 <= not w20092 and not w20522;
w20847 <= not w20521 and w20846;
w20848 <= not w20845 and not w20847;
w20849 <= not b(19) and not w20848;
w20850 <= not w20111 and w20326;
w20851 <= not w20322 and w20850;
w20852 <= not w20323 and not w20326;
w20853 <= not w20851 and not w20852;
w20854 <= not w20523 and not w20853;
w20855 <= not w20101 and not w20522;
w20856 <= not w20521 and w20855;
w20857 <= not w20854 and not w20856;
w20858 <= not b(18) and not w20857;
w20859 <= not w20120 and w20321;
w20860 <= not w20317 and w20859;
w20861 <= not w20318 and not w20321;
w20862 <= not w20860 and not w20861;
w20863 <= not w20523 and not w20862;
w20864 <= not w20110 and not w20522;
w20865 <= not w20521 and w20864;
w20866 <= not w20863 and not w20865;
w20867 <= not b(17) and not w20866;
w20868 <= not w20129 and w20316;
w20869 <= not w20312 and w20868;
w20870 <= not w20313 and not w20316;
w20871 <= not w20869 and not w20870;
w20872 <= not w20523 and not w20871;
w20873 <= not w20119 and not w20522;
w20874 <= not w20521 and w20873;
w20875 <= not w20872 and not w20874;
w20876 <= not b(16) and not w20875;
w20877 <= not w20138 and w20311;
w20878 <= not w20307 and w20877;
w20879 <= not w20308 and not w20311;
w20880 <= not w20878 and not w20879;
w20881 <= not w20523 and not w20880;
w20882 <= not w20128 and not w20522;
w20883 <= not w20521 and w20882;
w20884 <= not w20881 and not w20883;
w20885 <= not b(15) and not w20884;
w20886 <= not w20147 and w20306;
w20887 <= not w20302 and w20886;
w20888 <= not w20303 and not w20306;
w20889 <= not w20887 and not w20888;
w20890 <= not w20523 and not w20889;
w20891 <= not w20137 and not w20522;
w20892 <= not w20521 and w20891;
w20893 <= not w20890 and not w20892;
w20894 <= not b(14) and not w20893;
w20895 <= not w20156 and w20301;
w20896 <= not w20297 and w20895;
w20897 <= not w20298 and not w20301;
w20898 <= not w20896 and not w20897;
w20899 <= not w20523 and not w20898;
w20900 <= not w20146 and not w20522;
w20901 <= not w20521 and w20900;
w20902 <= not w20899 and not w20901;
w20903 <= not b(13) and not w20902;
w20904 <= not w20165 and w20296;
w20905 <= not w20292 and w20904;
w20906 <= not w20293 and not w20296;
w20907 <= not w20905 and not w20906;
w20908 <= not w20523 and not w20907;
w20909 <= not w20155 and not w20522;
w20910 <= not w20521 and w20909;
w20911 <= not w20908 and not w20910;
w20912 <= not b(12) and not w20911;
w20913 <= not w20174 and w20291;
w20914 <= not w20287 and w20913;
w20915 <= not w20288 and not w20291;
w20916 <= not w20914 and not w20915;
w20917 <= not w20523 and not w20916;
w20918 <= not w20164 and not w20522;
w20919 <= not w20521 and w20918;
w20920 <= not w20917 and not w20919;
w20921 <= not b(11) and not w20920;
w20922 <= not w20183 and w20286;
w20923 <= not w20282 and w20922;
w20924 <= not w20283 and not w20286;
w20925 <= not w20923 and not w20924;
w20926 <= not w20523 and not w20925;
w20927 <= not w20173 and not w20522;
w20928 <= not w20521 and w20927;
w20929 <= not w20926 and not w20928;
w20930 <= not b(10) and not w20929;
w20931 <= not w20192 and w20281;
w20932 <= not w20277 and w20931;
w20933 <= not w20278 and not w20281;
w20934 <= not w20932 and not w20933;
w20935 <= not w20523 and not w20934;
w20936 <= not w20182 and not w20522;
w20937 <= not w20521 and w20936;
w20938 <= not w20935 and not w20937;
w20939 <= not b(9) and not w20938;
w20940 <= not w20201 and w20276;
w20941 <= not w20272 and w20940;
w20942 <= not w20273 and not w20276;
w20943 <= not w20941 and not w20942;
w20944 <= not w20523 and not w20943;
w20945 <= not w20191 and not w20522;
w20946 <= not w20521 and w20945;
w20947 <= not w20944 and not w20946;
w20948 <= not b(8) and not w20947;
w20949 <= not w20210 and w20271;
w20950 <= not w20267 and w20949;
w20951 <= not w20268 and not w20271;
w20952 <= not w20950 and not w20951;
w20953 <= not w20523 and not w20952;
w20954 <= not w20200 and not w20522;
w20955 <= not w20521 and w20954;
w20956 <= not w20953 and not w20955;
w20957 <= not b(7) and not w20956;
w20958 <= not w20219 and w20266;
w20959 <= not w20262 and w20958;
w20960 <= not w20263 and not w20266;
w20961 <= not w20959 and not w20960;
w20962 <= not w20523 and not w20961;
w20963 <= not w20209 and not w20522;
w20964 <= not w20521 and w20963;
w20965 <= not w20962 and not w20964;
w20966 <= not b(6) and not w20965;
w20967 <= not w20228 and w20261;
w20968 <= not w20257 and w20967;
w20969 <= not w20258 and not w20261;
w20970 <= not w20968 and not w20969;
w20971 <= not w20523 and not w20970;
w20972 <= not w20218 and not w20522;
w20973 <= not w20521 and w20972;
w20974 <= not w20971 and not w20973;
w20975 <= not b(5) and not w20974;
w20976 <= not w20236 and w20256;
w20977 <= not w20252 and w20976;
w20978 <= not w20253 and not w20256;
w20979 <= not w20977 and not w20978;
w20980 <= not w20523 and not w20979;
w20981 <= not w20227 and not w20522;
w20982 <= not w20521 and w20981;
w20983 <= not w20980 and not w20982;
w20984 <= not b(4) and not w20983;
w20985 <= not w20247 and w20251;
w20986 <= not w20246 and w20985;
w20987 <= not w20248 and not w20251;
w20988 <= not w20986 and not w20987;
w20989 <= not w20523 and not w20988;
w20990 <= not w20235 and not w20522;
w20991 <= not w20521 and w20990;
w20992 <= not w20989 and not w20991;
w20993 <= not b(3) and not w20992;
w20994 <= not w20243 and w20245;
w20995 <= not w20241 and w20994;
w20996 <= not w20246 and not w20995;
w20997 <= not w20523 and w20996;
w20998 <= not w20240 and not w20522;
w20999 <= not w20521 and w20998;
w21000 <= not w20997 and not w20999;
w21001 <= not b(2) and not w21000;
w21002 <= b(0) and not w20523;
w21003 <= a(10) and not w21002;
w21004 <= w20245 and not w20523;
w21005 <= not w21003 and not w21004;
w21006 <= b(1) and not w21005;
w21007 <= not b(1) and not w21004;
w21008 <= not w21003 and w21007;
w21009 <= not w21006 and not w21008;
w21010 <= not a(9) and b(0);
w21011 <= not w21009 and not w21010;
w21012 <= not b(1) and not w21005;
w21013 <= not w21011 and not w21012;
w21014 <= b(2) and not w20999;
w21015 <= not w20997 and w21014;
w21016 <= not w21001 and not w21015;
w21017 <= not w21013 and w21016;
w21018 <= not w21001 and not w21017;
w21019 <= b(3) and not w20991;
w21020 <= not w20989 and w21019;
w21021 <= not w20993 and not w21020;
w21022 <= not w21018 and w21021;
w21023 <= not w20993 and not w21022;
w21024 <= b(4) and not w20982;
w21025 <= not w20980 and w21024;
w21026 <= not w20984 and not w21025;
w21027 <= not w21023 and w21026;
w21028 <= not w20984 and not w21027;
w21029 <= b(5) and not w20973;
w21030 <= not w20971 and w21029;
w21031 <= not w20975 and not w21030;
w21032 <= not w21028 and w21031;
w21033 <= not w20975 and not w21032;
w21034 <= b(6) and not w20964;
w21035 <= not w20962 and w21034;
w21036 <= not w20966 and not w21035;
w21037 <= not w21033 and w21036;
w21038 <= not w20966 and not w21037;
w21039 <= b(7) and not w20955;
w21040 <= not w20953 and w21039;
w21041 <= not w20957 and not w21040;
w21042 <= not w21038 and w21041;
w21043 <= not w20957 and not w21042;
w21044 <= b(8) and not w20946;
w21045 <= not w20944 and w21044;
w21046 <= not w20948 and not w21045;
w21047 <= not w21043 and w21046;
w21048 <= not w20948 and not w21047;
w21049 <= b(9) and not w20937;
w21050 <= not w20935 and w21049;
w21051 <= not w20939 and not w21050;
w21052 <= not w21048 and w21051;
w21053 <= not w20939 and not w21052;
w21054 <= b(10) and not w20928;
w21055 <= not w20926 and w21054;
w21056 <= not w20930 and not w21055;
w21057 <= not w21053 and w21056;
w21058 <= not w20930 and not w21057;
w21059 <= b(11) and not w20919;
w21060 <= not w20917 and w21059;
w21061 <= not w20921 and not w21060;
w21062 <= not w21058 and w21061;
w21063 <= not w20921 and not w21062;
w21064 <= b(12) and not w20910;
w21065 <= not w20908 and w21064;
w21066 <= not w20912 and not w21065;
w21067 <= not w21063 and w21066;
w21068 <= not w20912 and not w21067;
w21069 <= b(13) and not w20901;
w21070 <= not w20899 and w21069;
w21071 <= not w20903 and not w21070;
w21072 <= not w21068 and w21071;
w21073 <= not w20903 and not w21072;
w21074 <= b(14) and not w20892;
w21075 <= not w20890 and w21074;
w21076 <= not w20894 and not w21075;
w21077 <= not w21073 and w21076;
w21078 <= not w20894 and not w21077;
w21079 <= b(15) and not w20883;
w21080 <= not w20881 and w21079;
w21081 <= not w20885 and not w21080;
w21082 <= not w21078 and w21081;
w21083 <= not w20885 and not w21082;
w21084 <= b(16) and not w20874;
w21085 <= not w20872 and w21084;
w21086 <= not w20876 and not w21085;
w21087 <= not w21083 and w21086;
w21088 <= not w20876 and not w21087;
w21089 <= b(17) and not w20865;
w21090 <= not w20863 and w21089;
w21091 <= not w20867 and not w21090;
w21092 <= not w21088 and w21091;
w21093 <= not w20867 and not w21092;
w21094 <= b(18) and not w20856;
w21095 <= not w20854 and w21094;
w21096 <= not w20858 and not w21095;
w21097 <= not w21093 and w21096;
w21098 <= not w20858 and not w21097;
w21099 <= b(19) and not w20847;
w21100 <= not w20845 and w21099;
w21101 <= not w20849 and not w21100;
w21102 <= not w21098 and w21101;
w21103 <= not w20849 and not w21102;
w21104 <= b(20) and not w20838;
w21105 <= not w20836 and w21104;
w21106 <= not w20840 and not w21105;
w21107 <= not w21103 and w21106;
w21108 <= not w20840 and not w21107;
w21109 <= b(21) and not w20829;
w21110 <= not w20827 and w21109;
w21111 <= not w20831 and not w21110;
w21112 <= not w21108 and w21111;
w21113 <= not w20831 and not w21112;
w21114 <= b(22) and not w20820;
w21115 <= not w20818 and w21114;
w21116 <= not w20822 and not w21115;
w21117 <= not w21113 and w21116;
w21118 <= not w20822 and not w21117;
w21119 <= b(23) and not w20811;
w21120 <= not w20809 and w21119;
w21121 <= not w20813 and not w21120;
w21122 <= not w21118 and w21121;
w21123 <= not w20813 and not w21122;
w21124 <= b(24) and not w20802;
w21125 <= not w20800 and w21124;
w21126 <= not w20804 and not w21125;
w21127 <= not w21123 and w21126;
w21128 <= not w20804 and not w21127;
w21129 <= b(25) and not w20793;
w21130 <= not w20791 and w21129;
w21131 <= not w20795 and not w21130;
w21132 <= not w21128 and w21131;
w21133 <= not w20795 and not w21132;
w21134 <= b(26) and not w20784;
w21135 <= not w20782 and w21134;
w21136 <= not w20786 and not w21135;
w21137 <= not w21133 and w21136;
w21138 <= not w20786 and not w21137;
w21139 <= b(27) and not w20775;
w21140 <= not w20773 and w21139;
w21141 <= not w20777 and not w21140;
w21142 <= not w21138 and w21141;
w21143 <= not w20777 and not w21142;
w21144 <= b(28) and not w20766;
w21145 <= not w20764 and w21144;
w21146 <= not w20768 and not w21145;
w21147 <= not w21143 and w21146;
w21148 <= not w20768 and not w21147;
w21149 <= b(29) and not w20757;
w21150 <= not w20755 and w21149;
w21151 <= not w20759 and not w21150;
w21152 <= not w21148 and w21151;
w21153 <= not w20759 and not w21152;
w21154 <= b(30) and not w20748;
w21155 <= not w20746 and w21154;
w21156 <= not w20750 and not w21155;
w21157 <= not w21153 and w21156;
w21158 <= not w20750 and not w21157;
w21159 <= b(31) and not w20739;
w21160 <= not w20737 and w21159;
w21161 <= not w20741 and not w21160;
w21162 <= not w21158 and w21161;
w21163 <= not w20741 and not w21162;
w21164 <= b(32) and not w20730;
w21165 <= not w20728 and w21164;
w21166 <= not w20732 and not w21165;
w21167 <= not w21163 and w21166;
w21168 <= not w20732 and not w21167;
w21169 <= b(33) and not w20721;
w21170 <= not w20719 and w21169;
w21171 <= not w20723 and not w21170;
w21172 <= not w21168 and w21171;
w21173 <= not w20723 and not w21172;
w21174 <= b(34) and not w20712;
w21175 <= not w20710 and w21174;
w21176 <= not w20714 and not w21175;
w21177 <= not w21173 and w21176;
w21178 <= not w20714 and not w21177;
w21179 <= b(35) and not w20703;
w21180 <= not w20701 and w21179;
w21181 <= not w20705 and not w21180;
w21182 <= not w21178 and w21181;
w21183 <= not w20705 and not w21182;
w21184 <= b(36) and not w20694;
w21185 <= not w20692 and w21184;
w21186 <= not w20696 and not w21185;
w21187 <= not w21183 and w21186;
w21188 <= not w20696 and not w21187;
w21189 <= b(37) and not w20685;
w21190 <= not w20683 and w21189;
w21191 <= not w20687 and not w21190;
w21192 <= not w21188 and w21191;
w21193 <= not w20687 and not w21192;
w21194 <= b(38) and not w20676;
w21195 <= not w20674 and w21194;
w21196 <= not w20678 and not w21195;
w21197 <= not w21193 and w21196;
w21198 <= not w20678 and not w21197;
w21199 <= b(39) and not w20667;
w21200 <= not w20665 and w21199;
w21201 <= not w20669 and not w21200;
w21202 <= not w21198 and w21201;
w21203 <= not w20669 and not w21202;
w21204 <= b(40) and not w20658;
w21205 <= not w20656 and w21204;
w21206 <= not w20660 and not w21205;
w21207 <= not w21203 and w21206;
w21208 <= not w20660 and not w21207;
w21209 <= b(41) and not w20649;
w21210 <= not w20647 and w21209;
w21211 <= not w20651 and not w21210;
w21212 <= not w21208 and w21211;
w21213 <= not w20651 and not w21212;
w21214 <= b(42) and not w20640;
w21215 <= not w20638 and w21214;
w21216 <= not w20642 and not w21215;
w21217 <= not w21213 and w21216;
w21218 <= not w20642 and not w21217;
w21219 <= b(43) and not w20631;
w21220 <= not w20629 and w21219;
w21221 <= not w20633 and not w21220;
w21222 <= not w21218 and w21221;
w21223 <= not w20633 and not w21222;
w21224 <= b(44) and not w20622;
w21225 <= not w20620 and w21224;
w21226 <= not w20624 and not w21225;
w21227 <= not w21223 and w21226;
w21228 <= not w20624 and not w21227;
w21229 <= b(45) and not w20613;
w21230 <= not w20611 and w21229;
w21231 <= not w20615 and not w21230;
w21232 <= not w21228 and w21231;
w21233 <= not w20615 and not w21232;
w21234 <= b(46) and not w20604;
w21235 <= not w20602 and w21234;
w21236 <= not w20606 and not w21235;
w21237 <= not w21233 and w21236;
w21238 <= not w20606 and not w21237;
w21239 <= b(47) and not w20595;
w21240 <= not w20593 and w21239;
w21241 <= not w20597 and not w21240;
w21242 <= not w21238 and w21241;
w21243 <= not w20597 and not w21242;
w21244 <= b(48) and not w20586;
w21245 <= not w20584 and w21244;
w21246 <= not w20588 and not w21245;
w21247 <= not w21243 and w21246;
w21248 <= not w20588 and not w21247;
w21249 <= b(49) and not w20577;
w21250 <= not w20575 and w21249;
w21251 <= not w20579 and not w21250;
w21252 <= not w21248 and w21251;
w21253 <= not w20579 and not w21252;
w21254 <= b(50) and not w20568;
w21255 <= not w20566 and w21254;
w21256 <= not w20570 and not w21255;
w21257 <= not w21253 and w21256;
w21258 <= not w20570 and not w21257;
w21259 <= b(51) and not w20559;
w21260 <= not w20557 and w21259;
w21261 <= not w20561 and not w21260;
w21262 <= not w21258 and w21261;
w21263 <= not w20561 and not w21262;
w21264 <= b(52) and not w20550;
w21265 <= not w20548 and w21264;
w21266 <= not w20552 and not w21265;
w21267 <= not w21263 and w21266;
w21268 <= not w20552 and not w21267;
w21269 <= b(53) and not w20530;
w21270 <= not w20528 and w21269;
w21271 <= not w20543 and not w21270;
w21272 <= not w21268 and w21271;
w21273 <= not w20543 and not w21272;
w21274 <= b(54) and not w20540;
w21275 <= not w20538 and w21274;
w21276 <= not w20542 and not w21275;
w21277 <= not w21273 and w21276;
w21278 <= not w20542 and not w21277;
w21279 <= w139 and w149;
w21280 <= w146 and w21279;
w21281 <= not w21278 and w21280;
w21282 <= not w20531 and not w21281;
w21283 <= not w20552 and w21271;
w21284 <= not w21267 and w21283;
w21285 <= not w21268 and not w21271;
w21286 <= not w21284 and not w21285;
w21287 <= w21280 and not w21286;
w21288 <= not w21278 and w21287;
w21289 <= not w21282 and not w21288;
w21290 <= not b(54) and not w21289;
w21291 <= not w20551 and not w21281;
w21292 <= not w20561 and w21266;
w21293 <= not w21262 and w21292;
w21294 <= not w21263 and not w21266;
w21295 <= not w21293 and not w21294;
w21296 <= w21280 and not w21295;
w21297 <= not w21278 and w21296;
w21298 <= not w21291 and not w21297;
w21299 <= not b(53) and not w21298;
w21300 <= not w20560 and not w21281;
w21301 <= not w20570 and w21261;
w21302 <= not w21257 and w21301;
w21303 <= not w21258 and not w21261;
w21304 <= not w21302 and not w21303;
w21305 <= w21280 and not w21304;
w21306 <= not w21278 and w21305;
w21307 <= not w21300 and not w21306;
w21308 <= not b(52) and not w21307;
w21309 <= not w20569 and not w21281;
w21310 <= not w20579 and w21256;
w21311 <= not w21252 and w21310;
w21312 <= not w21253 and not w21256;
w21313 <= not w21311 and not w21312;
w21314 <= w21280 and not w21313;
w21315 <= not w21278 and w21314;
w21316 <= not w21309 and not w21315;
w21317 <= not b(51) and not w21316;
w21318 <= not w20578 and not w21281;
w21319 <= not w20588 and w21251;
w21320 <= not w21247 and w21319;
w21321 <= not w21248 and not w21251;
w21322 <= not w21320 and not w21321;
w21323 <= w21280 and not w21322;
w21324 <= not w21278 and w21323;
w21325 <= not w21318 and not w21324;
w21326 <= not b(50) and not w21325;
w21327 <= not w20587 and not w21281;
w21328 <= not w20597 and w21246;
w21329 <= not w21242 and w21328;
w21330 <= not w21243 and not w21246;
w21331 <= not w21329 and not w21330;
w21332 <= w21280 and not w21331;
w21333 <= not w21278 and w21332;
w21334 <= not w21327 and not w21333;
w21335 <= not b(49) and not w21334;
w21336 <= not w20596 and not w21281;
w21337 <= not w20606 and w21241;
w21338 <= not w21237 and w21337;
w21339 <= not w21238 and not w21241;
w21340 <= not w21338 and not w21339;
w21341 <= w21280 and not w21340;
w21342 <= not w21278 and w21341;
w21343 <= not w21336 and not w21342;
w21344 <= not b(48) and not w21343;
w21345 <= not w20605 and not w21281;
w21346 <= not w20615 and w21236;
w21347 <= not w21232 and w21346;
w21348 <= not w21233 and not w21236;
w21349 <= not w21347 and not w21348;
w21350 <= w21280 and not w21349;
w21351 <= not w21278 and w21350;
w21352 <= not w21345 and not w21351;
w21353 <= not b(47) and not w21352;
w21354 <= not w20614 and not w21281;
w21355 <= not w20624 and w21231;
w21356 <= not w21227 and w21355;
w21357 <= not w21228 and not w21231;
w21358 <= not w21356 and not w21357;
w21359 <= w21280 and not w21358;
w21360 <= not w21278 and w21359;
w21361 <= not w21354 and not w21360;
w21362 <= not b(46) and not w21361;
w21363 <= not w20623 and not w21281;
w21364 <= not w20633 and w21226;
w21365 <= not w21222 and w21364;
w21366 <= not w21223 and not w21226;
w21367 <= not w21365 and not w21366;
w21368 <= w21280 and not w21367;
w21369 <= not w21278 and w21368;
w21370 <= not w21363 and not w21369;
w21371 <= not b(45) and not w21370;
w21372 <= not w20632 and not w21281;
w21373 <= not w20642 and w21221;
w21374 <= not w21217 and w21373;
w21375 <= not w21218 and not w21221;
w21376 <= not w21374 and not w21375;
w21377 <= w21280 and not w21376;
w21378 <= not w21278 and w21377;
w21379 <= not w21372 and not w21378;
w21380 <= not b(44) and not w21379;
w21381 <= not w20641 and not w21281;
w21382 <= not w20651 and w21216;
w21383 <= not w21212 and w21382;
w21384 <= not w21213 and not w21216;
w21385 <= not w21383 and not w21384;
w21386 <= w21280 and not w21385;
w21387 <= not w21278 and w21386;
w21388 <= not w21381 and not w21387;
w21389 <= not b(43) and not w21388;
w21390 <= not w20650 and not w21281;
w21391 <= not w20660 and w21211;
w21392 <= not w21207 and w21391;
w21393 <= not w21208 and not w21211;
w21394 <= not w21392 and not w21393;
w21395 <= w21280 and not w21394;
w21396 <= not w21278 and w21395;
w21397 <= not w21390 and not w21396;
w21398 <= not b(42) and not w21397;
w21399 <= not w20659 and not w21281;
w21400 <= not w20669 and w21206;
w21401 <= not w21202 and w21400;
w21402 <= not w21203 and not w21206;
w21403 <= not w21401 and not w21402;
w21404 <= w21280 and not w21403;
w21405 <= not w21278 and w21404;
w21406 <= not w21399 and not w21405;
w21407 <= not b(41) and not w21406;
w21408 <= not w20668 and not w21281;
w21409 <= not w20678 and w21201;
w21410 <= not w21197 and w21409;
w21411 <= not w21198 and not w21201;
w21412 <= not w21410 and not w21411;
w21413 <= w21280 and not w21412;
w21414 <= not w21278 and w21413;
w21415 <= not w21408 and not w21414;
w21416 <= not b(40) and not w21415;
w21417 <= not w20677 and not w21281;
w21418 <= not w20687 and w21196;
w21419 <= not w21192 and w21418;
w21420 <= not w21193 and not w21196;
w21421 <= not w21419 and not w21420;
w21422 <= w21280 and not w21421;
w21423 <= not w21278 and w21422;
w21424 <= not w21417 and not w21423;
w21425 <= not b(39) and not w21424;
w21426 <= not w20686 and not w21281;
w21427 <= not w20696 and w21191;
w21428 <= not w21187 and w21427;
w21429 <= not w21188 and not w21191;
w21430 <= not w21428 and not w21429;
w21431 <= w21280 and not w21430;
w21432 <= not w21278 and w21431;
w21433 <= not w21426 and not w21432;
w21434 <= not b(38) and not w21433;
w21435 <= not w20695 and not w21281;
w21436 <= not w20705 and w21186;
w21437 <= not w21182 and w21436;
w21438 <= not w21183 and not w21186;
w21439 <= not w21437 and not w21438;
w21440 <= w21280 and not w21439;
w21441 <= not w21278 and w21440;
w21442 <= not w21435 and not w21441;
w21443 <= not b(37) and not w21442;
w21444 <= not w20704 and not w21281;
w21445 <= not w20714 and w21181;
w21446 <= not w21177 and w21445;
w21447 <= not w21178 and not w21181;
w21448 <= not w21446 and not w21447;
w21449 <= w21280 and not w21448;
w21450 <= not w21278 and w21449;
w21451 <= not w21444 and not w21450;
w21452 <= not b(36) and not w21451;
w21453 <= not w20713 and not w21281;
w21454 <= not w20723 and w21176;
w21455 <= not w21172 and w21454;
w21456 <= not w21173 and not w21176;
w21457 <= not w21455 and not w21456;
w21458 <= w21280 and not w21457;
w21459 <= not w21278 and w21458;
w21460 <= not w21453 and not w21459;
w21461 <= not b(35) and not w21460;
w21462 <= not w20722 and not w21281;
w21463 <= not w20732 and w21171;
w21464 <= not w21167 and w21463;
w21465 <= not w21168 and not w21171;
w21466 <= not w21464 and not w21465;
w21467 <= w21280 and not w21466;
w21468 <= not w21278 and w21467;
w21469 <= not w21462 and not w21468;
w21470 <= not b(34) and not w21469;
w21471 <= not w20731 and not w21281;
w21472 <= not w20741 and w21166;
w21473 <= not w21162 and w21472;
w21474 <= not w21163 and not w21166;
w21475 <= not w21473 and not w21474;
w21476 <= w21280 and not w21475;
w21477 <= not w21278 and w21476;
w21478 <= not w21471 and not w21477;
w21479 <= not b(33) and not w21478;
w21480 <= not w20740 and not w21281;
w21481 <= not w20750 and w21161;
w21482 <= not w21157 and w21481;
w21483 <= not w21158 and not w21161;
w21484 <= not w21482 and not w21483;
w21485 <= w21280 and not w21484;
w21486 <= not w21278 and w21485;
w21487 <= not w21480 and not w21486;
w21488 <= not b(32) and not w21487;
w21489 <= not w20749 and not w21281;
w21490 <= not w20759 and w21156;
w21491 <= not w21152 and w21490;
w21492 <= not w21153 and not w21156;
w21493 <= not w21491 and not w21492;
w21494 <= w21280 and not w21493;
w21495 <= not w21278 and w21494;
w21496 <= not w21489 and not w21495;
w21497 <= not b(31) and not w21496;
w21498 <= not w20758 and not w21281;
w21499 <= not w20768 and w21151;
w21500 <= not w21147 and w21499;
w21501 <= not w21148 and not w21151;
w21502 <= not w21500 and not w21501;
w21503 <= w21280 and not w21502;
w21504 <= not w21278 and w21503;
w21505 <= not w21498 and not w21504;
w21506 <= not b(30) and not w21505;
w21507 <= not w20767 and not w21281;
w21508 <= not w20777 and w21146;
w21509 <= not w21142 and w21508;
w21510 <= not w21143 and not w21146;
w21511 <= not w21509 and not w21510;
w21512 <= w21280 and not w21511;
w21513 <= not w21278 and w21512;
w21514 <= not w21507 and not w21513;
w21515 <= not b(29) and not w21514;
w21516 <= not w20776 and not w21281;
w21517 <= not w20786 and w21141;
w21518 <= not w21137 and w21517;
w21519 <= not w21138 and not w21141;
w21520 <= not w21518 and not w21519;
w21521 <= w21280 and not w21520;
w21522 <= not w21278 and w21521;
w21523 <= not w21516 and not w21522;
w21524 <= not b(28) and not w21523;
w21525 <= not w20785 and not w21281;
w21526 <= not w20795 and w21136;
w21527 <= not w21132 and w21526;
w21528 <= not w21133 and not w21136;
w21529 <= not w21527 and not w21528;
w21530 <= w21280 and not w21529;
w21531 <= not w21278 and w21530;
w21532 <= not w21525 and not w21531;
w21533 <= not b(27) and not w21532;
w21534 <= not w20794 and not w21281;
w21535 <= not w20804 and w21131;
w21536 <= not w21127 and w21535;
w21537 <= not w21128 and not w21131;
w21538 <= not w21536 and not w21537;
w21539 <= w21280 and not w21538;
w21540 <= not w21278 and w21539;
w21541 <= not w21534 and not w21540;
w21542 <= not b(26) and not w21541;
w21543 <= not w20803 and not w21281;
w21544 <= not w20813 and w21126;
w21545 <= not w21122 and w21544;
w21546 <= not w21123 and not w21126;
w21547 <= not w21545 and not w21546;
w21548 <= w21280 and not w21547;
w21549 <= not w21278 and w21548;
w21550 <= not w21543 and not w21549;
w21551 <= not b(25) and not w21550;
w21552 <= not w20812 and not w21281;
w21553 <= not w20822 and w21121;
w21554 <= not w21117 and w21553;
w21555 <= not w21118 and not w21121;
w21556 <= not w21554 and not w21555;
w21557 <= w21280 and not w21556;
w21558 <= not w21278 and w21557;
w21559 <= not w21552 and not w21558;
w21560 <= not b(24) and not w21559;
w21561 <= not w20821 and not w21281;
w21562 <= not w20831 and w21116;
w21563 <= not w21112 and w21562;
w21564 <= not w21113 and not w21116;
w21565 <= not w21563 and not w21564;
w21566 <= w21280 and not w21565;
w21567 <= not w21278 and w21566;
w21568 <= not w21561 and not w21567;
w21569 <= not b(23) and not w21568;
w21570 <= not w20830 and not w21281;
w21571 <= not w20840 and w21111;
w21572 <= not w21107 and w21571;
w21573 <= not w21108 and not w21111;
w21574 <= not w21572 and not w21573;
w21575 <= w21280 and not w21574;
w21576 <= not w21278 and w21575;
w21577 <= not w21570 and not w21576;
w21578 <= not b(22) and not w21577;
w21579 <= not w20839 and not w21281;
w21580 <= not w20849 and w21106;
w21581 <= not w21102 and w21580;
w21582 <= not w21103 and not w21106;
w21583 <= not w21581 and not w21582;
w21584 <= w21280 and not w21583;
w21585 <= not w21278 and w21584;
w21586 <= not w21579 and not w21585;
w21587 <= not b(21) and not w21586;
w21588 <= not w20848 and not w21281;
w21589 <= not w20858 and w21101;
w21590 <= not w21097 and w21589;
w21591 <= not w21098 and not w21101;
w21592 <= not w21590 and not w21591;
w21593 <= w21280 and not w21592;
w21594 <= not w21278 and w21593;
w21595 <= not w21588 and not w21594;
w21596 <= not b(20) and not w21595;
w21597 <= not w20857 and not w21281;
w21598 <= not w20867 and w21096;
w21599 <= not w21092 and w21598;
w21600 <= not w21093 and not w21096;
w21601 <= not w21599 and not w21600;
w21602 <= w21280 and not w21601;
w21603 <= not w21278 and w21602;
w21604 <= not w21597 and not w21603;
w21605 <= not b(19) and not w21604;
w21606 <= not w20866 and not w21281;
w21607 <= not w20876 and w21091;
w21608 <= not w21087 and w21607;
w21609 <= not w21088 and not w21091;
w21610 <= not w21608 and not w21609;
w21611 <= w21280 and not w21610;
w21612 <= not w21278 and w21611;
w21613 <= not w21606 and not w21612;
w21614 <= not b(18) and not w21613;
w21615 <= not w20875 and not w21281;
w21616 <= not w20885 and w21086;
w21617 <= not w21082 and w21616;
w21618 <= not w21083 and not w21086;
w21619 <= not w21617 and not w21618;
w21620 <= w21280 and not w21619;
w21621 <= not w21278 and w21620;
w21622 <= not w21615 and not w21621;
w21623 <= not b(17) and not w21622;
w21624 <= not w20884 and not w21281;
w21625 <= not w20894 and w21081;
w21626 <= not w21077 and w21625;
w21627 <= not w21078 and not w21081;
w21628 <= not w21626 and not w21627;
w21629 <= w21280 and not w21628;
w21630 <= not w21278 and w21629;
w21631 <= not w21624 and not w21630;
w21632 <= not b(16) and not w21631;
w21633 <= not w20893 and not w21281;
w21634 <= not w20903 and w21076;
w21635 <= not w21072 and w21634;
w21636 <= not w21073 and not w21076;
w21637 <= not w21635 and not w21636;
w21638 <= w21280 and not w21637;
w21639 <= not w21278 and w21638;
w21640 <= not w21633 and not w21639;
w21641 <= not b(15) and not w21640;
w21642 <= not w20902 and not w21281;
w21643 <= not w20912 and w21071;
w21644 <= not w21067 and w21643;
w21645 <= not w21068 and not w21071;
w21646 <= not w21644 and not w21645;
w21647 <= w21280 and not w21646;
w21648 <= not w21278 and w21647;
w21649 <= not w21642 and not w21648;
w21650 <= not b(14) and not w21649;
w21651 <= not w20911 and not w21281;
w21652 <= not w20921 and w21066;
w21653 <= not w21062 and w21652;
w21654 <= not w21063 and not w21066;
w21655 <= not w21653 and not w21654;
w21656 <= w21280 and not w21655;
w21657 <= not w21278 and w21656;
w21658 <= not w21651 and not w21657;
w21659 <= not b(13) and not w21658;
w21660 <= not w20920 and not w21281;
w21661 <= not w20930 and w21061;
w21662 <= not w21057 and w21661;
w21663 <= not w21058 and not w21061;
w21664 <= not w21662 and not w21663;
w21665 <= w21280 and not w21664;
w21666 <= not w21278 and w21665;
w21667 <= not w21660 and not w21666;
w21668 <= not b(12) and not w21667;
w21669 <= not w20929 and not w21281;
w21670 <= not w20939 and w21056;
w21671 <= not w21052 and w21670;
w21672 <= not w21053 and not w21056;
w21673 <= not w21671 and not w21672;
w21674 <= w21280 and not w21673;
w21675 <= not w21278 and w21674;
w21676 <= not w21669 and not w21675;
w21677 <= not b(11) and not w21676;
w21678 <= not w20938 and not w21281;
w21679 <= not w20948 and w21051;
w21680 <= not w21047 and w21679;
w21681 <= not w21048 and not w21051;
w21682 <= not w21680 and not w21681;
w21683 <= w21280 and not w21682;
w21684 <= not w21278 and w21683;
w21685 <= not w21678 and not w21684;
w21686 <= not b(10) and not w21685;
w21687 <= not w20947 and not w21281;
w21688 <= not w20957 and w21046;
w21689 <= not w21042 and w21688;
w21690 <= not w21043 and not w21046;
w21691 <= not w21689 and not w21690;
w21692 <= w21280 and not w21691;
w21693 <= not w21278 and w21692;
w21694 <= not w21687 and not w21693;
w21695 <= not b(9) and not w21694;
w21696 <= not w20956 and not w21281;
w21697 <= not w20966 and w21041;
w21698 <= not w21037 and w21697;
w21699 <= not w21038 and not w21041;
w21700 <= not w21698 and not w21699;
w21701 <= w21280 and not w21700;
w21702 <= not w21278 and w21701;
w21703 <= not w21696 and not w21702;
w21704 <= not b(8) and not w21703;
w21705 <= not w20965 and not w21281;
w21706 <= not w20975 and w21036;
w21707 <= not w21032 and w21706;
w21708 <= not w21033 and not w21036;
w21709 <= not w21707 and not w21708;
w21710 <= w21280 and not w21709;
w21711 <= not w21278 and w21710;
w21712 <= not w21705 and not w21711;
w21713 <= not b(7) and not w21712;
w21714 <= not w20974 and not w21281;
w21715 <= not w20984 and w21031;
w21716 <= not w21027 and w21715;
w21717 <= not w21028 and not w21031;
w21718 <= not w21716 and not w21717;
w21719 <= w21280 and not w21718;
w21720 <= not w21278 and w21719;
w21721 <= not w21714 and not w21720;
w21722 <= not b(6) and not w21721;
w21723 <= not w20983 and not w21281;
w21724 <= not w20993 and w21026;
w21725 <= not w21022 and w21724;
w21726 <= not w21023 and not w21026;
w21727 <= not w21725 and not w21726;
w21728 <= w21280 and not w21727;
w21729 <= not w21278 and w21728;
w21730 <= not w21723 and not w21729;
w21731 <= not b(5) and not w21730;
w21732 <= not w20992 and not w21281;
w21733 <= not w21001 and w21021;
w21734 <= not w21017 and w21733;
w21735 <= not w21018 and not w21021;
w21736 <= not w21734 and not w21735;
w21737 <= w21280 and not w21736;
w21738 <= not w21278 and w21737;
w21739 <= not w21732 and not w21738;
w21740 <= not b(4) and not w21739;
w21741 <= not w21000 and not w21281;
w21742 <= not w21012 and w21016;
w21743 <= not w21011 and w21742;
w21744 <= not w21013 and not w21016;
w21745 <= not w21743 and not w21744;
w21746 <= w21280 and not w21745;
w21747 <= not w21278 and w21746;
w21748 <= not w21741 and not w21747;
w21749 <= not b(3) and not w21748;
w21750 <= not w21005 and not w21281;
w21751 <= not w21008 and w21010;
w21752 <= not w21006 and w21751;
w21753 <= w21280 and not w21752;
w21754 <= not w21011 and w21753;
w21755 <= not w21278 and w21754;
w21756 <= not w21750 and not w21755;
w21757 <= not b(2) and not w21756;
w21758 <= b(0) and not b(55);
w21759 <= w26 and w21758;
w21760 <= w23 and w21759;
w21761 <= not w21278 and w21760;
w21762 <= a(9) and not w21761;
w21763 <= w139 and w21010;
w21764 <= w149 and w21763;
w21765 <= w146 and w21764;
w21766 <= not w21278 and w21765;
w21767 <= not w21762 and not w21766;
w21768 <= b(1) and not w21767;
w21769 <= not b(1) and not w21766;
w21770 <= not w21762 and w21769;
w21771 <= not w21768 and not w21770;
w21772 <= not a(8) and b(0);
w21773 <= not w21771 and not w21772;
w21774 <= not b(1) and not w21767;
w21775 <= not w21773 and not w21774;
w21776 <= b(2) and not w21755;
w21777 <= not w21750 and w21776;
w21778 <= not w21757 and not w21777;
w21779 <= not w21775 and w21778;
w21780 <= not w21757 and not w21779;
w21781 <= b(3) and not w21747;
w21782 <= not w21741 and w21781;
w21783 <= not w21749 and not w21782;
w21784 <= not w21780 and w21783;
w21785 <= not w21749 and not w21784;
w21786 <= b(4) and not w21738;
w21787 <= not w21732 and w21786;
w21788 <= not w21740 and not w21787;
w21789 <= not w21785 and w21788;
w21790 <= not w21740 and not w21789;
w21791 <= b(5) and not w21729;
w21792 <= not w21723 and w21791;
w21793 <= not w21731 and not w21792;
w21794 <= not w21790 and w21793;
w21795 <= not w21731 and not w21794;
w21796 <= b(6) and not w21720;
w21797 <= not w21714 and w21796;
w21798 <= not w21722 and not w21797;
w21799 <= not w21795 and w21798;
w21800 <= not w21722 and not w21799;
w21801 <= b(7) and not w21711;
w21802 <= not w21705 and w21801;
w21803 <= not w21713 and not w21802;
w21804 <= not w21800 and w21803;
w21805 <= not w21713 and not w21804;
w21806 <= b(8) and not w21702;
w21807 <= not w21696 and w21806;
w21808 <= not w21704 and not w21807;
w21809 <= not w21805 and w21808;
w21810 <= not w21704 and not w21809;
w21811 <= b(9) and not w21693;
w21812 <= not w21687 and w21811;
w21813 <= not w21695 and not w21812;
w21814 <= not w21810 and w21813;
w21815 <= not w21695 and not w21814;
w21816 <= b(10) and not w21684;
w21817 <= not w21678 and w21816;
w21818 <= not w21686 and not w21817;
w21819 <= not w21815 and w21818;
w21820 <= not w21686 and not w21819;
w21821 <= b(11) and not w21675;
w21822 <= not w21669 and w21821;
w21823 <= not w21677 and not w21822;
w21824 <= not w21820 and w21823;
w21825 <= not w21677 and not w21824;
w21826 <= b(12) and not w21666;
w21827 <= not w21660 and w21826;
w21828 <= not w21668 and not w21827;
w21829 <= not w21825 and w21828;
w21830 <= not w21668 and not w21829;
w21831 <= b(13) and not w21657;
w21832 <= not w21651 and w21831;
w21833 <= not w21659 and not w21832;
w21834 <= not w21830 and w21833;
w21835 <= not w21659 and not w21834;
w21836 <= b(14) and not w21648;
w21837 <= not w21642 and w21836;
w21838 <= not w21650 and not w21837;
w21839 <= not w21835 and w21838;
w21840 <= not w21650 and not w21839;
w21841 <= b(15) and not w21639;
w21842 <= not w21633 and w21841;
w21843 <= not w21641 and not w21842;
w21844 <= not w21840 and w21843;
w21845 <= not w21641 and not w21844;
w21846 <= b(16) and not w21630;
w21847 <= not w21624 and w21846;
w21848 <= not w21632 and not w21847;
w21849 <= not w21845 and w21848;
w21850 <= not w21632 and not w21849;
w21851 <= b(17) and not w21621;
w21852 <= not w21615 and w21851;
w21853 <= not w21623 and not w21852;
w21854 <= not w21850 and w21853;
w21855 <= not w21623 and not w21854;
w21856 <= b(18) and not w21612;
w21857 <= not w21606 and w21856;
w21858 <= not w21614 and not w21857;
w21859 <= not w21855 and w21858;
w21860 <= not w21614 and not w21859;
w21861 <= b(19) and not w21603;
w21862 <= not w21597 and w21861;
w21863 <= not w21605 and not w21862;
w21864 <= not w21860 and w21863;
w21865 <= not w21605 and not w21864;
w21866 <= b(20) and not w21594;
w21867 <= not w21588 and w21866;
w21868 <= not w21596 and not w21867;
w21869 <= not w21865 and w21868;
w21870 <= not w21596 and not w21869;
w21871 <= b(21) and not w21585;
w21872 <= not w21579 and w21871;
w21873 <= not w21587 and not w21872;
w21874 <= not w21870 and w21873;
w21875 <= not w21587 and not w21874;
w21876 <= b(22) and not w21576;
w21877 <= not w21570 and w21876;
w21878 <= not w21578 and not w21877;
w21879 <= not w21875 and w21878;
w21880 <= not w21578 and not w21879;
w21881 <= b(23) and not w21567;
w21882 <= not w21561 and w21881;
w21883 <= not w21569 and not w21882;
w21884 <= not w21880 and w21883;
w21885 <= not w21569 and not w21884;
w21886 <= b(24) and not w21558;
w21887 <= not w21552 and w21886;
w21888 <= not w21560 and not w21887;
w21889 <= not w21885 and w21888;
w21890 <= not w21560 and not w21889;
w21891 <= b(25) and not w21549;
w21892 <= not w21543 and w21891;
w21893 <= not w21551 and not w21892;
w21894 <= not w21890 and w21893;
w21895 <= not w21551 and not w21894;
w21896 <= b(26) and not w21540;
w21897 <= not w21534 and w21896;
w21898 <= not w21542 and not w21897;
w21899 <= not w21895 and w21898;
w21900 <= not w21542 and not w21899;
w21901 <= b(27) and not w21531;
w21902 <= not w21525 and w21901;
w21903 <= not w21533 and not w21902;
w21904 <= not w21900 and w21903;
w21905 <= not w21533 and not w21904;
w21906 <= b(28) and not w21522;
w21907 <= not w21516 and w21906;
w21908 <= not w21524 and not w21907;
w21909 <= not w21905 and w21908;
w21910 <= not w21524 and not w21909;
w21911 <= b(29) and not w21513;
w21912 <= not w21507 and w21911;
w21913 <= not w21515 and not w21912;
w21914 <= not w21910 and w21913;
w21915 <= not w21515 and not w21914;
w21916 <= b(30) and not w21504;
w21917 <= not w21498 and w21916;
w21918 <= not w21506 and not w21917;
w21919 <= not w21915 and w21918;
w21920 <= not w21506 and not w21919;
w21921 <= b(31) and not w21495;
w21922 <= not w21489 and w21921;
w21923 <= not w21497 and not w21922;
w21924 <= not w21920 and w21923;
w21925 <= not w21497 and not w21924;
w21926 <= b(32) and not w21486;
w21927 <= not w21480 and w21926;
w21928 <= not w21488 and not w21927;
w21929 <= not w21925 and w21928;
w21930 <= not w21488 and not w21929;
w21931 <= b(33) and not w21477;
w21932 <= not w21471 and w21931;
w21933 <= not w21479 and not w21932;
w21934 <= not w21930 and w21933;
w21935 <= not w21479 and not w21934;
w21936 <= b(34) and not w21468;
w21937 <= not w21462 and w21936;
w21938 <= not w21470 and not w21937;
w21939 <= not w21935 and w21938;
w21940 <= not w21470 and not w21939;
w21941 <= b(35) and not w21459;
w21942 <= not w21453 and w21941;
w21943 <= not w21461 and not w21942;
w21944 <= not w21940 and w21943;
w21945 <= not w21461 and not w21944;
w21946 <= b(36) and not w21450;
w21947 <= not w21444 and w21946;
w21948 <= not w21452 and not w21947;
w21949 <= not w21945 and w21948;
w21950 <= not w21452 and not w21949;
w21951 <= b(37) and not w21441;
w21952 <= not w21435 and w21951;
w21953 <= not w21443 and not w21952;
w21954 <= not w21950 and w21953;
w21955 <= not w21443 and not w21954;
w21956 <= b(38) and not w21432;
w21957 <= not w21426 and w21956;
w21958 <= not w21434 and not w21957;
w21959 <= not w21955 and w21958;
w21960 <= not w21434 and not w21959;
w21961 <= b(39) and not w21423;
w21962 <= not w21417 and w21961;
w21963 <= not w21425 and not w21962;
w21964 <= not w21960 and w21963;
w21965 <= not w21425 and not w21964;
w21966 <= b(40) and not w21414;
w21967 <= not w21408 and w21966;
w21968 <= not w21416 and not w21967;
w21969 <= not w21965 and w21968;
w21970 <= not w21416 and not w21969;
w21971 <= b(41) and not w21405;
w21972 <= not w21399 and w21971;
w21973 <= not w21407 and not w21972;
w21974 <= not w21970 and w21973;
w21975 <= not w21407 and not w21974;
w21976 <= b(42) and not w21396;
w21977 <= not w21390 and w21976;
w21978 <= not w21398 and not w21977;
w21979 <= not w21975 and w21978;
w21980 <= not w21398 and not w21979;
w21981 <= b(43) and not w21387;
w21982 <= not w21381 and w21981;
w21983 <= not w21389 and not w21982;
w21984 <= not w21980 and w21983;
w21985 <= not w21389 and not w21984;
w21986 <= b(44) and not w21378;
w21987 <= not w21372 and w21986;
w21988 <= not w21380 and not w21987;
w21989 <= not w21985 and w21988;
w21990 <= not w21380 and not w21989;
w21991 <= b(45) and not w21369;
w21992 <= not w21363 and w21991;
w21993 <= not w21371 and not w21992;
w21994 <= not w21990 and w21993;
w21995 <= not w21371 and not w21994;
w21996 <= b(46) and not w21360;
w21997 <= not w21354 and w21996;
w21998 <= not w21362 and not w21997;
w21999 <= not w21995 and w21998;
w22000 <= not w21362 and not w21999;
w22001 <= b(47) and not w21351;
w22002 <= not w21345 and w22001;
w22003 <= not w21353 and not w22002;
w22004 <= not w22000 and w22003;
w22005 <= not w21353 and not w22004;
w22006 <= b(48) and not w21342;
w22007 <= not w21336 and w22006;
w22008 <= not w21344 and not w22007;
w22009 <= not w22005 and w22008;
w22010 <= not w21344 and not w22009;
w22011 <= b(49) and not w21333;
w22012 <= not w21327 and w22011;
w22013 <= not w21335 and not w22012;
w22014 <= not w22010 and w22013;
w22015 <= not w21335 and not w22014;
w22016 <= b(50) and not w21324;
w22017 <= not w21318 and w22016;
w22018 <= not w21326 and not w22017;
w22019 <= not w22015 and w22018;
w22020 <= not w21326 and not w22019;
w22021 <= b(51) and not w21315;
w22022 <= not w21309 and w22021;
w22023 <= not w21317 and not w22022;
w22024 <= not w22020 and w22023;
w22025 <= not w21317 and not w22024;
w22026 <= b(52) and not w21306;
w22027 <= not w21300 and w22026;
w22028 <= not w21308 and not w22027;
w22029 <= not w22025 and w22028;
w22030 <= not w21308 and not w22029;
w22031 <= b(53) and not w21297;
w22032 <= not w21291 and w22031;
w22033 <= not w21299 and not w22032;
w22034 <= not w22030 and w22033;
w22035 <= not w21299 and not w22034;
w22036 <= b(54) and not w21288;
w22037 <= not w21282 and w22036;
w22038 <= not w21290 and not w22037;
w22039 <= not w22035 and w22038;
w22040 <= not w21290 and not w22039;
w22041 <= not w20541 and not w21281;
w22042 <= not w20543 and w21276;
w22043 <= not w21272 and w22042;
w22044 <= not w21273 and not w21276;
w22045 <= not w22043 and not w22044;
w22046 <= w21281 and not w22045;
w22047 <= not w22041 and not w22046;
w22048 <= not b(55) and not w22047;
w22049 <= b(55) and not w22041;
w22050 <= not w22046 and w22049;
w22051 <= w80 and not w22050;
w22052 <= not w22048 and w22051;
w22053 <= not w22040 and w22052;
w22054 <= w21280 and not w22047;
w22055 <= not w22053 and not w22054;
w22056 <= not w21299 and w22038;
w22057 <= not w22034 and w22056;
w22058 <= not w22035 and not w22038;
w22059 <= not w22057 and not w22058;
w22060 <= not w22055 and not w22059;
w22061 <= not w21289 and not w22054;
w22062 <= not w22053 and w22061;
w22063 <= not w22060 and not w22062;
w22064 <= not b(55) and not w22063;
w22065 <= not w21308 and w22033;
w22066 <= not w22029 and w22065;
w22067 <= not w22030 and not w22033;
w22068 <= not w22066 and not w22067;
w22069 <= not w22055 and not w22068;
w22070 <= not w21298 and not w22054;
w22071 <= not w22053 and w22070;
w22072 <= not w22069 and not w22071;
w22073 <= not b(54) and not w22072;
w22074 <= not w21317 and w22028;
w22075 <= not w22024 and w22074;
w22076 <= not w22025 and not w22028;
w22077 <= not w22075 and not w22076;
w22078 <= not w22055 and not w22077;
w22079 <= not w21307 and not w22054;
w22080 <= not w22053 and w22079;
w22081 <= not w22078 and not w22080;
w22082 <= not b(53) and not w22081;
w22083 <= not w21326 and w22023;
w22084 <= not w22019 and w22083;
w22085 <= not w22020 and not w22023;
w22086 <= not w22084 and not w22085;
w22087 <= not w22055 and not w22086;
w22088 <= not w21316 and not w22054;
w22089 <= not w22053 and w22088;
w22090 <= not w22087 and not w22089;
w22091 <= not b(52) and not w22090;
w22092 <= not w21335 and w22018;
w22093 <= not w22014 and w22092;
w22094 <= not w22015 and not w22018;
w22095 <= not w22093 and not w22094;
w22096 <= not w22055 and not w22095;
w22097 <= not w21325 and not w22054;
w22098 <= not w22053 and w22097;
w22099 <= not w22096 and not w22098;
w22100 <= not b(51) and not w22099;
w22101 <= not w21344 and w22013;
w22102 <= not w22009 and w22101;
w22103 <= not w22010 and not w22013;
w22104 <= not w22102 and not w22103;
w22105 <= not w22055 and not w22104;
w22106 <= not w21334 and not w22054;
w22107 <= not w22053 and w22106;
w22108 <= not w22105 and not w22107;
w22109 <= not b(50) and not w22108;
w22110 <= not w21353 and w22008;
w22111 <= not w22004 and w22110;
w22112 <= not w22005 and not w22008;
w22113 <= not w22111 and not w22112;
w22114 <= not w22055 and not w22113;
w22115 <= not w21343 and not w22054;
w22116 <= not w22053 and w22115;
w22117 <= not w22114 and not w22116;
w22118 <= not b(49) and not w22117;
w22119 <= not w21362 and w22003;
w22120 <= not w21999 and w22119;
w22121 <= not w22000 and not w22003;
w22122 <= not w22120 and not w22121;
w22123 <= not w22055 and not w22122;
w22124 <= not w21352 and not w22054;
w22125 <= not w22053 and w22124;
w22126 <= not w22123 and not w22125;
w22127 <= not b(48) and not w22126;
w22128 <= not w21371 and w21998;
w22129 <= not w21994 and w22128;
w22130 <= not w21995 and not w21998;
w22131 <= not w22129 and not w22130;
w22132 <= not w22055 and not w22131;
w22133 <= not w21361 and not w22054;
w22134 <= not w22053 and w22133;
w22135 <= not w22132 and not w22134;
w22136 <= not b(47) and not w22135;
w22137 <= not w21380 and w21993;
w22138 <= not w21989 and w22137;
w22139 <= not w21990 and not w21993;
w22140 <= not w22138 and not w22139;
w22141 <= not w22055 and not w22140;
w22142 <= not w21370 and not w22054;
w22143 <= not w22053 and w22142;
w22144 <= not w22141 and not w22143;
w22145 <= not b(46) and not w22144;
w22146 <= not w21389 and w21988;
w22147 <= not w21984 and w22146;
w22148 <= not w21985 and not w21988;
w22149 <= not w22147 and not w22148;
w22150 <= not w22055 and not w22149;
w22151 <= not w21379 and not w22054;
w22152 <= not w22053 and w22151;
w22153 <= not w22150 and not w22152;
w22154 <= not b(45) and not w22153;
w22155 <= not w21398 and w21983;
w22156 <= not w21979 and w22155;
w22157 <= not w21980 and not w21983;
w22158 <= not w22156 and not w22157;
w22159 <= not w22055 and not w22158;
w22160 <= not w21388 and not w22054;
w22161 <= not w22053 and w22160;
w22162 <= not w22159 and not w22161;
w22163 <= not b(44) and not w22162;
w22164 <= not w21407 and w21978;
w22165 <= not w21974 and w22164;
w22166 <= not w21975 and not w21978;
w22167 <= not w22165 and not w22166;
w22168 <= not w22055 and not w22167;
w22169 <= not w21397 and not w22054;
w22170 <= not w22053 and w22169;
w22171 <= not w22168 and not w22170;
w22172 <= not b(43) and not w22171;
w22173 <= not w21416 and w21973;
w22174 <= not w21969 and w22173;
w22175 <= not w21970 and not w21973;
w22176 <= not w22174 and not w22175;
w22177 <= not w22055 and not w22176;
w22178 <= not w21406 and not w22054;
w22179 <= not w22053 and w22178;
w22180 <= not w22177 and not w22179;
w22181 <= not b(42) and not w22180;
w22182 <= not w21425 and w21968;
w22183 <= not w21964 and w22182;
w22184 <= not w21965 and not w21968;
w22185 <= not w22183 and not w22184;
w22186 <= not w22055 and not w22185;
w22187 <= not w21415 and not w22054;
w22188 <= not w22053 and w22187;
w22189 <= not w22186 and not w22188;
w22190 <= not b(41) and not w22189;
w22191 <= not w21434 and w21963;
w22192 <= not w21959 and w22191;
w22193 <= not w21960 and not w21963;
w22194 <= not w22192 and not w22193;
w22195 <= not w22055 and not w22194;
w22196 <= not w21424 and not w22054;
w22197 <= not w22053 and w22196;
w22198 <= not w22195 and not w22197;
w22199 <= not b(40) and not w22198;
w22200 <= not w21443 and w21958;
w22201 <= not w21954 and w22200;
w22202 <= not w21955 and not w21958;
w22203 <= not w22201 and not w22202;
w22204 <= not w22055 and not w22203;
w22205 <= not w21433 and not w22054;
w22206 <= not w22053 and w22205;
w22207 <= not w22204 and not w22206;
w22208 <= not b(39) and not w22207;
w22209 <= not w21452 and w21953;
w22210 <= not w21949 and w22209;
w22211 <= not w21950 and not w21953;
w22212 <= not w22210 and not w22211;
w22213 <= not w22055 and not w22212;
w22214 <= not w21442 and not w22054;
w22215 <= not w22053 and w22214;
w22216 <= not w22213 and not w22215;
w22217 <= not b(38) and not w22216;
w22218 <= not w21461 and w21948;
w22219 <= not w21944 and w22218;
w22220 <= not w21945 and not w21948;
w22221 <= not w22219 and not w22220;
w22222 <= not w22055 and not w22221;
w22223 <= not w21451 and not w22054;
w22224 <= not w22053 and w22223;
w22225 <= not w22222 and not w22224;
w22226 <= not b(37) and not w22225;
w22227 <= not w21470 and w21943;
w22228 <= not w21939 and w22227;
w22229 <= not w21940 and not w21943;
w22230 <= not w22228 and not w22229;
w22231 <= not w22055 and not w22230;
w22232 <= not w21460 and not w22054;
w22233 <= not w22053 and w22232;
w22234 <= not w22231 and not w22233;
w22235 <= not b(36) and not w22234;
w22236 <= not w21479 and w21938;
w22237 <= not w21934 and w22236;
w22238 <= not w21935 and not w21938;
w22239 <= not w22237 and not w22238;
w22240 <= not w22055 and not w22239;
w22241 <= not w21469 and not w22054;
w22242 <= not w22053 and w22241;
w22243 <= not w22240 and not w22242;
w22244 <= not b(35) and not w22243;
w22245 <= not w21488 and w21933;
w22246 <= not w21929 and w22245;
w22247 <= not w21930 and not w21933;
w22248 <= not w22246 and not w22247;
w22249 <= not w22055 and not w22248;
w22250 <= not w21478 and not w22054;
w22251 <= not w22053 and w22250;
w22252 <= not w22249 and not w22251;
w22253 <= not b(34) and not w22252;
w22254 <= not w21497 and w21928;
w22255 <= not w21924 and w22254;
w22256 <= not w21925 and not w21928;
w22257 <= not w22255 and not w22256;
w22258 <= not w22055 and not w22257;
w22259 <= not w21487 and not w22054;
w22260 <= not w22053 and w22259;
w22261 <= not w22258 and not w22260;
w22262 <= not b(33) and not w22261;
w22263 <= not w21506 and w21923;
w22264 <= not w21919 and w22263;
w22265 <= not w21920 and not w21923;
w22266 <= not w22264 and not w22265;
w22267 <= not w22055 and not w22266;
w22268 <= not w21496 and not w22054;
w22269 <= not w22053 and w22268;
w22270 <= not w22267 and not w22269;
w22271 <= not b(32) and not w22270;
w22272 <= not w21515 and w21918;
w22273 <= not w21914 and w22272;
w22274 <= not w21915 and not w21918;
w22275 <= not w22273 and not w22274;
w22276 <= not w22055 and not w22275;
w22277 <= not w21505 and not w22054;
w22278 <= not w22053 and w22277;
w22279 <= not w22276 and not w22278;
w22280 <= not b(31) and not w22279;
w22281 <= not w21524 and w21913;
w22282 <= not w21909 and w22281;
w22283 <= not w21910 and not w21913;
w22284 <= not w22282 and not w22283;
w22285 <= not w22055 and not w22284;
w22286 <= not w21514 and not w22054;
w22287 <= not w22053 and w22286;
w22288 <= not w22285 and not w22287;
w22289 <= not b(30) and not w22288;
w22290 <= not w21533 and w21908;
w22291 <= not w21904 and w22290;
w22292 <= not w21905 and not w21908;
w22293 <= not w22291 and not w22292;
w22294 <= not w22055 and not w22293;
w22295 <= not w21523 and not w22054;
w22296 <= not w22053 and w22295;
w22297 <= not w22294 and not w22296;
w22298 <= not b(29) and not w22297;
w22299 <= not w21542 and w21903;
w22300 <= not w21899 and w22299;
w22301 <= not w21900 and not w21903;
w22302 <= not w22300 and not w22301;
w22303 <= not w22055 and not w22302;
w22304 <= not w21532 and not w22054;
w22305 <= not w22053 and w22304;
w22306 <= not w22303 and not w22305;
w22307 <= not b(28) and not w22306;
w22308 <= not w21551 and w21898;
w22309 <= not w21894 and w22308;
w22310 <= not w21895 and not w21898;
w22311 <= not w22309 and not w22310;
w22312 <= not w22055 and not w22311;
w22313 <= not w21541 and not w22054;
w22314 <= not w22053 and w22313;
w22315 <= not w22312 and not w22314;
w22316 <= not b(27) and not w22315;
w22317 <= not w21560 and w21893;
w22318 <= not w21889 and w22317;
w22319 <= not w21890 and not w21893;
w22320 <= not w22318 and not w22319;
w22321 <= not w22055 and not w22320;
w22322 <= not w21550 and not w22054;
w22323 <= not w22053 and w22322;
w22324 <= not w22321 and not w22323;
w22325 <= not b(26) and not w22324;
w22326 <= not w21569 and w21888;
w22327 <= not w21884 and w22326;
w22328 <= not w21885 and not w21888;
w22329 <= not w22327 and not w22328;
w22330 <= not w22055 and not w22329;
w22331 <= not w21559 and not w22054;
w22332 <= not w22053 and w22331;
w22333 <= not w22330 and not w22332;
w22334 <= not b(25) and not w22333;
w22335 <= not w21578 and w21883;
w22336 <= not w21879 and w22335;
w22337 <= not w21880 and not w21883;
w22338 <= not w22336 and not w22337;
w22339 <= not w22055 and not w22338;
w22340 <= not w21568 and not w22054;
w22341 <= not w22053 and w22340;
w22342 <= not w22339 and not w22341;
w22343 <= not b(24) and not w22342;
w22344 <= not w21587 and w21878;
w22345 <= not w21874 and w22344;
w22346 <= not w21875 and not w21878;
w22347 <= not w22345 and not w22346;
w22348 <= not w22055 and not w22347;
w22349 <= not w21577 and not w22054;
w22350 <= not w22053 and w22349;
w22351 <= not w22348 and not w22350;
w22352 <= not b(23) and not w22351;
w22353 <= not w21596 and w21873;
w22354 <= not w21869 and w22353;
w22355 <= not w21870 and not w21873;
w22356 <= not w22354 and not w22355;
w22357 <= not w22055 and not w22356;
w22358 <= not w21586 and not w22054;
w22359 <= not w22053 and w22358;
w22360 <= not w22357 and not w22359;
w22361 <= not b(22) and not w22360;
w22362 <= not w21605 and w21868;
w22363 <= not w21864 and w22362;
w22364 <= not w21865 and not w21868;
w22365 <= not w22363 and not w22364;
w22366 <= not w22055 and not w22365;
w22367 <= not w21595 and not w22054;
w22368 <= not w22053 and w22367;
w22369 <= not w22366 and not w22368;
w22370 <= not b(21) and not w22369;
w22371 <= not w21614 and w21863;
w22372 <= not w21859 and w22371;
w22373 <= not w21860 and not w21863;
w22374 <= not w22372 and not w22373;
w22375 <= not w22055 and not w22374;
w22376 <= not w21604 and not w22054;
w22377 <= not w22053 and w22376;
w22378 <= not w22375 and not w22377;
w22379 <= not b(20) and not w22378;
w22380 <= not w21623 and w21858;
w22381 <= not w21854 and w22380;
w22382 <= not w21855 and not w21858;
w22383 <= not w22381 and not w22382;
w22384 <= not w22055 and not w22383;
w22385 <= not w21613 and not w22054;
w22386 <= not w22053 and w22385;
w22387 <= not w22384 and not w22386;
w22388 <= not b(19) and not w22387;
w22389 <= not w21632 and w21853;
w22390 <= not w21849 and w22389;
w22391 <= not w21850 and not w21853;
w22392 <= not w22390 and not w22391;
w22393 <= not w22055 and not w22392;
w22394 <= not w21622 and not w22054;
w22395 <= not w22053 and w22394;
w22396 <= not w22393 and not w22395;
w22397 <= not b(18) and not w22396;
w22398 <= not w21641 and w21848;
w22399 <= not w21844 and w22398;
w22400 <= not w21845 and not w21848;
w22401 <= not w22399 and not w22400;
w22402 <= not w22055 and not w22401;
w22403 <= not w21631 and not w22054;
w22404 <= not w22053 and w22403;
w22405 <= not w22402 and not w22404;
w22406 <= not b(17) and not w22405;
w22407 <= not w21650 and w21843;
w22408 <= not w21839 and w22407;
w22409 <= not w21840 and not w21843;
w22410 <= not w22408 and not w22409;
w22411 <= not w22055 and not w22410;
w22412 <= not w21640 and not w22054;
w22413 <= not w22053 and w22412;
w22414 <= not w22411 and not w22413;
w22415 <= not b(16) and not w22414;
w22416 <= not w21659 and w21838;
w22417 <= not w21834 and w22416;
w22418 <= not w21835 and not w21838;
w22419 <= not w22417 and not w22418;
w22420 <= not w22055 and not w22419;
w22421 <= not w21649 and not w22054;
w22422 <= not w22053 and w22421;
w22423 <= not w22420 and not w22422;
w22424 <= not b(15) and not w22423;
w22425 <= not w21668 and w21833;
w22426 <= not w21829 and w22425;
w22427 <= not w21830 and not w21833;
w22428 <= not w22426 and not w22427;
w22429 <= not w22055 and not w22428;
w22430 <= not w21658 and not w22054;
w22431 <= not w22053 and w22430;
w22432 <= not w22429 and not w22431;
w22433 <= not b(14) and not w22432;
w22434 <= not w21677 and w21828;
w22435 <= not w21824 and w22434;
w22436 <= not w21825 and not w21828;
w22437 <= not w22435 and not w22436;
w22438 <= not w22055 and not w22437;
w22439 <= not w21667 and not w22054;
w22440 <= not w22053 and w22439;
w22441 <= not w22438 and not w22440;
w22442 <= not b(13) and not w22441;
w22443 <= not w21686 and w21823;
w22444 <= not w21819 and w22443;
w22445 <= not w21820 and not w21823;
w22446 <= not w22444 and not w22445;
w22447 <= not w22055 and not w22446;
w22448 <= not w21676 and not w22054;
w22449 <= not w22053 and w22448;
w22450 <= not w22447 and not w22449;
w22451 <= not b(12) and not w22450;
w22452 <= not w21695 and w21818;
w22453 <= not w21814 and w22452;
w22454 <= not w21815 and not w21818;
w22455 <= not w22453 and not w22454;
w22456 <= not w22055 and not w22455;
w22457 <= not w21685 and not w22054;
w22458 <= not w22053 and w22457;
w22459 <= not w22456 and not w22458;
w22460 <= not b(11) and not w22459;
w22461 <= not w21704 and w21813;
w22462 <= not w21809 and w22461;
w22463 <= not w21810 and not w21813;
w22464 <= not w22462 and not w22463;
w22465 <= not w22055 and not w22464;
w22466 <= not w21694 and not w22054;
w22467 <= not w22053 and w22466;
w22468 <= not w22465 and not w22467;
w22469 <= not b(10) and not w22468;
w22470 <= not w21713 and w21808;
w22471 <= not w21804 and w22470;
w22472 <= not w21805 and not w21808;
w22473 <= not w22471 and not w22472;
w22474 <= not w22055 and not w22473;
w22475 <= not w21703 and not w22054;
w22476 <= not w22053 and w22475;
w22477 <= not w22474 and not w22476;
w22478 <= not b(9) and not w22477;
w22479 <= not w21722 and w21803;
w22480 <= not w21799 and w22479;
w22481 <= not w21800 and not w21803;
w22482 <= not w22480 and not w22481;
w22483 <= not w22055 and not w22482;
w22484 <= not w21712 and not w22054;
w22485 <= not w22053 and w22484;
w22486 <= not w22483 and not w22485;
w22487 <= not b(8) and not w22486;
w22488 <= not w21731 and w21798;
w22489 <= not w21794 and w22488;
w22490 <= not w21795 and not w21798;
w22491 <= not w22489 and not w22490;
w22492 <= not w22055 and not w22491;
w22493 <= not w21721 and not w22054;
w22494 <= not w22053 and w22493;
w22495 <= not w22492 and not w22494;
w22496 <= not b(7) and not w22495;
w22497 <= not w21740 and w21793;
w22498 <= not w21789 and w22497;
w22499 <= not w21790 and not w21793;
w22500 <= not w22498 and not w22499;
w22501 <= not w22055 and not w22500;
w22502 <= not w21730 and not w22054;
w22503 <= not w22053 and w22502;
w22504 <= not w22501 and not w22503;
w22505 <= not b(6) and not w22504;
w22506 <= not w21749 and w21788;
w22507 <= not w21784 and w22506;
w22508 <= not w21785 and not w21788;
w22509 <= not w22507 and not w22508;
w22510 <= not w22055 and not w22509;
w22511 <= not w21739 and not w22054;
w22512 <= not w22053 and w22511;
w22513 <= not w22510 and not w22512;
w22514 <= not b(5) and not w22513;
w22515 <= not w21757 and w21783;
w22516 <= not w21779 and w22515;
w22517 <= not w21780 and not w21783;
w22518 <= not w22516 and not w22517;
w22519 <= not w22055 and not w22518;
w22520 <= not w21748 and not w22054;
w22521 <= not w22053 and w22520;
w22522 <= not w22519 and not w22521;
w22523 <= not b(4) and not w22522;
w22524 <= not w21774 and w21778;
w22525 <= not w21773 and w22524;
w22526 <= not w21775 and not w21778;
w22527 <= not w22525 and not w22526;
w22528 <= not w22055 and not w22527;
w22529 <= not w21756 and not w22054;
w22530 <= not w22053 and w22529;
w22531 <= not w22528 and not w22530;
w22532 <= not b(3) and not w22531;
w22533 <= not w21770 and w21772;
w22534 <= not w21768 and w22533;
w22535 <= not w21773 and not w22534;
w22536 <= not w22055 and w22535;
w22537 <= not w21767 and not w22054;
w22538 <= not w22053 and w22537;
w22539 <= not w22536 and not w22538;
w22540 <= not b(2) and not w22539;
w22541 <= b(0) and not w22055;
w22542 <= a(8) and not w22541;
w22543 <= w21772 and not w22055;
w22544 <= not w22542 and not w22543;
w22545 <= b(1) and not w22544;
w22546 <= not b(1) and not w22543;
w22547 <= not w22542 and w22546;
w22548 <= not w22545 and not w22547;
w22549 <= not a(7) and b(0);
w22550 <= not w22548 and not w22549;
w22551 <= not b(1) and not w22544;
w22552 <= not w22550 and not w22551;
w22553 <= b(2) and not w22538;
w22554 <= not w22536 and w22553;
w22555 <= not w22540 and not w22554;
w22556 <= not w22552 and w22555;
w22557 <= not w22540 and not w22556;
w22558 <= b(3) and not w22530;
w22559 <= not w22528 and w22558;
w22560 <= not w22532 and not w22559;
w22561 <= not w22557 and w22560;
w22562 <= not w22532 and not w22561;
w22563 <= b(4) and not w22521;
w22564 <= not w22519 and w22563;
w22565 <= not w22523 and not w22564;
w22566 <= not w22562 and w22565;
w22567 <= not w22523 and not w22566;
w22568 <= b(5) and not w22512;
w22569 <= not w22510 and w22568;
w22570 <= not w22514 and not w22569;
w22571 <= not w22567 and w22570;
w22572 <= not w22514 and not w22571;
w22573 <= b(6) and not w22503;
w22574 <= not w22501 and w22573;
w22575 <= not w22505 and not w22574;
w22576 <= not w22572 and w22575;
w22577 <= not w22505 and not w22576;
w22578 <= b(7) and not w22494;
w22579 <= not w22492 and w22578;
w22580 <= not w22496 and not w22579;
w22581 <= not w22577 and w22580;
w22582 <= not w22496 and not w22581;
w22583 <= b(8) and not w22485;
w22584 <= not w22483 and w22583;
w22585 <= not w22487 and not w22584;
w22586 <= not w22582 and w22585;
w22587 <= not w22487 and not w22586;
w22588 <= b(9) and not w22476;
w22589 <= not w22474 and w22588;
w22590 <= not w22478 and not w22589;
w22591 <= not w22587 and w22590;
w22592 <= not w22478 and not w22591;
w22593 <= b(10) and not w22467;
w22594 <= not w22465 and w22593;
w22595 <= not w22469 and not w22594;
w22596 <= not w22592 and w22595;
w22597 <= not w22469 and not w22596;
w22598 <= b(11) and not w22458;
w22599 <= not w22456 and w22598;
w22600 <= not w22460 and not w22599;
w22601 <= not w22597 and w22600;
w22602 <= not w22460 and not w22601;
w22603 <= b(12) and not w22449;
w22604 <= not w22447 and w22603;
w22605 <= not w22451 and not w22604;
w22606 <= not w22602 and w22605;
w22607 <= not w22451 and not w22606;
w22608 <= b(13) and not w22440;
w22609 <= not w22438 and w22608;
w22610 <= not w22442 and not w22609;
w22611 <= not w22607 and w22610;
w22612 <= not w22442 and not w22611;
w22613 <= b(14) and not w22431;
w22614 <= not w22429 and w22613;
w22615 <= not w22433 and not w22614;
w22616 <= not w22612 and w22615;
w22617 <= not w22433 and not w22616;
w22618 <= b(15) and not w22422;
w22619 <= not w22420 and w22618;
w22620 <= not w22424 and not w22619;
w22621 <= not w22617 and w22620;
w22622 <= not w22424 and not w22621;
w22623 <= b(16) and not w22413;
w22624 <= not w22411 and w22623;
w22625 <= not w22415 and not w22624;
w22626 <= not w22622 and w22625;
w22627 <= not w22415 and not w22626;
w22628 <= b(17) and not w22404;
w22629 <= not w22402 and w22628;
w22630 <= not w22406 and not w22629;
w22631 <= not w22627 and w22630;
w22632 <= not w22406 and not w22631;
w22633 <= b(18) and not w22395;
w22634 <= not w22393 and w22633;
w22635 <= not w22397 and not w22634;
w22636 <= not w22632 and w22635;
w22637 <= not w22397 and not w22636;
w22638 <= b(19) and not w22386;
w22639 <= not w22384 and w22638;
w22640 <= not w22388 and not w22639;
w22641 <= not w22637 and w22640;
w22642 <= not w22388 and not w22641;
w22643 <= b(20) and not w22377;
w22644 <= not w22375 and w22643;
w22645 <= not w22379 and not w22644;
w22646 <= not w22642 and w22645;
w22647 <= not w22379 and not w22646;
w22648 <= b(21) and not w22368;
w22649 <= not w22366 and w22648;
w22650 <= not w22370 and not w22649;
w22651 <= not w22647 and w22650;
w22652 <= not w22370 and not w22651;
w22653 <= b(22) and not w22359;
w22654 <= not w22357 and w22653;
w22655 <= not w22361 and not w22654;
w22656 <= not w22652 and w22655;
w22657 <= not w22361 and not w22656;
w22658 <= b(23) and not w22350;
w22659 <= not w22348 and w22658;
w22660 <= not w22352 and not w22659;
w22661 <= not w22657 and w22660;
w22662 <= not w22352 and not w22661;
w22663 <= b(24) and not w22341;
w22664 <= not w22339 and w22663;
w22665 <= not w22343 and not w22664;
w22666 <= not w22662 and w22665;
w22667 <= not w22343 and not w22666;
w22668 <= b(25) and not w22332;
w22669 <= not w22330 and w22668;
w22670 <= not w22334 and not w22669;
w22671 <= not w22667 and w22670;
w22672 <= not w22334 and not w22671;
w22673 <= b(26) and not w22323;
w22674 <= not w22321 and w22673;
w22675 <= not w22325 and not w22674;
w22676 <= not w22672 and w22675;
w22677 <= not w22325 and not w22676;
w22678 <= b(27) and not w22314;
w22679 <= not w22312 and w22678;
w22680 <= not w22316 and not w22679;
w22681 <= not w22677 and w22680;
w22682 <= not w22316 and not w22681;
w22683 <= b(28) and not w22305;
w22684 <= not w22303 and w22683;
w22685 <= not w22307 and not w22684;
w22686 <= not w22682 and w22685;
w22687 <= not w22307 and not w22686;
w22688 <= b(29) and not w22296;
w22689 <= not w22294 and w22688;
w22690 <= not w22298 and not w22689;
w22691 <= not w22687 and w22690;
w22692 <= not w22298 and not w22691;
w22693 <= b(30) and not w22287;
w22694 <= not w22285 and w22693;
w22695 <= not w22289 and not w22694;
w22696 <= not w22692 and w22695;
w22697 <= not w22289 and not w22696;
w22698 <= b(31) and not w22278;
w22699 <= not w22276 and w22698;
w22700 <= not w22280 and not w22699;
w22701 <= not w22697 and w22700;
w22702 <= not w22280 and not w22701;
w22703 <= b(32) and not w22269;
w22704 <= not w22267 and w22703;
w22705 <= not w22271 and not w22704;
w22706 <= not w22702 and w22705;
w22707 <= not w22271 and not w22706;
w22708 <= b(33) and not w22260;
w22709 <= not w22258 and w22708;
w22710 <= not w22262 and not w22709;
w22711 <= not w22707 and w22710;
w22712 <= not w22262 and not w22711;
w22713 <= b(34) and not w22251;
w22714 <= not w22249 and w22713;
w22715 <= not w22253 and not w22714;
w22716 <= not w22712 and w22715;
w22717 <= not w22253 and not w22716;
w22718 <= b(35) and not w22242;
w22719 <= not w22240 and w22718;
w22720 <= not w22244 and not w22719;
w22721 <= not w22717 and w22720;
w22722 <= not w22244 and not w22721;
w22723 <= b(36) and not w22233;
w22724 <= not w22231 and w22723;
w22725 <= not w22235 and not w22724;
w22726 <= not w22722 and w22725;
w22727 <= not w22235 and not w22726;
w22728 <= b(37) and not w22224;
w22729 <= not w22222 and w22728;
w22730 <= not w22226 and not w22729;
w22731 <= not w22727 and w22730;
w22732 <= not w22226 and not w22731;
w22733 <= b(38) and not w22215;
w22734 <= not w22213 and w22733;
w22735 <= not w22217 and not w22734;
w22736 <= not w22732 and w22735;
w22737 <= not w22217 and not w22736;
w22738 <= b(39) and not w22206;
w22739 <= not w22204 and w22738;
w22740 <= not w22208 and not w22739;
w22741 <= not w22737 and w22740;
w22742 <= not w22208 and not w22741;
w22743 <= b(40) and not w22197;
w22744 <= not w22195 and w22743;
w22745 <= not w22199 and not w22744;
w22746 <= not w22742 and w22745;
w22747 <= not w22199 and not w22746;
w22748 <= b(41) and not w22188;
w22749 <= not w22186 and w22748;
w22750 <= not w22190 and not w22749;
w22751 <= not w22747 and w22750;
w22752 <= not w22190 and not w22751;
w22753 <= b(42) and not w22179;
w22754 <= not w22177 and w22753;
w22755 <= not w22181 and not w22754;
w22756 <= not w22752 and w22755;
w22757 <= not w22181 and not w22756;
w22758 <= b(43) and not w22170;
w22759 <= not w22168 and w22758;
w22760 <= not w22172 and not w22759;
w22761 <= not w22757 and w22760;
w22762 <= not w22172 and not w22761;
w22763 <= b(44) and not w22161;
w22764 <= not w22159 and w22763;
w22765 <= not w22163 and not w22764;
w22766 <= not w22762 and w22765;
w22767 <= not w22163 and not w22766;
w22768 <= b(45) and not w22152;
w22769 <= not w22150 and w22768;
w22770 <= not w22154 and not w22769;
w22771 <= not w22767 and w22770;
w22772 <= not w22154 and not w22771;
w22773 <= b(46) and not w22143;
w22774 <= not w22141 and w22773;
w22775 <= not w22145 and not w22774;
w22776 <= not w22772 and w22775;
w22777 <= not w22145 and not w22776;
w22778 <= b(47) and not w22134;
w22779 <= not w22132 and w22778;
w22780 <= not w22136 and not w22779;
w22781 <= not w22777 and w22780;
w22782 <= not w22136 and not w22781;
w22783 <= b(48) and not w22125;
w22784 <= not w22123 and w22783;
w22785 <= not w22127 and not w22784;
w22786 <= not w22782 and w22785;
w22787 <= not w22127 and not w22786;
w22788 <= b(49) and not w22116;
w22789 <= not w22114 and w22788;
w22790 <= not w22118 and not w22789;
w22791 <= not w22787 and w22790;
w22792 <= not w22118 and not w22791;
w22793 <= b(50) and not w22107;
w22794 <= not w22105 and w22793;
w22795 <= not w22109 and not w22794;
w22796 <= not w22792 and w22795;
w22797 <= not w22109 and not w22796;
w22798 <= b(51) and not w22098;
w22799 <= not w22096 and w22798;
w22800 <= not w22100 and not w22799;
w22801 <= not w22797 and w22800;
w22802 <= not w22100 and not w22801;
w22803 <= b(52) and not w22089;
w22804 <= not w22087 and w22803;
w22805 <= not w22091 and not w22804;
w22806 <= not w22802 and w22805;
w22807 <= not w22091 and not w22806;
w22808 <= b(53) and not w22080;
w22809 <= not w22078 and w22808;
w22810 <= not w22082 and not w22809;
w22811 <= not w22807 and w22810;
w22812 <= not w22082 and not w22811;
w22813 <= b(54) and not w22071;
w22814 <= not w22069 and w22813;
w22815 <= not w22073 and not w22814;
w22816 <= not w22812 and w22815;
w22817 <= not w22073 and not w22816;
w22818 <= b(55) and not w22062;
w22819 <= not w22060 and w22818;
w22820 <= not w22064 and not w22819;
w22821 <= not w22817 and w22820;
w22822 <= not w22064 and not w22821;
w22823 <= not w21290 and not w22050;
w22824 <= not w22048 and w22823;
w22825 <= not w22039 and w22824;
w22826 <= not w22048 and not w22050;
w22827 <= not w22040 and not w22826;
w22828 <= not w22825 and not w22827;
w22829 <= not w22055 and not w22828;
w22830 <= not w22047 and not w22054;
w22831 <= not w22053 and w22830;
w22832 <= not w22829 and not w22831;
w22833 <= not b(56) and not w22832;
w22834 <= b(56) and not w22831;
w22835 <= not w22829 and w22834;
w22836 <= w150 and not w22835;
w22837 <= not w22833 and w22836;
w22838 <= not w22822 and w22837;
w22839 <= w80 and not w22832;
w22840 <= not w22838 and not w22839;
w22841 <= not w22073 and w22820;
w22842 <= not w22816 and w22841;
w22843 <= not w22817 and not w22820;
w22844 <= not w22842 and not w22843;
w22845 <= not w22840 and not w22844;
w22846 <= not w22063 and not w22839;
w22847 <= not w22838 and w22846;
w22848 <= not w22845 and not w22847;
w22849 <= not w22064 and not w22835;
w22850 <= not w22833 and w22849;
w22851 <= not w22821 and w22850;
w22852 <= not w22833 and not w22835;
w22853 <= not w22822 and not w22852;
w22854 <= not w22851 and not w22853;
w22855 <= not w22840 and not w22854;
w22856 <= not w22832 and not w22839;
w22857 <= not w22838 and w22856;
w22858 <= not w22855 and not w22857;
w22859 <= not b(57) and not w22858;
w22860 <= not b(56) and not w22848;
w22861 <= not w22082 and w22815;
w22862 <= not w22811 and w22861;
w22863 <= not w22812 and not w22815;
w22864 <= not w22862 and not w22863;
w22865 <= not w22840 and not w22864;
w22866 <= not w22072 and not w22839;
w22867 <= not w22838 and w22866;
w22868 <= not w22865 and not w22867;
w22869 <= not b(55) and not w22868;
w22870 <= not w22091 and w22810;
w22871 <= not w22806 and w22870;
w22872 <= not w22807 and not w22810;
w22873 <= not w22871 and not w22872;
w22874 <= not w22840 and not w22873;
w22875 <= not w22081 and not w22839;
w22876 <= not w22838 and w22875;
w22877 <= not w22874 and not w22876;
w22878 <= not b(54) and not w22877;
w22879 <= not w22100 and w22805;
w22880 <= not w22801 and w22879;
w22881 <= not w22802 and not w22805;
w22882 <= not w22880 and not w22881;
w22883 <= not w22840 and not w22882;
w22884 <= not w22090 and not w22839;
w22885 <= not w22838 and w22884;
w22886 <= not w22883 and not w22885;
w22887 <= not b(53) and not w22886;
w22888 <= not w22109 and w22800;
w22889 <= not w22796 and w22888;
w22890 <= not w22797 and not w22800;
w22891 <= not w22889 and not w22890;
w22892 <= not w22840 and not w22891;
w22893 <= not w22099 and not w22839;
w22894 <= not w22838 and w22893;
w22895 <= not w22892 and not w22894;
w22896 <= not b(52) and not w22895;
w22897 <= not w22118 and w22795;
w22898 <= not w22791 and w22897;
w22899 <= not w22792 and not w22795;
w22900 <= not w22898 and not w22899;
w22901 <= not w22840 and not w22900;
w22902 <= not w22108 and not w22839;
w22903 <= not w22838 and w22902;
w22904 <= not w22901 and not w22903;
w22905 <= not b(51) and not w22904;
w22906 <= not w22127 and w22790;
w22907 <= not w22786 and w22906;
w22908 <= not w22787 and not w22790;
w22909 <= not w22907 and not w22908;
w22910 <= not w22840 and not w22909;
w22911 <= not w22117 and not w22839;
w22912 <= not w22838 and w22911;
w22913 <= not w22910 and not w22912;
w22914 <= not b(50) and not w22913;
w22915 <= not w22136 and w22785;
w22916 <= not w22781 and w22915;
w22917 <= not w22782 and not w22785;
w22918 <= not w22916 and not w22917;
w22919 <= not w22840 and not w22918;
w22920 <= not w22126 and not w22839;
w22921 <= not w22838 and w22920;
w22922 <= not w22919 and not w22921;
w22923 <= not b(49) and not w22922;
w22924 <= not w22145 and w22780;
w22925 <= not w22776 and w22924;
w22926 <= not w22777 and not w22780;
w22927 <= not w22925 and not w22926;
w22928 <= not w22840 and not w22927;
w22929 <= not w22135 and not w22839;
w22930 <= not w22838 and w22929;
w22931 <= not w22928 and not w22930;
w22932 <= not b(48) and not w22931;
w22933 <= not w22154 and w22775;
w22934 <= not w22771 and w22933;
w22935 <= not w22772 and not w22775;
w22936 <= not w22934 and not w22935;
w22937 <= not w22840 and not w22936;
w22938 <= not w22144 and not w22839;
w22939 <= not w22838 and w22938;
w22940 <= not w22937 and not w22939;
w22941 <= not b(47) and not w22940;
w22942 <= not w22163 and w22770;
w22943 <= not w22766 and w22942;
w22944 <= not w22767 and not w22770;
w22945 <= not w22943 and not w22944;
w22946 <= not w22840 and not w22945;
w22947 <= not w22153 and not w22839;
w22948 <= not w22838 and w22947;
w22949 <= not w22946 and not w22948;
w22950 <= not b(46) and not w22949;
w22951 <= not w22172 and w22765;
w22952 <= not w22761 and w22951;
w22953 <= not w22762 and not w22765;
w22954 <= not w22952 and not w22953;
w22955 <= not w22840 and not w22954;
w22956 <= not w22162 and not w22839;
w22957 <= not w22838 and w22956;
w22958 <= not w22955 and not w22957;
w22959 <= not b(45) and not w22958;
w22960 <= not w22181 and w22760;
w22961 <= not w22756 and w22960;
w22962 <= not w22757 and not w22760;
w22963 <= not w22961 and not w22962;
w22964 <= not w22840 and not w22963;
w22965 <= not w22171 and not w22839;
w22966 <= not w22838 and w22965;
w22967 <= not w22964 and not w22966;
w22968 <= not b(44) and not w22967;
w22969 <= not w22190 and w22755;
w22970 <= not w22751 and w22969;
w22971 <= not w22752 and not w22755;
w22972 <= not w22970 and not w22971;
w22973 <= not w22840 and not w22972;
w22974 <= not w22180 and not w22839;
w22975 <= not w22838 and w22974;
w22976 <= not w22973 and not w22975;
w22977 <= not b(43) and not w22976;
w22978 <= not w22199 and w22750;
w22979 <= not w22746 and w22978;
w22980 <= not w22747 and not w22750;
w22981 <= not w22979 and not w22980;
w22982 <= not w22840 and not w22981;
w22983 <= not w22189 and not w22839;
w22984 <= not w22838 and w22983;
w22985 <= not w22982 and not w22984;
w22986 <= not b(42) and not w22985;
w22987 <= not w22208 and w22745;
w22988 <= not w22741 and w22987;
w22989 <= not w22742 and not w22745;
w22990 <= not w22988 and not w22989;
w22991 <= not w22840 and not w22990;
w22992 <= not w22198 and not w22839;
w22993 <= not w22838 and w22992;
w22994 <= not w22991 and not w22993;
w22995 <= not b(41) and not w22994;
w22996 <= not w22217 and w22740;
w22997 <= not w22736 and w22996;
w22998 <= not w22737 and not w22740;
w22999 <= not w22997 and not w22998;
w23000 <= not w22840 and not w22999;
w23001 <= not w22207 and not w22839;
w23002 <= not w22838 and w23001;
w23003 <= not w23000 and not w23002;
w23004 <= not b(40) and not w23003;
w23005 <= not w22226 and w22735;
w23006 <= not w22731 and w23005;
w23007 <= not w22732 and not w22735;
w23008 <= not w23006 and not w23007;
w23009 <= not w22840 and not w23008;
w23010 <= not w22216 and not w22839;
w23011 <= not w22838 and w23010;
w23012 <= not w23009 and not w23011;
w23013 <= not b(39) and not w23012;
w23014 <= not w22235 and w22730;
w23015 <= not w22726 and w23014;
w23016 <= not w22727 and not w22730;
w23017 <= not w23015 and not w23016;
w23018 <= not w22840 and not w23017;
w23019 <= not w22225 and not w22839;
w23020 <= not w22838 and w23019;
w23021 <= not w23018 and not w23020;
w23022 <= not b(38) and not w23021;
w23023 <= not w22244 and w22725;
w23024 <= not w22721 and w23023;
w23025 <= not w22722 and not w22725;
w23026 <= not w23024 and not w23025;
w23027 <= not w22840 and not w23026;
w23028 <= not w22234 and not w22839;
w23029 <= not w22838 and w23028;
w23030 <= not w23027 and not w23029;
w23031 <= not b(37) and not w23030;
w23032 <= not w22253 and w22720;
w23033 <= not w22716 and w23032;
w23034 <= not w22717 and not w22720;
w23035 <= not w23033 and not w23034;
w23036 <= not w22840 and not w23035;
w23037 <= not w22243 and not w22839;
w23038 <= not w22838 and w23037;
w23039 <= not w23036 and not w23038;
w23040 <= not b(36) and not w23039;
w23041 <= not w22262 and w22715;
w23042 <= not w22711 and w23041;
w23043 <= not w22712 and not w22715;
w23044 <= not w23042 and not w23043;
w23045 <= not w22840 and not w23044;
w23046 <= not w22252 and not w22839;
w23047 <= not w22838 and w23046;
w23048 <= not w23045 and not w23047;
w23049 <= not b(35) and not w23048;
w23050 <= not w22271 and w22710;
w23051 <= not w22706 and w23050;
w23052 <= not w22707 and not w22710;
w23053 <= not w23051 and not w23052;
w23054 <= not w22840 and not w23053;
w23055 <= not w22261 and not w22839;
w23056 <= not w22838 and w23055;
w23057 <= not w23054 and not w23056;
w23058 <= not b(34) and not w23057;
w23059 <= not w22280 and w22705;
w23060 <= not w22701 and w23059;
w23061 <= not w22702 and not w22705;
w23062 <= not w23060 and not w23061;
w23063 <= not w22840 and not w23062;
w23064 <= not w22270 and not w22839;
w23065 <= not w22838 and w23064;
w23066 <= not w23063 and not w23065;
w23067 <= not b(33) and not w23066;
w23068 <= not w22289 and w22700;
w23069 <= not w22696 and w23068;
w23070 <= not w22697 and not w22700;
w23071 <= not w23069 and not w23070;
w23072 <= not w22840 and not w23071;
w23073 <= not w22279 and not w22839;
w23074 <= not w22838 and w23073;
w23075 <= not w23072 and not w23074;
w23076 <= not b(32) and not w23075;
w23077 <= not w22298 and w22695;
w23078 <= not w22691 and w23077;
w23079 <= not w22692 and not w22695;
w23080 <= not w23078 and not w23079;
w23081 <= not w22840 and not w23080;
w23082 <= not w22288 and not w22839;
w23083 <= not w22838 and w23082;
w23084 <= not w23081 and not w23083;
w23085 <= not b(31) and not w23084;
w23086 <= not w22307 and w22690;
w23087 <= not w22686 and w23086;
w23088 <= not w22687 and not w22690;
w23089 <= not w23087 and not w23088;
w23090 <= not w22840 and not w23089;
w23091 <= not w22297 and not w22839;
w23092 <= not w22838 and w23091;
w23093 <= not w23090 and not w23092;
w23094 <= not b(30) and not w23093;
w23095 <= not w22316 and w22685;
w23096 <= not w22681 and w23095;
w23097 <= not w22682 and not w22685;
w23098 <= not w23096 and not w23097;
w23099 <= not w22840 and not w23098;
w23100 <= not w22306 and not w22839;
w23101 <= not w22838 and w23100;
w23102 <= not w23099 and not w23101;
w23103 <= not b(29) and not w23102;
w23104 <= not w22325 and w22680;
w23105 <= not w22676 and w23104;
w23106 <= not w22677 and not w22680;
w23107 <= not w23105 and not w23106;
w23108 <= not w22840 and not w23107;
w23109 <= not w22315 and not w22839;
w23110 <= not w22838 and w23109;
w23111 <= not w23108 and not w23110;
w23112 <= not b(28) and not w23111;
w23113 <= not w22334 and w22675;
w23114 <= not w22671 and w23113;
w23115 <= not w22672 and not w22675;
w23116 <= not w23114 and not w23115;
w23117 <= not w22840 and not w23116;
w23118 <= not w22324 and not w22839;
w23119 <= not w22838 and w23118;
w23120 <= not w23117 and not w23119;
w23121 <= not b(27) and not w23120;
w23122 <= not w22343 and w22670;
w23123 <= not w22666 and w23122;
w23124 <= not w22667 and not w22670;
w23125 <= not w23123 and not w23124;
w23126 <= not w22840 and not w23125;
w23127 <= not w22333 and not w22839;
w23128 <= not w22838 and w23127;
w23129 <= not w23126 and not w23128;
w23130 <= not b(26) and not w23129;
w23131 <= not w22352 and w22665;
w23132 <= not w22661 and w23131;
w23133 <= not w22662 and not w22665;
w23134 <= not w23132 and not w23133;
w23135 <= not w22840 and not w23134;
w23136 <= not w22342 and not w22839;
w23137 <= not w22838 and w23136;
w23138 <= not w23135 and not w23137;
w23139 <= not b(25) and not w23138;
w23140 <= not w22361 and w22660;
w23141 <= not w22656 and w23140;
w23142 <= not w22657 and not w22660;
w23143 <= not w23141 and not w23142;
w23144 <= not w22840 and not w23143;
w23145 <= not w22351 and not w22839;
w23146 <= not w22838 and w23145;
w23147 <= not w23144 and not w23146;
w23148 <= not b(24) and not w23147;
w23149 <= not w22370 and w22655;
w23150 <= not w22651 and w23149;
w23151 <= not w22652 and not w22655;
w23152 <= not w23150 and not w23151;
w23153 <= not w22840 and not w23152;
w23154 <= not w22360 and not w22839;
w23155 <= not w22838 and w23154;
w23156 <= not w23153 and not w23155;
w23157 <= not b(23) and not w23156;
w23158 <= not w22379 and w22650;
w23159 <= not w22646 and w23158;
w23160 <= not w22647 and not w22650;
w23161 <= not w23159 and not w23160;
w23162 <= not w22840 and not w23161;
w23163 <= not w22369 and not w22839;
w23164 <= not w22838 and w23163;
w23165 <= not w23162 and not w23164;
w23166 <= not b(22) and not w23165;
w23167 <= not w22388 and w22645;
w23168 <= not w22641 and w23167;
w23169 <= not w22642 and not w22645;
w23170 <= not w23168 and not w23169;
w23171 <= not w22840 and not w23170;
w23172 <= not w22378 and not w22839;
w23173 <= not w22838 and w23172;
w23174 <= not w23171 and not w23173;
w23175 <= not b(21) and not w23174;
w23176 <= not w22397 and w22640;
w23177 <= not w22636 and w23176;
w23178 <= not w22637 and not w22640;
w23179 <= not w23177 and not w23178;
w23180 <= not w22840 and not w23179;
w23181 <= not w22387 and not w22839;
w23182 <= not w22838 and w23181;
w23183 <= not w23180 and not w23182;
w23184 <= not b(20) and not w23183;
w23185 <= not w22406 and w22635;
w23186 <= not w22631 and w23185;
w23187 <= not w22632 and not w22635;
w23188 <= not w23186 and not w23187;
w23189 <= not w22840 and not w23188;
w23190 <= not w22396 and not w22839;
w23191 <= not w22838 and w23190;
w23192 <= not w23189 and not w23191;
w23193 <= not b(19) and not w23192;
w23194 <= not w22415 and w22630;
w23195 <= not w22626 and w23194;
w23196 <= not w22627 and not w22630;
w23197 <= not w23195 and not w23196;
w23198 <= not w22840 and not w23197;
w23199 <= not w22405 and not w22839;
w23200 <= not w22838 and w23199;
w23201 <= not w23198 and not w23200;
w23202 <= not b(18) and not w23201;
w23203 <= not w22424 and w22625;
w23204 <= not w22621 and w23203;
w23205 <= not w22622 and not w22625;
w23206 <= not w23204 and not w23205;
w23207 <= not w22840 and not w23206;
w23208 <= not w22414 and not w22839;
w23209 <= not w22838 and w23208;
w23210 <= not w23207 and not w23209;
w23211 <= not b(17) and not w23210;
w23212 <= not w22433 and w22620;
w23213 <= not w22616 and w23212;
w23214 <= not w22617 and not w22620;
w23215 <= not w23213 and not w23214;
w23216 <= not w22840 and not w23215;
w23217 <= not w22423 and not w22839;
w23218 <= not w22838 and w23217;
w23219 <= not w23216 and not w23218;
w23220 <= not b(16) and not w23219;
w23221 <= not w22442 and w22615;
w23222 <= not w22611 and w23221;
w23223 <= not w22612 and not w22615;
w23224 <= not w23222 and not w23223;
w23225 <= not w22840 and not w23224;
w23226 <= not w22432 and not w22839;
w23227 <= not w22838 and w23226;
w23228 <= not w23225 and not w23227;
w23229 <= not b(15) and not w23228;
w23230 <= not w22451 and w22610;
w23231 <= not w22606 and w23230;
w23232 <= not w22607 and not w22610;
w23233 <= not w23231 and not w23232;
w23234 <= not w22840 and not w23233;
w23235 <= not w22441 and not w22839;
w23236 <= not w22838 and w23235;
w23237 <= not w23234 and not w23236;
w23238 <= not b(14) and not w23237;
w23239 <= not w22460 and w22605;
w23240 <= not w22601 and w23239;
w23241 <= not w22602 and not w22605;
w23242 <= not w23240 and not w23241;
w23243 <= not w22840 and not w23242;
w23244 <= not w22450 and not w22839;
w23245 <= not w22838 and w23244;
w23246 <= not w23243 and not w23245;
w23247 <= not b(13) and not w23246;
w23248 <= not w22469 and w22600;
w23249 <= not w22596 and w23248;
w23250 <= not w22597 and not w22600;
w23251 <= not w23249 and not w23250;
w23252 <= not w22840 and not w23251;
w23253 <= not w22459 and not w22839;
w23254 <= not w22838 and w23253;
w23255 <= not w23252 and not w23254;
w23256 <= not b(12) and not w23255;
w23257 <= not w22478 and w22595;
w23258 <= not w22591 and w23257;
w23259 <= not w22592 and not w22595;
w23260 <= not w23258 and not w23259;
w23261 <= not w22840 and not w23260;
w23262 <= not w22468 and not w22839;
w23263 <= not w22838 and w23262;
w23264 <= not w23261 and not w23263;
w23265 <= not b(11) and not w23264;
w23266 <= not w22487 and w22590;
w23267 <= not w22586 and w23266;
w23268 <= not w22587 and not w22590;
w23269 <= not w23267 and not w23268;
w23270 <= not w22840 and not w23269;
w23271 <= not w22477 and not w22839;
w23272 <= not w22838 and w23271;
w23273 <= not w23270 and not w23272;
w23274 <= not b(10) and not w23273;
w23275 <= not w22496 and w22585;
w23276 <= not w22581 and w23275;
w23277 <= not w22582 and not w22585;
w23278 <= not w23276 and not w23277;
w23279 <= not w22840 and not w23278;
w23280 <= not w22486 and not w22839;
w23281 <= not w22838 and w23280;
w23282 <= not w23279 and not w23281;
w23283 <= not b(9) and not w23282;
w23284 <= not w22505 and w22580;
w23285 <= not w22576 and w23284;
w23286 <= not w22577 and not w22580;
w23287 <= not w23285 and not w23286;
w23288 <= not w22840 and not w23287;
w23289 <= not w22495 and not w22839;
w23290 <= not w22838 and w23289;
w23291 <= not w23288 and not w23290;
w23292 <= not b(8) and not w23291;
w23293 <= not w22514 and w22575;
w23294 <= not w22571 and w23293;
w23295 <= not w22572 and not w22575;
w23296 <= not w23294 and not w23295;
w23297 <= not w22840 and not w23296;
w23298 <= not w22504 and not w22839;
w23299 <= not w22838 and w23298;
w23300 <= not w23297 and not w23299;
w23301 <= not b(7) and not w23300;
w23302 <= not w22523 and w22570;
w23303 <= not w22566 and w23302;
w23304 <= not w22567 and not w22570;
w23305 <= not w23303 and not w23304;
w23306 <= not w22840 and not w23305;
w23307 <= not w22513 and not w22839;
w23308 <= not w22838 and w23307;
w23309 <= not w23306 and not w23308;
w23310 <= not b(6) and not w23309;
w23311 <= not w22532 and w22565;
w23312 <= not w22561 and w23311;
w23313 <= not w22562 and not w22565;
w23314 <= not w23312 and not w23313;
w23315 <= not w22840 and not w23314;
w23316 <= not w22522 and not w22839;
w23317 <= not w22838 and w23316;
w23318 <= not w23315 and not w23317;
w23319 <= not b(5) and not w23318;
w23320 <= not w22540 and w22560;
w23321 <= not w22556 and w23320;
w23322 <= not w22557 and not w22560;
w23323 <= not w23321 and not w23322;
w23324 <= not w22840 and not w23323;
w23325 <= not w22531 and not w22839;
w23326 <= not w22838 and w23325;
w23327 <= not w23324 and not w23326;
w23328 <= not b(4) and not w23327;
w23329 <= not w22551 and w22555;
w23330 <= not w22550 and w23329;
w23331 <= not w22552 and not w22555;
w23332 <= not w23330 and not w23331;
w23333 <= not w22840 and not w23332;
w23334 <= not w22539 and not w22839;
w23335 <= not w22838 and w23334;
w23336 <= not w23333 and not w23335;
w23337 <= not b(3) and not w23336;
w23338 <= not w22547 and w22549;
w23339 <= not w22545 and w23338;
w23340 <= not w22550 and not w23339;
w23341 <= not w22840 and w23340;
w23342 <= not w22544 and not w22839;
w23343 <= not w22838 and w23342;
w23344 <= not w23341 and not w23343;
w23345 <= not b(2) and not w23344;
w23346 <= b(0) and not w22840;
w23347 <= a(7) and not w23346;
w23348 <= w22549 and not w22840;
w23349 <= not w23347 and not w23348;
w23350 <= b(1) and not w23349;
w23351 <= not b(1) and not w23348;
w23352 <= not w23347 and w23351;
w23353 <= not w23350 and not w23352;
w23354 <= not a(6) and b(0);
w23355 <= not w23353 and not w23354;
w23356 <= not b(1) and not w23349;
w23357 <= not w23355 and not w23356;
w23358 <= b(2) and not w23343;
w23359 <= not w23341 and w23358;
w23360 <= not w23345 and not w23359;
w23361 <= not w23357 and w23360;
w23362 <= not w23345 and not w23361;
w23363 <= b(3) and not w23335;
w23364 <= not w23333 and w23363;
w23365 <= not w23337 and not w23364;
w23366 <= not w23362 and w23365;
w23367 <= not w23337 and not w23366;
w23368 <= b(4) and not w23326;
w23369 <= not w23324 and w23368;
w23370 <= not w23328 and not w23369;
w23371 <= not w23367 and w23370;
w23372 <= not w23328 and not w23371;
w23373 <= b(5) and not w23317;
w23374 <= not w23315 and w23373;
w23375 <= not w23319 and not w23374;
w23376 <= not w23372 and w23375;
w23377 <= not w23319 and not w23376;
w23378 <= b(6) and not w23308;
w23379 <= not w23306 and w23378;
w23380 <= not w23310 and not w23379;
w23381 <= not w23377 and w23380;
w23382 <= not w23310 and not w23381;
w23383 <= b(7) and not w23299;
w23384 <= not w23297 and w23383;
w23385 <= not w23301 and not w23384;
w23386 <= not w23382 and w23385;
w23387 <= not w23301 and not w23386;
w23388 <= b(8) and not w23290;
w23389 <= not w23288 and w23388;
w23390 <= not w23292 and not w23389;
w23391 <= not w23387 and w23390;
w23392 <= not w23292 and not w23391;
w23393 <= b(9) and not w23281;
w23394 <= not w23279 and w23393;
w23395 <= not w23283 and not w23394;
w23396 <= not w23392 and w23395;
w23397 <= not w23283 and not w23396;
w23398 <= b(10) and not w23272;
w23399 <= not w23270 and w23398;
w23400 <= not w23274 and not w23399;
w23401 <= not w23397 and w23400;
w23402 <= not w23274 and not w23401;
w23403 <= b(11) and not w23263;
w23404 <= not w23261 and w23403;
w23405 <= not w23265 and not w23404;
w23406 <= not w23402 and w23405;
w23407 <= not w23265 and not w23406;
w23408 <= b(12) and not w23254;
w23409 <= not w23252 and w23408;
w23410 <= not w23256 and not w23409;
w23411 <= not w23407 and w23410;
w23412 <= not w23256 and not w23411;
w23413 <= b(13) and not w23245;
w23414 <= not w23243 and w23413;
w23415 <= not w23247 and not w23414;
w23416 <= not w23412 and w23415;
w23417 <= not w23247 and not w23416;
w23418 <= b(14) and not w23236;
w23419 <= not w23234 and w23418;
w23420 <= not w23238 and not w23419;
w23421 <= not w23417 and w23420;
w23422 <= not w23238 and not w23421;
w23423 <= b(15) and not w23227;
w23424 <= not w23225 and w23423;
w23425 <= not w23229 and not w23424;
w23426 <= not w23422 and w23425;
w23427 <= not w23229 and not w23426;
w23428 <= b(16) and not w23218;
w23429 <= not w23216 and w23428;
w23430 <= not w23220 and not w23429;
w23431 <= not w23427 and w23430;
w23432 <= not w23220 and not w23431;
w23433 <= b(17) and not w23209;
w23434 <= not w23207 and w23433;
w23435 <= not w23211 and not w23434;
w23436 <= not w23432 and w23435;
w23437 <= not w23211 and not w23436;
w23438 <= b(18) and not w23200;
w23439 <= not w23198 and w23438;
w23440 <= not w23202 and not w23439;
w23441 <= not w23437 and w23440;
w23442 <= not w23202 and not w23441;
w23443 <= b(19) and not w23191;
w23444 <= not w23189 and w23443;
w23445 <= not w23193 and not w23444;
w23446 <= not w23442 and w23445;
w23447 <= not w23193 and not w23446;
w23448 <= b(20) and not w23182;
w23449 <= not w23180 and w23448;
w23450 <= not w23184 and not w23449;
w23451 <= not w23447 and w23450;
w23452 <= not w23184 and not w23451;
w23453 <= b(21) and not w23173;
w23454 <= not w23171 and w23453;
w23455 <= not w23175 and not w23454;
w23456 <= not w23452 and w23455;
w23457 <= not w23175 and not w23456;
w23458 <= b(22) and not w23164;
w23459 <= not w23162 and w23458;
w23460 <= not w23166 and not w23459;
w23461 <= not w23457 and w23460;
w23462 <= not w23166 and not w23461;
w23463 <= b(23) and not w23155;
w23464 <= not w23153 and w23463;
w23465 <= not w23157 and not w23464;
w23466 <= not w23462 and w23465;
w23467 <= not w23157 and not w23466;
w23468 <= b(24) and not w23146;
w23469 <= not w23144 and w23468;
w23470 <= not w23148 and not w23469;
w23471 <= not w23467 and w23470;
w23472 <= not w23148 and not w23471;
w23473 <= b(25) and not w23137;
w23474 <= not w23135 and w23473;
w23475 <= not w23139 and not w23474;
w23476 <= not w23472 and w23475;
w23477 <= not w23139 and not w23476;
w23478 <= b(26) and not w23128;
w23479 <= not w23126 and w23478;
w23480 <= not w23130 and not w23479;
w23481 <= not w23477 and w23480;
w23482 <= not w23130 and not w23481;
w23483 <= b(27) and not w23119;
w23484 <= not w23117 and w23483;
w23485 <= not w23121 and not w23484;
w23486 <= not w23482 and w23485;
w23487 <= not w23121 and not w23486;
w23488 <= b(28) and not w23110;
w23489 <= not w23108 and w23488;
w23490 <= not w23112 and not w23489;
w23491 <= not w23487 and w23490;
w23492 <= not w23112 and not w23491;
w23493 <= b(29) and not w23101;
w23494 <= not w23099 and w23493;
w23495 <= not w23103 and not w23494;
w23496 <= not w23492 and w23495;
w23497 <= not w23103 and not w23496;
w23498 <= b(30) and not w23092;
w23499 <= not w23090 and w23498;
w23500 <= not w23094 and not w23499;
w23501 <= not w23497 and w23500;
w23502 <= not w23094 and not w23501;
w23503 <= b(31) and not w23083;
w23504 <= not w23081 and w23503;
w23505 <= not w23085 and not w23504;
w23506 <= not w23502 and w23505;
w23507 <= not w23085 and not w23506;
w23508 <= b(32) and not w23074;
w23509 <= not w23072 and w23508;
w23510 <= not w23076 and not w23509;
w23511 <= not w23507 and w23510;
w23512 <= not w23076 and not w23511;
w23513 <= b(33) and not w23065;
w23514 <= not w23063 and w23513;
w23515 <= not w23067 and not w23514;
w23516 <= not w23512 and w23515;
w23517 <= not w23067 and not w23516;
w23518 <= b(34) and not w23056;
w23519 <= not w23054 and w23518;
w23520 <= not w23058 and not w23519;
w23521 <= not w23517 and w23520;
w23522 <= not w23058 and not w23521;
w23523 <= b(35) and not w23047;
w23524 <= not w23045 and w23523;
w23525 <= not w23049 and not w23524;
w23526 <= not w23522 and w23525;
w23527 <= not w23049 and not w23526;
w23528 <= b(36) and not w23038;
w23529 <= not w23036 and w23528;
w23530 <= not w23040 and not w23529;
w23531 <= not w23527 and w23530;
w23532 <= not w23040 and not w23531;
w23533 <= b(37) and not w23029;
w23534 <= not w23027 and w23533;
w23535 <= not w23031 and not w23534;
w23536 <= not w23532 and w23535;
w23537 <= not w23031 and not w23536;
w23538 <= b(38) and not w23020;
w23539 <= not w23018 and w23538;
w23540 <= not w23022 and not w23539;
w23541 <= not w23537 and w23540;
w23542 <= not w23022 and not w23541;
w23543 <= b(39) and not w23011;
w23544 <= not w23009 and w23543;
w23545 <= not w23013 and not w23544;
w23546 <= not w23542 and w23545;
w23547 <= not w23013 and not w23546;
w23548 <= b(40) and not w23002;
w23549 <= not w23000 and w23548;
w23550 <= not w23004 and not w23549;
w23551 <= not w23547 and w23550;
w23552 <= not w23004 and not w23551;
w23553 <= b(41) and not w22993;
w23554 <= not w22991 and w23553;
w23555 <= not w22995 and not w23554;
w23556 <= not w23552 and w23555;
w23557 <= not w22995 and not w23556;
w23558 <= b(42) and not w22984;
w23559 <= not w22982 and w23558;
w23560 <= not w22986 and not w23559;
w23561 <= not w23557 and w23560;
w23562 <= not w22986 and not w23561;
w23563 <= b(43) and not w22975;
w23564 <= not w22973 and w23563;
w23565 <= not w22977 and not w23564;
w23566 <= not w23562 and w23565;
w23567 <= not w22977 and not w23566;
w23568 <= b(44) and not w22966;
w23569 <= not w22964 and w23568;
w23570 <= not w22968 and not w23569;
w23571 <= not w23567 and w23570;
w23572 <= not w22968 and not w23571;
w23573 <= b(45) and not w22957;
w23574 <= not w22955 and w23573;
w23575 <= not w22959 and not w23574;
w23576 <= not w23572 and w23575;
w23577 <= not w22959 and not w23576;
w23578 <= b(46) and not w22948;
w23579 <= not w22946 and w23578;
w23580 <= not w22950 and not w23579;
w23581 <= not w23577 and w23580;
w23582 <= not w22950 and not w23581;
w23583 <= b(47) and not w22939;
w23584 <= not w22937 and w23583;
w23585 <= not w22941 and not w23584;
w23586 <= not w23582 and w23585;
w23587 <= not w22941 and not w23586;
w23588 <= b(48) and not w22930;
w23589 <= not w22928 and w23588;
w23590 <= not w22932 and not w23589;
w23591 <= not w23587 and w23590;
w23592 <= not w22932 and not w23591;
w23593 <= b(49) and not w22921;
w23594 <= not w22919 and w23593;
w23595 <= not w22923 and not w23594;
w23596 <= not w23592 and w23595;
w23597 <= not w22923 and not w23596;
w23598 <= b(50) and not w22912;
w23599 <= not w22910 and w23598;
w23600 <= not w22914 and not w23599;
w23601 <= not w23597 and w23600;
w23602 <= not w22914 and not w23601;
w23603 <= b(51) and not w22903;
w23604 <= not w22901 and w23603;
w23605 <= not w22905 and not w23604;
w23606 <= not w23602 and w23605;
w23607 <= not w22905 and not w23606;
w23608 <= b(52) and not w22894;
w23609 <= not w22892 and w23608;
w23610 <= not w22896 and not w23609;
w23611 <= not w23607 and w23610;
w23612 <= not w22896 and not w23611;
w23613 <= b(53) and not w22885;
w23614 <= not w22883 and w23613;
w23615 <= not w22887 and not w23614;
w23616 <= not w23612 and w23615;
w23617 <= not w22887 and not w23616;
w23618 <= b(54) and not w22876;
w23619 <= not w22874 and w23618;
w23620 <= not w22878 and not w23619;
w23621 <= not w23617 and w23620;
w23622 <= not w22878 and not w23621;
w23623 <= b(55) and not w22867;
w23624 <= not w22865 and w23623;
w23625 <= not w22869 and not w23624;
w23626 <= not w23622 and w23625;
w23627 <= not w22869 and not w23626;
w23628 <= b(56) and not w22847;
w23629 <= not w22845 and w23628;
w23630 <= not w22860 and not w23629;
w23631 <= not w23627 and w23630;
w23632 <= not w22860 and not w23631;
w23633 <= b(57) and not w22857;
w23634 <= not w22855 and w23633;
w23635 <= not w22859 and not w23634;
w23636 <= not w23632 and w23635;
w23637 <= not w22859 and not w23636;
w23638 <= w23 and w25;
w23639 <= not w23637 and w23638;
w23640 <= not w22848 and not w23639;
w23641 <= not w22869 and w23630;
w23642 <= not w23626 and w23641;
w23643 <= not w23627 and not w23630;
w23644 <= not w23642 and not w23643;
w23645 <= w23638 and not w23644;
w23646 <= not w23637 and w23645;
w23647 <= not w23640 and not w23646;
w23648 <= not b(57) and not w23647;
w23649 <= not w22868 and not w23639;
w23650 <= not w22878 and w23625;
w23651 <= not w23621 and w23650;
w23652 <= not w23622 and not w23625;
w23653 <= not w23651 and not w23652;
w23654 <= w23638 and not w23653;
w23655 <= not w23637 and w23654;
w23656 <= not w23649 and not w23655;
w23657 <= not b(56) and not w23656;
w23658 <= not w22877 and not w23639;
w23659 <= not w22887 and w23620;
w23660 <= not w23616 and w23659;
w23661 <= not w23617 and not w23620;
w23662 <= not w23660 and not w23661;
w23663 <= w23638 and not w23662;
w23664 <= not w23637 and w23663;
w23665 <= not w23658 and not w23664;
w23666 <= not b(55) and not w23665;
w23667 <= not w22886 and not w23639;
w23668 <= not w22896 and w23615;
w23669 <= not w23611 and w23668;
w23670 <= not w23612 and not w23615;
w23671 <= not w23669 and not w23670;
w23672 <= w23638 and not w23671;
w23673 <= not w23637 and w23672;
w23674 <= not w23667 and not w23673;
w23675 <= not b(54) and not w23674;
w23676 <= not w22895 and not w23639;
w23677 <= not w22905 and w23610;
w23678 <= not w23606 and w23677;
w23679 <= not w23607 and not w23610;
w23680 <= not w23678 and not w23679;
w23681 <= w23638 and not w23680;
w23682 <= not w23637 and w23681;
w23683 <= not w23676 and not w23682;
w23684 <= not b(53) and not w23683;
w23685 <= not w22904 and not w23639;
w23686 <= not w22914 and w23605;
w23687 <= not w23601 and w23686;
w23688 <= not w23602 and not w23605;
w23689 <= not w23687 and not w23688;
w23690 <= w23638 and not w23689;
w23691 <= not w23637 and w23690;
w23692 <= not w23685 and not w23691;
w23693 <= not b(52) and not w23692;
w23694 <= not w22913 and not w23639;
w23695 <= not w22923 and w23600;
w23696 <= not w23596 and w23695;
w23697 <= not w23597 and not w23600;
w23698 <= not w23696 and not w23697;
w23699 <= w23638 and not w23698;
w23700 <= not w23637 and w23699;
w23701 <= not w23694 and not w23700;
w23702 <= not b(51) and not w23701;
w23703 <= not w22922 and not w23639;
w23704 <= not w22932 and w23595;
w23705 <= not w23591 and w23704;
w23706 <= not w23592 and not w23595;
w23707 <= not w23705 and not w23706;
w23708 <= w23638 and not w23707;
w23709 <= not w23637 and w23708;
w23710 <= not w23703 and not w23709;
w23711 <= not b(50) and not w23710;
w23712 <= not w22931 and not w23639;
w23713 <= not w22941 and w23590;
w23714 <= not w23586 and w23713;
w23715 <= not w23587 and not w23590;
w23716 <= not w23714 and not w23715;
w23717 <= w23638 and not w23716;
w23718 <= not w23637 and w23717;
w23719 <= not w23712 and not w23718;
w23720 <= not b(49) and not w23719;
w23721 <= not w22940 and not w23639;
w23722 <= not w22950 and w23585;
w23723 <= not w23581 and w23722;
w23724 <= not w23582 and not w23585;
w23725 <= not w23723 and not w23724;
w23726 <= w23638 and not w23725;
w23727 <= not w23637 and w23726;
w23728 <= not w23721 and not w23727;
w23729 <= not b(48) and not w23728;
w23730 <= not w22949 and not w23639;
w23731 <= not w22959 and w23580;
w23732 <= not w23576 and w23731;
w23733 <= not w23577 and not w23580;
w23734 <= not w23732 and not w23733;
w23735 <= w23638 and not w23734;
w23736 <= not w23637 and w23735;
w23737 <= not w23730 and not w23736;
w23738 <= not b(47) and not w23737;
w23739 <= not w22958 and not w23639;
w23740 <= not w22968 and w23575;
w23741 <= not w23571 and w23740;
w23742 <= not w23572 and not w23575;
w23743 <= not w23741 and not w23742;
w23744 <= w23638 and not w23743;
w23745 <= not w23637 and w23744;
w23746 <= not w23739 and not w23745;
w23747 <= not b(46) and not w23746;
w23748 <= not w22967 and not w23639;
w23749 <= not w22977 and w23570;
w23750 <= not w23566 and w23749;
w23751 <= not w23567 and not w23570;
w23752 <= not w23750 and not w23751;
w23753 <= w23638 and not w23752;
w23754 <= not w23637 and w23753;
w23755 <= not w23748 and not w23754;
w23756 <= not b(45) and not w23755;
w23757 <= not w22976 and not w23639;
w23758 <= not w22986 and w23565;
w23759 <= not w23561 and w23758;
w23760 <= not w23562 and not w23565;
w23761 <= not w23759 and not w23760;
w23762 <= w23638 and not w23761;
w23763 <= not w23637 and w23762;
w23764 <= not w23757 and not w23763;
w23765 <= not b(44) and not w23764;
w23766 <= not w22985 and not w23639;
w23767 <= not w22995 and w23560;
w23768 <= not w23556 and w23767;
w23769 <= not w23557 and not w23560;
w23770 <= not w23768 and not w23769;
w23771 <= w23638 and not w23770;
w23772 <= not w23637 and w23771;
w23773 <= not w23766 and not w23772;
w23774 <= not b(43) and not w23773;
w23775 <= not w22994 and not w23639;
w23776 <= not w23004 and w23555;
w23777 <= not w23551 and w23776;
w23778 <= not w23552 and not w23555;
w23779 <= not w23777 and not w23778;
w23780 <= w23638 and not w23779;
w23781 <= not w23637 and w23780;
w23782 <= not w23775 and not w23781;
w23783 <= not b(42) and not w23782;
w23784 <= not w23003 and not w23639;
w23785 <= not w23013 and w23550;
w23786 <= not w23546 and w23785;
w23787 <= not w23547 and not w23550;
w23788 <= not w23786 and not w23787;
w23789 <= w23638 and not w23788;
w23790 <= not w23637 and w23789;
w23791 <= not w23784 and not w23790;
w23792 <= not b(41) and not w23791;
w23793 <= not w23012 and not w23639;
w23794 <= not w23022 and w23545;
w23795 <= not w23541 and w23794;
w23796 <= not w23542 and not w23545;
w23797 <= not w23795 and not w23796;
w23798 <= w23638 and not w23797;
w23799 <= not w23637 and w23798;
w23800 <= not w23793 and not w23799;
w23801 <= not b(40) and not w23800;
w23802 <= not w23021 and not w23639;
w23803 <= not w23031 and w23540;
w23804 <= not w23536 and w23803;
w23805 <= not w23537 and not w23540;
w23806 <= not w23804 and not w23805;
w23807 <= w23638 and not w23806;
w23808 <= not w23637 and w23807;
w23809 <= not w23802 and not w23808;
w23810 <= not b(39) and not w23809;
w23811 <= not w23030 and not w23639;
w23812 <= not w23040 and w23535;
w23813 <= not w23531 and w23812;
w23814 <= not w23532 and not w23535;
w23815 <= not w23813 and not w23814;
w23816 <= w23638 and not w23815;
w23817 <= not w23637 and w23816;
w23818 <= not w23811 and not w23817;
w23819 <= not b(38) and not w23818;
w23820 <= not w23039 and not w23639;
w23821 <= not w23049 and w23530;
w23822 <= not w23526 and w23821;
w23823 <= not w23527 and not w23530;
w23824 <= not w23822 and not w23823;
w23825 <= w23638 and not w23824;
w23826 <= not w23637 and w23825;
w23827 <= not w23820 and not w23826;
w23828 <= not b(37) and not w23827;
w23829 <= not w23048 and not w23639;
w23830 <= not w23058 and w23525;
w23831 <= not w23521 and w23830;
w23832 <= not w23522 and not w23525;
w23833 <= not w23831 and not w23832;
w23834 <= w23638 and not w23833;
w23835 <= not w23637 and w23834;
w23836 <= not w23829 and not w23835;
w23837 <= not b(36) and not w23836;
w23838 <= not w23057 and not w23639;
w23839 <= not w23067 and w23520;
w23840 <= not w23516 and w23839;
w23841 <= not w23517 and not w23520;
w23842 <= not w23840 and not w23841;
w23843 <= w23638 and not w23842;
w23844 <= not w23637 and w23843;
w23845 <= not w23838 and not w23844;
w23846 <= not b(35) and not w23845;
w23847 <= not w23066 and not w23639;
w23848 <= not w23076 and w23515;
w23849 <= not w23511 and w23848;
w23850 <= not w23512 and not w23515;
w23851 <= not w23849 and not w23850;
w23852 <= w23638 and not w23851;
w23853 <= not w23637 and w23852;
w23854 <= not w23847 and not w23853;
w23855 <= not b(34) and not w23854;
w23856 <= not w23075 and not w23639;
w23857 <= not w23085 and w23510;
w23858 <= not w23506 and w23857;
w23859 <= not w23507 and not w23510;
w23860 <= not w23858 and not w23859;
w23861 <= w23638 and not w23860;
w23862 <= not w23637 and w23861;
w23863 <= not w23856 and not w23862;
w23864 <= not b(33) and not w23863;
w23865 <= not w23084 and not w23639;
w23866 <= not w23094 and w23505;
w23867 <= not w23501 and w23866;
w23868 <= not w23502 and not w23505;
w23869 <= not w23867 and not w23868;
w23870 <= w23638 and not w23869;
w23871 <= not w23637 and w23870;
w23872 <= not w23865 and not w23871;
w23873 <= not b(32) and not w23872;
w23874 <= not w23093 and not w23639;
w23875 <= not w23103 and w23500;
w23876 <= not w23496 and w23875;
w23877 <= not w23497 and not w23500;
w23878 <= not w23876 and not w23877;
w23879 <= w23638 and not w23878;
w23880 <= not w23637 and w23879;
w23881 <= not w23874 and not w23880;
w23882 <= not b(31) and not w23881;
w23883 <= not w23102 and not w23639;
w23884 <= not w23112 and w23495;
w23885 <= not w23491 and w23884;
w23886 <= not w23492 and not w23495;
w23887 <= not w23885 and not w23886;
w23888 <= w23638 and not w23887;
w23889 <= not w23637 and w23888;
w23890 <= not w23883 and not w23889;
w23891 <= not b(30) and not w23890;
w23892 <= not w23111 and not w23639;
w23893 <= not w23121 and w23490;
w23894 <= not w23486 and w23893;
w23895 <= not w23487 and not w23490;
w23896 <= not w23894 and not w23895;
w23897 <= w23638 and not w23896;
w23898 <= not w23637 and w23897;
w23899 <= not w23892 and not w23898;
w23900 <= not b(29) and not w23899;
w23901 <= not w23120 and not w23639;
w23902 <= not w23130 and w23485;
w23903 <= not w23481 and w23902;
w23904 <= not w23482 and not w23485;
w23905 <= not w23903 and not w23904;
w23906 <= w23638 and not w23905;
w23907 <= not w23637 and w23906;
w23908 <= not w23901 and not w23907;
w23909 <= not b(28) and not w23908;
w23910 <= not w23129 and not w23639;
w23911 <= not w23139 and w23480;
w23912 <= not w23476 and w23911;
w23913 <= not w23477 and not w23480;
w23914 <= not w23912 and not w23913;
w23915 <= w23638 and not w23914;
w23916 <= not w23637 and w23915;
w23917 <= not w23910 and not w23916;
w23918 <= not b(27) and not w23917;
w23919 <= not w23138 and not w23639;
w23920 <= not w23148 and w23475;
w23921 <= not w23471 and w23920;
w23922 <= not w23472 and not w23475;
w23923 <= not w23921 and not w23922;
w23924 <= w23638 and not w23923;
w23925 <= not w23637 and w23924;
w23926 <= not w23919 and not w23925;
w23927 <= not b(26) and not w23926;
w23928 <= not w23147 and not w23639;
w23929 <= not w23157 and w23470;
w23930 <= not w23466 and w23929;
w23931 <= not w23467 and not w23470;
w23932 <= not w23930 and not w23931;
w23933 <= w23638 and not w23932;
w23934 <= not w23637 and w23933;
w23935 <= not w23928 and not w23934;
w23936 <= not b(25) and not w23935;
w23937 <= not w23156 and not w23639;
w23938 <= not w23166 and w23465;
w23939 <= not w23461 and w23938;
w23940 <= not w23462 and not w23465;
w23941 <= not w23939 and not w23940;
w23942 <= w23638 and not w23941;
w23943 <= not w23637 and w23942;
w23944 <= not w23937 and not w23943;
w23945 <= not b(24) and not w23944;
w23946 <= not w23165 and not w23639;
w23947 <= not w23175 and w23460;
w23948 <= not w23456 and w23947;
w23949 <= not w23457 and not w23460;
w23950 <= not w23948 and not w23949;
w23951 <= w23638 and not w23950;
w23952 <= not w23637 and w23951;
w23953 <= not w23946 and not w23952;
w23954 <= not b(23) and not w23953;
w23955 <= not w23174 and not w23639;
w23956 <= not w23184 and w23455;
w23957 <= not w23451 and w23956;
w23958 <= not w23452 and not w23455;
w23959 <= not w23957 and not w23958;
w23960 <= w23638 and not w23959;
w23961 <= not w23637 and w23960;
w23962 <= not w23955 and not w23961;
w23963 <= not b(22) and not w23962;
w23964 <= not w23183 and not w23639;
w23965 <= not w23193 and w23450;
w23966 <= not w23446 and w23965;
w23967 <= not w23447 and not w23450;
w23968 <= not w23966 and not w23967;
w23969 <= w23638 and not w23968;
w23970 <= not w23637 and w23969;
w23971 <= not w23964 and not w23970;
w23972 <= not b(21) and not w23971;
w23973 <= not w23192 and not w23639;
w23974 <= not w23202 and w23445;
w23975 <= not w23441 and w23974;
w23976 <= not w23442 and not w23445;
w23977 <= not w23975 and not w23976;
w23978 <= w23638 and not w23977;
w23979 <= not w23637 and w23978;
w23980 <= not w23973 and not w23979;
w23981 <= not b(20) and not w23980;
w23982 <= not w23201 and not w23639;
w23983 <= not w23211 and w23440;
w23984 <= not w23436 and w23983;
w23985 <= not w23437 and not w23440;
w23986 <= not w23984 and not w23985;
w23987 <= w23638 and not w23986;
w23988 <= not w23637 and w23987;
w23989 <= not w23982 and not w23988;
w23990 <= not b(19) and not w23989;
w23991 <= not w23210 and not w23639;
w23992 <= not w23220 and w23435;
w23993 <= not w23431 and w23992;
w23994 <= not w23432 and not w23435;
w23995 <= not w23993 and not w23994;
w23996 <= w23638 and not w23995;
w23997 <= not w23637 and w23996;
w23998 <= not w23991 and not w23997;
w23999 <= not b(18) and not w23998;
w24000 <= not w23219 and not w23639;
w24001 <= not w23229 and w23430;
w24002 <= not w23426 and w24001;
w24003 <= not w23427 and not w23430;
w24004 <= not w24002 and not w24003;
w24005 <= w23638 and not w24004;
w24006 <= not w23637 and w24005;
w24007 <= not w24000 and not w24006;
w24008 <= not b(17) and not w24007;
w24009 <= not w23228 and not w23639;
w24010 <= not w23238 and w23425;
w24011 <= not w23421 and w24010;
w24012 <= not w23422 and not w23425;
w24013 <= not w24011 and not w24012;
w24014 <= w23638 and not w24013;
w24015 <= not w23637 and w24014;
w24016 <= not w24009 and not w24015;
w24017 <= not b(16) and not w24016;
w24018 <= not w23237 and not w23639;
w24019 <= not w23247 and w23420;
w24020 <= not w23416 and w24019;
w24021 <= not w23417 and not w23420;
w24022 <= not w24020 and not w24021;
w24023 <= w23638 and not w24022;
w24024 <= not w23637 and w24023;
w24025 <= not w24018 and not w24024;
w24026 <= not b(15) and not w24025;
w24027 <= not w23246 and not w23639;
w24028 <= not w23256 and w23415;
w24029 <= not w23411 and w24028;
w24030 <= not w23412 and not w23415;
w24031 <= not w24029 and not w24030;
w24032 <= w23638 and not w24031;
w24033 <= not w23637 and w24032;
w24034 <= not w24027 and not w24033;
w24035 <= not b(14) and not w24034;
w24036 <= not w23255 and not w23639;
w24037 <= not w23265 and w23410;
w24038 <= not w23406 and w24037;
w24039 <= not w23407 and not w23410;
w24040 <= not w24038 and not w24039;
w24041 <= w23638 and not w24040;
w24042 <= not w23637 and w24041;
w24043 <= not w24036 and not w24042;
w24044 <= not b(13) and not w24043;
w24045 <= not w23264 and not w23639;
w24046 <= not w23274 and w23405;
w24047 <= not w23401 and w24046;
w24048 <= not w23402 and not w23405;
w24049 <= not w24047 and not w24048;
w24050 <= w23638 and not w24049;
w24051 <= not w23637 and w24050;
w24052 <= not w24045 and not w24051;
w24053 <= not b(12) and not w24052;
w24054 <= not w23273 and not w23639;
w24055 <= not w23283 and w23400;
w24056 <= not w23396 and w24055;
w24057 <= not w23397 and not w23400;
w24058 <= not w24056 and not w24057;
w24059 <= w23638 and not w24058;
w24060 <= not w23637 and w24059;
w24061 <= not w24054 and not w24060;
w24062 <= not b(11) and not w24061;
w24063 <= not w23282 and not w23639;
w24064 <= not w23292 and w23395;
w24065 <= not w23391 and w24064;
w24066 <= not w23392 and not w23395;
w24067 <= not w24065 and not w24066;
w24068 <= w23638 and not w24067;
w24069 <= not w23637 and w24068;
w24070 <= not w24063 and not w24069;
w24071 <= not b(10) and not w24070;
w24072 <= not w23291 and not w23639;
w24073 <= not w23301 and w23390;
w24074 <= not w23386 and w24073;
w24075 <= not w23387 and not w23390;
w24076 <= not w24074 and not w24075;
w24077 <= w23638 and not w24076;
w24078 <= not w23637 and w24077;
w24079 <= not w24072 and not w24078;
w24080 <= not b(9) and not w24079;
w24081 <= not w23300 and not w23639;
w24082 <= not w23310 and w23385;
w24083 <= not w23381 and w24082;
w24084 <= not w23382 and not w23385;
w24085 <= not w24083 and not w24084;
w24086 <= w23638 and not w24085;
w24087 <= not w23637 and w24086;
w24088 <= not w24081 and not w24087;
w24089 <= not b(8) and not w24088;
w24090 <= not w23309 and not w23639;
w24091 <= not w23319 and w23380;
w24092 <= not w23376 and w24091;
w24093 <= not w23377 and not w23380;
w24094 <= not w24092 and not w24093;
w24095 <= w23638 and not w24094;
w24096 <= not w23637 and w24095;
w24097 <= not w24090 and not w24096;
w24098 <= not b(7) and not w24097;
w24099 <= not w23318 and not w23639;
w24100 <= not w23328 and w23375;
w24101 <= not w23371 and w24100;
w24102 <= not w23372 and not w23375;
w24103 <= not w24101 and not w24102;
w24104 <= w23638 and not w24103;
w24105 <= not w23637 and w24104;
w24106 <= not w24099 and not w24105;
w24107 <= not b(6) and not w24106;
w24108 <= not w23327 and not w23639;
w24109 <= not w23337 and w23370;
w24110 <= not w23366 and w24109;
w24111 <= not w23367 and not w23370;
w24112 <= not w24110 and not w24111;
w24113 <= w23638 and not w24112;
w24114 <= not w23637 and w24113;
w24115 <= not w24108 and not w24114;
w24116 <= not b(5) and not w24115;
w24117 <= not w23336 and not w23639;
w24118 <= not w23345 and w23365;
w24119 <= not w23361 and w24118;
w24120 <= not w23362 and not w23365;
w24121 <= not w24119 and not w24120;
w24122 <= w23638 and not w24121;
w24123 <= not w23637 and w24122;
w24124 <= not w24117 and not w24123;
w24125 <= not b(4) and not w24124;
w24126 <= not w23344 and not w23639;
w24127 <= not w23356 and w23360;
w24128 <= not w23355 and w24127;
w24129 <= not w23357 and not w23360;
w24130 <= not w24128 and not w24129;
w24131 <= w23638 and not w24130;
w24132 <= not w23637 and w24131;
w24133 <= not w24126 and not w24132;
w24134 <= not b(3) and not w24133;
w24135 <= not w23349 and not w23639;
w24136 <= not w23352 and w23354;
w24137 <= not w23350 and w24136;
w24138 <= w23638 and not w24137;
w24139 <= not w23355 and w24138;
w24140 <= not w23637 and w24139;
w24141 <= not w24135 and not w24140;
w24142 <= not b(2) and not w24141;
w24143 <= b(0) and not b(58);
w24144 <= w148 and w24143;
w24145 <= w146 and w24144;
w24146 <= not w23637 and w24145;
w24147 <= a(6) and not w24146;
w24148 <= w25 and w23354;
w24149 <= w23 and w24148;
w24150 <= not w23637 and w24149;
w24151 <= not w24147 and not w24150;
w24152 <= b(1) and not w24151;
w24153 <= not b(1) and not w24150;
w24154 <= not w24147 and w24153;
w24155 <= not w24152 and not w24154;
w24156 <= not a(5) and b(0);
w24157 <= not w24155 and not w24156;
w24158 <= not b(1) and not w24151;
w24159 <= not w24157 and not w24158;
w24160 <= b(2) and not w24140;
w24161 <= not w24135 and w24160;
w24162 <= not w24142 and not w24161;
w24163 <= not w24159 and w24162;
w24164 <= not w24142 and not w24163;
w24165 <= b(3) and not w24132;
w24166 <= not w24126 and w24165;
w24167 <= not w24134 and not w24166;
w24168 <= not w24164 and w24167;
w24169 <= not w24134 and not w24168;
w24170 <= b(4) and not w24123;
w24171 <= not w24117 and w24170;
w24172 <= not w24125 and not w24171;
w24173 <= not w24169 and w24172;
w24174 <= not w24125 and not w24173;
w24175 <= b(5) and not w24114;
w24176 <= not w24108 and w24175;
w24177 <= not w24116 and not w24176;
w24178 <= not w24174 and w24177;
w24179 <= not w24116 and not w24178;
w24180 <= b(6) and not w24105;
w24181 <= not w24099 and w24180;
w24182 <= not w24107 and not w24181;
w24183 <= not w24179 and w24182;
w24184 <= not w24107 and not w24183;
w24185 <= b(7) and not w24096;
w24186 <= not w24090 and w24185;
w24187 <= not w24098 and not w24186;
w24188 <= not w24184 and w24187;
w24189 <= not w24098 and not w24188;
w24190 <= b(8) and not w24087;
w24191 <= not w24081 and w24190;
w24192 <= not w24089 and not w24191;
w24193 <= not w24189 and w24192;
w24194 <= not w24089 and not w24193;
w24195 <= b(9) and not w24078;
w24196 <= not w24072 and w24195;
w24197 <= not w24080 and not w24196;
w24198 <= not w24194 and w24197;
w24199 <= not w24080 and not w24198;
w24200 <= b(10) and not w24069;
w24201 <= not w24063 and w24200;
w24202 <= not w24071 and not w24201;
w24203 <= not w24199 and w24202;
w24204 <= not w24071 and not w24203;
w24205 <= b(11) and not w24060;
w24206 <= not w24054 and w24205;
w24207 <= not w24062 and not w24206;
w24208 <= not w24204 and w24207;
w24209 <= not w24062 and not w24208;
w24210 <= b(12) and not w24051;
w24211 <= not w24045 and w24210;
w24212 <= not w24053 and not w24211;
w24213 <= not w24209 and w24212;
w24214 <= not w24053 and not w24213;
w24215 <= b(13) and not w24042;
w24216 <= not w24036 and w24215;
w24217 <= not w24044 and not w24216;
w24218 <= not w24214 and w24217;
w24219 <= not w24044 and not w24218;
w24220 <= b(14) and not w24033;
w24221 <= not w24027 and w24220;
w24222 <= not w24035 and not w24221;
w24223 <= not w24219 and w24222;
w24224 <= not w24035 and not w24223;
w24225 <= b(15) and not w24024;
w24226 <= not w24018 and w24225;
w24227 <= not w24026 and not w24226;
w24228 <= not w24224 and w24227;
w24229 <= not w24026 and not w24228;
w24230 <= b(16) and not w24015;
w24231 <= not w24009 and w24230;
w24232 <= not w24017 and not w24231;
w24233 <= not w24229 and w24232;
w24234 <= not w24017 and not w24233;
w24235 <= b(17) and not w24006;
w24236 <= not w24000 and w24235;
w24237 <= not w24008 and not w24236;
w24238 <= not w24234 and w24237;
w24239 <= not w24008 and not w24238;
w24240 <= b(18) and not w23997;
w24241 <= not w23991 and w24240;
w24242 <= not w23999 and not w24241;
w24243 <= not w24239 and w24242;
w24244 <= not w23999 and not w24243;
w24245 <= b(19) and not w23988;
w24246 <= not w23982 and w24245;
w24247 <= not w23990 and not w24246;
w24248 <= not w24244 and w24247;
w24249 <= not w23990 and not w24248;
w24250 <= b(20) and not w23979;
w24251 <= not w23973 and w24250;
w24252 <= not w23981 and not w24251;
w24253 <= not w24249 and w24252;
w24254 <= not w23981 and not w24253;
w24255 <= b(21) and not w23970;
w24256 <= not w23964 and w24255;
w24257 <= not w23972 and not w24256;
w24258 <= not w24254 and w24257;
w24259 <= not w23972 and not w24258;
w24260 <= b(22) and not w23961;
w24261 <= not w23955 and w24260;
w24262 <= not w23963 and not w24261;
w24263 <= not w24259 and w24262;
w24264 <= not w23963 and not w24263;
w24265 <= b(23) and not w23952;
w24266 <= not w23946 and w24265;
w24267 <= not w23954 and not w24266;
w24268 <= not w24264 and w24267;
w24269 <= not w23954 and not w24268;
w24270 <= b(24) and not w23943;
w24271 <= not w23937 and w24270;
w24272 <= not w23945 and not w24271;
w24273 <= not w24269 and w24272;
w24274 <= not w23945 and not w24273;
w24275 <= b(25) and not w23934;
w24276 <= not w23928 and w24275;
w24277 <= not w23936 and not w24276;
w24278 <= not w24274 and w24277;
w24279 <= not w23936 and not w24278;
w24280 <= b(26) and not w23925;
w24281 <= not w23919 and w24280;
w24282 <= not w23927 and not w24281;
w24283 <= not w24279 and w24282;
w24284 <= not w23927 and not w24283;
w24285 <= b(27) and not w23916;
w24286 <= not w23910 and w24285;
w24287 <= not w23918 and not w24286;
w24288 <= not w24284 and w24287;
w24289 <= not w23918 and not w24288;
w24290 <= b(28) and not w23907;
w24291 <= not w23901 and w24290;
w24292 <= not w23909 and not w24291;
w24293 <= not w24289 and w24292;
w24294 <= not w23909 and not w24293;
w24295 <= b(29) and not w23898;
w24296 <= not w23892 and w24295;
w24297 <= not w23900 and not w24296;
w24298 <= not w24294 and w24297;
w24299 <= not w23900 and not w24298;
w24300 <= b(30) and not w23889;
w24301 <= not w23883 and w24300;
w24302 <= not w23891 and not w24301;
w24303 <= not w24299 and w24302;
w24304 <= not w23891 and not w24303;
w24305 <= b(31) and not w23880;
w24306 <= not w23874 and w24305;
w24307 <= not w23882 and not w24306;
w24308 <= not w24304 and w24307;
w24309 <= not w23882 and not w24308;
w24310 <= b(32) and not w23871;
w24311 <= not w23865 and w24310;
w24312 <= not w23873 and not w24311;
w24313 <= not w24309 and w24312;
w24314 <= not w23873 and not w24313;
w24315 <= b(33) and not w23862;
w24316 <= not w23856 and w24315;
w24317 <= not w23864 and not w24316;
w24318 <= not w24314 and w24317;
w24319 <= not w23864 and not w24318;
w24320 <= b(34) and not w23853;
w24321 <= not w23847 and w24320;
w24322 <= not w23855 and not w24321;
w24323 <= not w24319 and w24322;
w24324 <= not w23855 and not w24323;
w24325 <= b(35) and not w23844;
w24326 <= not w23838 and w24325;
w24327 <= not w23846 and not w24326;
w24328 <= not w24324 and w24327;
w24329 <= not w23846 and not w24328;
w24330 <= b(36) and not w23835;
w24331 <= not w23829 and w24330;
w24332 <= not w23837 and not w24331;
w24333 <= not w24329 and w24332;
w24334 <= not w23837 and not w24333;
w24335 <= b(37) and not w23826;
w24336 <= not w23820 and w24335;
w24337 <= not w23828 and not w24336;
w24338 <= not w24334 and w24337;
w24339 <= not w23828 and not w24338;
w24340 <= b(38) and not w23817;
w24341 <= not w23811 and w24340;
w24342 <= not w23819 and not w24341;
w24343 <= not w24339 and w24342;
w24344 <= not w23819 and not w24343;
w24345 <= b(39) and not w23808;
w24346 <= not w23802 and w24345;
w24347 <= not w23810 and not w24346;
w24348 <= not w24344 and w24347;
w24349 <= not w23810 and not w24348;
w24350 <= b(40) and not w23799;
w24351 <= not w23793 and w24350;
w24352 <= not w23801 and not w24351;
w24353 <= not w24349 and w24352;
w24354 <= not w23801 and not w24353;
w24355 <= b(41) and not w23790;
w24356 <= not w23784 and w24355;
w24357 <= not w23792 and not w24356;
w24358 <= not w24354 and w24357;
w24359 <= not w23792 and not w24358;
w24360 <= b(42) and not w23781;
w24361 <= not w23775 and w24360;
w24362 <= not w23783 and not w24361;
w24363 <= not w24359 and w24362;
w24364 <= not w23783 and not w24363;
w24365 <= b(43) and not w23772;
w24366 <= not w23766 and w24365;
w24367 <= not w23774 and not w24366;
w24368 <= not w24364 and w24367;
w24369 <= not w23774 and not w24368;
w24370 <= b(44) and not w23763;
w24371 <= not w23757 and w24370;
w24372 <= not w23765 and not w24371;
w24373 <= not w24369 and w24372;
w24374 <= not w23765 and not w24373;
w24375 <= b(45) and not w23754;
w24376 <= not w23748 and w24375;
w24377 <= not w23756 and not w24376;
w24378 <= not w24374 and w24377;
w24379 <= not w23756 and not w24378;
w24380 <= b(46) and not w23745;
w24381 <= not w23739 and w24380;
w24382 <= not w23747 and not w24381;
w24383 <= not w24379 and w24382;
w24384 <= not w23747 and not w24383;
w24385 <= b(47) and not w23736;
w24386 <= not w23730 and w24385;
w24387 <= not w23738 and not w24386;
w24388 <= not w24384 and w24387;
w24389 <= not w23738 and not w24388;
w24390 <= b(48) and not w23727;
w24391 <= not w23721 and w24390;
w24392 <= not w23729 and not w24391;
w24393 <= not w24389 and w24392;
w24394 <= not w23729 and not w24393;
w24395 <= b(49) and not w23718;
w24396 <= not w23712 and w24395;
w24397 <= not w23720 and not w24396;
w24398 <= not w24394 and w24397;
w24399 <= not w23720 and not w24398;
w24400 <= b(50) and not w23709;
w24401 <= not w23703 and w24400;
w24402 <= not w23711 and not w24401;
w24403 <= not w24399 and w24402;
w24404 <= not w23711 and not w24403;
w24405 <= b(51) and not w23700;
w24406 <= not w23694 and w24405;
w24407 <= not w23702 and not w24406;
w24408 <= not w24404 and w24407;
w24409 <= not w23702 and not w24408;
w24410 <= b(52) and not w23691;
w24411 <= not w23685 and w24410;
w24412 <= not w23693 and not w24411;
w24413 <= not w24409 and w24412;
w24414 <= not w23693 and not w24413;
w24415 <= b(53) and not w23682;
w24416 <= not w23676 and w24415;
w24417 <= not w23684 and not w24416;
w24418 <= not w24414 and w24417;
w24419 <= not w23684 and not w24418;
w24420 <= b(54) and not w23673;
w24421 <= not w23667 and w24420;
w24422 <= not w23675 and not w24421;
w24423 <= not w24419 and w24422;
w24424 <= not w23675 and not w24423;
w24425 <= b(55) and not w23664;
w24426 <= not w23658 and w24425;
w24427 <= not w23666 and not w24426;
w24428 <= not w24424 and w24427;
w24429 <= not w23666 and not w24428;
w24430 <= b(56) and not w23655;
w24431 <= not w23649 and w24430;
w24432 <= not w23657 and not w24431;
w24433 <= not w24429 and w24432;
w24434 <= not w23657 and not w24433;
w24435 <= b(57) and not w23646;
w24436 <= not w23640 and w24435;
w24437 <= not w23648 and not w24436;
w24438 <= not w24434 and w24437;
w24439 <= not w23648 and not w24438;
w24440 <= not w22858 and not w23639;
w24441 <= not w22860 and w23635;
w24442 <= not w23631 and w24441;
w24443 <= not w23632 and not w23635;
w24444 <= not w24442 and not w24443;
w24445 <= w23639 and not w24444;
w24446 <= not w24440 and not w24445;
w24447 <= not b(58) and not w24446;
w24448 <= b(58) and not w24440;
w24449 <= not w24445 and w24448;
w24450 <= w146 and w148;
w24451 <= not w24449 and w24450;
w24452 <= not w24447 and w24451;
w24453 <= not w24439 and w24452;
w24454 <= w23638 and not w24446;
w24455 <= not w24453 and not w24454;
w24456 <= not w23657 and w24437;
w24457 <= not w24433 and w24456;
w24458 <= not w24434 and not w24437;
w24459 <= not w24457 and not w24458;
w24460 <= not w24455 and not w24459;
w24461 <= not w23647 and not w24454;
w24462 <= not w24453 and w24461;
w24463 <= not w24460 and not w24462;
w24464 <= not b(58) and not w24463;
w24465 <= not w23666 and w24432;
w24466 <= not w24428 and w24465;
w24467 <= not w24429 and not w24432;
w24468 <= not w24466 and not w24467;
w24469 <= not w24455 and not w24468;
w24470 <= not w23656 and not w24454;
w24471 <= not w24453 and w24470;
w24472 <= not w24469 and not w24471;
w24473 <= not b(57) and not w24472;
w24474 <= not w23675 and w24427;
w24475 <= not w24423 and w24474;
w24476 <= not w24424 and not w24427;
w24477 <= not w24475 and not w24476;
w24478 <= not w24455 and not w24477;
w24479 <= not w23665 and not w24454;
w24480 <= not w24453 and w24479;
w24481 <= not w24478 and not w24480;
w24482 <= not b(56) and not w24481;
w24483 <= not w23684 and w24422;
w24484 <= not w24418 and w24483;
w24485 <= not w24419 and not w24422;
w24486 <= not w24484 and not w24485;
w24487 <= not w24455 and not w24486;
w24488 <= not w23674 and not w24454;
w24489 <= not w24453 and w24488;
w24490 <= not w24487 and not w24489;
w24491 <= not b(55) and not w24490;
w24492 <= not w23693 and w24417;
w24493 <= not w24413 and w24492;
w24494 <= not w24414 and not w24417;
w24495 <= not w24493 and not w24494;
w24496 <= not w24455 and not w24495;
w24497 <= not w23683 and not w24454;
w24498 <= not w24453 and w24497;
w24499 <= not w24496 and not w24498;
w24500 <= not b(54) and not w24499;
w24501 <= not w23702 and w24412;
w24502 <= not w24408 and w24501;
w24503 <= not w24409 and not w24412;
w24504 <= not w24502 and not w24503;
w24505 <= not w24455 and not w24504;
w24506 <= not w23692 and not w24454;
w24507 <= not w24453 and w24506;
w24508 <= not w24505 and not w24507;
w24509 <= not b(53) and not w24508;
w24510 <= not w23711 and w24407;
w24511 <= not w24403 and w24510;
w24512 <= not w24404 and not w24407;
w24513 <= not w24511 and not w24512;
w24514 <= not w24455 and not w24513;
w24515 <= not w23701 and not w24454;
w24516 <= not w24453 and w24515;
w24517 <= not w24514 and not w24516;
w24518 <= not b(52) and not w24517;
w24519 <= not w23720 and w24402;
w24520 <= not w24398 and w24519;
w24521 <= not w24399 and not w24402;
w24522 <= not w24520 and not w24521;
w24523 <= not w24455 and not w24522;
w24524 <= not w23710 and not w24454;
w24525 <= not w24453 and w24524;
w24526 <= not w24523 and not w24525;
w24527 <= not b(51) and not w24526;
w24528 <= not w23729 and w24397;
w24529 <= not w24393 and w24528;
w24530 <= not w24394 and not w24397;
w24531 <= not w24529 and not w24530;
w24532 <= not w24455 and not w24531;
w24533 <= not w23719 and not w24454;
w24534 <= not w24453 and w24533;
w24535 <= not w24532 and not w24534;
w24536 <= not b(50) and not w24535;
w24537 <= not w23738 and w24392;
w24538 <= not w24388 and w24537;
w24539 <= not w24389 and not w24392;
w24540 <= not w24538 and not w24539;
w24541 <= not w24455 and not w24540;
w24542 <= not w23728 and not w24454;
w24543 <= not w24453 and w24542;
w24544 <= not w24541 and not w24543;
w24545 <= not b(49) and not w24544;
w24546 <= not w23747 and w24387;
w24547 <= not w24383 and w24546;
w24548 <= not w24384 and not w24387;
w24549 <= not w24547 and not w24548;
w24550 <= not w24455 and not w24549;
w24551 <= not w23737 and not w24454;
w24552 <= not w24453 and w24551;
w24553 <= not w24550 and not w24552;
w24554 <= not b(48) and not w24553;
w24555 <= not w23756 and w24382;
w24556 <= not w24378 and w24555;
w24557 <= not w24379 and not w24382;
w24558 <= not w24556 and not w24557;
w24559 <= not w24455 and not w24558;
w24560 <= not w23746 and not w24454;
w24561 <= not w24453 and w24560;
w24562 <= not w24559 and not w24561;
w24563 <= not b(47) and not w24562;
w24564 <= not w23765 and w24377;
w24565 <= not w24373 and w24564;
w24566 <= not w24374 and not w24377;
w24567 <= not w24565 and not w24566;
w24568 <= not w24455 and not w24567;
w24569 <= not w23755 and not w24454;
w24570 <= not w24453 and w24569;
w24571 <= not w24568 and not w24570;
w24572 <= not b(46) and not w24571;
w24573 <= not w23774 and w24372;
w24574 <= not w24368 and w24573;
w24575 <= not w24369 and not w24372;
w24576 <= not w24574 and not w24575;
w24577 <= not w24455 and not w24576;
w24578 <= not w23764 and not w24454;
w24579 <= not w24453 and w24578;
w24580 <= not w24577 and not w24579;
w24581 <= not b(45) and not w24580;
w24582 <= not w23783 and w24367;
w24583 <= not w24363 and w24582;
w24584 <= not w24364 and not w24367;
w24585 <= not w24583 and not w24584;
w24586 <= not w24455 and not w24585;
w24587 <= not w23773 and not w24454;
w24588 <= not w24453 and w24587;
w24589 <= not w24586 and not w24588;
w24590 <= not b(44) and not w24589;
w24591 <= not w23792 and w24362;
w24592 <= not w24358 and w24591;
w24593 <= not w24359 and not w24362;
w24594 <= not w24592 and not w24593;
w24595 <= not w24455 and not w24594;
w24596 <= not w23782 and not w24454;
w24597 <= not w24453 and w24596;
w24598 <= not w24595 and not w24597;
w24599 <= not b(43) and not w24598;
w24600 <= not w23801 and w24357;
w24601 <= not w24353 and w24600;
w24602 <= not w24354 and not w24357;
w24603 <= not w24601 and not w24602;
w24604 <= not w24455 and not w24603;
w24605 <= not w23791 and not w24454;
w24606 <= not w24453 and w24605;
w24607 <= not w24604 and not w24606;
w24608 <= not b(42) and not w24607;
w24609 <= not w23810 and w24352;
w24610 <= not w24348 and w24609;
w24611 <= not w24349 and not w24352;
w24612 <= not w24610 and not w24611;
w24613 <= not w24455 and not w24612;
w24614 <= not w23800 and not w24454;
w24615 <= not w24453 and w24614;
w24616 <= not w24613 and not w24615;
w24617 <= not b(41) and not w24616;
w24618 <= not w23819 and w24347;
w24619 <= not w24343 and w24618;
w24620 <= not w24344 and not w24347;
w24621 <= not w24619 and not w24620;
w24622 <= not w24455 and not w24621;
w24623 <= not w23809 and not w24454;
w24624 <= not w24453 and w24623;
w24625 <= not w24622 and not w24624;
w24626 <= not b(40) and not w24625;
w24627 <= not w23828 and w24342;
w24628 <= not w24338 and w24627;
w24629 <= not w24339 and not w24342;
w24630 <= not w24628 and not w24629;
w24631 <= not w24455 and not w24630;
w24632 <= not w23818 and not w24454;
w24633 <= not w24453 and w24632;
w24634 <= not w24631 and not w24633;
w24635 <= not b(39) and not w24634;
w24636 <= not w23837 and w24337;
w24637 <= not w24333 and w24636;
w24638 <= not w24334 and not w24337;
w24639 <= not w24637 and not w24638;
w24640 <= not w24455 and not w24639;
w24641 <= not w23827 and not w24454;
w24642 <= not w24453 and w24641;
w24643 <= not w24640 and not w24642;
w24644 <= not b(38) and not w24643;
w24645 <= not w23846 and w24332;
w24646 <= not w24328 and w24645;
w24647 <= not w24329 and not w24332;
w24648 <= not w24646 and not w24647;
w24649 <= not w24455 and not w24648;
w24650 <= not w23836 and not w24454;
w24651 <= not w24453 and w24650;
w24652 <= not w24649 and not w24651;
w24653 <= not b(37) and not w24652;
w24654 <= not w23855 and w24327;
w24655 <= not w24323 and w24654;
w24656 <= not w24324 and not w24327;
w24657 <= not w24655 and not w24656;
w24658 <= not w24455 and not w24657;
w24659 <= not w23845 and not w24454;
w24660 <= not w24453 and w24659;
w24661 <= not w24658 and not w24660;
w24662 <= not b(36) and not w24661;
w24663 <= not w23864 and w24322;
w24664 <= not w24318 and w24663;
w24665 <= not w24319 and not w24322;
w24666 <= not w24664 and not w24665;
w24667 <= not w24455 and not w24666;
w24668 <= not w23854 and not w24454;
w24669 <= not w24453 and w24668;
w24670 <= not w24667 and not w24669;
w24671 <= not b(35) and not w24670;
w24672 <= not w23873 and w24317;
w24673 <= not w24313 and w24672;
w24674 <= not w24314 and not w24317;
w24675 <= not w24673 and not w24674;
w24676 <= not w24455 and not w24675;
w24677 <= not w23863 and not w24454;
w24678 <= not w24453 and w24677;
w24679 <= not w24676 and not w24678;
w24680 <= not b(34) and not w24679;
w24681 <= not w23882 and w24312;
w24682 <= not w24308 and w24681;
w24683 <= not w24309 and not w24312;
w24684 <= not w24682 and not w24683;
w24685 <= not w24455 and not w24684;
w24686 <= not w23872 and not w24454;
w24687 <= not w24453 and w24686;
w24688 <= not w24685 and not w24687;
w24689 <= not b(33) and not w24688;
w24690 <= not w23891 and w24307;
w24691 <= not w24303 and w24690;
w24692 <= not w24304 and not w24307;
w24693 <= not w24691 and not w24692;
w24694 <= not w24455 and not w24693;
w24695 <= not w23881 and not w24454;
w24696 <= not w24453 and w24695;
w24697 <= not w24694 and not w24696;
w24698 <= not b(32) and not w24697;
w24699 <= not w23900 and w24302;
w24700 <= not w24298 and w24699;
w24701 <= not w24299 and not w24302;
w24702 <= not w24700 and not w24701;
w24703 <= not w24455 and not w24702;
w24704 <= not w23890 and not w24454;
w24705 <= not w24453 and w24704;
w24706 <= not w24703 and not w24705;
w24707 <= not b(31) and not w24706;
w24708 <= not w23909 and w24297;
w24709 <= not w24293 and w24708;
w24710 <= not w24294 and not w24297;
w24711 <= not w24709 and not w24710;
w24712 <= not w24455 and not w24711;
w24713 <= not w23899 and not w24454;
w24714 <= not w24453 and w24713;
w24715 <= not w24712 and not w24714;
w24716 <= not b(30) and not w24715;
w24717 <= not w23918 and w24292;
w24718 <= not w24288 and w24717;
w24719 <= not w24289 and not w24292;
w24720 <= not w24718 and not w24719;
w24721 <= not w24455 and not w24720;
w24722 <= not w23908 and not w24454;
w24723 <= not w24453 and w24722;
w24724 <= not w24721 and not w24723;
w24725 <= not b(29) and not w24724;
w24726 <= not w23927 and w24287;
w24727 <= not w24283 and w24726;
w24728 <= not w24284 and not w24287;
w24729 <= not w24727 and not w24728;
w24730 <= not w24455 and not w24729;
w24731 <= not w23917 and not w24454;
w24732 <= not w24453 and w24731;
w24733 <= not w24730 and not w24732;
w24734 <= not b(28) and not w24733;
w24735 <= not w23936 and w24282;
w24736 <= not w24278 and w24735;
w24737 <= not w24279 and not w24282;
w24738 <= not w24736 and not w24737;
w24739 <= not w24455 and not w24738;
w24740 <= not w23926 and not w24454;
w24741 <= not w24453 and w24740;
w24742 <= not w24739 and not w24741;
w24743 <= not b(27) and not w24742;
w24744 <= not w23945 and w24277;
w24745 <= not w24273 and w24744;
w24746 <= not w24274 and not w24277;
w24747 <= not w24745 and not w24746;
w24748 <= not w24455 and not w24747;
w24749 <= not w23935 and not w24454;
w24750 <= not w24453 and w24749;
w24751 <= not w24748 and not w24750;
w24752 <= not b(26) and not w24751;
w24753 <= not w23954 and w24272;
w24754 <= not w24268 and w24753;
w24755 <= not w24269 and not w24272;
w24756 <= not w24754 and not w24755;
w24757 <= not w24455 and not w24756;
w24758 <= not w23944 and not w24454;
w24759 <= not w24453 and w24758;
w24760 <= not w24757 and not w24759;
w24761 <= not b(25) and not w24760;
w24762 <= not w23963 and w24267;
w24763 <= not w24263 and w24762;
w24764 <= not w24264 and not w24267;
w24765 <= not w24763 and not w24764;
w24766 <= not w24455 and not w24765;
w24767 <= not w23953 and not w24454;
w24768 <= not w24453 and w24767;
w24769 <= not w24766 and not w24768;
w24770 <= not b(24) and not w24769;
w24771 <= not w23972 and w24262;
w24772 <= not w24258 and w24771;
w24773 <= not w24259 and not w24262;
w24774 <= not w24772 and not w24773;
w24775 <= not w24455 and not w24774;
w24776 <= not w23962 and not w24454;
w24777 <= not w24453 and w24776;
w24778 <= not w24775 and not w24777;
w24779 <= not b(23) and not w24778;
w24780 <= not w23981 and w24257;
w24781 <= not w24253 and w24780;
w24782 <= not w24254 and not w24257;
w24783 <= not w24781 and not w24782;
w24784 <= not w24455 and not w24783;
w24785 <= not w23971 and not w24454;
w24786 <= not w24453 and w24785;
w24787 <= not w24784 and not w24786;
w24788 <= not b(22) and not w24787;
w24789 <= not w23990 and w24252;
w24790 <= not w24248 and w24789;
w24791 <= not w24249 and not w24252;
w24792 <= not w24790 and not w24791;
w24793 <= not w24455 and not w24792;
w24794 <= not w23980 and not w24454;
w24795 <= not w24453 and w24794;
w24796 <= not w24793 and not w24795;
w24797 <= not b(21) and not w24796;
w24798 <= not w23999 and w24247;
w24799 <= not w24243 and w24798;
w24800 <= not w24244 and not w24247;
w24801 <= not w24799 and not w24800;
w24802 <= not w24455 and not w24801;
w24803 <= not w23989 and not w24454;
w24804 <= not w24453 and w24803;
w24805 <= not w24802 and not w24804;
w24806 <= not b(20) and not w24805;
w24807 <= not w24008 and w24242;
w24808 <= not w24238 and w24807;
w24809 <= not w24239 and not w24242;
w24810 <= not w24808 and not w24809;
w24811 <= not w24455 and not w24810;
w24812 <= not w23998 and not w24454;
w24813 <= not w24453 and w24812;
w24814 <= not w24811 and not w24813;
w24815 <= not b(19) and not w24814;
w24816 <= not w24017 and w24237;
w24817 <= not w24233 and w24816;
w24818 <= not w24234 and not w24237;
w24819 <= not w24817 and not w24818;
w24820 <= not w24455 and not w24819;
w24821 <= not w24007 and not w24454;
w24822 <= not w24453 and w24821;
w24823 <= not w24820 and not w24822;
w24824 <= not b(18) and not w24823;
w24825 <= not w24026 and w24232;
w24826 <= not w24228 and w24825;
w24827 <= not w24229 and not w24232;
w24828 <= not w24826 and not w24827;
w24829 <= not w24455 and not w24828;
w24830 <= not w24016 and not w24454;
w24831 <= not w24453 and w24830;
w24832 <= not w24829 and not w24831;
w24833 <= not b(17) and not w24832;
w24834 <= not w24035 and w24227;
w24835 <= not w24223 and w24834;
w24836 <= not w24224 and not w24227;
w24837 <= not w24835 and not w24836;
w24838 <= not w24455 and not w24837;
w24839 <= not w24025 and not w24454;
w24840 <= not w24453 and w24839;
w24841 <= not w24838 and not w24840;
w24842 <= not b(16) and not w24841;
w24843 <= not w24044 and w24222;
w24844 <= not w24218 and w24843;
w24845 <= not w24219 and not w24222;
w24846 <= not w24844 and not w24845;
w24847 <= not w24455 and not w24846;
w24848 <= not w24034 and not w24454;
w24849 <= not w24453 and w24848;
w24850 <= not w24847 and not w24849;
w24851 <= not b(15) and not w24850;
w24852 <= not w24053 and w24217;
w24853 <= not w24213 and w24852;
w24854 <= not w24214 and not w24217;
w24855 <= not w24853 and not w24854;
w24856 <= not w24455 and not w24855;
w24857 <= not w24043 and not w24454;
w24858 <= not w24453 and w24857;
w24859 <= not w24856 and not w24858;
w24860 <= not b(14) and not w24859;
w24861 <= not w24062 and w24212;
w24862 <= not w24208 and w24861;
w24863 <= not w24209 and not w24212;
w24864 <= not w24862 and not w24863;
w24865 <= not w24455 and not w24864;
w24866 <= not w24052 and not w24454;
w24867 <= not w24453 and w24866;
w24868 <= not w24865 and not w24867;
w24869 <= not b(13) and not w24868;
w24870 <= not w24071 and w24207;
w24871 <= not w24203 and w24870;
w24872 <= not w24204 and not w24207;
w24873 <= not w24871 and not w24872;
w24874 <= not w24455 and not w24873;
w24875 <= not w24061 and not w24454;
w24876 <= not w24453 and w24875;
w24877 <= not w24874 and not w24876;
w24878 <= not b(12) and not w24877;
w24879 <= not w24080 and w24202;
w24880 <= not w24198 and w24879;
w24881 <= not w24199 and not w24202;
w24882 <= not w24880 and not w24881;
w24883 <= not w24455 and not w24882;
w24884 <= not w24070 and not w24454;
w24885 <= not w24453 and w24884;
w24886 <= not w24883 and not w24885;
w24887 <= not b(11) and not w24886;
w24888 <= not w24089 and w24197;
w24889 <= not w24193 and w24888;
w24890 <= not w24194 and not w24197;
w24891 <= not w24889 and not w24890;
w24892 <= not w24455 and not w24891;
w24893 <= not w24079 and not w24454;
w24894 <= not w24453 and w24893;
w24895 <= not w24892 and not w24894;
w24896 <= not b(10) and not w24895;
w24897 <= not w24098 and w24192;
w24898 <= not w24188 and w24897;
w24899 <= not w24189 and not w24192;
w24900 <= not w24898 and not w24899;
w24901 <= not w24455 and not w24900;
w24902 <= not w24088 and not w24454;
w24903 <= not w24453 and w24902;
w24904 <= not w24901 and not w24903;
w24905 <= not b(9) and not w24904;
w24906 <= not w24107 and w24187;
w24907 <= not w24183 and w24906;
w24908 <= not w24184 and not w24187;
w24909 <= not w24907 and not w24908;
w24910 <= not w24455 and not w24909;
w24911 <= not w24097 and not w24454;
w24912 <= not w24453 and w24911;
w24913 <= not w24910 and not w24912;
w24914 <= not b(8) and not w24913;
w24915 <= not w24116 and w24182;
w24916 <= not w24178 and w24915;
w24917 <= not w24179 and not w24182;
w24918 <= not w24916 and not w24917;
w24919 <= not w24455 and not w24918;
w24920 <= not w24106 and not w24454;
w24921 <= not w24453 and w24920;
w24922 <= not w24919 and not w24921;
w24923 <= not b(7) and not w24922;
w24924 <= not w24125 and w24177;
w24925 <= not w24173 and w24924;
w24926 <= not w24174 and not w24177;
w24927 <= not w24925 and not w24926;
w24928 <= not w24455 and not w24927;
w24929 <= not w24115 and not w24454;
w24930 <= not w24453 and w24929;
w24931 <= not w24928 and not w24930;
w24932 <= not b(6) and not w24931;
w24933 <= not w24134 and w24172;
w24934 <= not w24168 and w24933;
w24935 <= not w24169 and not w24172;
w24936 <= not w24934 and not w24935;
w24937 <= not w24455 and not w24936;
w24938 <= not w24124 and not w24454;
w24939 <= not w24453 and w24938;
w24940 <= not w24937 and not w24939;
w24941 <= not b(5) and not w24940;
w24942 <= not w24142 and w24167;
w24943 <= not w24163 and w24942;
w24944 <= not w24164 and not w24167;
w24945 <= not w24943 and not w24944;
w24946 <= not w24455 and not w24945;
w24947 <= not w24133 and not w24454;
w24948 <= not w24453 and w24947;
w24949 <= not w24946 and not w24948;
w24950 <= not b(4) and not w24949;
w24951 <= not w24158 and w24162;
w24952 <= not w24157 and w24951;
w24953 <= not w24159 and not w24162;
w24954 <= not w24952 and not w24953;
w24955 <= not w24455 and not w24954;
w24956 <= not w24141 and not w24454;
w24957 <= not w24453 and w24956;
w24958 <= not w24955 and not w24957;
w24959 <= not b(3) and not w24958;
w24960 <= not w24154 and w24156;
w24961 <= not w24152 and w24960;
w24962 <= not w24157 and not w24961;
w24963 <= not w24455 and w24962;
w24964 <= not w24151 and not w24454;
w24965 <= not w24453 and w24964;
w24966 <= not w24963 and not w24965;
w24967 <= not b(2) and not w24966;
w24968 <= b(0) and not w24455;
w24969 <= a(5) and not w24968;
w24970 <= w24156 and not w24455;
w24971 <= not w24969 and not w24970;
w24972 <= b(1) and not w24971;
w24973 <= not b(1) and not w24970;
w24974 <= not w24969 and w24973;
w24975 <= not w24972 and not w24974;
w24976 <= not a(4) and b(0);
w24977 <= not w24975 and not w24976;
w24978 <= not b(1) and not w24971;
w24979 <= not w24977 and not w24978;
w24980 <= b(2) and not w24965;
w24981 <= not w24963 and w24980;
w24982 <= not w24967 and not w24981;
w24983 <= not w24979 and w24982;
w24984 <= not w24967 and not w24983;
w24985 <= b(3) and not w24957;
w24986 <= not w24955 and w24985;
w24987 <= not w24959 and not w24986;
w24988 <= not w24984 and w24987;
w24989 <= not w24959 and not w24988;
w24990 <= b(4) and not w24948;
w24991 <= not w24946 and w24990;
w24992 <= not w24950 and not w24991;
w24993 <= not w24989 and w24992;
w24994 <= not w24950 and not w24993;
w24995 <= b(5) and not w24939;
w24996 <= not w24937 and w24995;
w24997 <= not w24941 and not w24996;
w24998 <= not w24994 and w24997;
w24999 <= not w24941 and not w24998;
w25000 <= b(6) and not w24930;
w25001 <= not w24928 and w25000;
w25002 <= not w24932 and not w25001;
w25003 <= not w24999 and w25002;
w25004 <= not w24932 and not w25003;
w25005 <= b(7) and not w24921;
w25006 <= not w24919 and w25005;
w25007 <= not w24923 and not w25006;
w25008 <= not w25004 and w25007;
w25009 <= not w24923 and not w25008;
w25010 <= b(8) and not w24912;
w25011 <= not w24910 and w25010;
w25012 <= not w24914 and not w25011;
w25013 <= not w25009 and w25012;
w25014 <= not w24914 and not w25013;
w25015 <= b(9) and not w24903;
w25016 <= not w24901 and w25015;
w25017 <= not w24905 and not w25016;
w25018 <= not w25014 and w25017;
w25019 <= not w24905 and not w25018;
w25020 <= b(10) and not w24894;
w25021 <= not w24892 and w25020;
w25022 <= not w24896 and not w25021;
w25023 <= not w25019 and w25022;
w25024 <= not w24896 and not w25023;
w25025 <= b(11) and not w24885;
w25026 <= not w24883 and w25025;
w25027 <= not w24887 and not w25026;
w25028 <= not w25024 and w25027;
w25029 <= not w24887 and not w25028;
w25030 <= b(12) and not w24876;
w25031 <= not w24874 and w25030;
w25032 <= not w24878 and not w25031;
w25033 <= not w25029 and w25032;
w25034 <= not w24878 and not w25033;
w25035 <= b(13) and not w24867;
w25036 <= not w24865 and w25035;
w25037 <= not w24869 and not w25036;
w25038 <= not w25034 and w25037;
w25039 <= not w24869 and not w25038;
w25040 <= b(14) and not w24858;
w25041 <= not w24856 and w25040;
w25042 <= not w24860 and not w25041;
w25043 <= not w25039 and w25042;
w25044 <= not w24860 and not w25043;
w25045 <= b(15) and not w24849;
w25046 <= not w24847 and w25045;
w25047 <= not w24851 and not w25046;
w25048 <= not w25044 and w25047;
w25049 <= not w24851 and not w25048;
w25050 <= b(16) and not w24840;
w25051 <= not w24838 and w25050;
w25052 <= not w24842 and not w25051;
w25053 <= not w25049 and w25052;
w25054 <= not w24842 and not w25053;
w25055 <= b(17) and not w24831;
w25056 <= not w24829 and w25055;
w25057 <= not w24833 and not w25056;
w25058 <= not w25054 and w25057;
w25059 <= not w24833 and not w25058;
w25060 <= b(18) and not w24822;
w25061 <= not w24820 and w25060;
w25062 <= not w24824 and not w25061;
w25063 <= not w25059 and w25062;
w25064 <= not w24824 and not w25063;
w25065 <= b(19) and not w24813;
w25066 <= not w24811 and w25065;
w25067 <= not w24815 and not w25066;
w25068 <= not w25064 and w25067;
w25069 <= not w24815 and not w25068;
w25070 <= b(20) and not w24804;
w25071 <= not w24802 and w25070;
w25072 <= not w24806 and not w25071;
w25073 <= not w25069 and w25072;
w25074 <= not w24806 and not w25073;
w25075 <= b(21) and not w24795;
w25076 <= not w24793 and w25075;
w25077 <= not w24797 and not w25076;
w25078 <= not w25074 and w25077;
w25079 <= not w24797 and not w25078;
w25080 <= b(22) and not w24786;
w25081 <= not w24784 and w25080;
w25082 <= not w24788 and not w25081;
w25083 <= not w25079 and w25082;
w25084 <= not w24788 and not w25083;
w25085 <= b(23) and not w24777;
w25086 <= not w24775 and w25085;
w25087 <= not w24779 and not w25086;
w25088 <= not w25084 and w25087;
w25089 <= not w24779 and not w25088;
w25090 <= b(24) and not w24768;
w25091 <= not w24766 and w25090;
w25092 <= not w24770 and not w25091;
w25093 <= not w25089 and w25092;
w25094 <= not w24770 and not w25093;
w25095 <= b(25) and not w24759;
w25096 <= not w24757 and w25095;
w25097 <= not w24761 and not w25096;
w25098 <= not w25094 and w25097;
w25099 <= not w24761 and not w25098;
w25100 <= b(26) and not w24750;
w25101 <= not w24748 and w25100;
w25102 <= not w24752 and not w25101;
w25103 <= not w25099 and w25102;
w25104 <= not w24752 and not w25103;
w25105 <= b(27) and not w24741;
w25106 <= not w24739 and w25105;
w25107 <= not w24743 and not w25106;
w25108 <= not w25104 and w25107;
w25109 <= not w24743 and not w25108;
w25110 <= b(28) and not w24732;
w25111 <= not w24730 and w25110;
w25112 <= not w24734 and not w25111;
w25113 <= not w25109 and w25112;
w25114 <= not w24734 and not w25113;
w25115 <= b(29) and not w24723;
w25116 <= not w24721 and w25115;
w25117 <= not w24725 and not w25116;
w25118 <= not w25114 and w25117;
w25119 <= not w24725 and not w25118;
w25120 <= b(30) and not w24714;
w25121 <= not w24712 and w25120;
w25122 <= not w24716 and not w25121;
w25123 <= not w25119 and w25122;
w25124 <= not w24716 and not w25123;
w25125 <= b(31) and not w24705;
w25126 <= not w24703 and w25125;
w25127 <= not w24707 and not w25126;
w25128 <= not w25124 and w25127;
w25129 <= not w24707 and not w25128;
w25130 <= b(32) and not w24696;
w25131 <= not w24694 and w25130;
w25132 <= not w24698 and not w25131;
w25133 <= not w25129 and w25132;
w25134 <= not w24698 and not w25133;
w25135 <= b(33) and not w24687;
w25136 <= not w24685 and w25135;
w25137 <= not w24689 and not w25136;
w25138 <= not w25134 and w25137;
w25139 <= not w24689 and not w25138;
w25140 <= b(34) and not w24678;
w25141 <= not w24676 and w25140;
w25142 <= not w24680 and not w25141;
w25143 <= not w25139 and w25142;
w25144 <= not w24680 and not w25143;
w25145 <= b(35) and not w24669;
w25146 <= not w24667 and w25145;
w25147 <= not w24671 and not w25146;
w25148 <= not w25144 and w25147;
w25149 <= not w24671 and not w25148;
w25150 <= b(36) and not w24660;
w25151 <= not w24658 and w25150;
w25152 <= not w24662 and not w25151;
w25153 <= not w25149 and w25152;
w25154 <= not w24662 and not w25153;
w25155 <= b(37) and not w24651;
w25156 <= not w24649 and w25155;
w25157 <= not w24653 and not w25156;
w25158 <= not w25154 and w25157;
w25159 <= not w24653 and not w25158;
w25160 <= b(38) and not w24642;
w25161 <= not w24640 and w25160;
w25162 <= not w24644 and not w25161;
w25163 <= not w25159 and w25162;
w25164 <= not w24644 and not w25163;
w25165 <= b(39) and not w24633;
w25166 <= not w24631 and w25165;
w25167 <= not w24635 and not w25166;
w25168 <= not w25164 and w25167;
w25169 <= not w24635 and not w25168;
w25170 <= b(40) and not w24624;
w25171 <= not w24622 and w25170;
w25172 <= not w24626 and not w25171;
w25173 <= not w25169 and w25172;
w25174 <= not w24626 and not w25173;
w25175 <= b(41) and not w24615;
w25176 <= not w24613 and w25175;
w25177 <= not w24617 and not w25176;
w25178 <= not w25174 and w25177;
w25179 <= not w24617 and not w25178;
w25180 <= b(42) and not w24606;
w25181 <= not w24604 and w25180;
w25182 <= not w24608 and not w25181;
w25183 <= not w25179 and w25182;
w25184 <= not w24608 and not w25183;
w25185 <= b(43) and not w24597;
w25186 <= not w24595 and w25185;
w25187 <= not w24599 and not w25186;
w25188 <= not w25184 and w25187;
w25189 <= not w24599 and not w25188;
w25190 <= b(44) and not w24588;
w25191 <= not w24586 and w25190;
w25192 <= not w24590 and not w25191;
w25193 <= not w25189 and w25192;
w25194 <= not w24590 and not w25193;
w25195 <= b(45) and not w24579;
w25196 <= not w24577 and w25195;
w25197 <= not w24581 and not w25196;
w25198 <= not w25194 and w25197;
w25199 <= not w24581 and not w25198;
w25200 <= b(46) and not w24570;
w25201 <= not w24568 and w25200;
w25202 <= not w24572 and not w25201;
w25203 <= not w25199 and w25202;
w25204 <= not w24572 and not w25203;
w25205 <= b(47) and not w24561;
w25206 <= not w24559 and w25205;
w25207 <= not w24563 and not w25206;
w25208 <= not w25204 and w25207;
w25209 <= not w24563 and not w25208;
w25210 <= b(48) and not w24552;
w25211 <= not w24550 and w25210;
w25212 <= not w24554 and not w25211;
w25213 <= not w25209 and w25212;
w25214 <= not w24554 and not w25213;
w25215 <= b(49) and not w24543;
w25216 <= not w24541 and w25215;
w25217 <= not w24545 and not w25216;
w25218 <= not w25214 and w25217;
w25219 <= not w24545 and not w25218;
w25220 <= b(50) and not w24534;
w25221 <= not w24532 and w25220;
w25222 <= not w24536 and not w25221;
w25223 <= not w25219 and w25222;
w25224 <= not w24536 and not w25223;
w25225 <= b(51) and not w24525;
w25226 <= not w24523 and w25225;
w25227 <= not w24527 and not w25226;
w25228 <= not w25224 and w25227;
w25229 <= not w24527 and not w25228;
w25230 <= b(52) and not w24516;
w25231 <= not w24514 and w25230;
w25232 <= not w24518 and not w25231;
w25233 <= not w25229 and w25232;
w25234 <= not w24518 and not w25233;
w25235 <= b(53) and not w24507;
w25236 <= not w24505 and w25235;
w25237 <= not w24509 and not w25236;
w25238 <= not w25234 and w25237;
w25239 <= not w24509 and not w25238;
w25240 <= b(54) and not w24498;
w25241 <= not w24496 and w25240;
w25242 <= not w24500 and not w25241;
w25243 <= not w25239 and w25242;
w25244 <= not w24500 and not w25243;
w25245 <= b(55) and not w24489;
w25246 <= not w24487 and w25245;
w25247 <= not w24491 and not w25246;
w25248 <= not w25244 and w25247;
w25249 <= not w24491 and not w25248;
w25250 <= b(56) and not w24480;
w25251 <= not w24478 and w25250;
w25252 <= not w24482 and not w25251;
w25253 <= not w25249 and w25252;
w25254 <= not w24482 and not w25253;
w25255 <= b(57) and not w24471;
w25256 <= not w24469 and w25255;
w25257 <= not w24473 and not w25256;
w25258 <= not w25254 and w25257;
w25259 <= not w24473 and not w25258;
w25260 <= b(58) and not w24462;
w25261 <= not w24460 and w25260;
w25262 <= not w24464 and not w25261;
w25263 <= not w25259 and w25262;
w25264 <= not w24464 and not w25263;
w25265 <= not w23648 and not w24449;
w25266 <= not w24447 and w25265;
w25267 <= not w24438 and w25266;
w25268 <= not w24447 and not w24449;
w25269 <= not w24439 and not w25268;
w25270 <= not w25267 and not w25269;
w25271 <= not w24455 and not w25270;
w25272 <= not w24446 and not w24454;
w25273 <= not w24453 and w25272;
w25274 <= not w25271 and not w25273;
w25275 <= not b(59) and not w25274;
w25276 <= b(59) and not w25273;
w25277 <= not w25271 and w25276;
w25278 <= w23 and not w25277;
w25279 <= not w25275 and w25278;
w25280 <= not w25264 and w25279;
w25281 <= w24450 and not w25274;
w25282 <= not w25280 and not w25281;
w25283 <= not w24473 and w25262;
w25284 <= not w25258 and w25283;
w25285 <= not w25259 and not w25262;
w25286 <= not w25284 and not w25285;
w25287 <= not w25282 and not w25286;
w25288 <= not w24463 and not w25281;
w25289 <= not w25280 and w25288;
w25290 <= not w25287 and not w25289;
w25291 <= not b(59) and not w25290;
w25292 <= not w24482 and w25257;
w25293 <= not w25253 and w25292;
w25294 <= not w25254 and not w25257;
w25295 <= not w25293 and not w25294;
w25296 <= not w25282 and not w25295;
w25297 <= not w24472 and not w25281;
w25298 <= not w25280 and w25297;
w25299 <= not w25296 and not w25298;
w25300 <= not b(58) and not w25299;
w25301 <= not w24491 and w25252;
w25302 <= not w25248 and w25301;
w25303 <= not w25249 and not w25252;
w25304 <= not w25302 and not w25303;
w25305 <= not w25282 and not w25304;
w25306 <= not w24481 and not w25281;
w25307 <= not w25280 and w25306;
w25308 <= not w25305 and not w25307;
w25309 <= not b(57) and not w25308;
w25310 <= not w24500 and w25247;
w25311 <= not w25243 and w25310;
w25312 <= not w25244 and not w25247;
w25313 <= not w25311 and not w25312;
w25314 <= not w25282 and not w25313;
w25315 <= not w24490 and not w25281;
w25316 <= not w25280 and w25315;
w25317 <= not w25314 and not w25316;
w25318 <= not b(56) and not w25317;
w25319 <= not w24509 and w25242;
w25320 <= not w25238 and w25319;
w25321 <= not w25239 and not w25242;
w25322 <= not w25320 and not w25321;
w25323 <= not w25282 and not w25322;
w25324 <= not w24499 and not w25281;
w25325 <= not w25280 and w25324;
w25326 <= not w25323 and not w25325;
w25327 <= not b(55) and not w25326;
w25328 <= not w24518 and w25237;
w25329 <= not w25233 and w25328;
w25330 <= not w25234 and not w25237;
w25331 <= not w25329 and not w25330;
w25332 <= not w25282 and not w25331;
w25333 <= not w24508 and not w25281;
w25334 <= not w25280 and w25333;
w25335 <= not w25332 and not w25334;
w25336 <= not b(54) and not w25335;
w25337 <= not w24527 and w25232;
w25338 <= not w25228 and w25337;
w25339 <= not w25229 and not w25232;
w25340 <= not w25338 and not w25339;
w25341 <= not w25282 and not w25340;
w25342 <= not w24517 and not w25281;
w25343 <= not w25280 and w25342;
w25344 <= not w25341 and not w25343;
w25345 <= not b(53) and not w25344;
w25346 <= not w24536 and w25227;
w25347 <= not w25223 and w25346;
w25348 <= not w25224 and not w25227;
w25349 <= not w25347 and not w25348;
w25350 <= not w25282 and not w25349;
w25351 <= not w24526 and not w25281;
w25352 <= not w25280 and w25351;
w25353 <= not w25350 and not w25352;
w25354 <= not b(52) and not w25353;
w25355 <= not w24545 and w25222;
w25356 <= not w25218 and w25355;
w25357 <= not w25219 and not w25222;
w25358 <= not w25356 and not w25357;
w25359 <= not w25282 and not w25358;
w25360 <= not w24535 and not w25281;
w25361 <= not w25280 and w25360;
w25362 <= not w25359 and not w25361;
w25363 <= not b(51) and not w25362;
w25364 <= not w24554 and w25217;
w25365 <= not w25213 and w25364;
w25366 <= not w25214 and not w25217;
w25367 <= not w25365 and not w25366;
w25368 <= not w25282 and not w25367;
w25369 <= not w24544 and not w25281;
w25370 <= not w25280 and w25369;
w25371 <= not w25368 and not w25370;
w25372 <= not b(50) and not w25371;
w25373 <= not w24563 and w25212;
w25374 <= not w25208 and w25373;
w25375 <= not w25209 and not w25212;
w25376 <= not w25374 and not w25375;
w25377 <= not w25282 and not w25376;
w25378 <= not w24553 and not w25281;
w25379 <= not w25280 and w25378;
w25380 <= not w25377 and not w25379;
w25381 <= not b(49) and not w25380;
w25382 <= not w24572 and w25207;
w25383 <= not w25203 and w25382;
w25384 <= not w25204 and not w25207;
w25385 <= not w25383 and not w25384;
w25386 <= not w25282 and not w25385;
w25387 <= not w24562 and not w25281;
w25388 <= not w25280 and w25387;
w25389 <= not w25386 and not w25388;
w25390 <= not b(48) and not w25389;
w25391 <= not w24581 and w25202;
w25392 <= not w25198 and w25391;
w25393 <= not w25199 and not w25202;
w25394 <= not w25392 and not w25393;
w25395 <= not w25282 and not w25394;
w25396 <= not w24571 and not w25281;
w25397 <= not w25280 and w25396;
w25398 <= not w25395 and not w25397;
w25399 <= not b(47) and not w25398;
w25400 <= not w24590 and w25197;
w25401 <= not w25193 and w25400;
w25402 <= not w25194 and not w25197;
w25403 <= not w25401 and not w25402;
w25404 <= not w25282 and not w25403;
w25405 <= not w24580 and not w25281;
w25406 <= not w25280 and w25405;
w25407 <= not w25404 and not w25406;
w25408 <= not b(46) and not w25407;
w25409 <= not w24599 and w25192;
w25410 <= not w25188 and w25409;
w25411 <= not w25189 and not w25192;
w25412 <= not w25410 and not w25411;
w25413 <= not w25282 and not w25412;
w25414 <= not w24589 and not w25281;
w25415 <= not w25280 and w25414;
w25416 <= not w25413 and not w25415;
w25417 <= not b(45) and not w25416;
w25418 <= not w24608 and w25187;
w25419 <= not w25183 and w25418;
w25420 <= not w25184 and not w25187;
w25421 <= not w25419 and not w25420;
w25422 <= not w25282 and not w25421;
w25423 <= not w24598 and not w25281;
w25424 <= not w25280 and w25423;
w25425 <= not w25422 and not w25424;
w25426 <= not b(44) and not w25425;
w25427 <= not w24617 and w25182;
w25428 <= not w25178 and w25427;
w25429 <= not w25179 and not w25182;
w25430 <= not w25428 and not w25429;
w25431 <= not w25282 and not w25430;
w25432 <= not w24607 and not w25281;
w25433 <= not w25280 and w25432;
w25434 <= not w25431 and not w25433;
w25435 <= not b(43) and not w25434;
w25436 <= not w24626 and w25177;
w25437 <= not w25173 and w25436;
w25438 <= not w25174 and not w25177;
w25439 <= not w25437 and not w25438;
w25440 <= not w25282 and not w25439;
w25441 <= not w24616 and not w25281;
w25442 <= not w25280 and w25441;
w25443 <= not w25440 and not w25442;
w25444 <= not b(42) and not w25443;
w25445 <= not w24635 and w25172;
w25446 <= not w25168 and w25445;
w25447 <= not w25169 and not w25172;
w25448 <= not w25446 and not w25447;
w25449 <= not w25282 and not w25448;
w25450 <= not w24625 and not w25281;
w25451 <= not w25280 and w25450;
w25452 <= not w25449 and not w25451;
w25453 <= not b(41) and not w25452;
w25454 <= not w24644 and w25167;
w25455 <= not w25163 and w25454;
w25456 <= not w25164 and not w25167;
w25457 <= not w25455 and not w25456;
w25458 <= not w25282 and not w25457;
w25459 <= not w24634 and not w25281;
w25460 <= not w25280 and w25459;
w25461 <= not w25458 and not w25460;
w25462 <= not b(40) and not w25461;
w25463 <= not w24653 and w25162;
w25464 <= not w25158 and w25463;
w25465 <= not w25159 and not w25162;
w25466 <= not w25464 and not w25465;
w25467 <= not w25282 and not w25466;
w25468 <= not w24643 and not w25281;
w25469 <= not w25280 and w25468;
w25470 <= not w25467 and not w25469;
w25471 <= not b(39) and not w25470;
w25472 <= not w24662 and w25157;
w25473 <= not w25153 and w25472;
w25474 <= not w25154 and not w25157;
w25475 <= not w25473 and not w25474;
w25476 <= not w25282 and not w25475;
w25477 <= not w24652 and not w25281;
w25478 <= not w25280 and w25477;
w25479 <= not w25476 and not w25478;
w25480 <= not b(38) and not w25479;
w25481 <= not w24671 and w25152;
w25482 <= not w25148 and w25481;
w25483 <= not w25149 and not w25152;
w25484 <= not w25482 and not w25483;
w25485 <= not w25282 and not w25484;
w25486 <= not w24661 and not w25281;
w25487 <= not w25280 and w25486;
w25488 <= not w25485 and not w25487;
w25489 <= not b(37) and not w25488;
w25490 <= not w24680 and w25147;
w25491 <= not w25143 and w25490;
w25492 <= not w25144 and not w25147;
w25493 <= not w25491 and not w25492;
w25494 <= not w25282 and not w25493;
w25495 <= not w24670 and not w25281;
w25496 <= not w25280 and w25495;
w25497 <= not w25494 and not w25496;
w25498 <= not b(36) and not w25497;
w25499 <= not w24689 and w25142;
w25500 <= not w25138 and w25499;
w25501 <= not w25139 and not w25142;
w25502 <= not w25500 and not w25501;
w25503 <= not w25282 and not w25502;
w25504 <= not w24679 and not w25281;
w25505 <= not w25280 and w25504;
w25506 <= not w25503 and not w25505;
w25507 <= not b(35) and not w25506;
w25508 <= not w24698 and w25137;
w25509 <= not w25133 and w25508;
w25510 <= not w25134 and not w25137;
w25511 <= not w25509 and not w25510;
w25512 <= not w25282 and not w25511;
w25513 <= not w24688 and not w25281;
w25514 <= not w25280 and w25513;
w25515 <= not w25512 and not w25514;
w25516 <= not b(34) and not w25515;
w25517 <= not w24707 and w25132;
w25518 <= not w25128 and w25517;
w25519 <= not w25129 and not w25132;
w25520 <= not w25518 and not w25519;
w25521 <= not w25282 and not w25520;
w25522 <= not w24697 and not w25281;
w25523 <= not w25280 and w25522;
w25524 <= not w25521 and not w25523;
w25525 <= not b(33) and not w25524;
w25526 <= not w24716 and w25127;
w25527 <= not w25123 and w25526;
w25528 <= not w25124 and not w25127;
w25529 <= not w25527 and not w25528;
w25530 <= not w25282 and not w25529;
w25531 <= not w24706 and not w25281;
w25532 <= not w25280 and w25531;
w25533 <= not w25530 and not w25532;
w25534 <= not b(32) and not w25533;
w25535 <= not w24725 and w25122;
w25536 <= not w25118 and w25535;
w25537 <= not w25119 and not w25122;
w25538 <= not w25536 and not w25537;
w25539 <= not w25282 and not w25538;
w25540 <= not w24715 and not w25281;
w25541 <= not w25280 and w25540;
w25542 <= not w25539 and not w25541;
w25543 <= not b(31) and not w25542;
w25544 <= not w24734 and w25117;
w25545 <= not w25113 and w25544;
w25546 <= not w25114 and not w25117;
w25547 <= not w25545 and not w25546;
w25548 <= not w25282 and not w25547;
w25549 <= not w24724 and not w25281;
w25550 <= not w25280 and w25549;
w25551 <= not w25548 and not w25550;
w25552 <= not b(30) and not w25551;
w25553 <= not w24743 and w25112;
w25554 <= not w25108 and w25553;
w25555 <= not w25109 and not w25112;
w25556 <= not w25554 and not w25555;
w25557 <= not w25282 and not w25556;
w25558 <= not w24733 and not w25281;
w25559 <= not w25280 and w25558;
w25560 <= not w25557 and not w25559;
w25561 <= not b(29) and not w25560;
w25562 <= not w24752 and w25107;
w25563 <= not w25103 and w25562;
w25564 <= not w25104 and not w25107;
w25565 <= not w25563 and not w25564;
w25566 <= not w25282 and not w25565;
w25567 <= not w24742 and not w25281;
w25568 <= not w25280 and w25567;
w25569 <= not w25566 and not w25568;
w25570 <= not b(28) and not w25569;
w25571 <= not w24761 and w25102;
w25572 <= not w25098 and w25571;
w25573 <= not w25099 and not w25102;
w25574 <= not w25572 and not w25573;
w25575 <= not w25282 and not w25574;
w25576 <= not w24751 and not w25281;
w25577 <= not w25280 and w25576;
w25578 <= not w25575 and not w25577;
w25579 <= not b(27) and not w25578;
w25580 <= not w24770 and w25097;
w25581 <= not w25093 and w25580;
w25582 <= not w25094 and not w25097;
w25583 <= not w25581 and not w25582;
w25584 <= not w25282 and not w25583;
w25585 <= not w24760 and not w25281;
w25586 <= not w25280 and w25585;
w25587 <= not w25584 and not w25586;
w25588 <= not b(26) and not w25587;
w25589 <= not w24779 and w25092;
w25590 <= not w25088 and w25589;
w25591 <= not w25089 and not w25092;
w25592 <= not w25590 and not w25591;
w25593 <= not w25282 and not w25592;
w25594 <= not w24769 and not w25281;
w25595 <= not w25280 and w25594;
w25596 <= not w25593 and not w25595;
w25597 <= not b(25) and not w25596;
w25598 <= not w24788 and w25087;
w25599 <= not w25083 and w25598;
w25600 <= not w25084 and not w25087;
w25601 <= not w25599 and not w25600;
w25602 <= not w25282 and not w25601;
w25603 <= not w24778 and not w25281;
w25604 <= not w25280 and w25603;
w25605 <= not w25602 and not w25604;
w25606 <= not b(24) and not w25605;
w25607 <= not w24797 and w25082;
w25608 <= not w25078 and w25607;
w25609 <= not w25079 and not w25082;
w25610 <= not w25608 and not w25609;
w25611 <= not w25282 and not w25610;
w25612 <= not w24787 and not w25281;
w25613 <= not w25280 and w25612;
w25614 <= not w25611 and not w25613;
w25615 <= not b(23) and not w25614;
w25616 <= not w24806 and w25077;
w25617 <= not w25073 and w25616;
w25618 <= not w25074 and not w25077;
w25619 <= not w25617 and not w25618;
w25620 <= not w25282 and not w25619;
w25621 <= not w24796 and not w25281;
w25622 <= not w25280 and w25621;
w25623 <= not w25620 and not w25622;
w25624 <= not b(22) and not w25623;
w25625 <= not w24815 and w25072;
w25626 <= not w25068 and w25625;
w25627 <= not w25069 and not w25072;
w25628 <= not w25626 and not w25627;
w25629 <= not w25282 and not w25628;
w25630 <= not w24805 and not w25281;
w25631 <= not w25280 and w25630;
w25632 <= not w25629 and not w25631;
w25633 <= not b(21) and not w25632;
w25634 <= not w24824 and w25067;
w25635 <= not w25063 and w25634;
w25636 <= not w25064 and not w25067;
w25637 <= not w25635 and not w25636;
w25638 <= not w25282 and not w25637;
w25639 <= not w24814 and not w25281;
w25640 <= not w25280 and w25639;
w25641 <= not w25638 and not w25640;
w25642 <= not b(20) and not w25641;
w25643 <= not w24833 and w25062;
w25644 <= not w25058 and w25643;
w25645 <= not w25059 and not w25062;
w25646 <= not w25644 and not w25645;
w25647 <= not w25282 and not w25646;
w25648 <= not w24823 and not w25281;
w25649 <= not w25280 and w25648;
w25650 <= not w25647 and not w25649;
w25651 <= not b(19) and not w25650;
w25652 <= not w24842 and w25057;
w25653 <= not w25053 and w25652;
w25654 <= not w25054 and not w25057;
w25655 <= not w25653 and not w25654;
w25656 <= not w25282 and not w25655;
w25657 <= not w24832 and not w25281;
w25658 <= not w25280 and w25657;
w25659 <= not w25656 and not w25658;
w25660 <= not b(18) and not w25659;
w25661 <= not w24851 and w25052;
w25662 <= not w25048 and w25661;
w25663 <= not w25049 and not w25052;
w25664 <= not w25662 and not w25663;
w25665 <= not w25282 and not w25664;
w25666 <= not w24841 and not w25281;
w25667 <= not w25280 and w25666;
w25668 <= not w25665 and not w25667;
w25669 <= not b(17) and not w25668;
w25670 <= not w24860 and w25047;
w25671 <= not w25043 and w25670;
w25672 <= not w25044 and not w25047;
w25673 <= not w25671 and not w25672;
w25674 <= not w25282 and not w25673;
w25675 <= not w24850 and not w25281;
w25676 <= not w25280 and w25675;
w25677 <= not w25674 and not w25676;
w25678 <= not b(16) and not w25677;
w25679 <= not w24869 and w25042;
w25680 <= not w25038 and w25679;
w25681 <= not w25039 and not w25042;
w25682 <= not w25680 and not w25681;
w25683 <= not w25282 and not w25682;
w25684 <= not w24859 and not w25281;
w25685 <= not w25280 and w25684;
w25686 <= not w25683 and not w25685;
w25687 <= not b(15) and not w25686;
w25688 <= not w24878 and w25037;
w25689 <= not w25033 and w25688;
w25690 <= not w25034 and not w25037;
w25691 <= not w25689 and not w25690;
w25692 <= not w25282 and not w25691;
w25693 <= not w24868 and not w25281;
w25694 <= not w25280 and w25693;
w25695 <= not w25692 and not w25694;
w25696 <= not b(14) and not w25695;
w25697 <= not w24887 and w25032;
w25698 <= not w25028 and w25697;
w25699 <= not w25029 and not w25032;
w25700 <= not w25698 and not w25699;
w25701 <= not w25282 and not w25700;
w25702 <= not w24877 and not w25281;
w25703 <= not w25280 and w25702;
w25704 <= not w25701 and not w25703;
w25705 <= not b(13) and not w25704;
w25706 <= not w24896 and w25027;
w25707 <= not w25023 and w25706;
w25708 <= not w25024 and not w25027;
w25709 <= not w25707 and not w25708;
w25710 <= not w25282 and not w25709;
w25711 <= not w24886 and not w25281;
w25712 <= not w25280 and w25711;
w25713 <= not w25710 and not w25712;
w25714 <= not b(12) and not w25713;
w25715 <= not w24905 and w25022;
w25716 <= not w25018 and w25715;
w25717 <= not w25019 and not w25022;
w25718 <= not w25716 and not w25717;
w25719 <= not w25282 and not w25718;
w25720 <= not w24895 and not w25281;
w25721 <= not w25280 and w25720;
w25722 <= not w25719 and not w25721;
w25723 <= not b(11) and not w25722;
w25724 <= not w24914 and w25017;
w25725 <= not w25013 and w25724;
w25726 <= not w25014 and not w25017;
w25727 <= not w25725 and not w25726;
w25728 <= not w25282 and not w25727;
w25729 <= not w24904 and not w25281;
w25730 <= not w25280 and w25729;
w25731 <= not w25728 and not w25730;
w25732 <= not b(10) and not w25731;
w25733 <= not w24923 and w25012;
w25734 <= not w25008 and w25733;
w25735 <= not w25009 and not w25012;
w25736 <= not w25734 and not w25735;
w25737 <= not w25282 and not w25736;
w25738 <= not w24913 and not w25281;
w25739 <= not w25280 and w25738;
w25740 <= not w25737 and not w25739;
w25741 <= not b(9) and not w25740;
w25742 <= not w24932 and w25007;
w25743 <= not w25003 and w25742;
w25744 <= not w25004 and not w25007;
w25745 <= not w25743 and not w25744;
w25746 <= not w25282 and not w25745;
w25747 <= not w24922 and not w25281;
w25748 <= not w25280 and w25747;
w25749 <= not w25746 and not w25748;
w25750 <= not b(8) and not w25749;
w25751 <= not w24941 and w25002;
w25752 <= not w24998 and w25751;
w25753 <= not w24999 and not w25002;
w25754 <= not w25752 and not w25753;
w25755 <= not w25282 and not w25754;
w25756 <= not w24931 and not w25281;
w25757 <= not w25280 and w25756;
w25758 <= not w25755 and not w25757;
w25759 <= not b(7) and not w25758;
w25760 <= not w24950 and w24997;
w25761 <= not w24993 and w25760;
w25762 <= not w24994 and not w24997;
w25763 <= not w25761 and not w25762;
w25764 <= not w25282 and not w25763;
w25765 <= not w24940 and not w25281;
w25766 <= not w25280 and w25765;
w25767 <= not w25764 and not w25766;
w25768 <= not b(6) and not w25767;
w25769 <= not w24959 and w24992;
w25770 <= not w24988 and w25769;
w25771 <= not w24989 and not w24992;
w25772 <= not w25770 and not w25771;
w25773 <= not w25282 and not w25772;
w25774 <= not w24949 and not w25281;
w25775 <= not w25280 and w25774;
w25776 <= not w25773 and not w25775;
w25777 <= not b(5) and not w25776;
w25778 <= not w24967 and w24987;
w25779 <= not w24983 and w25778;
w25780 <= not w24984 and not w24987;
w25781 <= not w25779 and not w25780;
w25782 <= not w25282 and not w25781;
w25783 <= not w24958 and not w25281;
w25784 <= not w25280 and w25783;
w25785 <= not w25782 and not w25784;
w25786 <= not b(4) and not w25785;
w25787 <= not w24978 and w24982;
w25788 <= not w24977 and w25787;
w25789 <= not w24979 and not w24982;
w25790 <= not w25788 and not w25789;
w25791 <= not w25282 and not w25790;
w25792 <= not w24966 and not w25281;
w25793 <= not w25280 and w25792;
w25794 <= not w25791 and not w25793;
w25795 <= not b(3) and not w25794;
w25796 <= not w24974 and w24976;
w25797 <= not w24972 and w25796;
w25798 <= not w24977 and not w25797;
w25799 <= not w25282 and w25798;
w25800 <= not w24971 and not w25281;
w25801 <= not w25280 and w25800;
w25802 <= not w25799 and not w25801;
w25803 <= not b(2) and not w25802;
w25804 <= b(0) and not w25282;
w25805 <= a(4) and not w25804;
w25806 <= w24976 and not w25282;
w25807 <= not w25805 and not w25806;
w25808 <= b(1) and not w25807;
w25809 <= not b(1) and not w25806;
w25810 <= not w25805 and w25809;
w25811 <= not w25808 and not w25810;
w25812 <= not a(3) and b(0);
w25813 <= not w25811 and not w25812;
w25814 <= not b(1) and not w25807;
w25815 <= not w25813 and not w25814;
w25816 <= b(2) and not w25801;
w25817 <= not w25799 and w25816;
w25818 <= not w25803 and not w25817;
w25819 <= not w25815 and w25818;
w25820 <= not w25803 and not w25819;
w25821 <= b(3) and not w25793;
w25822 <= not w25791 and w25821;
w25823 <= not w25795 and not w25822;
w25824 <= not w25820 and w25823;
w25825 <= not w25795 and not w25824;
w25826 <= b(4) and not w25784;
w25827 <= not w25782 and w25826;
w25828 <= not w25786 and not w25827;
w25829 <= not w25825 and w25828;
w25830 <= not w25786 and not w25829;
w25831 <= b(5) and not w25775;
w25832 <= not w25773 and w25831;
w25833 <= not w25777 and not w25832;
w25834 <= not w25830 and w25833;
w25835 <= not w25777 and not w25834;
w25836 <= b(6) and not w25766;
w25837 <= not w25764 and w25836;
w25838 <= not w25768 and not w25837;
w25839 <= not w25835 and w25838;
w25840 <= not w25768 and not w25839;
w25841 <= b(7) and not w25757;
w25842 <= not w25755 and w25841;
w25843 <= not w25759 and not w25842;
w25844 <= not w25840 and w25843;
w25845 <= not w25759 and not w25844;
w25846 <= b(8) and not w25748;
w25847 <= not w25746 and w25846;
w25848 <= not w25750 and not w25847;
w25849 <= not w25845 and w25848;
w25850 <= not w25750 and not w25849;
w25851 <= b(9) and not w25739;
w25852 <= not w25737 and w25851;
w25853 <= not w25741 and not w25852;
w25854 <= not w25850 and w25853;
w25855 <= not w25741 and not w25854;
w25856 <= b(10) and not w25730;
w25857 <= not w25728 and w25856;
w25858 <= not w25732 and not w25857;
w25859 <= not w25855 and w25858;
w25860 <= not w25732 and not w25859;
w25861 <= b(11) and not w25721;
w25862 <= not w25719 and w25861;
w25863 <= not w25723 and not w25862;
w25864 <= not w25860 and w25863;
w25865 <= not w25723 and not w25864;
w25866 <= b(12) and not w25712;
w25867 <= not w25710 and w25866;
w25868 <= not w25714 and not w25867;
w25869 <= not w25865 and w25868;
w25870 <= not w25714 and not w25869;
w25871 <= b(13) and not w25703;
w25872 <= not w25701 and w25871;
w25873 <= not w25705 and not w25872;
w25874 <= not w25870 and w25873;
w25875 <= not w25705 and not w25874;
w25876 <= b(14) and not w25694;
w25877 <= not w25692 and w25876;
w25878 <= not w25696 and not w25877;
w25879 <= not w25875 and w25878;
w25880 <= not w25696 and not w25879;
w25881 <= b(15) and not w25685;
w25882 <= not w25683 and w25881;
w25883 <= not w25687 and not w25882;
w25884 <= not w25880 and w25883;
w25885 <= not w25687 and not w25884;
w25886 <= b(16) and not w25676;
w25887 <= not w25674 and w25886;
w25888 <= not w25678 and not w25887;
w25889 <= not w25885 and w25888;
w25890 <= not w25678 and not w25889;
w25891 <= b(17) and not w25667;
w25892 <= not w25665 and w25891;
w25893 <= not w25669 and not w25892;
w25894 <= not w25890 and w25893;
w25895 <= not w25669 and not w25894;
w25896 <= b(18) and not w25658;
w25897 <= not w25656 and w25896;
w25898 <= not w25660 and not w25897;
w25899 <= not w25895 and w25898;
w25900 <= not w25660 and not w25899;
w25901 <= b(19) and not w25649;
w25902 <= not w25647 and w25901;
w25903 <= not w25651 and not w25902;
w25904 <= not w25900 and w25903;
w25905 <= not w25651 and not w25904;
w25906 <= b(20) and not w25640;
w25907 <= not w25638 and w25906;
w25908 <= not w25642 and not w25907;
w25909 <= not w25905 and w25908;
w25910 <= not w25642 and not w25909;
w25911 <= b(21) and not w25631;
w25912 <= not w25629 and w25911;
w25913 <= not w25633 and not w25912;
w25914 <= not w25910 and w25913;
w25915 <= not w25633 and not w25914;
w25916 <= b(22) and not w25622;
w25917 <= not w25620 and w25916;
w25918 <= not w25624 and not w25917;
w25919 <= not w25915 and w25918;
w25920 <= not w25624 and not w25919;
w25921 <= b(23) and not w25613;
w25922 <= not w25611 and w25921;
w25923 <= not w25615 and not w25922;
w25924 <= not w25920 and w25923;
w25925 <= not w25615 and not w25924;
w25926 <= b(24) and not w25604;
w25927 <= not w25602 and w25926;
w25928 <= not w25606 and not w25927;
w25929 <= not w25925 and w25928;
w25930 <= not w25606 and not w25929;
w25931 <= b(25) and not w25595;
w25932 <= not w25593 and w25931;
w25933 <= not w25597 and not w25932;
w25934 <= not w25930 and w25933;
w25935 <= not w25597 and not w25934;
w25936 <= b(26) and not w25586;
w25937 <= not w25584 and w25936;
w25938 <= not w25588 and not w25937;
w25939 <= not w25935 and w25938;
w25940 <= not w25588 and not w25939;
w25941 <= b(27) and not w25577;
w25942 <= not w25575 and w25941;
w25943 <= not w25579 and not w25942;
w25944 <= not w25940 and w25943;
w25945 <= not w25579 and not w25944;
w25946 <= b(28) and not w25568;
w25947 <= not w25566 and w25946;
w25948 <= not w25570 and not w25947;
w25949 <= not w25945 and w25948;
w25950 <= not w25570 and not w25949;
w25951 <= b(29) and not w25559;
w25952 <= not w25557 and w25951;
w25953 <= not w25561 and not w25952;
w25954 <= not w25950 and w25953;
w25955 <= not w25561 and not w25954;
w25956 <= b(30) and not w25550;
w25957 <= not w25548 and w25956;
w25958 <= not w25552 and not w25957;
w25959 <= not w25955 and w25958;
w25960 <= not w25552 and not w25959;
w25961 <= b(31) and not w25541;
w25962 <= not w25539 and w25961;
w25963 <= not w25543 and not w25962;
w25964 <= not w25960 and w25963;
w25965 <= not w25543 and not w25964;
w25966 <= b(32) and not w25532;
w25967 <= not w25530 and w25966;
w25968 <= not w25534 and not w25967;
w25969 <= not w25965 and w25968;
w25970 <= not w25534 and not w25969;
w25971 <= b(33) and not w25523;
w25972 <= not w25521 and w25971;
w25973 <= not w25525 and not w25972;
w25974 <= not w25970 and w25973;
w25975 <= not w25525 and not w25974;
w25976 <= b(34) and not w25514;
w25977 <= not w25512 and w25976;
w25978 <= not w25516 and not w25977;
w25979 <= not w25975 and w25978;
w25980 <= not w25516 and not w25979;
w25981 <= b(35) and not w25505;
w25982 <= not w25503 and w25981;
w25983 <= not w25507 and not w25982;
w25984 <= not w25980 and w25983;
w25985 <= not w25507 and not w25984;
w25986 <= b(36) and not w25496;
w25987 <= not w25494 and w25986;
w25988 <= not w25498 and not w25987;
w25989 <= not w25985 and w25988;
w25990 <= not w25498 and not w25989;
w25991 <= b(37) and not w25487;
w25992 <= not w25485 and w25991;
w25993 <= not w25489 and not w25992;
w25994 <= not w25990 and w25993;
w25995 <= not w25489 and not w25994;
w25996 <= b(38) and not w25478;
w25997 <= not w25476 and w25996;
w25998 <= not w25480 and not w25997;
w25999 <= not w25995 and w25998;
w26000 <= not w25480 and not w25999;
w26001 <= b(39) and not w25469;
w26002 <= not w25467 and w26001;
w26003 <= not w25471 and not w26002;
w26004 <= not w26000 and w26003;
w26005 <= not w25471 and not w26004;
w26006 <= b(40) and not w25460;
w26007 <= not w25458 and w26006;
w26008 <= not w25462 and not w26007;
w26009 <= not w26005 and w26008;
w26010 <= not w25462 and not w26009;
w26011 <= b(41) and not w25451;
w26012 <= not w25449 and w26011;
w26013 <= not w25453 and not w26012;
w26014 <= not w26010 and w26013;
w26015 <= not w25453 and not w26014;
w26016 <= b(42) and not w25442;
w26017 <= not w25440 and w26016;
w26018 <= not w25444 and not w26017;
w26019 <= not w26015 and w26018;
w26020 <= not w25444 and not w26019;
w26021 <= b(43) and not w25433;
w26022 <= not w25431 and w26021;
w26023 <= not w25435 and not w26022;
w26024 <= not w26020 and w26023;
w26025 <= not w25435 and not w26024;
w26026 <= b(44) and not w25424;
w26027 <= not w25422 and w26026;
w26028 <= not w25426 and not w26027;
w26029 <= not w26025 and w26028;
w26030 <= not w25426 and not w26029;
w26031 <= b(45) and not w25415;
w26032 <= not w25413 and w26031;
w26033 <= not w25417 and not w26032;
w26034 <= not w26030 and w26033;
w26035 <= not w25417 and not w26034;
w26036 <= b(46) and not w25406;
w26037 <= not w25404 and w26036;
w26038 <= not w25408 and not w26037;
w26039 <= not w26035 and w26038;
w26040 <= not w25408 and not w26039;
w26041 <= b(47) and not w25397;
w26042 <= not w25395 and w26041;
w26043 <= not w25399 and not w26042;
w26044 <= not w26040 and w26043;
w26045 <= not w25399 and not w26044;
w26046 <= b(48) and not w25388;
w26047 <= not w25386 and w26046;
w26048 <= not w25390 and not w26047;
w26049 <= not w26045 and w26048;
w26050 <= not w25390 and not w26049;
w26051 <= b(49) and not w25379;
w26052 <= not w25377 and w26051;
w26053 <= not w25381 and not w26052;
w26054 <= not w26050 and w26053;
w26055 <= not w25381 and not w26054;
w26056 <= b(50) and not w25370;
w26057 <= not w25368 and w26056;
w26058 <= not w25372 and not w26057;
w26059 <= not w26055 and w26058;
w26060 <= not w25372 and not w26059;
w26061 <= b(51) and not w25361;
w26062 <= not w25359 and w26061;
w26063 <= not w25363 and not w26062;
w26064 <= not w26060 and w26063;
w26065 <= not w25363 and not w26064;
w26066 <= b(52) and not w25352;
w26067 <= not w25350 and w26066;
w26068 <= not w25354 and not w26067;
w26069 <= not w26065 and w26068;
w26070 <= not w25354 and not w26069;
w26071 <= b(53) and not w25343;
w26072 <= not w25341 and w26071;
w26073 <= not w25345 and not w26072;
w26074 <= not w26070 and w26073;
w26075 <= not w25345 and not w26074;
w26076 <= b(54) and not w25334;
w26077 <= not w25332 and w26076;
w26078 <= not w25336 and not w26077;
w26079 <= not w26075 and w26078;
w26080 <= not w25336 and not w26079;
w26081 <= b(55) and not w25325;
w26082 <= not w25323 and w26081;
w26083 <= not w25327 and not w26082;
w26084 <= not w26080 and w26083;
w26085 <= not w25327 and not w26084;
w26086 <= b(56) and not w25316;
w26087 <= not w25314 and w26086;
w26088 <= not w25318 and not w26087;
w26089 <= not w26085 and w26088;
w26090 <= not w25318 and not w26089;
w26091 <= b(57) and not w25307;
w26092 <= not w25305 and w26091;
w26093 <= not w25309 and not w26092;
w26094 <= not w26090 and w26093;
w26095 <= not w25309 and not w26094;
w26096 <= b(58) and not w25298;
w26097 <= not w25296 and w26096;
w26098 <= not w25300 and not w26097;
w26099 <= not w26095 and w26098;
w26100 <= not w25300 and not w26099;
w26101 <= b(59) and not w25289;
w26102 <= not w25287 and w26101;
w26103 <= not w25291 and not w26102;
w26104 <= not w26100 and w26103;
w26105 <= not w25291 and not w26104;
w26106 <= not w24464 and not w25277;
w26107 <= not w25275 and w26106;
w26108 <= not w25263 and w26107;
w26109 <= not w25275 and not w25277;
w26110 <= not w25264 and not w26109;
w26111 <= not w26108 and not w26110;
w26112 <= not w25282 and not w26111;
w26113 <= not w25274 and not w25281;
w26114 <= not w25280 and w26113;
w26115 <= not w26112 and not w26114;
w26116 <= not b(60) and not w26115;
w26117 <= b(60) and not w26114;
w26118 <= not w26112 and w26117;
w26119 <= w146 and not w26118;
w26120 <= not w26116 and w26119;
w26121 <= not w26105 and w26120;
w26122 <= w23 and not w26115;
w26123 <= not w26121 and not w26122;
w26124 <= not w25300 and w26103;
w26125 <= not w26099 and w26124;
w26126 <= not w26100 and not w26103;
w26127 <= not w26125 and not w26126;
w26128 <= not w26123 and not w26127;
w26129 <= not w25290 and not w26122;
w26130 <= not w26121 and w26129;
w26131 <= not w26128 and not w26130;
w26132 <= not b(60) and not w26131;
w26133 <= not w25309 and w26098;
w26134 <= not w26094 and w26133;
w26135 <= not w26095 and not w26098;
w26136 <= not w26134 and not w26135;
w26137 <= not w26123 and not w26136;
w26138 <= not w25299 and not w26122;
w26139 <= not w26121 and w26138;
w26140 <= not w26137 and not w26139;
w26141 <= not b(59) and not w26140;
w26142 <= not w25318 and w26093;
w26143 <= not w26089 and w26142;
w26144 <= not w26090 and not w26093;
w26145 <= not w26143 and not w26144;
w26146 <= not w26123 and not w26145;
w26147 <= not w25308 and not w26122;
w26148 <= not w26121 and w26147;
w26149 <= not w26146 and not w26148;
w26150 <= not b(58) and not w26149;
w26151 <= not w25327 and w26088;
w26152 <= not w26084 and w26151;
w26153 <= not w26085 and not w26088;
w26154 <= not w26152 and not w26153;
w26155 <= not w26123 and not w26154;
w26156 <= not w25317 and not w26122;
w26157 <= not w26121 and w26156;
w26158 <= not w26155 and not w26157;
w26159 <= not b(57) and not w26158;
w26160 <= not w25336 and w26083;
w26161 <= not w26079 and w26160;
w26162 <= not w26080 and not w26083;
w26163 <= not w26161 and not w26162;
w26164 <= not w26123 and not w26163;
w26165 <= not w25326 and not w26122;
w26166 <= not w26121 and w26165;
w26167 <= not w26164 and not w26166;
w26168 <= not b(56) and not w26167;
w26169 <= not w25345 and w26078;
w26170 <= not w26074 and w26169;
w26171 <= not w26075 and not w26078;
w26172 <= not w26170 and not w26171;
w26173 <= not w26123 and not w26172;
w26174 <= not w25335 and not w26122;
w26175 <= not w26121 and w26174;
w26176 <= not w26173 and not w26175;
w26177 <= not b(55) and not w26176;
w26178 <= not w25354 and w26073;
w26179 <= not w26069 and w26178;
w26180 <= not w26070 and not w26073;
w26181 <= not w26179 and not w26180;
w26182 <= not w26123 and not w26181;
w26183 <= not w25344 and not w26122;
w26184 <= not w26121 and w26183;
w26185 <= not w26182 and not w26184;
w26186 <= not b(54) and not w26185;
w26187 <= not w25363 and w26068;
w26188 <= not w26064 and w26187;
w26189 <= not w26065 and not w26068;
w26190 <= not w26188 and not w26189;
w26191 <= not w26123 and not w26190;
w26192 <= not w25353 and not w26122;
w26193 <= not w26121 and w26192;
w26194 <= not w26191 and not w26193;
w26195 <= not b(53) and not w26194;
w26196 <= not w25372 and w26063;
w26197 <= not w26059 and w26196;
w26198 <= not w26060 and not w26063;
w26199 <= not w26197 and not w26198;
w26200 <= not w26123 and not w26199;
w26201 <= not w25362 and not w26122;
w26202 <= not w26121 and w26201;
w26203 <= not w26200 and not w26202;
w26204 <= not b(52) and not w26203;
w26205 <= not w25381 and w26058;
w26206 <= not w26054 and w26205;
w26207 <= not w26055 and not w26058;
w26208 <= not w26206 and not w26207;
w26209 <= not w26123 and not w26208;
w26210 <= not w25371 and not w26122;
w26211 <= not w26121 and w26210;
w26212 <= not w26209 and not w26211;
w26213 <= not b(51) and not w26212;
w26214 <= not w25390 and w26053;
w26215 <= not w26049 and w26214;
w26216 <= not w26050 and not w26053;
w26217 <= not w26215 and not w26216;
w26218 <= not w26123 and not w26217;
w26219 <= not w25380 and not w26122;
w26220 <= not w26121 and w26219;
w26221 <= not w26218 and not w26220;
w26222 <= not b(50) and not w26221;
w26223 <= not w25399 and w26048;
w26224 <= not w26044 and w26223;
w26225 <= not w26045 and not w26048;
w26226 <= not w26224 and not w26225;
w26227 <= not w26123 and not w26226;
w26228 <= not w25389 and not w26122;
w26229 <= not w26121 and w26228;
w26230 <= not w26227 and not w26229;
w26231 <= not b(49) and not w26230;
w26232 <= not w25408 and w26043;
w26233 <= not w26039 and w26232;
w26234 <= not w26040 and not w26043;
w26235 <= not w26233 and not w26234;
w26236 <= not w26123 and not w26235;
w26237 <= not w25398 and not w26122;
w26238 <= not w26121 and w26237;
w26239 <= not w26236 and not w26238;
w26240 <= not b(48) and not w26239;
w26241 <= not w25417 and w26038;
w26242 <= not w26034 and w26241;
w26243 <= not w26035 and not w26038;
w26244 <= not w26242 and not w26243;
w26245 <= not w26123 and not w26244;
w26246 <= not w25407 and not w26122;
w26247 <= not w26121 and w26246;
w26248 <= not w26245 and not w26247;
w26249 <= not b(47) and not w26248;
w26250 <= not w25426 and w26033;
w26251 <= not w26029 and w26250;
w26252 <= not w26030 and not w26033;
w26253 <= not w26251 and not w26252;
w26254 <= not w26123 and not w26253;
w26255 <= not w25416 and not w26122;
w26256 <= not w26121 and w26255;
w26257 <= not w26254 and not w26256;
w26258 <= not b(46) and not w26257;
w26259 <= not w25435 and w26028;
w26260 <= not w26024 and w26259;
w26261 <= not w26025 and not w26028;
w26262 <= not w26260 and not w26261;
w26263 <= not w26123 and not w26262;
w26264 <= not w25425 and not w26122;
w26265 <= not w26121 and w26264;
w26266 <= not w26263 and not w26265;
w26267 <= not b(45) and not w26266;
w26268 <= not w25444 and w26023;
w26269 <= not w26019 and w26268;
w26270 <= not w26020 and not w26023;
w26271 <= not w26269 and not w26270;
w26272 <= not w26123 and not w26271;
w26273 <= not w25434 and not w26122;
w26274 <= not w26121 and w26273;
w26275 <= not w26272 and not w26274;
w26276 <= not b(44) and not w26275;
w26277 <= not w25453 and w26018;
w26278 <= not w26014 and w26277;
w26279 <= not w26015 and not w26018;
w26280 <= not w26278 and not w26279;
w26281 <= not w26123 and not w26280;
w26282 <= not w25443 and not w26122;
w26283 <= not w26121 and w26282;
w26284 <= not w26281 and not w26283;
w26285 <= not b(43) and not w26284;
w26286 <= not w25462 and w26013;
w26287 <= not w26009 and w26286;
w26288 <= not w26010 and not w26013;
w26289 <= not w26287 and not w26288;
w26290 <= not w26123 and not w26289;
w26291 <= not w25452 and not w26122;
w26292 <= not w26121 and w26291;
w26293 <= not w26290 and not w26292;
w26294 <= not b(42) and not w26293;
w26295 <= not w25471 and w26008;
w26296 <= not w26004 and w26295;
w26297 <= not w26005 and not w26008;
w26298 <= not w26296 and not w26297;
w26299 <= not w26123 and not w26298;
w26300 <= not w25461 and not w26122;
w26301 <= not w26121 and w26300;
w26302 <= not w26299 and not w26301;
w26303 <= not b(41) and not w26302;
w26304 <= not w25480 and w26003;
w26305 <= not w25999 and w26304;
w26306 <= not w26000 and not w26003;
w26307 <= not w26305 and not w26306;
w26308 <= not w26123 and not w26307;
w26309 <= not w25470 and not w26122;
w26310 <= not w26121 and w26309;
w26311 <= not w26308 and not w26310;
w26312 <= not b(40) and not w26311;
w26313 <= not w25489 and w25998;
w26314 <= not w25994 and w26313;
w26315 <= not w25995 and not w25998;
w26316 <= not w26314 and not w26315;
w26317 <= not w26123 and not w26316;
w26318 <= not w25479 and not w26122;
w26319 <= not w26121 and w26318;
w26320 <= not w26317 and not w26319;
w26321 <= not b(39) and not w26320;
w26322 <= not w25498 and w25993;
w26323 <= not w25989 and w26322;
w26324 <= not w25990 and not w25993;
w26325 <= not w26323 and not w26324;
w26326 <= not w26123 and not w26325;
w26327 <= not w25488 and not w26122;
w26328 <= not w26121 and w26327;
w26329 <= not w26326 and not w26328;
w26330 <= not b(38) and not w26329;
w26331 <= not w25507 and w25988;
w26332 <= not w25984 and w26331;
w26333 <= not w25985 and not w25988;
w26334 <= not w26332 and not w26333;
w26335 <= not w26123 and not w26334;
w26336 <= not w25497 and not w26122;
w26337 <= not w26121 and w26336;
w26338 <= not w26335 and not w26337;
w26339 <= not b(37) and not w26338;
w26340 <= not w25516 and w25983;
w26341 <= not w25979 and w26340;
w26342 <= not w25980 and not w25983;
w26343 <= not w26341 and not w26342;
w26344 <= not w26123 and not w26343;
w26345 <= not w25506 and not w26122;
w26346 <= not w26121 and w26345;
w26347 <= not w26344 and not w26346;
w26348 <= not b(36) and not w26347;
w26349 <= not w25525 and w25978;
w26350 <= not w25974 and w26349;
w26351 <= not w25975 and not w25978;
w26352 <= not w26350 and not w26351;
w26353 <= not w26123 and not w26352;
w26354 <= not w25515 and not w26122;
w26355 <= not w26121 and w26354;
w26356 <= not w26353 and not w26355;
w26357 <= not b(35) and not w26356;
w26358 <= not w25534 and w25973;
w26359 <= not w25969 and w26358;
w26360 <= not w25970 and not w25973;
w26361 <= not w26359 and not w26360;
w26362 <= not w26123 and not w26361;
w26363 <= not w25524 and not w26122;
w26364 <= not w26121 and w26363;
w26365 <= not w26362 and not w26364;
w26366 <= not b(34) and not w26365;
w26367 <= not w25543 and w25968;
w26368 <= not w25964 and w26367;
w26369 <= not w25965 and not w25968;
w26370 <= not w26368 and not w26369;
w26371 <= not w26123 and not w26370;
w26372 <= not w25533 and not w26122;
w26373 <= not w26121 and w26372;
w26374 <= not w26371 and not w26373;
w26375 <= not b(33) and not w26374;
w26376 <= not w25552 and w25963;
w26377 <= not w25959 and w26376;
w26378 <= not w25960 and not w25963;
w26379 <= not w26377 and not w26378;
w26380 <= not w26123 and not w26379;
w26381 <= not w25542 and not w26122;
w26382 <= not w26121 and w26381;
w26383 <= not w26380 and not w26382;
w26384 <= not b(32) and not w26383;
w26385 <= not w25561 and w25958;
w26386 <= not w25954 and w26385;
w26387 <= not w25955 and not w25958;
w26388 <= not w26386 and not w26387;
w26389 <= not w26123 and not w26388;
w26390 <= not w25551 and not w26122;
w26391 <= not w26121 and w26390;
w26392 <= not w26389 and not w26391;
w26393 <= not b(31) and not w26392;
w26394 <= not w25570 and w25953;
w26395 <= not w25949 and w26394;
w26396 <= not w25950 and not w25953;
w26397 <= not w26395 and not w26396;
w26398 <= not w26123 and not w26397;
w26399 <= not w25560 and not w26122;
w26400 <= not w26121 and w26399;
w26401 <= not w26398 and not w26400;
w26402 <= not b(30) and not w26401;
w26403 <= not w25579 and w25948;
w26404 <= not w25944 and w26403;
w26405 <= not w25945 and not w25948;
w26406 <= not w26404 and not w26405;
w26407 <= not w26123 and not w26406;
w26408 <= not w25569 and not w26122;
w26409 <= not w26121 and w26408;
w26410 <= not w26407 and not w26409;
w26411 <= not b(29) and not w26410;
w26412 <= not w25588 and w25943;
w26413 <= not w25939 and w26412;
w26414 <= not w25940 and not w25943;
w26415 <= not w26413 and not w26414;
w26416 <= not w26123 and not w26415;
w26417 <= not w25578 and not w26122;
w26418 <= not w26121 and w26417;
w26419 <= not w26416 and not w26418;
w26420 <= not b(28) and not w26419;
w26421 <= not w25597 and w25938;
w26422 <= not w25934 and w26421;
w26423 <= not w25935 and not w25938;
w26424 <= not w26422 and not w26423;
w26425 <= not w26123 and not w26424;
w26426 <= not w25587 and not w26122;
w26427 <= not w26121 and w26426;
w26428 <= not w26425 and not w26427;
w26429 <= not b(27) and not w26428;
w26430 <= not w25606 and w25933;
w26431 <= not w25929 and w26430;
w26432 <= not w25930 and not w25933;
w26433 <= not w26431 and not w26432;
w26434 <= not w26123 and not w26433;
w26435 <= not w25596 and not w26122;
w26436 <= not w26121 and w26435;
w26437 <= not w26434 and not w26436;
w26438 <= not b(26) and not w26437;
w26439 <= not w25615 and w25928;
w26440 <= not w25924 and w26439;
w26441 <= not w25925 and not w25928;
w26442 <= not w26440 and not w26441;
w26443 <= not w26123 and not w26442;
w26444 <= not w25605 and not w26122;
w26445 <= not w26121 and w26444;
w26446 <= not w26443 and not w26445;
w26447 <= not b(25) and not w26446;
w26448 <= not w25624 and w25923;
w26449 <= not w25919 and w26448;
w26450 <= not w25920 and not w25923;
w26451 <= not w26449 and not w26450;
w26452 <= not w26123 and not w26451;
w26453 <= not w25614 and not w26122;
w26454 <= not w26121 and w26453;
w26455 <= not w26452 and not w26454;
w26456 <= not b(24) and not w26455;
w26457 <= not w25633 and w25918;
w26458 <= not w25914 and w26457;
w26459 <= not w25915 and not w25918;
w26460 <= not w26458 and not w26459;
w26461 <= not w26123 and not w26460;
w26462 <= not w25623 and not w26122;
w26463 <= not w26121 and w26462;
w26464 <= not w26461 and not w26463;
w26465 <= not b(23) and not w26464;
w26466 <= not w25642 and w25913;
w26467 <= not w25909 and w26466;
w26468 <= not w25910 and not w25913;
w26469 <= not w26467 and not w26468;
w26470 <= not w26123 and not w26469;
w26471 <= not w25632 and not w26122;
w26472 <= not w26121 and w26471;
w26473 <= not w26470 and not w26472;
w26474 <= not b(22) and not w26473;
w26475 <= not w25651 and w25908;
w26476 <= not w25904 and w26475;
w26477 <= not w25905 and not w25908;
w26478 <= not w26476 and not w26477;
w26479 <= not w26123 and not w26478;
w26480 <= not w25641 and not w26122;
w26481 <= not w26121 and w26480;
w26482 <= not w26479 and not w26481;
w26483 <= not b(21) and not w26482;
w26484 <= not w25660 and w25903;
w26485 <= not w25899 and w26484;
w26486 <= not w25900 and not w25903;
w26487 <= not w26485 and not w26486;
w26488 <= not w26123 and not w26487;
w26489 <= not w25650 and not w26122;
w26490 <= not w26121 and w26489;
w26491 <= not w26488 and not w26490;
w26492 <= not b(20) and not w26491;
w26493 <= not w25669 and w25898;
w26494 <= not w25894 and w26493;
w26495 <= not w25895 and not w25898;
w26496 <= not w26494 and not w26495;
w26497 <= not w26123 and not w26496;
w26498 <= not w25659 and not w26122;
w26499 <= not w26121 and w26498;
w26500 <= not w26497 and not w26499;
w26501 <= not b(19) and not w26500;
w26502 <= not w25678 and w25893;
w26503 <= not w25889 and w26502;
w26504 <= not w25890 and not w25893;
w26505 <= not w26503 and not w26504;
w26506 <= not w26123 and not w26505;
w26507 <= not w25668 and not w26122;
w26508 <= not w26121 and w26507;
w26509 <= not w26506 and not w26508;
w26510 <= not b(18) and not w26509;
w26511 <= not w25687 and w25888;
w26512 <= not w25884 and w26511;
w26513 <= not w25885 and not w25888;
w26514 <= not w26512 and not w26513;
w26515 <= not w26123 and not w26514;
w26516 <= not w25677 and not w26122;
w26517 <= not w26121 and w26516;
w26518 <= not w26515 and not w26517;
w26519 <= not b(17) and not w26518;
w26520 <= not w25696 and w25883;
w26521 <= not w25879 and w26520;
w26522 <= not w25880 and not w25883;
w26523 <= not w26521 and not w26522;
w26524 <= not w26123 and not w26523;
w26525 <= not w25686 and not w26122;
w26526 <= not w26121 and w26525;
w26527 <= not w26524 and not w26526;
w26528 <= not b(16) and not w26527;
w26529 <= not w25705 and w25878;
w26530 <= not w25874 and w26529;
w26531 <= not w25875 and not w25878;
w26532 <= not w26530 and not w26531;
w26533 <= not w26123 and not w26532;
w26534 <= not w25695 and not w26122;
w26535 <= not w26121 and w26534;
w26536 <= not w26533 and not w26535;
w26537 <= not b(15) and not w26536;
w26538 <= not w25714 and w25873;
w26539 <= not w25869 and w26538;
w26540 <= not w25870 and not w25873;
w26541 <= not w26539 and not w26540;
w26542 <= not w26123 and not w26541;
w26543 <= not w25704 and not w26122;
w26544 <= not w26121 and w26543;
w26545 <= not w26542 and not w26544;
w26546 <= not b(14) and not w26545;
w26547 <= not w25723 and w25868;
w26548 <= not w25864 and w26547;
w26549 <= not w25865 and not w25868;
w26550 <= not w26548 and not w26549;
w26551 <= not w26123 and not w26550;
w26552 <= not w25713 and not w26122;
w26553 <= not w26121 and w26552;
w26554 <= not w26551 and not w26553;
w26555 <= not b(13) and not w26554;
w26556 <= not w25732 and w25863;
w26557 <= not w25859 and w26556;
w26558 <= not w25860 and not w25863;
w26559 <= not w26557 and not w26558;
w26560 <= not w26123 and not w26559;
w26561 <= not w25722 and not w26122;
w26562 <= not w26121 and w26561;
w26563 <= not w26560 and not w26562;
w26564 <= not b(12) and not w26563;
w26565 <= not w25741 and w25858;
w26566 <= not w25854 and w26565;
w26567 <= not w25855 and not w25858;
w26568 <= not w26566 and not w26567;
w26569 <= not w26123 and not w26568;
w26570 <= not w25731 and not w26122;
w26571 <= not w26121 and w26570;
w26572 <= not w26569 and not w26571;
w26573 <= not b(11) and not w26572;
w26574 <= not w25750 and w25853;
w26575 <= not w25849 and w26574;
w26576 <= not w25850 and not w25853;
w26577 <= not w26575 and not w26576;
w26578 <= not w26123 and not w26577;
w26579 <= not w25740 and not w26122;
w26580 <= not w26121 and w26579;
w26581 <= not w26578 and not w26580;
w26582 <= not b(10) and not w26581;
w26583 <= not w25759 and w25848;
w26584 <= not w25844 and w26583;
w26585 <= not w25845 and not w25848;
w26586 <= not w26584 and not w26585;
w26587 <= not w26123 and not w26586;
w26588 <= not w25749 and not w26122;
w26589 <= not w26121 and w26588;
w26590 <= not w26587 and not w26589;
w26591 <= not b(9) and not w26590;
w26592 <= not w25768 and w25843;
w26593 <= not w25839 and w26592;
w26594 <= not w25840 and not w25843;
w26595 <= not w26593 and not w26594;
w26596 <= not w26123 and not w26595;
w26597 <= not w25758 and not w26122;
w26598 <= not w26121 and w26597;
w26599 <= not w26596 and not w26598;
w26600 <= not b(8) and not w26599;
w26601 <= not w25777 and w25838;
w26602 <= not w25834 and w26601;
w26603 <= not w25835 and not w25838;
w26604 <= not w26602 and not w26603;
w26605 <= not w26123 and not w26604;
w26606 <= not w25767 and not w26122;
w26607 <= not w26121 and w26606;
w26608 <= not w26605 and not w26607;
w26609 <= not b(7) and not w26608;
w26610 <= not w25786 and w25833;
w26611 <= not w25829 and w26610;
w26612 <= not w25830 and not w25833;
w26613 <= not w26611 and not w26612;
w26614 <= not w26123 and not w26613;
w26615 <= not w25776 and not w26122;
w26616 <= not w26121 and w26615;
w26617 <= not w26614 and not w26616;
w26618 <= not b(6) and not w26617;
w26619 <= not w25795 and w25828;
w26620 <= not w25824 and w26619;
w26621 <= not w25825 and not w25828;
w26622 <= not w26620 and not w26621;
w26623 <= not w26123 and not w26622;
w26624 <= not w25785 and not w26122;
w26625 <= not w26121 and w26624;
w26626 <= not w26623 and not w26625;
w26627 <= not b(5) and not w26626;
w26628 <= not w25803 and w25823;
w26629 <= not w25819 and w26628;
w26630 <= not w25820 and not w25823;
w26631 <= not w26629 and not w26630;
w26632 <= not w26123 and not w26631;
w26633 <= not w25794 and not w26122;
w26634 <= not w26121 and w26633;
w26635 <= not w26632 and not w26634;
w26636 <= not b(4) and not w26635;
w26637 <= not w25814 and w25818;
w26638 <= not w25813 and w26637;
w26639 <= not w25815 and not w25818;
w26640 <= not w26638 and not w26639;
w26641 <= not w26123 and not w26640;
w26642 <= not w25802 and not w26122;
w26643 <= not w26121 and w26642;
w26644 <= not w26641 and not w26643;
w26645 <= not b(3) and not w26644;
w26646 <= not w25810 and w25812;
w26647 <= not w25808 and w26646;
w26648 <= not w25813 and not w26647;
w26649 <= not w26123 and w26648;
w26650 <= not w25807 and not w26122;
w26651 <= not w26121 and w26650;
w26652 <= not w26649 and not w26651;
w26653 <= not b(2) and not w26652;
w26654 <= b(0) and not w26123;
w26655 <= a(3) and not w26654;
w26656 <= w25812 and not w26123;
w26657 <= not w26655 and not w26656;
w26658 <= b(1) and not w26657;
w26659 <= not b(1) and not w26656;
w26660 <= not w26655 and w26659;
w26661 <= not w26658 and not w26660;
w26662 <= not a(2) and b(0);
w26663 <= not w26661 and not w26662;
w26664 <= not b(1) and not w26657;
w26665 <= not w26663 and not w26664;
w26666 <= b(2) and not w26651;
w26667 <= not w26649 and w26666;
w26668 <= not w26653 and not w26667;
w26669 <= not w26665 and w26668;
w26670 <= not w26653 and not w26669;
w26671 <= b(3) and not w26643;
w26672 <= not w26641 and w26671;
w26673 <= not w26645 and not w26672;
w26674 <= not w26670 and w26673;
w26675 <= not w26645 and not w26674;
w26676 <= b(4) and not w26634;
w26677 <= not w26632 and w26676;
w26678 <= not w26636 and not w26677;
w26679 <= not w26675 and w26678;
w26680 <= not w26636 and not w26679;
w26681 <= b(5) and not w26625;
w26682 <= not w26623 and w26681;
w26683 <= not w26627 and not w26682;
w26684 <= not w26680 and w26683;
w26685 <= not w26627 and not w26684;
w26686 <= b(6) and not w26616;
w26687 <= not w26614 and w26686;
w26688 <= not w26618 and not w26687;
w26689 <= not w26685 and w26688;
w26690 <= not w26618 and not w26689;
w26691 <= b(7) and not w26607;
w26692 <= not w26605 and w26691;
w26693 <= not w26609 and not w26692;
w26694 <= not w26690 and w26693;
w26695 <= not w26609 and not w26694;
w26696 <= b(8) and not w26598;
w26697 <= not w26596 and w26696;
w26698 <= not w26600 and not w26697;
w26699 <= not w26695 and w26698;
w26700 <= not w26600 and not w26699;
w26701 <= b(9) and not w26589;
w26702 <= not w26587 and w26701;
w26703 <= not w26591 and not w26702;
w26704 <= not w26700 and w26703;
w26705 <= not w26591 and not w26704;
w26706 <= b(10) and not w26580;
w26707 <= not w26578 and w26706;
w26708 <= not w26582 and not w26707;
w26709 <= not w26705 and w26708;
w26710 <= not w26582 and not w26709;
w26711 <= b(11) and not w26571;
w26712 <= not w26569 and w26711;
w26713 <= not w26573 and not w26712;
w26714 <= not w26710 and w26713;
w26715 <= not w26573 and not w26714;
w26716 <= b(12) and not w26562;
w26717 <= not w26560 and w26716;
w26718 <= not w26564 and not w26717;
w26719 <= not w26715 and w26718;
w26720 <= not w26564 and not w26719;
w26721 <= b(13) and not w26553;
w26722 <= not w26551 and w26721;
w26723 <= not w26555 and not w26722;
w26724 <= not w26720 and w26723;
w26725 <= not w26555 and not w26724;
w26726 <= b(14) and not w26544;
w26727 <= not w26542 and w26726;
w26728 <= not w26546 and not w26727;
w26729 <= not w26725 and w26728;
w26730 <= not w26546 and not w26729;
w26731 <= b(15) and not w26535;
w26732 <= not w26533 and w26731;
w26733 <= not w26537 and not w26732;
w26734 <= not w26730 and w26733;
w26735 <= not w26537 and not w26734;
w26736 <= b(16) and not w26526;
w26737 <= not w26524 and w26736;
w26738 <= not w26528 and not w26737;
w26739 <= not w26735 and w26738;
w26740 <= not w26528 and not w26739;
w26741 <= b(17) and not w26517;
w26742 <= not w26515 and w26741;
w26743 <= not w26519 and not w26742;
w26744 <= not w26740 and w26743;
w26745 <= not w26519 and not w26744;
w26746 <= b(18) and not w26508;
w26747 <= not w26506 and w26746;
w26748 <= not w26510 and not w26747;
w26749 <= not w26745 and w26748;
w26750 <= not w26510 and not w26749;
w26751 <= b(19) and not w26499;
w26752 <= not w26497 and w26751;
w26753 <= not w26501 and not w26752;
w26754 <= not w26750 and w26753;
w26755 <= not w26501 and not w26754;
w26756 <= b(20) and not w26490;
w26757 <= not w26488 and w26756;
w26758 <= not w26492 and not w26757;
w26759 <= not w26755 and w26758;
w26760 <= not w26492 and not w26759;
w26761 <= b(21) and not w26481;
w26762 <= not w26479 and w26761;
w26763 <= not w26483 and not w26762;
w26764 <= not w26760 and w26763;
w26765 <= not w26483 and not w26764;
w26766 <= b(22) and not w26472;
w26767 <= not w26470 and w26766;
w26768 <= not w26474 and not w26767;
w26769 <= not w26765 and w26768;
w26770 <= not w26474 and not w26769;
w26771 <= b(23) and not w26463;
w26772 <= not w26461 and w26771;
w26773 <= not w26465 and not w26772;
w26774 <= not w26770 and w26773;
w26775 <= not w26465 and not w26774;
w26776 <= b(24) and not w26454;
w26777 <= not w26452 and w26776;
w26778 <= not w26456 and not w26777;
w26779 <= not w26775 and w26778;
w26780 <= not w26456 and not w26779;
w26781 <= b(25) and not w26445;
w26782 <= not w26443 and w26781;
w26783 <= not w26447 and not w26782;
w26784 <= not w26780 and w26783;
w26785 <= not w26447 and not w26784;
w26786 <= b(26) and not w26436;
w26787 <= not w26434 and w26786;
w26788 <= not w26438 and not w26787;
w26789 <= not w26785 and w26788;
w26790 <= not w26438 and not w26789;
w26791 <= b(27) and not w26427;
w26792 <= not w26425 and w26791;
w26793 <= not w26429 and not w26792;
w26794 <= not w26790 and w26793;
w26795 <= not w26429 and not w26794;
w26796 <= b(28) and not w26418;
w26797 <= not w26416 and w26796;
w26798 <= not w26420 and not w26797;
w26799 <= not w26795 and w26798;
w26800 <= not w26420 and not w26799;
w26801 <= b(29) and not w26409;
w26802 <= not w26407 and w26801;
w26803 <= not w26411 and not w26802;
w26804 <= not w26800 and w26803;
w26805 <= not w26411 and not w26804;
w26806 <= b(30) and not w26400;
w26807 <= not w26398 and w26806;
w26808 <= not w26402 and not w26807;
w26809 <= not w26805 and w26808;
w26810 <= not w26402 and not w26809;
w26811 <= b(31) and not w26391;
w26812 <= not w26389 and w26811;
w26813 <= not w26393 and not w26812;
w26814 <= not w26810 and w26813;
w26815 <= not w26393 and not w26814;
w26816 <= b(32) and not w26382;
w26817 <= not w26380 and w26816;
w26818 <= not w26384 and not w26817;
w26819 <= not w26815 and w26818;
w26820 <= not w26384 and not w26819;
w26821 <= b(33) and not w26373;
w26822 <= not w26371 and w26821;
w26823 <= not w26375 and not w26822;
w26824 <= not w26820 and w26823;
w26825 <= not w26375 and not w26824;
w26826 <= b(34) and not w26364;
w26827 <= not w26362 and w26826;
w26828 <= not w26366 and not w26827;
w26829 <= not w26825 and w26828;
w26830 <= not w26366 and not w26829;
w26831 <= b(35) and not w26355;
w26832 <= not w26353 and w26831;
w26833 <= not w26357 and not w26832;
w26834 <= not w26830 and w26833;
w26835 <= not w26357 and not w26834;
w26836 <= b(36) and not w26346;
w26837 <= not w26344 and w26836;
w26838 <= not w26348 and not w26837;
w26839 <= not w26835 and w26838;
w26840 <= not w26348 and not w26839;
w26841 <= b(37) and not w26337;
w26842 <= not w26335 and w26841;
w26843 <= not w26339 and not w26842;
w26844 <= not w26840 and w26843;
w26845 <= not w26339 and not w26844;
w26846 <= b(38) and not w26328;
w26847 <= not w26326 and w26846;
w26848 <= not w26330 and not w26847;
w26849 <= not w26845 and w26848;
w26850 <= not w26330 and not w26849;
w26851 <= b(39) and not w26319;
w26852 <= not w26317 and w26851;
w26853 <= not w26321 and not w26852;
w26854 <= not w26850 and w26853;
w26855 <= not w26321 and not w26854;
w26856 <= b(40) and not w26310;
w26857 <= not w26308 and w26856;
w26858 <= not w26312 and not w26857;
w26859 <= not w26855 and w26858;
w26860 <= not w26312 and not w26859;
w26861 <= b(41) and not w26301;
w26862 <= not w26299 and w26861;
w26863 <= not w26303 and not w26862;
w26864 <= not w26860 and w26863;
w26865 <= not w26303 and not w26864;
w26866 <= b(42) and not w26292;
w26867 <= not w26290 and w26866;
w26868 <= not w26294 and not w26867;
w26869 <= not w26865 and w26868;
w26870 <= not w26294 and not w26869;
w26871 <= b(43) and not w26283;
w26872 <= not w26281 and w26871;
w26873 <= not w26285 and not w26872;
w26874 <= not w26870 and w26873;
w26875 <= not w26285 and not w26874;
w26876 <= b(44) and not w26274;
w26877 <= not w26272 and w26876;
w26878 <= not w26276 and not w26877;
w26879 <= not w26875 and w26878;
w26880 <= not w26276 and not w26879;
w26881 <= b(45) and not w26265;
w26882 <= not w26263 and w26881;
w26883 <= not w26267 and not w26882;
w26884 <= not w26880 and w26883;
w26885 <= not w26267 and not w26884;
w26886 <= b(46) and not w26256;
w26887 <= not w26254 and w26886;
w26888 <= not w26258 and not w26887;
w26889 <= not w26885 and w26888;
w26890 <= not w26258 and not w26889;
w26891 <= b(47) and not w26247;
w26892 <= not w26245 and w26891;
w26893 <= not w26249 and not w26892;
w26894 <= not w26890 and w26893;
w26895 <= not w26249 and not w26894;
w26896 <= b(48) and not w26238;
w26897 <= not w26236 and w26896;
w26898 <= not w26240 and not w26897;
w26899 <= not w26895 and w26898;
w26900 <= not w26240 and not w26899;
w26901 <= b(49) and not w26229;
w26902 <= not w26227 and w26901;
w26903 <= not w26231 and not w26902;
w26904 <= not w26900 and w26903;
w26905 <= not w26231 and not w26904;
w26906 <= b(50) and not w26220;
w26907 <= not w26218 and w26906;
w26908 <= not w26222 and not w26907;
w26909 <= not w26905 and w26908;
w26910 <= not w26222 and not w26909;
w26911 <= b(51) and not w26211;
w26912 <= not w26209 and w26911;
w26913 <= not w26213 and not w26912;
w26914 <= not w26910 and w26913;
w26915 <= not w26213 and not w26914;
w26916 <= b(52) and not w26202;
w26917 <= not w26200 and w26916;
w26918 <= not w26204 and not w26917;
w26919 <= not w26915 and w26918;
w26920 <= not w26204 and not w26919;
w26921 <= b(53) and not w26193;
w26922 <= not w26191 and w26921;
w26923 <= not w26195 and not w26922;
w26924 <= not w26920 and w26923;
w26925 <= not w26195 and not w26924;
w26926 <= b(54) and not w26184;
w26927 <= not w26182 and w26926;
w26928 <= not w26186 and not w26927;
w26929 <= not w26925 and w26928;
w26930 <= not w26186 and not w26929;
w26931 <= b(55) and not w26175;
w26932 <= not w26173 and w26931;
w26933 <= not w26177 and not w26932;
w26934 <= not w26930 and w26933;
w26935 <= not w26177 and not w26934;
w26936 <= b(56) and not w26166;
w26937 <= not w26164 and w26936;
w26938 <= not w26168 and not w26937;
w26939 <= not w26935 and w26938;
w26940 <= not w26168 and not w26939;
w26941 <= b(57) and not w26157;
w26942 <= not w26155 and w26941;
w26943 <= not w26159 and not w26942;
w26944 <= not w26940 and w26943;
w26945 <= not w26159 and not w26944;
w26946 <= b(58) and not w26148;
w26947 <= not w26146 and w26946;
w26948 <= not w26150 and not w26947;
w26949 <= not w26945 and w26948;
w26950 <= not w26150 and not w26949;
w26951 <= b(59) and not w26139;
w26952 <= not w26137 and w26951;
w26953 <= not w26141 and not w26952;
w26954 <= not w26950 and w26953;
w26955 <= not w26141 and not w26954;
w26956 <= b(60) and not w26130;
w26957 <= not w26128 and w26956;
w26958 <= not w26132 and not w26957;
w26959 <= not w26955 and w26958;
w26960 <= not w26132 and not w26959;
w26961 <= not w25291 and not w26118;
w26962 <= not w26116 and w26961;
w26963 <= not w26104 and w26962;
w26964 <= not w26116 and not w26118;
w26965 <= not w26105 and not w26964;
w26966 <= not w26963 and not w26965;
w26967 <= not w26123 and not w26966;
w26968 <= not w26115 and not w26122;
w26969 <= not w26121 and w26968;
w26970 <= not w26967 and not w26969;
w26971 <= not b(61) and not w26970;
w26972 <= b(61) and not w26969;
w26973 <= not w26967 and w26972;
w26974 <= w22 and not w26973;
w26975 <= not w26971 and w26974;
w26976 <= not w26960 and w26975;
w26977 <= w146 and not w26970;
w26978 <= not w26976 and not w26977;
w26979 <= not w26141 and w26958;
w26980 <= not w26954 and w26979;
w26981 <= not w26955 and not w26958;
w26982 <= not w26980 and not w26981;
w26983 <= not w26978 and not w26982;
w26984 <= not w26131 and not w26977;
w26985 <= not w26976 and w26984;
w26986 <= not w26983 and not w26985;
w26987 <= not b(61) and not w26986;
w26988 <= not w26150 and w26953;
w26989 <= not w26949 and w26988;
w26990 <= not w26950 and not w26953;
w26991 <= not w26989 and not w26990;
w26992 <= not w26978 and not w26991;
w26993 <= not w26140 and not w26977;
w26994 <= not w26976 and w26993;
w26995 <= not w26992 and not w26994;
w26996 <= not b(60) and not w26995;
w26997 <= not w26159 and w26948;
w26998 <= not w26944 and w26997;
w26999 <= not w26945 and not w26948;
w27000 <= not w26998 and not w26999;
w27001 <= not w26978 and not w27000;
w27002 <= not w26149 and not w26977;
w27003 <= not w26976 and w27002;
w27004 <= not w27001 and not w27003;
w27005 <= not b(59) and not w27004;
w27006 <= not w26168 and w26943;
w27007 <= not w26939 and w27006;
w27008 <= not w26940 and not w26943;
w27009 <= not w27007 and not w27008;
w27010 <= not w26978 and not w27009;
w27011 <= not w26158 and not w26977;
w27012 <= not w26976 and w27011;
w27013 <= not w27010 and not w27012;
w27014 <= not b(58) and not w27013;
w27015 <= not w26177 and w26938;
w27016 <= not w26934 and w27015;
w27017 <= not w26935 and not w26938;
w27018 <= not w27016 and not w27017;
w27019 <= not w26978 and not w27018;
w27020 <= not w26167 and not w26977;
w27021 <= not w26976 and w27020;
w27022 <= not w27019 and not w27021;
w27023 <= not b(57) and not w27022;
w27024 <= not w26186 and w26933;
w27025 <= not w26929 and w27024;
w27026 <= not w26930 and not w26933;
w27027 <= not w27025 and not w27026;
w27028 <= not w26978 and not w27027;
w27029 <= not w26176 and not w26977;
w27030 <= not w26976 and w27029;
w27031 <= not w27028 and not w27030;
w27032 <= not b(56) and not w27031;
w27033 <= not w26195 and w26928;
w27034 <= not w26924 and w27033;
w27035 <= not w26925 and not w26928;
w27036 <= not w27034 and not w27035;
w27037 <= not w26978 and not w27036;
w27038 <= not w26185 and not w26977;
w27039 <= not w26976 and w27038;
w27040 <= not w27037 and not w27039;
w27041 <= not b(55) and not w27040;
w27042 <= not w26204 and w26923;
w27043 <= not w26919 and w27042;
w27044 <= not w26920 and not w26923;
w27045 <= not w27043 and not w27044;
w27046 <= not w26978 and not w27045;
w27047 <= not w26194 and not w26977;
w27048 <= not w26976 and w27047;
w27049 <= not w27046 and not w27048;
w27050 <= not b(54) and not w27049;
w27051 <= not w26213 and w26918;
w27052 <= not w26914 and w27051;
w27053 <= not w26915 and not w26918;
w27054 <= not w27052 and not w27053;
w27055 <= not w26978 and not w27054;
w27056 <= not w26203 and not w26977;
w27057 <= not w26976 and w27056;
w27058 <= not w27055 and not w27057;
w27059 <= not b(53) and not w27058;
w27060 <= not w26222 and w26913;
w27061 <= not w26909 and w27060;
w27062 <= not w26910 and not w26913;
w27063 <= not w27061 and not w27062;
w27064 <= not w26978 and not w27063;
w27065 <= not w26212 and not w26977;
w27066 <= not w26976 and w27065;
w27067 <= not w27064 and not w27066;
w27068 <= not b(52) and not w27067;
w27069 <= not w26231 and w26908;
w27070 <= not w26904 and w27069;
w27071 <= not w26905 and not w26908;
w27072 <= not w27070 and not w27071;
w27073 <= not w26978 and not w27072;
w27074 <= not w26221 and not w26977;
w27075 <= not w26976 and w27074;
w27076 <= not w27073 and not w27075;
w27077 <= not b(51) and not w27076;
w27078 <= not w26240 and w26903;
w27079 <= not w26899 and w27078;
w27080 <= not w26900 and not w26903;
w27081 <= not w27079 and not w27080;
w27082 <= not w26978 and not w27081;
w27083 <= not w26230 and not w26977;
w27084 <= not w26976 and w27083;
w27085 <= not w27082 and not w27084;
w27086 <= not b(50) and not w27085;
w27087 <= not w26249 and w26898;
w27088 <= not w26894 and w27087;
w27089 <= not w26895 and not w26898;
w27090 <= not w27088 and not w27089;
w27091 <= not w26978 and not w27090;
w27092 <= not w26239 and not w26977;
w27093 <= not w26976 and w27092;
w27094 <= not w27091 and not w27093;
w27095 <= not b(49) and not w27094;
w27096 <= not w26258 and w26893;
w27097 <= not w26889 and w27096;
w27098 <= not w26890 and not w26893;
w27099 <= not w27097 and not w27098;
w27100 <= not w26978 and not w27099;
w27101 <= not w26248 and not w26977;
w27102 <= not w26976 and w27101;
w27103 <= not w27100 and not w27102;
w27104 <= not b(48) and not w27103;
w27105 <= not w26267 and w26888;
w27106 <= not w26884 and w27105;
w27107 <= not w26885 and not w26888;
w27108 <= not w27106 and not w27107;
w27109 <= not w26978 and not w27108;
w27110 <= not w26257 and not w26977;
w27111 <= not w26976 and w27110;
w27112 <= not w27109 and not w27111;
w27113 <= not b(47) and not w27112;
w27114 <= not w26276 and w26883;
w27115 <= not w26879 and w27114;
w27116 <= not w26880 and not w26883;
w27117 <= not w27115 and not w27116;
w27118 <= not w26978 and not w27117;
w27119 <= not w26266 and not w26977;
w27120 <= not w26976 and w27119;
w27121 <= not w27118 and not w27120;
w27122 <= not b(46) and not w27121;
w27123 <= not w26285 and w26878;
w27124 <= not w26874 and w27123;
w27125 <= not w26875 and not w26878;
w27126 <= not w27124 and not w27125;
w27127 <= not w26978 and not w27126;
w27128 <= not w26275 and not w26977;
w27129 <= not w26976 and w27128;
w27130 <= not w27127 and not w27129;
w27131 <= not b(45) and not w27130;
w27132 <= not w26294 and w26873;
w27133 <= not w26869 and w27132;
w27134 <= not w26870 and not w26873;
w27135 <= not w27133 and not w27134;
w27136 <= not w26978 and not w27135;
w27137 <= not w26284 and not w26977;
w27138 <= not w26976 and w27137;
w27139 <= not w27136 and not w27138;
w27140 <= not b(44) and not w27139;
w27141 <= not w26303 and w26868;
w27142 <= not w26864 and w27141;
w27143 <= not w26865 and not w26868;
w27144 <= not w27142 and not w27143;
w27145 <= not w26978 and not w27144;
w27146 <= not w26293 and not w26977;
w27147 <= not w26976 and w27146;
w27148 <= not w27145 and not w27147;
w27149 <= not b(43) and not w27148;
w27150 <= not w26312 and w26863;
w27151 <= not w26859 and w27150;
w27152 <= not w26860 and not w26863;
w27153 <= not w27151 and not w27152;
w27154 <= not w26978 and not w27153;
w27155 <= not w26302 and not w26977;
w27156 <= not w26976 and w27155;
w27157 <= not w27154 and not w27156;
w27158 <= not b(42) and not w27157;
w27159 <= not w26321 and w26858;
w27160 <= not w26854 and w27159;
w27161 <= not w26855 and not w26858;
w27162 <= not w27160 and not w27161;
w27163 <= not w26978 and not w27162;
w27164 <= not w26311 and not w26977;
w27165 <= not w26976 and w27164;
w27166 <= not w27163 and not w27165;
w27167 <= not b(41) and not w27166;
w27168 <= not w26330 and w26853;
w27169 <= not w26849 and w27168;
w27170 <= not w26850 and not w26853;
w27171 <= not w27169 and not w27170;
w27172 <= not w26978 and not w27171;
w27173 <= not w26320 and not w26977;
w27174 <= not w26976 and w27173;
w27175 <= not w27172 and not w27174;
w27176 <= not b(40) and not w27175;
w27177 <= not w26339 and w26848;
w27178 <= not w26844 and w27177;
w27179 <= not w26845 and not w26848;
w27180 <= not w27178 and not w27179;
w27181 <= not w26978 and not w27180;
w27182 <= not w26329 and not w26977;
w27183 <= not w26976 and w27182;
w27184 <= not w27181 and not w27183;
w27185 <= not b(39) and not w27184;
w27186 <= not w26348 and w26843;
w27187 <= not w26839 and w27186;
w27188 <= not w26840 and not w26843;
w27189 <= not w27187 and not w27188;
w27190 <= not w26978 and not w27189;
w27191 <= not w26338 and not w26977;
w27192 <= not w26976 and w27191;
w27193 <= not w27190 and not w27192;
w27194 <= not b(38) and not w27193;
w27195 <= not w26357 and w26838;
w27196 <= not w26834 and w27195;
w27197 <= not w26835 and not w26838;
w27198 <= not w27196 and not w27197;
w27199 <= not w26978 and not w27198;
w27200 <= not w26347 and not w26977;
w27201 <= not w26976 and w27200;
w27202 <= not w27199 and not w27201;
w27203 <= not b(37) and not w27202;
w27204 <= not w26366 and w26833;
w27205 <= not w26829 and w27204;
w27206 <= not w26830 and not w26833;
w27207 <= not w27205 and not w27206;
w27208 <= not w26978 and not w27207;
w27209 <= not w26356 and not w26977;
w27210 <= not w26976 and w27209;
w27211 <= not w27208 and not w27210;
w27212 <= not b(36) and not w27211;
w27213 <= not w26375 and w26828;
w27214 <= not w26824 and w27213;
w27215 <= not w26825 and not w26828;
w27216 <= not w27214 and not w27215;
w27217 <= not w26978 and not w27216;
w27218 <= not w26365 and not w26977;
w27219 <= not w26976 and w27218;
w27220 <= not w27217 and not w27219;
w27221 <= not b(35) and not w27220;
w27222 <= not w26384 and w26823;
w27223 <= not w26819 and w27222;
w27224 <= not w26820 and not w26823;
w27225 <= not w27223 and not w27224;
w27226 <= not w26978 and not w27225;
w27227 <= not w26374 and not w26977;
w27228 <= not w26976 and w27227;
w27229 <= not w27226 and not w27228;
w27230 <= not b(34) and not w27229;
w27231 <= not w26393 and w26818;
w27232 <= not w26814 and w27231;
w27233 <= not w26815 and not w26818;
w27234 <= not w27232 and not w27233;
w27235 <= not w26978 and not w27234;
w27236 <= not w26383 and not w26977;
w27237 <= not w26976 and w27236;
w27238 <= not w27235 and not w27237;
w27239 <= not b(33) and not w27238;
w27240 <= not w26402 and w26813;
w27241 <= not w26809 and w27240;
w27242 <= not w26810 and not w26813;
w27243 <= not w27241 and not w27242;
w27244 <= not w26978 and not w27243;
w27245 <= not w26392 and not w26977;
w27246 <= not w26976 and w27245;
w27247 <= not w27244 and not w27246;
w27248 <= not b(32) and not w27247;
w27249 <= not w26411 and w26808;
w27250 <= not w26804 and w27249;
w27251 <= not w26805 and not w26808;
w27252 <= not w27250 and not w27251;
w27253 <= not w26978 and not w27252;
w27254 <= not w26401 and not w26977;
w27255 <= not w26976 and w27254;
w27256 <= not w27253 and not w27255;
w27257 <= not b(31) and not w27256;
w27258 <= not w26420 and w26803;
w27259 <= not w26799 and w27258;
w27260 <= not w26800 and not w26803;
w27261 <= not w27259 and not w27260;
w27262 <= not w26978 and not w27261;
w27263 <= not w26410 and not w26977;
w27264 <= not w26976 and w27263;
w27265 <= not w27262 and not w27264;
w27266 <= not b(30) and not w27265;
w27267 <= not w26429 and w26798;
w27268 <= not w26794 and w27267;
w27269 <= not w26795 and not w26798;
w27270 <= not w27268 and not w27269;
w27271 <= not w26978 and not w27270;
w27272 <= not w26419 and not w26977;
w27273 <= not w26976 and w27272;
w27274 <= not w27271 and not w27273;
w27275 <= not b(29) and not w27274;
w27276 <= not w26438 and w26793;
w27277 <= not w26789 and w27276;
w27278 <= not w26790 and not w26793;
w27279 <= not w27277 and not w27278;
w27280 <= not w26978 and not w27279;
w27281 <= not w26428 and not w26977;
w27282 <= not w26976 and w27281;
w27283 <= not w27280 and not w27282;
w27284 <= not b(28) and not w27283;
w27285 <= not w26447 and w26788;
w27286 <= not w26784 and w27285;
w27287 <= not w26785 and not w26788;
w27288 <= not w27286 and not w27287;
w27289 <= not w26978 and not w27288;
w27290 <= not w26437 and not w26977;
w27291 <= not w26976 and w27290;
w27292 <= not w27289 and not w27291;
w27293 <= not b(27) and not w27292;
w27294 <= not w26456 and w26783;
w27295 <= not w26779 and w27294;
w27296 <= not w26780 and not w26783;
w27297 <= not w27295 and not w27296;
w27298 <= not w26978 and not w27297;
w27299 <= not w26446 and not w26977;
w27300 <= not w26976 and w27299;
w27301 <= not w27298 and not w27300;
w27302 <= not b(26) and not w27301;
w27303 <= not w26465 and w26778;
w27304 <= not w26774 and w27303;
w27305 <= not w26775 and not w26778;
w27306 <= not w27304 and not w27305;
w27307 <= not w26978 and not w27306;
w27308 <= not w26455 and not w26977;
w27309 <= not w26976 and w27308;
w27310 <= not w27307 and not w27309;
w27311 <= not b(25) and not w27310;
w27312 <= not w26474 and w26773;
w27313 <= not w26769 and w27312;
w27314 <= not w26770 and not w26773;
w27315 <= not w27313 and not w27314;
w27316 <= not w26978 and not w27315;
w27317 <= not w26464 and not w26977;
w27318 <= not w26976 and w27317;
w27319 <= not w27316 and not w27318;
w27320 <= not b(24) and not w27319;
w27321 <= not w26483 and w26768;
w27322 <= not w26764 and w27321;
w27323 <= not w26765 and not w26768;
w27324 <= not w27322 and not w27323;
w27325 <= not w26978 and not w27324;
w27326 <= not w26473 and not w26977;
w27327 <= not w26976 and w27326;
w27328 <= not w27325 and not w27327;
w27329 <= not b(23) and not w27328;
w27330 <= not w26492 and w26763;
w27331 <= not w26759 and w27330;
w27332 <= not w26760 and not w26763;
w27333 <= not w27331 and not w27332;
w27334 <= not w26978 and not w27333;
w27335 <= not w26482 and not w26977;
w27336 <= not w26976 and w27335;
w27337 <= not w27334 and not w27336;
w27338 <= not b(22) and not w27337;
w27339 <= not w26501 and w26758;
w27340 <= not w26754 and w27339;
w27341 <= not w26755 and not w26758;
w27342 <= not w27340 and not w27341;
w27343 <= not w26978 and not w27342;
w27344 <= not w26491 and not w26977;
w27345 <= not w26976 and w27344;
w27346 <= not w27343 and not w27345;
w27347 <= not b(21) and not w27346;
w27348 <= not w26510 and w26753;
w27349 <= not w26749 and w27348;
w27350 <= not w26750 and not w26753;
w27351 <= not w27349 and not w27350;
w27352 <= not w26978 and not w27351;
w27353 <= not w26500 and not w26977;
w27354 <= not w26976 and w27353;
w27355 <= not w27352 and not w27354;
w27356 <= not b(20) and not w27355;
w27357 <= not w26519 and w26748;
w27358 <= not w26744 and w27357;
w27359 <= not w26745 and not w26748;
w27360 <= not w27358 and not w27359;
w27361 <= not w26978 and not w27360;
w27362 <= not w26509 and not w26977;
w27363 <= not w26976 and w27362;
w27364 <= not w27361 and not w27363;
w27365 <= not b(19) and not w27364;
w27366 <= not w26528 and w26743;
w27367 <= not w26739 and w27366;
w27368 <= not w26740 and not w26743;
w27369 <= not w27367 and not w27368;
w27370 <= not w26978 and not w27369;
w27371 <= not w26518 and not w26977;
w27372 <= not w26976 and w27371;
w27373 <= not w27370 and not w27372;
w27374 <= not b(18) and not w27373;
w27375 <= not w26537 and w26738;
w27376 <= not w26734 and w27375;
w27377 <= not w26735 and not w26738;
w27378 <= not w27376 and not w27377;
w27379 <= not w26978 and not w27378;
w27380 <= not w26527 and not w26977;
w27381 <= not w26976 and w27380;
w27382 <= not w27379 and not w27381;
w27383 <= not b(17) and not w27382;
w27384 <= not w26546 and w26733;
w27385 <= not w26729 and w27384;
w27386 <= not w26730 and not w26733;
w27387 <= not w27385 and not w27386;
w27388 <= not w26978 and not w27387;
w27389 <= not w26536 and not w26977;
w27390 <= not w26976 and w27389;
w27391 <= not w27388 and not w27390;
w27392 <= not b(16) and not w27391;
w27393 <= not w26555 and w26728;
w27394 <= not w26724 and w27393;
w27395 <= not w26725 and not w26728;
w27396 <= not w27394 and not w27395;
w27397 <= not w26978 and not w27396;
w27398 <= not w26545 and not w26977;
w27399 <= not w26976 and w27398;
w27400 <= not w27397 and not w27399;
w27401 <= not b(15) and not w27400;
w27402 <= not w26564 and w26723;
w27403 <= not w26719 and w27402;
w27404 <= not w26720 and not w26723;
w27405 <= not w27403 and not w27404;
w27406 <= not w26978 and not w27405;
w27407 <= not w26554 and not w26977;
w27408 <= not w26976 and w27407;
w27409 <= not w27406 and not w27408;
w27410 <= not b(14) and not w27409;
w27411 <= not w26573 and w26718;
w27412 <= not w26714 and w27411;
w27413 <= not w26715 and not w26718;
w27414 <= not w27412 and not w27413;
w27415 <= not w26978 and not w27414;
w27416 <= not w26563 and not w26977;
w27417 <= not w26976 and w27416;
w27418 <= not w27415 and not w27417;
w27419 <= not b(13) and not w27418;
w27420 <= not w26582 and w26713;
w27421 <= not w26709 and w27420;
w27422 <= not w26710 and not w26713;
w27423 <= not w27421 and not w27422;
w27424 <= not w26978 and not w27423;
w27425 <= not w26572 and not w26977;
w27426 <= not w26976 and w27425;
w27427 <= not w27424 and not w27426;
w27428 <= not b(12) and not w27427;
w27429 <= not w26591 and w26708;
w27430 <= not w26704 and w27429;
w27431 <= not w26705 and not w26708;
w27432 <= not w27430 and not w27431;
w27433 <= not w26978 and not w27432;
w27434 <= not w26581 and not w26977;
w27435 <= not w26976 and w27434;
w27436 <= not w27433 and not w27435;
w27437 <= not b(11) and not w27436;
w27438 <= not w26600 and w26703;
w27439 <= not w26699 and w27438;
w27440 <= not w26700 and not w26703;
w27441 <= not w27439 and not w27440;
w27442 <= not w26978 and not w27441;
w27443 <= not w26590 and not w26977;
w27444 <= not w26976 and w27443;
w27445 <= not w27442 and not w27444;
w27446 <= not b(10) and not w27445;
w27447 <= not w26609 and w26698;
w27448 <= not w26694 and w27447;
w27449 <= not w26695 and not w26698;
w27450 <= not w27448 and not w27449;
w27451 <= not w26978 and not w27450;
w27452 <= not w26599 and not w26977;
w27453 <= not w26976 and w27452;
w27454 <= not w27451 and not w27453;
w27455 <= not b(9) and not w27454;
w27456 <= not w26618 and w26693;
w27457 <= not w26689 and w27456;
w27458 <= not w26690 and not w26693;
w27459 <= not w27457 and not w27458;
w27460 <= not w26978 and not w27459;
w27461 <= not w26608 and not w26977;
w27462 <= not w26976 and w27461;
w27463 <= not w27460 and not w27462;
w27464 <= not b(8) and not w27463;
w27465 <= not w26627 and w26688;
w27466 <= not w26684 and w27465;
w27467 <= not w26685 and not w26688;
w27468 <= not w27466 and not w27467;
w27469 <= not w26978 and not w27468;
w27470 <= not w26617 and not w26977;
w27471 <= not w26976 and w27470;
w27472 <= not w27469 and not w27471;
w27473 <= not b(7) and not w27472;
w27474 <= not w26636 and w26683;
w27475 <= not w26679 and w27474;
w27476 <= not w26680 and not w26683;
w27477 <= not w27475 and not w27476;
w27478 <= not w26978 and not w27477;
w27479 <= not w26626 and not w26977;
w27480 <= not w26976 and w27479;
w27481 <= not w27478 and not w27480;
w27482 <= not b(6) and not w27481;
w27483 <= not w26645 and w26678;
w27484 <= not w26674 and w27483;
w27485 <= not w26675 and not w26678;
w27486 <= not w27484 and not w27485;
w27487 <= not w26978 and not w27486;
w27488 <= not w26635 and not w26977;
w27489 <= not w26976 and w27488;
w27490 <= not w27487 and not w27489;
w27491 <= not b(5) and not w27490;
w27492 <= not w26653 and w26673;
w27493 <= not w26669 and w27492;
w27494 <= not w26670 and not w26673;
w27495 <= not w27493 and not w27494;
w27496 <= not w26978 and not w27495;
w27497 <= not w26644 and not w26977;
w27498 <= not w26976 and w27497;
w27499 <= not w27496 and not w27498;
w27500 <= not b(4) and not w27499;
w27501 <= not w26664 and w26668;
w27502 <= not w26663 and w27501;
w27503 <= not w26665 and not w26668;
w27504 <= not w27502 and not w27503;
w27505 <= not w26978 and not w27504;
w27506 <= not w26652 and not w26977;
w27507 <= not w26976 and w27506;
w27508 <= not w27505 and not w27507;
w27509 <= not b(3) and not w27508;
w27510 <= not w26660 and w26662;
w27511 <= not w26658 and w27510;
w27512 <= not w26663 and not w27511;
w27513 <= not w26978 and w27512;
w27514 <= not w26657 and not w26977;
w27515 <= not w26976 and w27514;
w27516 <= not w27513 and not w27515;
w27517 <= not b(2) and not w27516;
w27518 <= b(0) and not w26978;
w27519 <= a(2) and not w27518;
w27520 <= w26662 and not w26978;
w27521 <= not w27519 and not w27520;
w27522 <= b(1) and not w27521;
w27523 <= not b(1) and not w27520;
w27524 <= not w27519 and w27523;
w27525 <= not w27522 and not w27524;
w27526 <= not a(1) and b(0);
w27527 <= not w27525 and not w27526;
w27528 <= not b(1) and not w27521;
w27529 <= not w27527 and not w27528;
w27530 <= b(2) and not w27515;
w27531 <= not w27513 and w27530;
w27532 <= not w27517 and not w27531;
w27533 <= not w27529 and w27532;
w27534 <= not w27517 and not w27533;
w27535 <= b(3) and not w27507;
w27536 <= not w27505 and w27535;
w27537 <= not w27509 and not w27536;
w27538 <= not w27534 and w27537;
w27539 <= not w27509 and not w27538;
w27540 <= b(4) and not w27498;
w27541 <= not w27496 and w27540;
w27542 <= not w27500 and not w27541;
w27543 <= not w27539 and w27542;
w27544 <= not w27500 and not w27543;
w27545 <= b(5) and not w27489;
w27546 <= not w27487 and w27545;
w27547 <= not w27491 and not w27546;
w27548 <= not w27544 and w27547;
w27549 <= not w27491 and not w27548;
w27550 <= b(6) and not w27480;
w27551 <= not w27478 and w27550;
w27552 <= not w27482 and not w27551;
w27553 <= not w27549 and w27552;
w27554 <= not w27482 and not w27553;
w27555 <= b(7) and not w27471;
w27556 <= not w27469 and w27555;
w27557 <= not w27473 and not w27556;
w27558 <= not w27554 and w27557;
w27559 <= not w27473 and not w27558;
w27560 <= b(8) and not w27462;
w27561 <= not w27460 and w27560;
w27562 <= not w27464 and not w27561;
w27563 <= not w27559 and w27562;
w27564 <= not w27464 and not w27563;
w27565 <= b(9) and not w27453;
w27566 <= not w27451 and w27565;
w27567 <= not w27455 and not w27566;
w27568 <= not w27564 and w27567;
w27569 <= not w27455 and not w27568;
w27570 <= b(10) and not w27444;
w27571 <= not w27442 and w27570;
w27572 <= not w27446 and not w27571;
w27573 <= not w27569 and w27572;
w27574 <= not w27446 and not w27573;
w27575 <= b(11) and not w27435;
w27576 <= not w27433 and w27575;
w27577 <= not w27437 and not w27576;
w27578 <= not w27574 and w27577;
w27579 <= not w27437 and not w27578;
w27580 <= b(12) and not w27426;
w27581 <= not w27424 and w27580;
w27582 <= not w27428 and not w27581;
w27583 <= not w27579 and w27582;
w27584 <= not w27428 and not w27583;
w27585 <= b(13) and not w27417;
w27586 <= not w27415 and w27585;
w27587 <= not w27419 and not w27586;
w27588 <= not w27584 and w27587;
w27589 <= not w27419 and not w27588;
w27590 <= b(14) and not w27408;
w27591 <= not w27406 and w27590;
w27592 <= not w27410 and not w27591;
w27593 <= not w27589 and w27592;
w27594 <= not w27410 and not w27593;
w27595 <= b(15) and not w27399;
w27596 <= not w27397 and w27595;
w27597 <= not w27401 and not w27596;
w27598 <= not w27594 and w27597;
w27599 <= not w27401 and not w27598;
w27600 <= b(16) and not w27390;
w27601 <= not w27388 and w27600;
w27602 <= not w27392 and not w27601;
w27603 <= not w27599 and w27602;
w27604 <= not w27392 and not w27603;
w27605 <= b(17) and not w27381;
w27606 <= not w27379 and w27605;
w27607 <= not w27383 and not w27606;
w27608 <= not w27604 and w27607;
w27609 <= not w27383 and not w27608;
w27610 <= b(18) and not w27372;
w27611 <= not w27370 and w27610;
w27612 <= not w27374 and not w27611;
w27613 <= not w27609 and w27612;
w27614 <= not w27374 and not w27613;
w27615 <= b(19) and not w27363;
w27616 <= not w27361 and w27615;
w27617 <= not w27365 and not w27616;
w27618 <= not w27614 and w27617;
w27619 <= not w27365 and not w27618;
w27620 <= b(20) and not w27354;
w27621 <= not w27352 and w27620;
w27622 <= not w27356 and not w27621;
w27623 <= not w27619 and w27622;
w27624 <= not w27356 and not w27623;
w27625 <= b(21) and not w27345;
w27626 <= not w27343 and w27625;
w27627 <= not w27347 and not w27626;
w27628 <= not w27624 and w27627;
w27629 <= not w27347 and not w27628;
w27630 <= b(22) and not w27336;
w27631 <= not w27334 and w27630;
w27632 <= not w27338 and not w27631;
w27633 <= not w27629 and w27632;
w27634 <= not w27338 and not w27633;
w27635 <= b(23) and not w27327;
w27636 <= not w27325 and w27635;
w27637 <= not w27329 and not w27636;
w27638 <= not w27634 and w27637;
w27639 <= not w27329 and not w27638;
w27640 <= b(24) and not w27318;
w27641 <= not w27316 and w27640;
w27642 <= not w27320 and not w27641;
w27643 <= not w27639 and w27642;
w27644 <= not w27320 and not w27643;
w27645 <= b(25) and not w27309;
w27646 <= not w27307 and w27645;
w27647 <= not w27311 and not w27646;
w27648 <= not w27644 and w27647;
w27649 <= not w27311 and not w27648;
w27650 <= b(26) and not w27300;
w27651 <= not w27298 and w27650;
w27652 <= not w27302 and not w27651;
w27653 <= not w27649 and w27652;
w27654 <= not w27302 and not w27653;
w27655 <= b(27) and not w27291;
w27656 <= not w27289 and w27655;
w27657 <= not w27293 and not w27656;
w27658 <= not w27654 and w27657;
w27659 <= not w27293 and not w27658;
w27660 <= b(28) and not w27282;
w27661 <= not w27280 and w27660;
w27662 <= not w27284 and not w27661;
w27663 <= not w27659 and w27662;
w27664 <= not w27284 and not w27663;
w27665 <= b(29) and not w27273;
w27666 <= not w27271 and w27665;
w27667 <= not w27275 and not w27666;
w27668 <= not w27664 and w27667;
w27669 <= not w27275 and not w27668;
w27670 <= b(30) and not w27264;
w27671 <= not w27262 and w27670;
w27672 <= not w27266 and not w27671;
w27673 <= not w27669 and w27672;
w27674 <= not w27266 and not w27673;
w27675 <= b(31) and not w27255;
w27676 <= not w27253 and w27675;
w27677 <= not w27257 and not w27676;
w27678 <= not w27674 and w27677;
w27679 <= not w27257 and not w27678;
w27680 <= b(32) and not w27246;
w27681 <= not w27244 and w27680;
w27682 <= not w27248 and not w27681;
w27683 <= not w27679 and w27682;
w27684 <= not w27248 and not w27683;
w27685 <= b(33) and not w27237;
w27686 <= not w27235 and w27685;
w27687 <= not w27239 and not w27686;
w27688 <= not w27684 and w27687;
w27689 <= not w27239 and not w27688;
w27690 <= b(34) and not w27228;
w27691 <= not w27226 and w27690;
w27692 <= not w27230 and not w27691;
w27693 <= not w27689 and w27692;
w27694 <= not w27230 and not w27693;
w27695 <= b(35) and not w27219;
w27696 <= not w27217 and w27695;
w27697 <= not w27221 and not w27696;
w27698 <= not w27694 and w27697;
w27699 <= not w27221 and not w27698;
w27700 <= b(36) and not w27210;
w27701 <= not w27208 and w27700;
w27702 <= not w27212 and not w27701;
w27703 <= not w27699 and w27702;
w27704 <= not w27212 and not w27703;
w27705 <= b(37) and not w27201;
w27706 <= not w27199 and w27705;
w27707 <= not w27203 and not w27706;
w27708 <= not w27704 and w27707;
w27709 <= not w27203 and not w27708;
w27710 <= b(38) and not w27192;
w27711 <= not w27190 and w27710;
w27712 <= not w27194 and not w27711;
w27713 <= not w27709 and w27712;
w27714 <= not w27194 and not w27713;
w27715 <= b(39) and not w27183;
w27716 <= not w27181 and w27715;
w27717 <= not w27185 and not w27716;
w27718 <= not w27714 and w27717;
w27719 <= not w27185 and not w27718;
w27720 <= b(40) and not w27174;
w27721 <= not w27172 and w27720;
w27722 <= not w27176 and not w27721;
w27723 <= not w27719 and w27722;
w27724 <= not w27176 and not w27723;
w27725 <= b(41) and not w27165;
w27726 <= not w27163 and w27725;
w27727 <= not w27167 and not w27726;
w27728 <= not w27724 and w27727;
w27729 <= not w27167 and not w27728;
w27730 <= b(42) and not w27156;
w27731 <= not w27154 and w27730;
w27732 <= not w27158 and not w27731;
w27733 <= not w27729 and w27732;
w27734 <= not w27158 and not w27733;
w27735 <= b(43) and not w27147;
w27736 <= not w27145 and w27735;
w27737 <= not w27149 and not w27736;
w27738 <= not w27734 and w27737;
w27739 <= not w27149 and not w27738;
w27740 <= b(44) and not w27138;
w27741 <= not w27136 and w27740;
w27742 <= not w27140 and not w27741;
w27743 <= not w27739 and w27742;
w27744 <= not w27140 and not w27743;
w27745 <= b(45) and not w27129;
w27746 <= not w27127 and w27745;
w27747 <= not w27131 and not w27746;
w27748 <= not w27744 and w27747;
w27749 <= not w27131 and not w27748;
w27750 <= b(46) and not w27120;
w27751 <= not w27118 and w27750;
w27752 <= not w27122 and not w27751;
w27753 <= not w27749 and w27752;
w27754 <= not w27122 and not w27753;
w27755 <= b(47) and not w27111;
w27756 <= not w27109 and w27755;
w27757 <= not w27113 and not w27756;
w27758 <= not w27754 and w27757;
w27759 <= not w27113 and not w27758;
w27760 <= b(48) and not w27102;
w27761 <= not w27100 and w27760;
w27762 <= not w27104 and not w27761;
w27763 <= not w27759 and w27762;
w27764 <= not w27104 and not w27763;
w27765 <= b(49) and not w27093;
w27766 <= not w27091 and w27765;
w27767 <= not w27095 and not w27766;
w27768 <= not w27764 and w27767;
w27769 <= not w27095 and not w27768;
w27770 <= b(50) and not w27084;
w27771 <= not w27082 and w27770;
w27772 <= not w27086 and not w27771;
w27773 <= not w27769 and w27772;
w27774 <= not w27086 and not w27773;
w27775 <= b(51) and not w27075;
w27776 <= not w27073 and w27775;
w27777 <= not w27077 and not w27776;
w27778 <= not w27774 and w27777;
w27779 <= not w27077 and not w27778;
w27780 <= b(52) and not w27066;
w27781 <= not w27064 and w27780;
w27782 <= not w27068 and not w27781;
w27783 <= not w27779 and w27782;
w27784 <= not w27068 and not w27783;
w27785 <= b(53) and not w27057;
w27786 <= not w27055 and w27785;
w27787 <= not w27059 and not w27786;
w27788 <= not w27784 and w27787;
w27789 <= not w27059 and not w27788;
w27790 <= b(54) and not w27048;
w27791 <= not w27046 and w27790;
w27792 <= not w27050 and not w27791;
w27793 <= not w27789 and w27792;
w27794 <= not w27050 and not w27793;
w27795 <= b(55) and not w27039;
w27796 <= not w27037 and w27795;
w27797 <= not w27041 and not w27796;
w27798 <= not w27794 and w27797;
w27799 <= not w27041 and not w27798;
w27800 <= b(56) and not w27030;
w27801 <= not w27028 and w27800;
w27802 <= not w27032 and not w27801;
w27803 <= not w27799 and w27802;
w27804 <= not w27032 and not w27803;
w27805 <= b(57) and not w27021;
w27806 <= not w27019 and w27805;
w27807 <= not w27023 and not w27806;
w27808 <= not w27804 and w27807;
w27809 <= not w27023 and not w27808;
w27810 <= b(58) and not w27012;
w27811 <= not w27010 and w27810;
w27812 <= not w27014 and not w27811;
w27813 <= not w27809 and w27812;
w27814 <= not w27014 and not w27813;
w27815 <= b(59) and not w27003;
w27816 <= not w27001 and w27815;
w27817 <= not w27005 and not w27816;
w27818 <= not w27814 and w27817;
w27819 <= not w27005 and not w27818;
w27820 <= b(60) and not w26994;
w27821 <= not w26992 and w27820;
w27822 <= not w26996 and not w27821;
w27823 <= not w27819 and w27822;
w27824 <= not w26996 and not w27823;
w27825 <= b(61) and not w26985;
w27826 <= not w26983 and w27825;
w27827 <= not w26987 and not w27826;
w27828 <= not w27824 and w27827;
w27829 <= not w26987 and not w27828;
w27830 <= not w26132 and not w26973;
w27831 <= not w26971 and w27830;
w27832 <= not w26959 and w27831;
w27833 <= not w26971 and not w26973;
w27834 <= not w26960 and not w27833;
w27835 <= not w27832 and not w27834;
w27836 <= not w26978 and not w27835;
w27837 <= not w26970 and not w26977;
w27838 <= not w26976 and w27837;
w27839 <= not w27836 and not w27838;
w27840 <= not b(62) and not w27839;
w27841 <= b(62) and not w27838;
w27842 <= not w27836 and w27841;
w27843 <= not b(63) and not w27842;
w27844 <= not w27840 and w27843;
w27845 <= not w27829 and w27844;
w27846 <= w22 and not w27839;
w27847 <= not w27845 and not w27846;
w27848 <= not w27005 and w27822;
w27849 <= not w27818 and w27848;
w27850 <= not w27819 and not w27822;
w27851 <= not w27849 and not w27850;
w27852 <= not w27847 and not w27851;
w27853 <= not w26995 and not w27846;
w27854 <= not w27845 and w27853;
w27855 <= not w27852 and not w27854;
w27856 <= not w27023 and w27812;
w27857 <= not w27808 and w27856;
w27858 <= not w27809 and not w27812;
w27859 <= not w27857 and not w27858;
w27860 <= not w27847 and not w27859;
w27861 <= not w27013 and not w27846;
w27862 <= not w27845 and w27861;
w27863 <= not w27860 and not w27862;
w27864 <= not w27041 and w27802;
w27865 <= not w27798 and w27864;
w27866 <= not w27799 and not w27802;
w27867 <= not w27865 and not w27866;
w27868 <= not w27847 and not w27867;
w27869 <= not w27031 and not w27846;
w27870 <= not w27845 and w27869;
w27871 <= not w27868 and not w27870;
w27872 <= not w27059 and w27792;
w27873 <= not w27788 and w27872;
w27874 <= not w27789 and not w27792;
w27875 <= not w27873 and not w27874;
w27876 <= not w27847 and not w27875;
w27877 <= not w27049 and not w27846;
w27878 <= not w27845 and w27877;
w27879 <= not w27876 and not w27878;
w27880 <= not w27077 and w27782;
w27881 <= not w27778 and w27880;
w27882 <= not w27779 and not w27782;
w27883 <= not w27881 and not w27882;
w27884 <= not w27847 and not w27883;
w27885 <= not w27067 and not w27846;
w27886 <= not w27845 and w27885;
w27887 <= not w27884 and not w27886;
w27888 <= not w27095 and w27772;
w27889 <= not w27768 and w27888;
w27890 <= not w27769 and not w27772;
w27891 <= not w27889 and not w27890;
w27892 <= not w27847 and not w27891;
w27893 <= not w27085 and not w27846;
w27894 <= not w27845 and w27893;
w27895 <= not w27892 and not w27894;
w27896 <= not w27113 and w27762;
w27897 <= not w27758 and w27896;
w27898 <= not w27759 and not w27762;
w27899 <= not w27897 and not w27898;
w27900 <= not w27847 and not w27899;
w27901 <= not w27103 and not w27846;
w27902 <= not w27845 and w27901;
w27903 <= not w27900 and not w27902;
w27904 <= not w27131 and w27752;
w27905 <= not w27748 and w27904;
w27906 <= not w27749 and not w27752;
w27907 <= not w27905 and not w27906;
w27908 <= not w27847 and not w27907;
w27909 <= not w27121 and not w27846;
w27910 <= not w27845 and w27909;
w27911 <= not w27908 and not w27910;
w27912 <= not w27149 and w27742;
w27913 <= not w27738 and w27912;
w27914 <= not w27739 and not w27742;
w27915 <= not w27913 and not w27914;
w27916 <= not w27847 and not w27915;
w27917 <= not w27139 and not w27846;
w27918 <= not w27845 and w27917;
w27919 <= not w27916 and not w27918;
w27920 <= not w27167 and w27732;
w27921 <= not w27728 and w27920;
w27922 <= not w27729 and not w27732;
w27923 <= not w27921 and not w27922;
w27924 <= not w27847 and not w27923;
w27925 <= not w27157 and not w27846;
w27926 <= not w27845 and w27925;
w27927 <= not w27924 and not w27926;
w27928 <= not w27185 and w27722;
w27929 <= not w27718 and w27928;
w27930 <= not w27719 and not w27722;
w27931 <= not w27929 and not w27930;
w27932 <= not w27847 and not w27931;
w27933 <= not w27175 and not w27846;
w27934 <= not w27845 and w27933;
w27935 <= not w27932 and not w27934;
w27936 <= not w27203 and w27712;
w27937 <= not w27708 and w27936;
w27938 <= not w27709 and not w27712;
w27939 <= not w27937 and not w27938;
w27940 <= not w27847 and not w27939;
w27941 <= not w27193 and not w27846;
w27942 <= not w27845 and w27941;
w27943 <= not w27940 and not w27942;
w27944 <= not w27221 and w27702;
w27945 <= not w27698 and w27944;
w27946 <= not w27699 and not w27702;
w27947 <= not w27945 and not w27946;
w27948 <= not w27847 and not w27947;
w27949 <= not w27211 and not w27846;
w27950 <= not w27845 and w27949;
w27951 <= not w27948 and not w27950;
w27952 <= not w27239 and w27692;
w27953 <= not w27688 and w27952;
w27954 <= not w27689 and not w27692;
w27955 <= not w27953 and not w27954;
w27956 <= not w27847 and not w27955;
w27957 <= not w27229 and not w27846;
w27958 <= not w27845 and w27957;
w27959 <= not w27956 and not w27958;
w27960 <= not w27257 and w27682;
w27961 <= not w27678 and w27960;
w27962 <= not w27679 and not w27682;
w27963 <= not w27961 and not w27962;
w27964 <= not w27847 and not w27963;
w27965 <= not w27247 and not w27846;
w27966 <= not w27845 and w27965;
w27967 <= not w27964 and not w27966;
w27968 <= not w27275 and w27672;
w27969 <= not w27668 and w27968;
w27970 <= not w27669 and not w27672;
w27971 <= not w27969 and not w27970;
w27972 <= not w27847 and not w27971;
w27973 <= not w27265 and not w27846;
w27974 <= not w27845 and w27973;
w27975 <= not w27972 and not w27974;
w27976 <= not w27293 and w27662;
w27977 <= not w27658 and w27976;
w27978 <= not w27659 and not w27662;
w27979 <= not w27977 and not w27978;
w27980 <= not w27847 and not w27979;
w27981 <= not w27283 and not w27846;
w27982 <= not w27845 and w27981;
w27983 <= not w27980 and not w27982;
w27984 <= not w27311 and w27652;
w27985 <= not w27648 and w27984;
w27986 <= not w27649 and not w27652;
w27987 <= not w27985 and not w27986;
w27988 <= not w27847 and not w27987;
w27989 <= not w27301 and not w27846;
w27990 <= not w27845 and w27989;
w27991 <= not w27988 and not w27990;
w27992 <= not w27329 and w27642;
w27993 <= not w27638 and w27992;
w27994 <= not w27639 and not w27642;
w27995 <= not w27993 and not w27994;
w27996 <= not w27847 and not w27995;
w27997 <= not w27319 and not w27846;
w27998 <= not w27845 and w27997;
w27999 <= not w27996 and not w27998;
w28000 <= not w27347 and w27632;
w28001 <= not w27628 and w28000;
w28002 <= not w27629 and not w27632;
w28003 <= not w28001 and not w28002;
w28004 <= not w27847 and not w28003;
w28005 <= not w27337 and not w27846;
w28006 <= not w27845 and w28005;
w28007 <= not w28004 and not w28006;
w28008 <= not w27365 and w27622;
w28009 <= not w27618 and w28008;
w28010 <= not w27619 and not w27622;
w28011 <= not w28009 and not w28010;
w28012 <= not w27847 and not w28011;
w28013 <= not w27355 and not w27846;
w28014 <= not w27845 and w28013;
w28015 <= not w28012 and not w28014;
w28016 <= not w27383 and w27612;
w28017 <= not w27608 and w28016;
w28018 <= not w27609 and not w27612;
w28019 <= not w28017 and not w28018;
w28020 <= not w27847 and not w28019;
w28021 <= not w27373 and not w27846;
w28022 <= not w27845 and w28021;
w28023 <= not w28020 and not w28022;
w28024 <= not w27401 and w27602;
w28025 <= not w27598 and w28024;
w28026 <= not w27599 and not w27602;
w28027 <= not w28025 and not w28026;
w28028 <= not w27847 and not w28027;
w28029 <= not w27391 and not w27846;
w28030 <= not w27845 and w28029;
w28031 <= not w28028 and not w28030;
w28032 <= not w27419 and w27592;
w28033 <= not w27588 and w28032;
w28034 <= not w27589 and not w27592;
w28035 <= not w28033 and not w28034;
w28036 <= not w27847 and not w28035;
w28037 <= not w27409 and not w27846;
w28038 <= not w27845 and w28037;
w28039 <= not w28036 and not w28038;
w28040 <= not w27437 and w27582;
w28041 <= not w27578 and w28040;
w28042 <= not w27579 and not w27582;
w28043 <= not w28041 and not w28042;
w28044 <= not w27847 and not w28043;
w28045 <= not w27427 and not w27846;
w28046 <= not w27845 and w28045;
w28047 <= not w28044 and not w28046;
w28048 <= not w27455 and w27572;
w28049 <= not w27568 and w28048;
w28050 <= not w27569 and not w27572;
w28051 <= not w28049 and not w28050;
w28052 <= not w27847 and not w28051;
w28053 <= not w27445 and not w27846;
w28054 <= not w27845 and w28053;
w28055 <= not w28052 and not w28054;
w28056 <= not w27473 and w27562;
w28057 <= not w27558 and w28056;
w28058 <= not w27559 and not w27562;
w28059 <= not w28057 and not w28058;
w28060 <= not w27847 and not w28059;
w28061 <= not w27463 and not w27846;
w28062 <= not w27845 and w28061;
w28063 <= not w28060 and not w28062;
w28064 <= not w27491 and w27552;
w28065 <= not w27548 and w28064;
w28066 <= not w27549 and not w27552;
w28067 <= not w28065 and not w28066;
w28068 <= not w27847 and not w28067;
w28069 <= not w27481 and not w27846;
w28070 <= not w27845 and w28069;
w28071 <= not w28068 and not w28070;
w28072 <= not w27509 and w27542;
w28073 <= not w27538 and w28072;
w28074 <= not w27539 and not w27542;
w28075 <= not w28073 and not w28074;
w28076 <= not w27847 and not w28075;
w28077 <= not w27499 and not w27846;
w28078 <= not w27845 and w28077;
w28079 <= not w28076 and not w28078;
w28080 <= not w27528 and w27532;
w28081 <= not w27527 and w28080;
w28082 <= not w27529 and not w27532;
w28083 <= not w28081 and not w28082;
w28084 <= not w27847 and not w28083;
w28085 <= not w27516 and not w27846;
w28086 <= not w27845 and w28085;
w28087 <= not w28084 and not w28086;
w28088 <= not a(0) and b(0);
w28089 <= b(0) and not w27847;
w28090 <= a(1) and not w28089;
w28091 <= w27526 and not w27847;
w28092 <= not w28090 and not w28091;
w28093 <= not w28088 and not w28092;
w28094 <= w28088 and not w28091;
w28095 <= not w28090 and w28094;
w28096 <= not b(1) and not w28095;
w28097 <= not w27524 and w27526;
w28098 <= not w27522 and w28097;
w28099 <= not w27527 and not w28098;
w28100 <= not w27847 and w28099;
w28101 <= not w27521 and not w27846;
w28102 <= not w27845 and w28101;
w28103 <= not w28100 and not w28102;
w28104 <= not w28096 and w28103;
w28105 <= not w28093 and w28104;
w28106 <= not b(2) and not w28105;
w28107 <= not w28093 and not w28096;
w28108 <= not w28103 and not w28107;
w28109 <= not w28106 and not w28108;
w28110 <= not w28087 and not w28109;
w28111 <= w28087 and not w28108;
w28112 <= not w28106 and w28111;
w28113 <= not b(3) and not w28112;
w28114 <= not w27517 and w27537;
w28115 <= not w27533 and w28114;
w28116 <= not w27534 and not w27537;
w28117 <= not w28115 and not w28116;
w28118 <= not w27847 and not w28117;
w28119 <= not w27508 and not w27846;
w28120 <= not w27845 and w28119;
w28121 <= not w28118 and not w28120;
w28122 <= not w28113 and w28121;
w28123 <= not w28110 and w28122;
w28124 <= not b(4) and not w28123;
w28125 <= not w28110 and not w28113;
w28126 <= not w28121 and not w28125;
w28127 <= not w28124 and not w28126;
w28128 <= not w28079 and not w28127;
w28129 <= w28079 and not w28126;
w28130 <= not w28124 and w28129;
w28131 <= not b(5) and not w28130;
w28132 <= not w27500 and w27547;
w28133 <= not w27543 and w28132;
w28134 <= not w27544 and not w27547;
w28135 <= not w28133 and not w28134;
w28136 <= not w27847 and not w28135;
w28137 <= not w27490 and not w27846;
w28138 <= not w27845 and w28137;
w28139 <= not w28136 and not w28138;
w28140 <= not w28131 and w28139;
w28141 <= not w28128 and w28140;
w28142 <= not b(6) and not w28141;
w28143 <= not w28128 and not w28131;
w28144 <= not w28139 and not w28143;
w28145 <= not w28142 and not w28144;
w28146 <= not w28071 and not w28145;
w28147 <= w28071 and not w28144;
w28148 <= not w28142 and w28147;
w28149 <= not b(7) and not w28148;
w28150 <= not w27482 and w27557;
w28151 <= not w27553 and w28150;
w28152 <= not w27554 and not w27557;
w28153 <= not w28151 and not w28152;
w28154 <= not w27847 and not w28153;
w28155 <= not w27472 and not w27846;
w28156 <= not w27845 and w28155;
w28157 <= not w28154 and not w28156;
w28158 <= not w28149 and w28157;
w28159 <= not w28146 and w28158;
w28160 <= not b(8) and not w28159;
w28161 <= not w28146 and not w28149;
w28162 <= not w28157 and not w28161;
w28163 <= not w28160 and not w28162;
w28164 <= not w28063 and not w28163;
w28165 <= w28063 and not w28162;
w28166 <= not w28160 and w28165;
w28167 <= not b(9) and not w28166;
w28168 <= not w27464 and w27567;
w28169 <= not w27563 and w28168;
w28170 <= not w27564 and not w27567;
w28171 <= not w28169 and not w28170;
w28172 <= not w27847 and not w28171;
w28173 <= not w27454 and not w27846;
w28174 <= not w27845 and w28173;
w28175 <= not w28172 and not w28174;
w28176 <= not w28167 and w28175;
w28177 <= not w28164 and w28176;
w28178 <= not b(10) and not w28177;
w28179 <= not w28164 and not w28167;
w28180 <= not w28175 and not w28179;
w28181 <= not w28178 and not w28180;
w28182 <= not w28055 and not w28181;
w28183 <= w28055 and not w28180;
w28184 <= not w28178 and w28183;
w28185 <= not b(11) and not w28184;
w28186 <= not w27446 and w27577;
w28187 <= not w27573 and w28186;
w28188 <= not w27574 and not w27577;
w28189 <= not w28187 and not w28188;
w28190 <= not w27847 and not w28189;
w28191 <= not w27436 and not w27846;
w28192 <= not w27845 and w28191;
w28193 <= not w28190 and not w28192;
w28194 <= not w28185 and w28193;
w28195 <= not w28182 and w28194;
w28196 <= not b(12) and not w28195;
w28197 <= not w28182 and not w28185;
w28198 <= not w28193 and not w28197;
w28199 <= not w28196 and not w28198;
w28200 <= not w28047 and not w28199;
w28201 <= w28047 and not w28198;
w28202 <= not w28196 and w28201;
w28203 <= not b(13) and not w28202;
w28204 <= not w27428 and w27587;
w28205 <= not w27583 and w28204;
w28206 <= not w27584 and not w27587;
w28207 <= not w28205 and not w28206;
w28208 <= not w27847 and not w28207;
w28209 <= not w27418 and not w27846;
w28210 <= not w27845 and w28209;
w28211 <= not w28208 and not w28210;
w28212 <= not w28203 and w28211;
w28213 <= not w28200 and w28212;
w28214 <= not b(14) and not w28213;
w28215 <= not w28200 and not w28203;
w28216 <= not w28211 and not w28215;
w28217 <= not w28214 and not w28216;
w28218 <= not w28039 and not w28217;
w28219 <= w28039 and not w28216;
w28220 <= not w28214 and w28219;
w28221 <= not b(15) and not w28220;
w28222 <= not w27410 and w27597;
w28223 <= not w27593 and w28222;
w28224 <= not w27594 and not w27597;
w28225 <= not w28223 and not w28224;
w28226 <= not w27847 and not w28225;
w28227 <= not w27400 and not w27846;
w28228 <= not w27845 and w28227;
w28229 <= not w28226 and not w28228;
w28230 <= not w28221 and w28229;
w28231 <= not w28218 and w28230;
w28232 <= not b(16) and not w28231;
w28233 <= not w28218 and not w28221;
w28234 <= not w28229 and not w28233;
w28235 <= not w28232 and not w28234;
w28236 <= not w28031 and not w28235;
w28237 <= w28031 and not w28234;
w28238 <= not w28232 and w28237;
w28239 <= not b(17) and not w28238;
w28240 <= not w27392 and w27607;
w28241 <= not w27603 and w28240;
w28242 <= not w27604 and not w27607;
w28243 <= not w28241 and not w28242;
w28244 <= not w27847 and not w28243;
w28245 <= not w27382 and not w27846;
w28246 <= not w27845 and w28245;
w28247 <= not w28244 and not w28246;
w28248 <= not w28239 and w28247;
w28249 <= not w28236 and w28248;
w28250 <= not b(18) and not w28249;
w28251 <= not w28236 and not w28239;
w28252 <= not w28247 and not w28251;
w28253 <= not w28250 and not w28252;
w28254 <= not w28023 and not w28253;
w28255 <= w28023 and not w28252;
w28256 <= not w28250 and w28255;
w28257 <= not b(19) and not w28256;
w28258 <= not w27374 and w27617;
w28259 <= not w27613 and w28258;
w28260 <= not w27614 and not w27617;
w28261 <= not w28259 and not w28260;
w28262 <= not w27847 and not w28261;
w28263 <= not w27364 and not w27846;
w28264 <= not w27845 and w28263;
w28265 <= not w28262 and not w28264;
w28266 <= not w28257 and w28265;
w28267 <= not w28254 and w28266;
w28268 <= not b(20) and not w28267;
w28269 <= not w28254 and not w28257;
w28270 <= not w28265 and not w28269;
w28271 <= not w28268 and not w28270;
w28272 <= not w28015 and not w28271;
w28273 <= w28015 and not w28270;
w28274 <= not w28268 and w28273;
w28275 <= not b(21) and not w28274;
w28276 <= not w27356 and w27627;
w28277 <= not w27623 and w28276;
w28278 <= not w27624 and not w27627;
w28279 <= not w28277 and not w28278;
w28280 <= not w27847 and not w28279;
w28281 <= not w27346 and not w27846;
w28282 <= not w27845 and w28281;
w28283 <= not w28280 and not w28282;
w28284 <= not w28275 and w28283;
w28285 <= not w28272 and w28284;
w28286 <= not b(22) and not w28285;
w28287 <= not w28272 and not w28275;
w28288 <= not w28283 and not w28287;
w28289 <= not w28286 and not w28288;
w28290 <= not w28007 and not w28289;
w28291 <= w28007 and not w28288;
w28292 <= not w28286 and w28291;
w28293 <= not b(23) and not w28292;
w28294 <= not w27338 and w27637;
w28295 <= not w27633 and w28294;
w28296 <= not w27634 and not w27637;
w28297 <= not w28295 and not w28296;
w28298 <= not w27847 and not w28297;
w28299 <= not w27328 and not w27846;
w28300 <= not w27845 and w28299;
w28301 <= not w28298 and not w28300;
w28302 <= not w28293 and w28301;
w28303 <= not w28290 and w28302;
w28304 <= not b(24) and not w28303;
w28305 <= not w28290 and not w28293;
w28306 <= not w28301 and not w28305;
w28307 <= not w28304 and not w28306;
w28308 <= not w27999 and not w28307;
w28309 <= w27999 and not w28306;
w28310 <= not w28304 and w28309;
w28311 <= not b(25) and not w28310;
w28312 <= not w27320 and w27647;
w28313 <= not w27643 and w28312;
w28314 <= not w27644 and not w27647;
w28315 <= not w28313 and not w28314;
w28316 <= not w27847 and not w28315;
w28317 <= not w27310 and not w27846;
w28318 <= not w27845 and w28317;
w28319 <= not w28316 and not w28318;
w28320 <= not w28311 and w28319;
w28321 <= not w28308 and w28320;
w28322 <= not b(26) and not w28321;
w28323 <= not w28308 and not w28311;
w28324 <= not w28319 and not w28323;
w28325 <= not w28322 and not w28324;
w28326 <= not w27991 and not w28325;
w28327 <= w27991 and not w28324;
w28328 <= not w28322 and w28327;
w28329 <= not b(27) and not w28328;
w28330 <= not w27302 and w27657;
w28331 <= not w27653 and w28330;
w28332 <= not w27654 and not w27657;
w28333 <= not w28331 and not w28332;
w28334 <= not w27847 and not w28333;
w28335 <= not w27292 and not w27846;
w28336 <= not w27845 and w28335;
w28337 <= not w28334 and not w28336;
w28338 <= not w28329 and w28337;
w28339 <= not w28326 and w28338;
w28340 <= not b(28) and not w28339;
w28341 <= not w28326 and not w28329;
w28342 <= not w28337 and not w28341;
w28343 <= not w28340 and not w28342;
w28344 <= not w27983 and not w28343;
w28345 <= w27983 and not w28342;
w28346 <= not w28340 and w28345;
w28347 <= not b(29) and not w28346;
w28348 <= not w27284 and w27667;
w28349 <= not w27663 and w28348;
w28350 <= not w27664 and not w27667;
w28351 <= not w28349 and not w28350;
w28352 <= not w27847 and not w28351;
w28353 <= not w27274 and not w27846;
w28354 <= not w27845 and w28353;
w28355 <= not w28352 and not w28354;
w28356 <= not w28347 and w28355;
w28357 <= not w28344 and w28356;
w28358 <= not b(30) and not w28357;
w28359 <= not w28344 and not w28347;
w28360 <= not w28355 and not w28359;
w28361 <= not w28358 and not w28360;
w28362 <= not w27975 and not w28361;
w28363 <= w27975 and not w28360;
w28364 <= not w28358 and w28363;
w28365 <= not b(31) and not w28364;
w28366 <= not w27266 and w27677;
w28367 <= not w27673 and w28366;
w28368 <= not w27674 and not w27677;
w28369 <= not w28367 and not w28368;
w28370 <= not w27847 and not w28369;
w28371 <= not w27256 and not w27846;
w28372 <= not w27845 and w28371;
w28373 <= not w28370 and not w28372;
w28374 <= not w28365 and w28373;
w28375 <= not w28362 and w28374;
w28376 <= not b(32) and not w28375;
w28377 <= not w28362 and not w28365;
w28378 <= not w28373 and not w28377;
w28379 <= not w28376 and not w28378;
w28380 <= not w27967 and not w28379;
w28381 <= w27967 and not w28378;
w28382 <= not w28376 and w28381;
w28383 <= not b(33) and not w28382;
w28384 <= not w27248 and w27687;
w28385 <= not w27683 and w28384;
w28386 <= not w27684 and not w27687;
w28387 <= not w28385 and not w28386;
w28388 <= not w27847 and not w28387;
w28389 <= not w27238 and not w27846;
w28390 <= not w27845 and w28389;
w28391 <= not w28388 and not w28390;
w28392 <= not w28383 and w28391;
w28393 <= not w28380 and w28392;
w28394 <= not b(34) and not w28393;
w28395 <= not w28380 and not w28383;
w28396 <= not w28391 and not w28395;
w28397 <= not w28394 and not w28396;
w28398 <= not w27959 and not w28397;
w28399 <= w27959 and not w28396;
w28400 <= not w28394 and w28399;
w28401 <= not b(35) and not w28400;
w28402 <= not w27230 and w27697;
w28403 <= not w27693 and w28402;
w28404 <= not w27694 and not w27697;
w28405 <= not w28403 and not w28404;
w28406 <= not w27847 and not w28405;
w28407 <= not w27220 and not w27846;
w28408 <= not w27845 and w28407;
w28409 <= not w28406 and not w28408;
w28410 <= not w28401 and w28409;
w28411 <= not w28398 and w28410;
w28412 <= not b(36) and not w28411;
w28413 <= not w28398 and not w28401;
w28414 <= not w28409 and not w28413;
w28415 <= not w28412 and not w28414;
w28416 <= not w27951 and not w28415;
w28417 <= w27951 and not w28414;
w28418 <= not w28412 and w28417;
w28419 <= not b(37) and not w28418;
w28420 <= not w27212 and w27707;
w28421 <= not w27703 and w28420;
w28422 <= not w27704 and not w27707;
w28423 <= not w28421 and not w28422;
w28424 <= not w27847 and not w28423;
w28425 <= not w27202 and not w27846;
w28426 <= not w27845 and w28425;
w28427 <= not w28424 and not w28426;
w28428 <= not w28419 and w28427;
w28429 <= not w28416 and w28428;
w28430 <= not b(38) and not w28429;
w28431 <= not w28416 and not w28419;
w28432 <= not w28427 and not w28431;
w28433 <= not w28430 and not w28432;
w28434 <= not w27943 and not w28433;
w28435 <= w27943 and not w28432;
w28436 <= not w28430 and w28435;
w28437 <= not b(39) and not w28436;
w28438 <= not w27194 and w27717;
w28439 <= not w27713 and w28438;
w28440 <= not w27714 and not w27717;
w28441 <= not w28439 and not w28440;
w28442 <= not w27847 and not w28441;
w28443 <= not w27184 and not w27846;
w28444 <= not w27845 and w28443;
w28445 <= not w28442 and not w28444;
w28446 <= not w28437 and w28445;
w28447 <= not w28434 and w28446;
w28448 <= not b(40) and not w28447;
w28449 <= not w28434 and not w28437;
w28450 <= not w28445 and not w28449;
w28451 <= not w28448 and not w28450;
w28452 <= not w27935 and not w28451;
w28453 <= w27935 and not w28450;
w28454 <= not w28448 and w28453;
w28455 <= not b(41) and not w28454;
w28456 <= not w27176 and w27727;
w28457 <= not w27723 and w28456;
w28458 <= not w27724 and not w27727;
w28459 <= not w28457 and not w28458;
w28460 <= not w27847 and not w28459;
w28461 <= not w27166 and not w27846;
w28462 <= not w27845 and w28461;
w28463 <= not w28460 and not w28462;
w28464 <= not w28455 and w28463;
w28465 <= not w28452 and w28464;
w28466 <= not b(42) and not w28465;
w28467 <= not w28452 and not w28455;
w28468 <= not w28463 and not w28467;
w28469 <= not w28466 and not w28468;
w28470 <= not w27927 and not w28469;
w28471 <= w27927 and not w28468;
w28472 <= not w28466 and w28471;
w28473 <= not b(43) and not w28472;
w28474 <= not w27158 and w27737;
w28475 <= not w27733 and w28474;
w28476 <= not w27734 and not w27737;
w28477 <= not w28475 and not w28476;
w28478 <= not w27847 and not w28477;
w28479 <= not w27148 and not w27846;
w28480 <= not w27845 and w28479;
w28481 <= not w28478 and not w28480;
w28482 <= not w28473 and w28481;
w28483 <= not w28470 and w28482;
w28484 <= not b(44) and not w28483;
w28485 <= not w28470 and not w28473;
w28486 <= not w28481 and not w28485;
w28487 <= not w28484 and not w28486;
w28488 <= not w27919 and not w28487;
w28489 <= w27919 and not w28486;
w28490 <= not w28484 and w28489;
w28491 <= not b(45) and not w28490;
w28492 <= not w27140 and w27747;
w28493 <= not w27743 and w28492;
w28494 <= not w27744 and not w27747;
w28495 <= not w28493 and not w28494;
w28496 <= not w27847 and not w28495;
w28497 <= not w27130 and not w27846;
w28498 <= not w27845 and w28497;
w28499 <= not w28496 and not w28498;
w28500 <= not w28491 and w28499;
w28501 <= not w28488 and w28500;
w28502 <= not b(46) and not w28501;
w28503 <= not w28488 and not w28491;
w28504 <= not w28499 and not w28503;
w28505 <= not w28502 and not w28504;
w28506 <= not w27911 and not w28505;
w28507 <= w27911 and not w28504;
w28508 <= not w28502 and w28507;
w28509 <= not b(47) and not w28508;
w28510 <= not w27122 and w27757;
w28511 <= not w27753 and w28510;
w28512 <= not w27754 and not w27757;
w28513 <= not w28511 and not w28512;
w28514 <= not w27847 and not w28513;
w28515 <= not w27112 and not w27846;
w28516 <= not w27845 and w28515;
w28517 <= not w28514 and not w28516;
w28518 <= not w28509 and w28517;
w28519 <= not w28506 and w28518;
w28520 <= not b(48) and not w28519;
w28521 <= not w28506 and not w28509;
w28522 <= not w28517 and not w28521;
w28523 <= not w28520 and not w28522;
w28524 <= not w27903 and not w28523;
w28525 <= w27903 and not w28522;
w28526 <= not w28520 and w28525;
w28527 <= not b(49) and not w28526;
w28528 <= not w27104 and w27767;
w28529 <= not w27763 and w28528;
w28530 <= not w27764 and not w27767;
w28531 <= not w28529 and not w28530;
w28532 <= not w27847 and not w28531;
w28533 <= not w27094 and not w27846;
w28534 <= not w27845 and w28533;
w28535 <= not w28532 and not w28534;
w28536 <= not w28527 and w28535;
w28537 <= not w28524 and w28536;
w28538 <= not b(50) and not w28537;
w28539 <= not w28524 and not w28527;
w28540 <= not w28535 and not w28539;
w28541 <= not w28538 and not w28540;
w28542 <= not w27895 and not w28541;
w28543 <= w27895 and not w28540;
w28544 <= not w28538 and w28543;
w28545 <= not b(51) and not w28544;
w28546 <= not w27086 and w27777;
w28547 <= not w27773 and w28546;
w28548 <= not w27774 and not w27777;
w28549 <= not w28547 and not w28548;
w28550 <= not w27847 and not w28549;
w28551 <= not w27076 and not w27846;
w28552 <= not w27845 and w28551;
w28553 <= not w28550 and not w28552;
w28554 <= not w28545 and w28553;
w28555 <= not w28542 and w28554;
w28556 <= not b(52) and not w28555;
w28557 <= not w28542 and not w28545;
w28558 <= not w28553 and not w28557;
w28559 <= not w28556 and not w28558;
w28560 <= not w27887 and not w28559;
w28561 <= w27887 and not w28558;
w28562 <= not w28556 and w28561;
w28563 <= not b(53) and not w28562;
w28564 <= not w27068 and w27787;
w28565 <= not w27783 and w28564;
w28566 <= not w27784 and not w27787;
w28567 <= not w28565 and not w28566;
w28568 <= not w27847 and not w28567;
w28569 <= not w27058 and not w27846;
w28570 <= not w27845 and w28569;
w28571 <= not w28568 and not w28570;
w28572 <= not w28563 and w28571;
w28573 <= not w28560 and w28572;
w28574 <= not b(54) and not w28573;
w28575 <= not w28560 and not w28563;
w28576 <= not w28571 and not w28575;
w28577 <= not w28574 and not w28576;
w28578 <= not w27879 and not w28577;
w28579 <= w27879 and not w28576;
w28580 <= not w28574 and w28579;
w28581 <= not b(55) and not w28580;
w28582 <= not w27050 and w27797;
w28583 <= not w27793 and w28582;
w28584 <= not w27794 and not w27797;
w28585 <= not w28583 and not w28584;
w28586 <= not w27847 and not w28585;
w28587 <= not w27040 and not w27846;
w28588 <= not w27845 and w28587;
w28589 <= not w28586 and not w28588;
w28590 <= not w28581 and w28589;
w28591 <= not w28578 and w28590;
w28592 <= not b(56) and not w28591;
w28593 <= not w28578 and not w28581;
w28594 <= not w28589 and not w28593;
w28595 <= not w28592 and not w28594;
w28596 <= not w27871 and not w28595;
w28597 <= w27871 and not w28594;
w28598 <= not w28592 and w28597;
w28599 <= not b(57) and not w28598;
w28600 <= not w27032 and w27807;
w28601 <= not w27803 and w28600;
w28602 <= not w27804 and not w27807;
w28603 <= not w28601 and not w28602;
w28604 <= not w27847 and not w28603;
w28605 <= not w27022 and not w27846;
w28606 <= not w27845 and w28605;
w28607 <= not w28604 and not w28606;
w28608 <= not w28599 and w28607;
w28609 <= not w28596 and w28608;
w28610 <= not b(58) and not w28609;
w28611 <= not w28596 and not w28599;
w28612 <= not w28607 and not w28611;
w28613 <= not w28610 and not w28612;
w28614 <= not w27863 and not w28613;
w28615 <= w27863 and not w28612;
w28616 <= not w28610 and w28615;
w28617 <= not b(59) and not w28616;
w28618 <= not w27014 and w27817;
w28619 <= not w27813 and w28618;
w28620 <= not w27814 and not w27817;
w28621 <= not w28619 and not w28620;
w28622 <= not w27847 and not w28621;
w28623 <= not w27004 and not w27846;
w28624 <= not w27845 and w28623;
w28625 <= not w28622 and not w28624;
w28626 <= not w28617 and w28625;
w28627 <= not w28614 and w28626;
w28628 <= not b(60) and not w28627;
w28629 <= not w28614 and not w28617;
w28630 <= not w28625 and not w28629;
w28631 <= not w28628 and not w28630;
w28632 <= not w27855 and not w28631;
w28633 <= w27855 and not w28630;
w28634 <= not w28628 and w28633;
w28635 <= not b(61) and not w28634;
w28636 <= not w26996 and w27827;
w28637 <= not w27823 and w28636;
w28638 <= not w27824 and not w27827;
w28639 <= not w28637 and not w28638;
w28640 <= not w27847 and not w28639;
w28641 <= not w26986 and not w27846;
w28642 <= not w27845 and w28641;
w28643 <= not w28640 and not w28642;
w28644 <= not w28635 and w28643;
w28645 <= not w28632 and w28644;
w28646 <= not b(62) and not w28645;
w28647 <= not w28632 and not w28635;
w28648 <= not w28643 and not w28647;
w28649 <= not w26987 and not w27842;
w28650 <= not w27840 and w28649;
w28651 <= not w27828 and w28650;
w28652 <= not w27840 and not w27842;
w28653 <= not w27829 and not w28652;
w28654 <= not w28651 and not w28653;
w28655 <= not w27847 and not w28654;
w28656 <= not w27839 and not w27846;
w28657 <= not w27845 and w28656;
w28658 <= not w28655 and not w28657;
w28659 <= not w28648 and w28658;
w28660 <= not w28646 and w28659;
w28661 <= not b(63) and not w28660;
w28662 <= not w28646 and not w28648;
w28663 <= not w28658 and not w28662;
w28664 <= not w28661 and not w28663;
w28665 <= not w326 and w343;
w28666 <= w77 and w87;
w28667 <= w175 and w28666;
w28668 <= not w70 and w28667;
w28669 <= not b(1) and not b(2);
w28670 <= w126 and w28669;
w28671 <= not w0 and w28670;
w28672 <= w335 and w28671;
w28673 <= w386 and w28672;
w28674 <= w3 and w10;
w28675 <= w76 and w28674;
w28676 <= w87 and w28675;
w28677 <= w175 and w28676;
w28678 <= w67 and not w28677;
w28679 <= not w69 and not w28678;
w28680 <= a(63) and not w28677;
w28681 <= w90 and not w28680;
w28682 <= not w28679 and w28681;
w28683 <= w101 and not w28679;
w28684 <= w28680 and not w28683;
w28685 <= not w28682 and not w28684;
w28686 <= w168 and not w28679;
w28687 <= a(62) and not w28686;
w28688 <= w176 and not w28679;
w28689 <= not w28687 and not w28688;
w28690 <= not w106 and not w28689;
w28691 <= not w180 and not w28690;
w28692 <= b(2) and not w28682;
w28693 <= not w28684 and w28692;
w28694 <= not b(2) and not w28685;
w28695 <= not w28693 and not w28694;
w28696 <= w28691 and not w28695;
w28697 <= not b(2) and not w28696;
w28698 <= not w28691 and not w28693;
w28699 <= not w28694 and not w28698;
w28700 <= w193 and not w28699;
w28701 <= not w28697 and w28700;
w28702 <= not w28685 and not w28701;
w28703 <= w193 and not w28698;
w28704 <= not w28696 and w28703;
w28705 <= not w28699 and w28704;
w28706 <= b(3) and not w28705;
w28707 <= not w28702 and w28706;
w28708 <= w210 and not w28699;
w28709 <= not w28689 and not w28708;
w28710 <= w219 and not w28688;
w28711 <= not w28687 and w28710;
w28712 <= not w28699 and w28711;
w28713 <= not w28709 and not w28712;
w28714 <= not b(2) and not w28713;
w28715 <= b(2) and not w28712;
w28716 <= not w28709 and w28715;
w28717 <= w231 and not w28699;
w28718 <= a(61) and not w28717;
w28719 <= w238 and not w28699;
w28720 <= not w28718 and not w28719;
w28721 <= not w242 and not w28720;
w28722 <= not w244 and not w28721;
w28723 <= not w28716 and not w28722;
w28724 <= not w28714 and not w28723;
w28725 <= not w28707 and not w28724;
w28726 <= not w28702 and not w28705;
w28727 <= not b(3) and not w28726;
w28728 <= not w28725 and not w28727;
w28729 <= not w28707 and not w28727;
w28730 <= not w28724 and w28729;
w28731 <= w28724 and not w28729;
w28732 <= w256 and not w28731;
w28733 <= not w28730 and w28732;
w28734 <= not w28728 and w28733;
w28735 <= w256 and not w28728;
w28736 <= not w28726 and not w28735;
w28737 <= b(4) and not w28736;
w28738 <= not w28734 and w28737;
w28739 <= not w28714 and not w28716;
w28740 <= w28722 and not w28739;
w28741 <= w256 and not w28723;
w28742 <= not w28740 and w28741;
w28743 <= not w28728 and w28742;
w28744 <= not b(2) and not w28740;
w28745 <= w256 and not w28744;
w28746 <= not w28728 and w28745;
w28747 <= not w28713 and not w28746;
w28748 <= not w28743 and not w28747;
w28749 <= not b(3) and not w28748;
w28750 <= b(3) and not w28743;
w28751 <= not w28747 and w28750;
w28752 <= w286 and not w28728;
w28753 <= not w28720 and not w28752;
w28754 <= w293 and not w28719;
w28755 <= not w28718 and w28754;
w28756 <= not w28728 and w28755;
w28757 <= not w28753 and not w28756;
w28758 <= not b(2) and not w28757;
w28759 <= b(2) and not w28756;
w28760 <= not w28753 and w28759;
w28761 <= w307 and not w28728;
w28762 <= a(60) and not w28761;
w28763 <= w313 and not w28728;
w28764 <= not w28762 and not w28763;
w28765 <= not w302 and not w28764;
w28766 <= not w317 and not w28765;
w28767 <= not w28760 and not w28766;
w28768 <= not w28758 and not w28767;
w28769 <= not w28751 and not w28768;
w28770 <= not w28749 and not w28769;
w28771 <= not w28738 and not w28770;
w28772 <= not w28734 and not w28736;
w28773 <= not b(4) and not w28772;
w28774 <= not w28771 and not w28773;
w28775 <= not w28749 and not w28751;
w28776 <= not w28758 and not w28775;
w28777 <= not w28767 and w28776;
w28778 <= w343 and not w28777;
w28779 <= not w28769 and w28778;
w28780 <= not w28774 and w28779;
w28781 <= not b(3) and not w28777;
w28782 <= w343 and not w28781;
w28783 <= not w28774 and w28782;
w28784 <= not w28748 and not w28783;
w28785 <= not w28780 and not w28784;
w28786 <= b(4) and not w28785;
w28787 <= not b(4) and not w28780;
w28788 <= not w28784 and w28787;
w28789 <= not w28786 and not w28788;
w28790 <= not w28758 and not w28760;
w28791 <= w28766 and not w28790;
w28792 <= w343 and not w28767;
w28793 <= not w28791 and w28792;
w28794 <= not w28774 and w28793;
w28795 <= not b(2) and not w28791;
w28796 <= w343 and not w28795;
w28797 <= not w28774 and w28796;
w28798 <= not w28757 and not w28797;
w28799 <= not w28794 and not w28798;
w28800 <= b(3) and not w28799;
w28801 <= not b(3) and not w28794;
w28802 <= not w28798 and w28801;
w28803 <= not w28800 and not w28802;
w28804 <= w378 and not w28774;
w28805 <= not w28764 and not w28804;
w28806 <= w387 and not w28763;
w28807 <= not w28762 and w28806;
w28808 <= not w28774 and w28807;
w28809 <= not w28805 and not w28808;
w28810 <= not b(2) and not w28809;
w28811 <= w398 and not w28774;
w28812 <= a(59) and not w28811;
w28813 <= w404 and not w28774;
w28814 <= not w28812 and not w28813;
w28815 <= b(1) and not w28814;
w28816 <= not b(1) and not w28813;
w28817 <= not w28812 and w28816;
w28818 <= not w28815 and not w28817;
w28819 <= not w411 and not w28818;
w28820 <= not b(1) and not w28814;
w28821 <= not w28819 and not w28820;
w28822 <= b(2) and not w28808;
w28823 <= not w28805 and w28822;
w28824 <= not w28810 and not w28823;
w28825 <= not w28821 and w28824;
w28826 <= not w28810 and not w28825;
w28827 <= not w28803 and not w28826;
w28828 <= not b(3) and not w28799;
w28829 <= not w28827 and not w28828;
w28830 <= not w28789 and not w28829;
w28831 <= not b(4) and not w28785;
w28832 <= not w28830 and not w28831;
w28833 <= not w28738 and not w28773;
w28834 <= not w28749 and not w28833;
w28835 <= not w28769 and w28834;
w28836 <= w343 and not w28835;
w28837 <= not w28771 and w28836;
w28838 <= not w28774 and w28837;
w28839 <= not b(4) and not w28835;
w28840 <= w343 and not w28839;
w28841 <= not w28774 and w28840;
w28842 <= not w28772 and not w28841;
w28843 <= not w28838 and not w28842;
w28844 <= b(5) and not w28843;
w28845 <= not b(5) and not w28838;
w28846 <= not w28842 and w28845;
w28847 <= not w28844 and not w28846;
w28848 <= w444 and not w28847;
w28849 <= not w28832 and w28848;
w28850 <= w343 and not w28843;
w28851 <= not w28849 and not w28850;
w28852 <= w28789 and not w28828;
w28853 <= not w28827 and w28852;
w28854 <= not w28830 and not w28853;
w28855 <= not w28851 and w28854;
w28856 <= not w28785 and not w28850;
w28857 <= not w28849 and w28856;
w28858 <= not w28855 and not w28857;
w28859 <= not w28832 and not w28847;
w28860 <= not w28831 and w28847;
w28861 <= not w28830 and w28860;
w28862 <= not w28859 and not w28861;
w28863 <= not w28851 and w28862;
w28864 <= not w28843 and not w28850;
w28865 <= not w28849 and w28864;
w28866 <= not w28863 and not w28865;
w28867 <= not b(6) and not w28866;
w28868 <= not b(5) and not w28858;
w28869 <= w28803 and not w28810;
w28870 <= not w28825 and w28869;
w28871 <= not w28827 and not w28870;
w28872 <= not w28851 and w28871;
w28873 <= not w28799 and not w28850;
w28874 <= not w28849 and w28873;
w28875 <= not w28872 and not w28874;
w28876 <= not b(4) and not w28875;
w28877 <= not w28820 and w28824;
w28878 <= not w28819 and w28877;
w28879 <= not w28821 and not w28824;
w28880 <= not w28878 and not w28879;
w28881 <= not w28851 and not w28880;
w28882 <= not w28809 and not w28850;
w28883 <= not w28849 and w28882;
w28884 <= not w28881 and not w28883;
w28885 <= not b(3) and not w28884;
w28886 <= w411 and not w28817;
w28887 <= not w28815 and w28886;
w28888 <= not w28819 and not w28887;
w28889 <= not w28851 and w28888;
w28890 <= not w28814 and not w28850;
w28891 <= not w28849 and w28890;
w28892 <= not w28889 and not w28891;
w28893 <= not b(2) and not w28892;
w28894 <= b(0) and not w28851;
w28895 <= a(58) and not w28894;
w28896 <= w411 and not w28851;
w28897 <= not w28895 and not w28896;
w28898 <= b(1) and not w28897;
w28899 <= not b(1) and not w28896;
w28900 <= not w28895 and w28899;
w28901 <= not w28898 and not w28900;
w28902 <= not w499 and not w28901;
w28903 <= not b(1) and not w28897;
w28904 <= not w28902 and not w28903;
w28905 <= b(2) and not w28891;
w28906 <= not w28889 and w28905;
w28907 <= not w28893 and not w28906;
w28908 <= not w28904 and w28907;
w28909 <= not w28893 and not w28908;
w28910 <= b(3) and not w28883;
w28911 <= not w28881 and w28910;
w28912 <= not w28885 and not w28911;
w28913 <= not w28909 and w28912;
w28914 <= not w28885 and not w28913;
w28915 <= b(4) and not w28874;
w28916 <= not w28872 and w28915;
w28917 <= not w28876 and not w28916;
w28918 <= not w28914 and w28917;
w28919 <= not w28876 and not w28918;
w28920 <= b(5) and not w28857;
w28921 <= not w28855 and w28920;
w28922 <= not w28868 and not w28921;
w28923 <= not w28919 and w28922;
w28924 <= not w28868 and not w28923;
w28925 <= b(6) and not w28865;
w28926 <= not w28863 and w28925;
w28927 <= not w28867 and not w28926;
w28928 <= not w28924 and w28927;
w28929 <= not w28867 and not w28928;
w28930 <= w531 and not w28929;
w28931 <= not w28858 and not w28930;
w28932 <= not w28876 and w28922;
w28933 <= not w28918 and w28932;
w28934 <= not w28919 and not w28922;
w28935 <= not w28933 and not w28934;
w28936 <= w531 and not w28935;
w28937 <= not w28929 and w28936;
w28938 <= not w28931 and not w28937;
w28939 <= not w28866 and not w28930;
w28940 <= not w28868 and w28927;
w28941 <= not w28923 and w28940;
w28942 <= not w28924 and not w28927;
w28943 <= not w28941 and not w28942;
w28944 <= w28930 and not w28943;
w28945 <= not w28939 and not w28944;
w28946 <= not b(7) and not w28945;
w28947 <= not b(6) and not w28938;
w28948 <= not w28875 and not w28930;
w28949 <= not w28885 and w28917;
w28950 <= not w28913 and w28949;
w28951 <= not w28914 and not w28917;
w28952 <= not w28950 and not w28951;
w28953 <= w531 and not w28952;
w28954 <= not w28929 and w28953;
w28955 <= not w28948 and not w28954;
w28956 <= not b(5) and not w28955;
w28957 <= not w28884 and not w28930;
w28958 <= not w28893 and w28912;
w28959 <= not w28908 and w28958;
w28960 <= not w28909 and not w28912;
w28961 <= not w28959 and not w28960;
w28962 <= w531 and not w28961;
w28963 <= not w28929 and w28962;
w28964 <= not w28957 and not w28963;
w28965 <= not b(4) and not w28964;
w28966 <= not w28892 and not w28930;
w28967 <= not w28903 and w28907;
w28968 <= not w28902 and w28967;
w28969 <= not w28904 and not w28907;
w28970 <= not w28968 and not w28969;
w28971 <= w531 and not w28970;
w28972 <= not w28929 and w28971;
w28973 <= not w28966 and not w28972;
w28974 <= not b(3) and not w28973;
w28975 <= not w28897 and not w28930;
w28976 <= w499 and not w28900;
w28977 <= not w28898 and w28976;
w28978 <= w531 and not w28977;
w28979 <= not w28902 and w28978;
w28980 <= not w28929 and w28979;
w28981 <= not w28975 and not w28980;
w28982 <= not b(2) and not w28981;
w28983 <= w589 and not w28929;
w28984 <= a(57) and not w28983;
w28985 <= w596 and not w28929;
w28986 <= not w28984 and not w28985;
w28987 <= b(1) and not w28986;
w28988 <= not b(1) and not w28985;
w28989 <= not w28984 and w28988;
w28990 <= not w28987 and not w28989;
w28991 <= not w603 and not w28990;
w28992 <= not b(1) and not w28986;
w28993 <= not w28991 and not w28992;
w28994 <= b(2) and not w28980;
w28995 <= not w28975 and w28994;
w28996 <= not w28982 and not w28995;
w28997 <= not w28993 and w28996;
w28998 <= not w28982 and not w28997;
w28999 <= b(3) and not w28972;
w29000 <= not w28966 and w28999;
w29001 <= not w28974 and not w29000;
w29002 <= not w28998 and w29001;
w29003 <= not w28974 and not w29002;
w29004 <= b(4) and not w28963;
w29005 <= not w28957 and w29004;
w29006 <= not w28965 and not w29005;
w29007 <= not w29003 and w29006;
w29008 <= not w28965 and not w29007;
w29009 <= b(5) and not w28954;
w29010 <= not w28948 and w29009;
w29011 <= not w28956 and not w29010;
w29012 <= not w29008 and w29011;
w29013 <= not w28956 and not w29012;
w29014 <= b(6) and not w28937;
w29015 <= not w28931 and w29014;
w29016 <= not w28947 and not w29015;
w29017 <= not w29013 and w29016;
w29018 <= not w28947 and not w29017;
w29019 <= b(7) and not w28939;
w29020 <= not w28944 and w29019;
w29021 <= not w28946 and not w29020;
w29022 <= not w29018 and w29021;
w29023 <= not w28946 and not w29022;
w29024 <= w638 and not w29023;
w29025 <= not w28938 and not w29024;
w29026 <= not w28956 and w29016;
w29027 <= not w29012 and w29026;
w29028 <= not w29013 and not w29016;
w29029 <= not w29027 and not w29028;
w29030 <= w638 and not w29029;
w29031 <= not w29023 and w29030;
w29032 <= not w29025 and not w29031;
w29033 <= not b(7) and not w29032;
w29034 <= not w28955 and not w29024;
w29035 <= not w28965 and w29011;
w29036 <= not w29007 and w29035;
w29037 <= not w29008 and not w29011;
w29038 <= not w29036 and not w29037;
w29039 <= w638 and not w29038;
w29040 <= not w29023 and w29039;
w29041 <= not w29034 and not w29040;
w29042 <= not b(6) and not w29041;
w29043 <= not w28964 and not w29024;
w29044 <= not w28974 and w29006;
w29045 <= not w29002 and w29044;
w29046 <= not w29003 and not w29006;
w29047 <= not w29045 and not w29046;
w29048 <= w638 and not w29047;
w29049 <= not w29023 and w29048;
w29050 <= not w29043 and not w29049;
w29051 <= not b(5) and not w29050;
w29052 <= not w28973 and not w29024;
w29053 <= not w28982 and w29001;
w29054 <= not w28997 and w29053;
w29055 <= not w28998 and not w29001;
w29056 <= not w29054 and not w29055;
w29057 <= w638 and not w29056;
w29058 <= not w29023 and w29057;
w29059 <= not w29052 and not w29058;
w29060 <= not b(4) and not w29059;
w29061 <= not w28981 and not w29024;
w29062 <= not w28992 and w28996;
w29063 <= not w28991 and w29062;
w29064 <= not w28993 and not w28996;
w29065 <= not w29063 and not w29064;
w29066 <= w638 and not w29065;
w29067 <= not w29023 and w29066;
w29068 <= not w29061 and not w29067;
w29069 <= not b(3) and not w29068;
w29070 <= not w28986 and not w29024;
w29071 <= w603 and not w28989;
w29072 <= not w28987 and w29071;
w29073 <= w638 and not w29072;
w29074 <= not w28991 and w29073;
w29075 <= not w29023 and w29074;
w29076 <= not w29070 and not w29075;
w29077 <= not b(2) and not w29076;
w29078 <= w697 and not w29023;
w29079 <= a(56) and not w29078;
w29080 <= w703 and not w29023;
w29081 <= not w29079 and not w29080;
w29082 <= b(1) and not w29081;
w29083 <= not b(1) and not w29080;
w29084 <= not w29079 and w29083;
w29085 <= not w29082 and not w29084;
w29086 <= not w710 and not w29085;
w29087 <= not b(1) and not w29081;
w29088 <= not w29086 and not w29087;
w29089 <= b(2) and not w29075;
w29090 <= not w29070 and w29089;
w29091 <= not w29077 and not w29090;
w29092 <= not w29088 and w29091;
w29093 <= not w29077 and not w29092;
w29094 <= b(3) and not w29067;
w29095 <= not w29061 and w29094;
w29096 <= not w29069 and not w29095;
w29097 <= not w29093 and w29096;
w29098 <= not w29069 and not w29097;
w29099 <= b(4) and not w29058;
w29100 <= not w29052 and w29099;
w29101 <= not w29060 and not w29100;
w29102 <= not w29098 and w29101;
w29103 <= not w29060 and not w29102;
w29104 <= b(5) and not w29049;
w29105 <= not w29043 and w29104;
w29106 <= not w29051 and not w29105;
w29107 <= not w29103 and w29106;
w29108 <= not w29051 and not w29107;
w29109 <= b(6) and not w29040;
w29110 <= not w29034 and w29109;
w29111 <= not w29042 and not w29110;
w29112 <= not w29108 and w29111;
w29113 <= not w29042 and not w29112;
w29114 <= b(7) and not w29031;
w29115 <= not w29025 and w29114;
w29116 <= not w29033 and not w29115;
w29117 <= not w29113 and w29116;
w29118 <= not w29033 and not w29117;
w29119 <= not w28945 and not w29024;
w29120 <= not w28947 and w29021;
w29121 <= not w29017 and w29120;
w29122 <= not w29018 and not w29021;
w29123 <= not w29121 and not w29122;
w29124 <= w29024 and not w29123;
w29125 <= not w29119 and not w29124;
w29126 <= not b(8) and not w29125;
w29127 <= b(8) and not w29119;
w29128 <= not w29124 and w29127;
w29129 <= w755 and not w29128;
w29130 <= not w29126 and w29129;
w29131 <= not w29118 and w29130;
w29132 <= w638 and not w29125;
w29133 <= not w29131 and not w29132;
w29134 <= not w29042 and w29116;
w29135 <= not w29112 and w29134;
w29136 <= not w29113 and not w29116;
w29137 <= not w29135 and not w29136;
w29138 <= not w29133 and not w29137;
w29139 <= not w29032 and not w29132;
w29140 <= not w29131 and w29139;
w29141 <= not w29138 and not w29140;
w29142 <= not w29033 and not w29128;
w29143 <= not w29126 and w29142;
w29144 <= not w29117 and w29143;
w29145 <= not w29126 and not w29128;
w29146 <= not w29118 and not w29145;
w29147 <= not w29144 and not w29146;
w29148 <= not w29133 and not w29147;
w29149 <= not w29125 and not w29132;
w29150 <= not w29131 and w29149;
w29151 <= not w29148 and not w29150;
w29152 <= not b(9) and not w29151;
w29153 <= not b(8) and not w29141;
w29154 <= not w29051 and w29111;
w29155 <= not w29107 and w29154;
w29156 <= not w29108 and not w29111;
w29157 <= not w29155 and not w29156;
w29158 <= not w29133 and not w29157;
w29159 <= not w29041 and not w29132;
w29160 <= not w29131 and w29159;
w29161 <= not w29158 and not w29160;
w29162 <= not b(7) and not w29161;
w29163 <= not w29060 and w29106;
w29164 <= not w29102 and w29163;
w29165 <= not w29103 and not w29106;
w29166 <= not w29164 and not w29165;
w29167 <= not w29133 and not w29166;
w29168 <= not w29050 and not w29132;
w29169 <= not w29131 and w29168;
w29170 <= not w29167 and not w29169;
w29171 <= not b(6) and not w29170;
w29172 <= not w29069 and w29101;
w29173 <= not w29097 and w29172;
w29174 <= not w29098 and not w29101;
w29175 <= not w29173 and not w29174;
w29176 <= not w29133 and not w29175;
w29177 <= not w29059 and not w29132;
w29178 <= not w29131 and w29177;
w29179 <= not w29176 and not w29178;
w29180 <= not b(5) and not w29179;
w29181 <= not w29077 and w29096;
w29182 <= not w29092 and w29181;
w29183 <= not w29093 and not w29096;
w29184 <= not w29182 and not w29183;
w29185 <= not w29133 and not w29184;
w29186 <= not w29068 and not w29132;
w29187 <= not w29131 and w29186;
w29188 <= not w29185 and not w29187;
w29189 <= not b(4) and not w29188;
w29190 <= not w29087 and w29091;
w29191 <= not w29086 and w29190;
w29192 <= not w29088 and not w29091;
w29193 <= not w29191 and not w29192;
w29194 <= not w29133 and not w29193;
w29195 <= not w29076 and not w29132;
w29196 <= not w29131 and w29195;
w29197 <= not w29194 and not w29196;
w29198 <= not b(3) and not w29197;
w29199 <= w710 and not w29084;
w29200 <= not w29082 and w29199;
w29201 <= not w29086 and not w29200;
w29202 <= not w29133 and w29201;
w29203 <= not w29081 and not w29132;
w29204 <= not w29131 and w29203;
w29205 <= not w29202 and not w29204;
w29206 <= not b(2) and not w29205;
w29207 <= b(0) and not w29133;
w29208 <= a(55) and not w29207;
w29209 <= w710 and not w29133;
w29210 <= not w29208 and not w29209;
w29211 <= b(1) and not w29210;
w29212 <= not b(1) and not w29209;
w29213 <= not w29208 and w29212;
w29214 <= not w29211 and not w29213;
w29215 <= not w842 and not w29214;
w29216 <= not b(1) and not w29210;
w29217 <= not w29215 and not w29216;
w29218 <= b(2) and not w29204;
w29219 <= not w29202 and w29218;
w29220 <= not w29206 and not w29219;
w29221 <= not w29217 and w29220;
w29222 <= not w29206 and not w29221;
w29223 <= b(3) and not w29196;
w29224 <= not w29194 and w29223;
w29225 <= not w29198 and not w29224;
w29226 <= not w29222 and w29225;
w29227 <= not w29198 and not w29226;
w29228 <= b(4) and not w29187;
w29229 <= not w29185 and w29228;
w29230 <= not w29189 and not w29229;
w29231 <= not w29227 and w29230;
w29232 <= not w29189 and not w29231;
w29233 <= b(5) and not w29178;
w29234 <= not w29176 and w29233;
w29235 <= not w29180 and not w29234;
w29236 <= not w29232 and w29235;
w29237 <= not w29180 and not w29236;
w29238 <= b(6) and not w29169;
w29239 <= not w29167 and w29238;
w29240 <= not w29171 and not w29239;
w29241 <= not w29237 and w29240;
w29242 <= not w29171 and not w29241;
w29243 <= b(7) and not w29160;
w29244 <= not w29158 and w29243;
w29245 <= not w29162 and not w29244;
w29246 <= not w29242 and w29245;
w29247 <= not w29162 and not w29246;
w29248 <= b(8) and not w29140;
w29249 <= not w29138 and w29248;
w29250 <= not w29153 and not w29249;
w29251 <= not w29247 and w29250;
w29252 <= not w29153 and not w29251;
w29253 <= b(9) and not w29150;
w29254 <= not w29148 and w29253;
w29255 <= not w29152 and not w29254;
w29256 <= not w29252 and w29255;
w29257 <= not w29152 and not w29256;
w29258 <= w888 and not w29257;
w29259 <= not w29141 and not w29258;
w29260 <= not w29162 and w29250;
w29261 <= not w29246 and w29260;
w29262 <= not w29247 and not w29250;
w29263 <= not w29261 and not w29262;
w29264 <= w888 and not w29263;
w29265 <= not w29257 and w29264;
w29266 <= not w29259 and not w29265;
w29267 <= not w29151 and not w29258;
w29268 <= not w29153 and w29255;
w29269 <= not w29251 and w29268;
w29270 <= not w29252 and not w29255;
w29271 <= not w29269 and not w29270;
w29272 <= w29258 and not w29271;
w29273 <= not w29267 and not w29272;
w29274 <= not b(10) and not w29273;
w29275 <= not b(9) and not w29266;
w29276 <= not w29161 and not w29258;
w29277 <= not w29171 and w29245;
w29278 <= not w29241 and w29277;
w29279 <= not w29242 and not w29245;
w29280 <= not w29278 and not w29279;
w29281 <= w888 and not w29280;
w29282 <= not w29257 and w29281;
w29283 <= not w29276 and not w29282;
w29284 <= not b(8) and not w29283;
w29285 <= not w29170 and not w29258;
w29286 <= not w29180 and w29240;
w29287 <= not w29236 and w29286;
w29288 <= not w29237 and not w29240;
w29289 <= not w29287 and not w29288;
w29290 <= w888 and not w29289;
w29291 <= not w29257 and w29290;
w29292 <= not w29285 and not w29291;
w29293 <= not b(7) and not w29292;
w29294 <= not w29179 and not w29258;
w29295 <= not w29189 and w29235;
w29296 <= not w29231 and w29295;
w29297 <= not w29232 and not w29235;
w29298 <= not w29296 and not w29297;
w29299 <= w888 and not w29298;
w29300 <= not w29257 and w29299;
w29301 <= not w29294 and not w29300;
w29302 <= not b(6) and not w29301;
w29303 <= not w29188 and not w29258;
w29304 <= not w29198 and w29230;
w29305 <= not w29226 and w29304;
w29306 <= not w29227 and not w29230;
w29307 <= not w29305 and not w29306;
w29308 <= w888 and not w29307;
w29309 <= not w29257 and w29308;
w29310 <= not w29303 and not w29309;
w29311 <= not b(5) and not w29310;
w29312 <= not w29197 and not w29258;
w29313 <= not w29206 and w29225;
w29314 <= not w29221 and w29313;
w29315 <= not w29222 and not w29225;
w29316 <= not w29314 and not w29315;
w29317 <= w888 and not w29316;
w29318 <= not w29257 and w29317;
w29319 <= not w29312 and not w29318;
w29320 <= not b(4) and not w29319;
w29321 <= not w29205 and not w29258;
w29322 <= not w29216 and w29220;
w29323 <= not w29215 and w29322;
w29324 <= not w29217 and not w29220;
w29325 <= not w29323 and not w29324;
w29326 <= w888 and not w29325;
w29327 <= not w29257 and w29326;
w29328 <= not w29321 and not w29327;
w29329 <= not b(3) and not w29328;
w29330 <= not w29210 and not w29258;
w29331 <= w842 and not w29213;
w29332 <= not w29211 and w29331;
w29333 <= w888 and not w29332;
w29334 <= not w29215 and w29333;
w29335 <= not w29257 and w29334;
w29336 <= not w29330 and not w29335;
w29337 <= not b(2) and not w29336;
w29338 <= w973 and not w29257;
w29339 <= a(54) and not w29338;
w29340 <= w979 and not w29257;
w29341 <= not w29339 and not w29340;
w29342 <= b(1) and not w29341;
w29343 <= not b(1) and not w29340;
w29344 <= not w29339 and w29343;
w29345 <= not w29342 and not w29344;
w29346 <= not w986 and not w29345;
w29347 <= not b(1) and not w29341;
w29348 <= not w29346 and not w29347;
w29349 <= b(2) and not w29335;
w29350 <= not w29330 and w29349;
w29351 <= not w29337 and not w29350;
w29352 <= not w29348 and w29351;
w29353 <= not w29337 and not w29352;
w29354 <= b(3) and not w29327;
w29355 <= not w29321 and w29354;
w29356 <= not w29329 and not w29355;
w29357 <= not w29353 and w29356;
w29358 <= not w29329 and not w29357;
w29359 <= b(4) and not w29318;
w29360 <= not w29312 and w29359;
w29361 <= not w29320 and not w29360;
w29362 <= not w29358 and w29361;
w29363 <= not w29320 and not w29362;
w29364 <= b(5) and not w29309;
w29365 <= not w29303 and w29364;
w29366 <= not w29311 and not w29365;
w29367 <= not w29363 and w29366;
w29368 <= not w29311 and not w29367;
w29369 <= b(6) and not w29300;
w29370 <= not w29294 and w29369;
w29371 <= not w29302 and not w29370;
w29372 <= not w29368 and w29371;
w29373 <= not w29302 and not w29372;
w29374 <= b(7) and not w29291;
w29375 <= not w29285 and w29374;
w29376 <= not w29293 and not w29375;
w29377 <= not w29373 and w29376;
w29378 <= not w29293 and not w29377;
w29379 <= b(8) and not w29282;
w29380 <= not w29276 and w29379;
w29381 <= not w29284 and not w29380;
w29382 <= not w29378 and w29381;
w29383 <= not w29284 and not w29382;
w29384 <= b(9) and not w29265;
w29385 <= not w29259 and w29384;
w29386 <= not w29275 and not w29385;
w29387 <= not w29383 and w29386;
w29388 <= not w29275 and not w29387;
w29389 <= b(10) and not w29267;
w29390 <= not w29272 and w29389;
w29391 <= not w29274 and not w29390;
w29392 <= not w29388 and w29391;
w29393 <= not w29274 and not w29392;
w29394 <= w1037 and not w29393;
w29395 <= not w29266 and not w29394;
w29396 <= not w29284 and w29386;
w29397 <= not w29382 and w29396;
w29398 <= not w29383 and not w29386;
w29399 <= not w29397 and not w29398;
w29400 <= w1037 and not w29399;
w29401 <= not w29393 and w29400;
w29402 <= not w29395 and not w29401;
w29403 <= not b(10) and not w29402;
w29404 <= not w29283 and not w29394;
w29405 <= not w29293 and w29381;
w29406 <= not w29377 and w29405;
w29407 <= not w29378 and not w29381;
w29408 <= not w29406 and not w29407;
w29409 <= w1037 and not w29408;
w29410 <= not w29393 and w29409;
w29411 <= not w29404 and not w29410;
w29412 <= not b(9) and not w29411;
w29413 <= not w29292 and not w29394;
w29414 <= not w29302 and w29376;
w29415 <= not w29372 and w29414;
w29416 <= not w29373 and not w29376;
w29417 <= not w29415 and not w29416;
w29418 <= w1037 and not w29417;
w29419 <= not w29393 and w29418;
w29420 <= not w29413 and not w29419;
w29421 <= not b(8) and not w29420;
w29422 <= not w29301 and not w29394;
w29423 <= not w29311 and w29371;
w29424 <= not w29367 and w29423;
w29425 <= not w29368 and not w29371;
w29426 <= not w29424 and not w29425;
w29427 <= w1037 and not w29426;
w29428 <= not w29393 and w29427;
w29429 <= not w29422 and not w29428;
w29430 <= not b(7) and not w29429;
w29431 <= not w29310 and not w29394;
w29432 <= not w29320 and w29366;
w29433 <= not w29362 and w29432;
w29434 <= not w29363 and not w29366;
w29435 <= not w29433 and not w29434;
w29436 <= w1037 and not w29435;
w29437 <= not w29393 and w29436;
w29438 <= not w29431 and not w29437;
w29439 <= not b(6) and not w29438;
w29440 <= not w29319 and not w29394;
w29441 <= not w29329 and w29361;
w29442 <= not w29357 and w29441;
w29443 <= not w29358 and not w29361;
w29444 <= not w29442 and not w29443;
w29445 <= w1037 and not w29444;
w29446 <= not w29393 and w29445;
w29447 <= not w29440 and not w29446;
w29448 <= not b(5) and not w29447;
w29449 <= not w29328 and not w29394;
w29450 <= not w29337 and w29356;
w29451 <= not w29352 and w29450;
w29452 <= not w29353 and not w29356;
w29453 <= not w29451 and not w29452;
w29454 <= w1037 and not w29453;
w29455 <= not w29393 and w29454;
w29456 <= not w29449 and not w29455;
w29457 <= not b(4) and not w29456;
w29458 <= not w29336 and not w29394;
w29459 <= not w29347 and w29351;
w29460 <= not w29346 and w29459;
w29461 <= not w29348 and not w29351;
w29462 <= not w29460 and not w29461;
w29463 <= w1037 and not w29462;
w29464 <= not w29393 and w29463;
w29465 <= not w29458 and not w29464;
w29466 <= not b(3) and not w29465;
w29467 <= not w29341 and not w29394;
w29468 <= w986 and not w29344;
w29469 <= not w29342 and w29468;
w29470 <= w1037 and not w29469;
w29471 <= not w29346 and w29470;
w29472 <= not w29393 and w29471;
w29473 <= not w29467 and not w29472;
w29474 <= not b(2) and not w29473;
w29475 <= w1122 and not w29393;
w29476 <= a(53) and not w29475;
w29477 <= w1128 and not w29393;
w29478 <= not w29476 and not w29477;
w29479 <= b(1) and not w29478;
w29480 <= not b(1) and not w29477;
w29481 <= not w29476 and w29480;
w29482 <= not w29479 and not w29481;
w29483 <= not w1135 and not w29482;
w29484 <= not b(1) and not w29478;
w29485 <= not w29483 and not w29484;
w29486 <= b(2) and not w29472;
w29487 <= not w29467 and w29486;
w29488 <= not w29474 and not w29487;
w29489 <= not w29485 and w29488;
w29490 <= not w29474 and not w29489;
w29491 <= b(3) and not w29464;
w29492 <= not w29458 and w29491;
w29493 <= not w29466 and not w29492;
w29494 <= not w29490 and w29493;
w29495 <= not w29466 and not w29494;
w29496 <= b(4) and not w29455;
w29497 <= not w29449 and w29496;
w29498 <= not w29457 and not w29497;
w29499 <= not w29495 and w29498;
w29500 <= not w29457 and not w29499;
w29501 <= b(5) and not w29446;
w29502 <= not w29440 and w29501;
w29503 <= not w29448 and not w29502;
w29504 <= not w29500 and w29503;
w29505 <= not w29448 and not w29504;
w29506 <= b(6) and not w29437;
w29507 <= not w29431 and w29506;
w29508 <= not w29439 and not w29507;
w29509 <= not w29505 and w29508;
w29510 <= not w29439 and not w29509;
w29511 <= b(7) and not w29428;
w29512 <= not w29422 and w29511;
w29513 <= not w29430 and not w29512;
w29514 <= not w29510 and w29513;
w29515 <= not w29430 and not w29514;
w29516 <= b(8) and not w29419;
w29517 <= not w29413 and w29516;
w29518 <= not w29421 and not w29517;
w29519 <= not w29515 and w29518;
w29520 <= not w29421 and not w29519;
w29521 <= b(9) and not w29410;
w29522 <= not w29404 and w29521;
w29523 <= not w29412 and not w29522;
w29524 <= not w29520 and w29523;
w29525 <= not w29412 and not w29524;
w29526 <= b(10) and not w29401;
w29527 <= not w29395 and w29526;
w29528 <= not w29403 and not w29527;
w29529 <= not w29525 and w29528;
w29530 <= not w29403 and not w29529;
w29531 <= not w29273 and not w29394;
w29532 <= not w29275 and w29391;
w29533 <= not w29387 and w29532;
w29534 <= not w29388 and not w29391;
w29535 <= not w29533 and not w29534;
w29536 <= w29394 and not w29535;
w29537 <= not w29531 and not w29536;
w29538 <= not b(11) and not w29537;
w29539 <= b(11) and not w29531;
w29540 <= not w29536 and w29539;
w29541 <= w1195 and not w29540;
w29542 <= not w29538 and w29541;
w29543 <= not w29530 and w29542;
w29544 <= w1037 and not w29537;
w29545 <= not w29543 and not w29544;
w29546 <= not w29412 and w29528;
w29547 <= not w29524 and w29546;
w29548 <= not w29525 and not w29528;
w29549 <= not w29547 and not w29548;
w29550 <= not w29545 and not w29549;
w29551 <= not w29402 and not w29544;
w29552 <= not w29543 and w29551;
w29553 <= not w29550 and not w29552;
w29554 <= not w29403 and not w29540;
w29555 <= not w29538 and w29554;
w29556 <= not w29529 and w29555;
w29557 <= not w29538 and not w29540;
w29558 <= not w29530 and not w29557;
w29559 <= not w29556 and not w29558;
w29560 <= not w29545 and not w29559;
w29561 <= not w29537 and not w29544;
w29562 <= not w29543 and w29561;
w29563 <= not w29560 and not w29562;
w29564 <= not b(12) and not w29563;
w29565 <= not b(11) and not w29553;
w29566 <= not w29421 and w29523;
w29567 <= not w29519 and w29566;
w29568 <= not w29520 and not w29523;
w29569 <= not w29567 and not w29568;
w29570 <= not w29545 and not w29569;
w29571 <= not w29411 and not w29544;
w29572 <= not w29543 and w29571;
w29573 <= not w29570 and not w29572;
w29574 <= not b(10) and not w29573;
w29575 <= not w29430 and w29518;
w29576 <= not w29514 and w29575;
w29577 <= not w29515 and not w29518;
w29578 <= not w29576 and not w29577;
w29579 <= not w29545 and not w29578;
w29580 <= not w29420 and not w29544;
w29581 <= not w29543 and w29580;
w29582 <= not w29579 and not w29581;
w29583 <= not b(9) and not w29582;
w29584 <= not w29439 and w29513;
w29585 <= not w29509 and w29584;
w29586 <= not w29510 and not w29513;
w29587 <= not w29585 and not w29586;
w29588 <= not w29545 and not w29587;
w29589 <= not w29429 and not w29544;
w29590 <= not w29543 and w29589;
w29591 <= not w29588 and not w29590;
w29592 <= not b(8) and not w29591;
w29593 <= not w29448 and w29508;
w29594 <= not w29504 and w29593;
w29595 <= not w29505 and not w29508;
w29596 <= not w29594 and not w29595;
w29597 <= not w29545 and not w29596;
w29598 <= not w29438 and not w29544;
w29599 <= not w29543 and w29598;
w29600 <= not w29597 and not w29599;
w29601 <= not b(7) and not w29600;
w29602 <= not w29457 and w29503;
w29603 <= not w29499 and w29602;
w29604 <= not w29500 and not w29503;
w29605 <= not w29603 and not w29604;
w29606 <= not w29545 and not w29605;
w29607 <= not w29447 and not w29544;
w29608 <= not w29543 and w29607;
w29609 <= not w29606 and not w29608;
w29610 <= not b(6) and not w29609;
w29611 <= not w29466 and w29498;
w29612 <= not w29494 and w29611;
w29613 <= not w29495 and not w29498;
w29614 <= not w29612 and not w29613;
w29615 <= not w29545 and not w29614;
w29616 <= not w29456 and not w29544;
w29617 <= not w29543 and w29616;
w29618 <= not w29615 and not w29617;
w29619 <= not b(5) and not w29618;
w29620 <= not w29474 and w29493;
w29621 <= not w29489 and w29620;
w29622 <= not w29490 and not w29493;
w29623 <= not w29621 and not w29622;
w29624 <= not w29545 and not w29623;
w29625 <= not w29465 and not w29544;
w29626 <= not w29543 and w29625;
w29627 <= not w29624 and not w29626;
w29628 <= not b(4) and not w29627;
w29629 <= not w29484 and w29488;
w29630 <= not w29483 and w29629;
w29631 <= not w29485 and not w29488;
w29632 <= not w29630 and not w29631;
w29633 <= not w29545 and not w29632;
w29634 <= not w29473 and not w29544;
w29635 <= not w29543 and w29634;
w29636 <= not w29633 and not w29635;
w29637 <= not b(3) and not w29636;
w29638 <= w1135 and not w29481;
w29639 <= not w29479 and w29638;
w29640 <= not w29483 and not w29639;
w29641 <= not w29545 and w29640;
w29642 <= not w29478 and not w29544;
w29643 <= not w29543 and w29642;
w29644 <= not w29641 and not w29643;
w29645 <= not b(2) and not w29644;
w29646 <= b(0) and not w29545;
w29647 <= a(52) and not w29646;
w29648 <= w1135 and not w29545;
w29649 <= not w29647 and not w29648;
w29650 <= b(1) and not w29649;
w29651 <= not b(1) and not w29648;
w29652 <= not w29647 and w29651;
w29653 <= not w29650 and not w29652;
w29654 <= not w1309 and not w29653;
w29655 <= not b(1) and not w29649;
w29656 <= not w29654 and not w29655;
w29657 <= b(2) and not w29643;
w29658 <= not w29641 and w29657;
w29659 <= not w29645 and not w29658;
w29660 <= not w29656 and w29659;
w29661 <= not w29645 and not w29660;
w29662 <= b(3) and not w29635;
w29663 <= not w29633 and w29662;
w29664 <= not w29637 and not w29663;
w29665 <= not w29661 and w29664;
w29666 <= not w29637 and not w29665;
w29667 <= b(4) and not w29626;
w29668 <= not w29624 and w29667;
w29669 <= not w29628 and not w29668;
w29670 <= not w29666 and w29669;
w29671 <= not w29628 and not w29670;
w29672 <= b(5) and not w29617;
w29673 <= not w29615 and w29672;
w29674 <= not w29619 and not w29673;
w29675 <= not w29671 and w29674;
w29676 <= not w29619 and not w29675;
w29677 <= b(6) and not w29608;
w29678 <= not w29606 and w29677;
w29679 <= not w29610 and not w29678;
w29680 <= not w29676 and w29679;
w29681 <= not w29610 and not w29680;
w29682 <= b(7) and not w29599;
w29683 <= not w29597 and w29682;
w29684 <= not w29601 and not w29683;
w29685 <= not w29681 and w29684;
w29686 <= not w29601 and not w29685;
w29687 <= b(8) and not w29590;
w29688 <= not w29588 and w29687;
w29689 <= not w29592 and not w29688;
w29690 <= not w29686 and w29689;
w29691 <= not w29592 and not w29690;
w29692 <= b(9) and not w29581;
w29693 <= not w29579 and w29692;
w29694 <= not w29583 and not w29693;
w29695 <= not w29691 and w29694;
w29696 <= not w29583 and not w29695;
w29697 <= b(10) and not w29572;
w29698 <= not w29570 and w29697;
w29699 <= not w29574 and not w29698;
w29700 <= not w29696 and w29699;
w29701 <= not w29574 and not w29700;
w29702 <= b(11) and not w29552;
w29703 <= not w29550 and w29702;
w29704 <= not w29565 and not w29703;
w29705 <= not w29701 and w29704;
w29706 <= not w29565 and not w29705;
w29707 <= b(12) and not w29562;
w29708 <= not w29560 and w29707;
w29709 <= not w29564 and not w29708;
w29710 <= not w29706 and w29709;
w29711 <= not w29564 and not w29710;
w29712 <= w1369 and not w29711;
w29713 <= not w29553 and not w29712;
w29714 <= not w29574 and w29704;
w29715 <= not w29700 and w29714;
w29716 <= not w29701 and not w29704;
w29717 <= not w29715 and not w29716;
w29718 <= w1369 and not w29717;
w29719 <= not w29711 and w29718;
w29720 <= not w29713 and not w29719;
w29721 <= not w29563 and not w29712;
w29722 <= not w29565 and w29709;
w29723 <= not w29705 and w29722;
w29724 <= not w29706 and not w29709;
w29725 <= not w29723 and not w29724;
w29726 <= w29712 and not w29725;
w29727 <= not w29721 and not w29726;
w29728 <= not b(13) and not w29727;
w29729 <= not b(12) and not w29720;
w29730 <= not w29573 and not w29712;
w29731 <= not w29583 and w29699;
w29732 <= not w29695 and w29731;
w29733 <= not w29696 and not w29699;
w29734 <= not w29732 and not w29733;
w29735 <= w1369 and not w29734;
w29736 <= not w29711 and w29735;
w29737 <= not w29730 and not w29736;
w29738 <= not b(11) and not w29737;
w29739 <= not w29582 and not w29712;
w29740 <= not w29592 and w29694;
w29741 <= not w29690 and w29740;
w29742 <= not w29691 and not w29694;
w29743 <= not w29741 and not w29742;
w29744 <= w1369 and not w29743;
w29745 <= not w29711 and w29744;
w29746 <= not w29739 and not w29745;
w29747 <= not b(10) and not w29746;
w29748 <= not w29591 and not w29712;
w29749 <= not w29601 and w29689;
w29750 <= not w29685 and w29749;
w29751 <= not w29686 and not w29689;
w29752 <= not w29750 and not w29751;
w29753 <= w1369 and not w29752;
w29754 <= not w29711 and w29753;
w29755 <= not w29748 and not w29754;
w29756 <= not b(9) and not w29755;
w29757 <= not w29600 and not w29712;
w29758 <= not w29610 and w29684;
w29759 <= not w29680 and w29758;
w29760 <= not w29681 and not w29684;
w29761 <= not w29759 and not w29760;
w29762 <= w1369 and not w29761;
w29763 <= not w29711 and w29762;
w29764 <= not w29757 and not w29763;
w29765 <= not b(8) and not w29764;
w29766 <= not w29609 and not w29712;
w29767 <= not w29619 and w29679;
w29768 <= not w29675 and w29767;
w29769 <= not w29676 and not w29679;
w29770 <= not w29768 and not w29769;
w29771 <= w1369 and not w29770;
w29772 <= not w29711 and w29771;
w29773 <= not w29766 and not w29772;
w29774 <= not b(7) and not w29773;
w29775 <= not w29618 and not w29712;
w29776 <= not w29628 and w29674;
w29777 <= not w29670 and w29776;
w29778 <= not w29671 and not w29674;
w29779 <= not w29777 and not w29778;
w29780 <= w1369 and not w29779;
w29781 <= not w29711 and w29780;
w29782 <= not w29775 and not w29781;
w29783 <= not b(6) and not w29782;
w29784 <= not w29627 and not w29712;
w29785 <= not w29637 and w29669;
w29786 <= not w29665 and w29785;
w29787 <= not w29666 and not w29669;
w29788 <= not w29786 and not w29787;
w29789 <= w1369 and not w29788;
w29790 <= not w29711 and w29789;
w29791 <= not w29784 and not w29790;
w29792 <= not b(5) and not w29791;
w29793 <= not w29636 and not w29712;
w29794 <= not w29645 and w29664;
w29795 <= not w29660 and w29794;
w29796 <= not w29661 and not w29664;
w29797 <= not w29795 and not w29796;
w29798 <= w1369 and not w29797;
w29799 <= not w29711 and w29798;
w29800 <= not w29793 and not w29799;
w29801 <= not b(4) and not w29800;
w29802 <= not w29644 and not w29712;
w29803 <= not w29655 and w29659;
w29804 <= not w29654 and w29803;
w29805 <= not w29656 and not w29659;
w29806 <= not w29804 and not w29805;
w29807 <= w1369 and not w29806;
w29808 <= not w29711 and w29807;
w29809 <= not w29802 and not w29808;
w29810 <= not b(3) and not w29809;
w29811 <= not w29649 and not w29712;
w29812 <= w1309 and not w29652;
w29813 <= not w29650 and w29812;
w29814 <= w1369 and not w29813;
w29815 <= not w29654 and w29814;
w29816 <= not w29711 and w29815;
w29817 <= not w29811 and not w29816;
w29818 <= not b(2) and not w29817;
w29819 <= w1481 and not w29711;
w29820 <= a(51) and not w29819;
w29821 <= w1486 and not w29711;
w29822 <= not w29820 and not w29821;
w29823 <= b(1) and not w29822;
w29824 <= not b(1) and not w29821;
w29825 <= not w29820 and w29824;
w29826 <= not w29823 and not w29825;
w29827 <= not w1493 and not w29826;
w29828 <= not b(1) and not w29822;
w29829 <= not w29827 and not w29828;
w29830 <= b(2) and not w29816;
w29831 <= not w29811 and w29830;
w29832 <= not w29818 and not w29831;
w29833 <= not w29829 and w29832;
w29834 <= not w29818 and not w29833;
w29835 <= b(3) and not w29808;
w29836 <= not w29802 and w29835;
w29837 <= not w29810 and not w29836;
w29838 <= not w29834 and w29837;
w29839 <= not w29810 and not w29838;
w29840 <= b(4) and not w29799;
w29841 <= not w29793 and w29840;
w29842 <= not w29801 and not w29841;
w29843 <= not w29839 and w29842;
w29844 <= not w29801 and not w29843;
w29845 <= b(5) and not w29790;
w29846 <= not w29784 and w29845;
w29847 <= not w29792 and not w29846;
w29848 <= not w29844 and w29847;
w29849 <= not w29792 and not w29848;
w29850 <= b(6) and not w29781;
w29851 <= not w29775 and w29850;
w29852 <= not w29783 and not w29851;
w29853 <= not w29849 and w29852;
w29854 <= not w29783 and not w29853;
w29855 <= b(7) and not w29772;
w29856 <= not w29766 and w29855;
w29857 <= not w29774 and not w29856;
w29858 <= not w29854 and w29857;
w29859 <= not w29774 and not w29858;
w29860 <= b(8) and not w29763;
w29861 <= not w29757 and w29860;
w29862 <= not w29765 and not w29861;
w29863 <= not w29859 and w29862;
w29864 <= not w29765 and not w29863;
w29865 <= b(9) and not w29754;
w29866 <= not w29748 and w29865;
w29867 <= not w29756 and not w29866;
w29868 <= not w29864 and w29867;
w29869 <= not w29756 and not w29868;
w29870 <= b(10) and not w29745;
w29871 <= not w29739 and w29870;
w29872 <= not w29747 and not w29871;
w29873 <= not w29869 and w29872;
w29874 <= not w29747 and not w29873;
w29875 <= b(11) and not w29736;
w29876 <= not w29730 and w29875;
w29877 <= not w29738 and not w29876;
w29878 <= not w29874 and w29877;
w29879 <= not w29738 and not w29878;
w29880 <= b(12) and not w29719;
w29881 <= not w29713 and w29880;
w29882 <= not w29729 and not w29881;
w29883 <= not w29879 and w29882;
w29884 <= not w29729 and not w29883;
w29885 <= b(13) and not w29721;
w29886 <= not w29726 and w29885;
w29887 <= not w29728 and not w29886;
w29888 <= not w29884 and w29887;
w29889 <= not w29728 and not w29888;
w29890 <= w1559 and not w29889;
w29891 <= not w29720 and not w29890;
w29892 <= not w29738 and w29882;
w29893 <= not w29878 and w29892;
w29894 <= not w29879 and not w29882;
w29895 <= not w29893 and not w29894;
w29896 <= w1559 and not w29895;
w29897 <= not w29889 and w29896;
w29898 <= not w29891 and not w29897;
w29899 <= not b(13) and not w29898;
w29900 <= not w29737 and not w29890;
w29901 <= not w29747 and w29877;
w29902 <= not w29873 and w29901;
w29903 <= not w29874 and not w29877;
w29904 <= not w29902 and not w29903;
w29905 <= w1559 and not w29904;
w29906 <= not w29889 and w29905;
w29907 <= not w29900 and not w29906;
w29908 <= not b(12) and not w29907;
w29909 <= not w29746 and not w29890;
w29910 <= not w29756 and w29872;
w29911 <= not w29868 and w29910;
w29912 <= not w29869 and not w29872;
w29913 <= not w29911 and not w29912;
w29914 <= w1559 and not w29913;
w29915 <= not w29889 and w29914;
w29916 <= not w29909 and not w29915;
w29917 <= not b(11) and not w29916;
w29918 <= not w29755 and not w29890;
w29919 <= not w29765 and w29867;
w29920 <= not w29863 and w29919;
w29921 <= not w29864 and not w29867;
w29922 <= not w29920 and not w29921;
w29923 <= w1559 and not w29922;
w29924 <= not w29889 and w29923;
w29925 <= not w29918 and not w29924;
w29926 <= not b(10) and not w29925;
w29927 <= not w29764 and not w29890;
w29928 <= not w29774 and w29862;
w29929 <= not w29858 and w29928;
w29930 <= not w29859 and not w29862;
w29931 <= not w29929 and not w29930;
w29932 <= w1559 and not w29931;
w29933 <= not w29889 and w29932;
w29934 <= not w29927 and not w29933;
w29935 <= not b(9) and not w29934;
w29936 <= not w29773 and not w29890;
w29937 <= not w29783 and w29857;
w29938 <= not w29853 and w29937;
w29939 <= not w29854 and not w29857;
w29940 <= not w29938 and not w29939;
w29941 <= w1559 and not w29940;
w29942 <= not w29889 and w29941;
w29943 <= not w29936 and not w29942;
w29944 <= not b(8) and not w29943;
w29945 <= not w29782 and not w29890;
w29946 <= not w29792 and w29852;
w29947 <= not w29848 and w29946;
w29948 <= not w29849 and not w29852;
w29949 <= not w29947 and not w29948;
w29950 <= w1559 and not w29949;
w29951 <= not w29889 and w29950;
w29952 <= not w29945 and not w29951;
w29953 <= not b(7) and not w29952;
w29954 <= not w29791 and not w29890;
w29955 <= not w29801 and w29847;
w29956 <= not w29843 and w29955;
w29957 <= not w29844 and not w29847;
w29958 <= not w29956 and not w29957;
w29959 <= w1559 and not w29958;
w29960 <= not w29889 and w29959;
w29961 <= not w29954 and not w29960;
w29962 <= not b(6) and not w29961;
w29963 <= not w29800 and not w29890;
w29964 <= not w29810 and w29842;
w29965 <= not w29838 and w29964;
w29966 <= not w29839 and not w29842;
w29967 <= not w29965 and not w29966;
w29968 <= w1559 and not w29967;
w29969 <= not w29889 and w29968;
w29970 <= not w29963 and not w29969;
w29971 <= not b(5) and not w29970;
w29972 <= not w29809 and not w29890;
w29973 <= not w29818 and w29837;
w29974 <= not w29833 and w29973;
w29975 <= not w29834 and not w29837;
w29976 <= not w29974 and not w29975;
w29977 <= w1559 and not w29976;
w29978 <= not w29889 and w29977;
w29979 <= not w29972 and not w29978;
w29980 <= not b(4) and not w29979;
w29981 <= not w29817 and not w29890;
w29982 <= not w29828 and w29832;
w29983 <= not w29827 and w29982;
w29984 <= not w29829 and not w29832;
w29985 <= not w29983 and not w29984;
w29986 <= w1559 and not w29985;
w29987 <= not w29889 and w29986;
w29988 <= not w29981 and not w29987;
w29989 <= not b(3) and not w29988;
w29990 <= not w29822 and not w29890;
w29991 <= w1493 and not w29825;
w29992 <= not w29823 and w29991;
w29993 <= w1559 and not w29992;
w29994 <= not w29827 and w29993;
w29995 <= not w29889 and w29994;
w29996 <= not w29990 and not w29995;
w29997 <= not b(2) and not w29996;
w29998 <= w1672 and not w29889;
w29999 <= a(50) and not w29998;
w30000 <= w1678 and not w29889;
w30001 <= not w29999 and not w30000;
w30002 <= b(1) and not w30001;
w30003 <= not b(1) and not w30000;
w30004 <= not w29999 and w30003;
w30005 <= not w30002 and not w30004;
w30006 <= not w1685 and not w30005;
w30007 <= not b(1) and not w30001;
w30008 <= not w30006 and not w30007;
w30009 <= b(2) and not w29995;
w30010 <= not w29990 and w30009;
w30011 <= not w29997 and not w30010;
w30012 <= not w30008 and w30011;
w30013 <= not w29997 and not w30012;
w30014 <= b(3) and not w29987;
w30015 <= not w29981 and w30014;
w30016 <= not w29989 and not w30015;
w30017 <= not w30013 and w30016;
w30018 <= not w29989 and not w30017;
w30019 <= b(4) and not w29978;
w30020 <= not w29972 and w30019;
w30021 <= not w29980 and not w30020;
w30022 <= not w30018 and w30021;
w30023 <= not w29980 and not w30022;
w30024 <= b(5) and not w29969;
w30025 <= not w29963 and w30024;
w30026 <= not w29971 and not w30025;
w30027 <= not w30023 and w30026;
w30028 <= not w29971 and not w30027;
w30029 <= b(6) and not w29960;
w30030 <= not w29954 and w30029;
w30031 <= not w29962 and not w30030;
w30032 <= not w30028 and w30031;
w30033 <= not w29962 and not w30032;
w30034 <= b(7) and not w29951;
w30035 <= not w29945 and w30034;
w30036 <= not w29953 and not w30035;
w30037 <= not w30033 and w30036;
w30038 <= not w29953 and not w30037;
w30039 <= b(8) and not w29942;
w30040 <= not w29936 and w30039;
w30041 <= not w29944 and not w30040;
w30042 <= not w30038 and w30041;
w30043 <= not w29944 and not w30042;
w30044 <= b(9) and not w29933;
w30045 <= not w29927 and w30044;
w30046 <= not w29935 and not w30045;
w30047 <= not w30043 and w30046;
w30048 <= not w29935 and not w30047;
w30049 <= b(10) and not w29924;
w30050 <= not w29918 and w30049;
w30051 <= not w29926 and not w30050;
w30052 <= not w30048 and w30051;
w30053 <= not w29926 and not w30052;
w30054 <= b(11) and not w29915;
w30055 <= not w29909 and w30054;
w30056 <= not w29917 and not w30055;
w30057 <= not w30053 and w30056;
w30058 <= not w29917 and not w30057;
w30059 <= b(12) and not w29906;
w30060 <= not w29900 and w30059;
w30061 <= not w29908 and not w30060;
w30062 <= not w30058 and w30061;
w30063 <= not w29908 and not w30062;
w30064 <= b(13) and not w29897;
w30065 <= not w29891 and w30064;
w30066 <= not w29899 and not w30065;
w30067 <= not w30063 and w30066;
w30068 <= not w29899 and not w30067;
w30069 <= not w29727 and not w29890;
w30070 <= not w29729 and w29887;
w30071 <= not w29883 and w30070;
w30072 <= not w29884 and not w29887;
w30073 <= not w30071 and not w30072;
w30074 <= w29890 and not w30073;
w30075 <= not w30069 and not w30074;
w30076 <= not b(14) and not w30075;
w30077 <= b(14) and not w30069;
w30078 <= not w30074 and w30077;
w30079 <= w1761 and not w30078;
w30080 <= not w30076 and w30079;
w30081 <= not w30068 and w30080;
w30082 <= w1559 and not w30075;
w30083 <= not w30081 and not w30082;
w30084 <= not w29908 and w30066;
w30085 <= not w30062 and w30084;
w30086 <= not w30063 and not w30066;
w30087 <= not w30085 and not w30086;
w30088 <= not w30083 and not w30087;
w30089 <= not w29898 and not w30082;
w30090 <= not w30081 and w30089;
w30091 <= not w30088 and not w30090;
w30092 <= not w29899 and not w30078;
w30093 <= not w30076 and w30092;
w30094 <= not w30067 and w30093;
w30095 <= not w30076 and not w30078;
w30096 <= not w30068 and not w30095;
w30097 <= not w30094 and not w30096;
w30098 <= not w30083 and not w30097;
w30099 <= not w30075 and not w30082;
w30100 <= not w30081 and w30099;
w30101 <= not w30098 and not w30100;
w30102 <= not b(15) and not w30101;
w30103 <= not b(14) and not w30091;
w30104 <= not w29917 and w30061;
w30105 <= not w30057 and w30104;
w30106 <= not w30058 and not w30061;
w30107 <= not w30105 and not w30106;
w30108 <= not w30083 and not w30107;
w30109 <= not w29907 and not w30082;
w30110 <= not w30081 and w30109;
w30111 <= not w30108 and not w30110;
w30112 <= not b(13) and not w30111;
w30113 <= not w29926 and w30056;
w30114 <= not w30052 and w30113;
w30115 <= not w30053 and not w30056;
w30116 <= not w30114 and not w30115;
w30117 <= not w30083 and not w30116;
w30118 <= not w29916 and not w30082;
w30119 <= not w30081 and w30118;
w30120 <= not w30117 and not w30119;
w30121 <= not b(12) and not w30120;
w30122 <= not w29935 and w30051;
w30123 <= not w30047 and w30122;
w30124 <= not w30048 and not w30051;
w30125 <= not w30123 and not w30124;
w30126 <= not w30083 and not w30125;
w30127 <= not w29925 and not w30082;
w30128 <= not w30081 and w30127;
w30129 <= not w30126 and not w30128;
w30130 <= not b(11) and not w30129;
w30131 <= not w29944 and w30046;
w30132 <= not w30042 and w30131;
w30133 <= not w30043 and not w30046;
w30134 <= not w30132 and not w30133;
w30135 <= not w30083 and not w30134;
w30136 <= not w29934 and not w30082;
w30137 <= not w30081 and w30136;
w30138 <= not w30135 and not w30137;
w30139 <= not b(10) and not w30138;
w30140 <= not w29953 and w30041;
w30141 <= not w30037 and w30140;
w30142 <= not w30038 and not w30041;
w30143 <= not w30141 and not w30142;
w30144 <= not w30083 and not w30143;
w30145 <= not w29943 and not w30082;
w30146 <= not w30081 and w30145;
w30147 <= not w30144 and not w30146;
w30148 <= not b(9) and not w30147;
w30149 <= not w29962 and w30036;
w30150 <= not w30032 and w30149;
w30151 <= not w30033 and not w30036;
w30152 <= not w30150 and not w30151;
w30153 <= not w30083 and not w30152;
w30154 <= not w29952 and not w30082;
w30155 <= not w30081 and w30154;
w30156 <= not w30153 and not w30155;
w30157 <= not b(8) and not w30156;
w30158 <= not w29971 and w30031;
w30159 <= not w30027 and w30158;
w30160 <= not w30028 and not w30031;
w30161 <= not w30159 and not w30160;
w30162 <= not w30083 and not w30161;
w30163 <= not w29961 and not w30082;
w30164 <= not w30081 and w30163;
w30165 <= not w30162 and not w30164;
w30166 <= not b(7) and not w30165;
w30167 <= not w29980 and w30026;
w30168 <= not w30022 and w30167;
w30169 <= not w30023 and not w30026;
w30170 <= not w30168 and not w30169;
w30171 <= not w30083 and not w30170;
w30172 <= not w29970 and not w30082;
w30173 <= not w30081 and w30172;
w30174 <= not w30171 and not w30173;
w30175 <= not b(6) and not w30174;
w30176 <= not w29989 and w30021;
w30177 <= not w30017 and w30176;
w30178 <= not w30018 and not w30021;
w30179 <= not w30177 and not w30178;
w30180 <= not w30083 and not w30179;
w30181 <= not w29979 and not w30082;
w30182 <= not w30081 and w30181;
w30183 <= not w30180 and not w30182;
w30184 <= not b(5) and not w30183;
w30185 <= not w29997 and w30016;
w30186 <= not w30012 and w30185;
w30187 <= not w30013 and not w30016;
w30188 <= not w30186 and not w30187;
w30189 <= not w30083 and not w30188;
w30190 <= not w29988 and not w30082;
w30191 <= not w30081 and w30190;
w30192 <= not w30189 and not w30191;
w30193 <= not b(4) and not w30192;
w30194 <= not w30007 and w30011;
w30195 <= not w30006 and w30194;
w30196 <= not w30008 and not w30011;
w30197 <= not w30195 and not w30196;
w30198 <= not w30083 and not w30197;
w30199 <= not w29996 and not w30082;
w30200 <= not w30081 and w30199;
w30201 <= not w30198 and not w30200;
w30202 <= not b(3) and not w30201;
w30203 <= w1685 and not w30004;
w30204 <= not w30002 and w30203;
w30205 <= not w30006 and not w30204;
w30206 <= not w30083 and w30205;
w30207 <= not w30001 and not w30082;
w30208 <= not w30081 and w30207;
w30209 <= not w30206 and not w30208;
w30210 <= not b(2) and not w30209;
w30211 <= b(0) and not w30083;
w30212 <= a(49) and not w30211;
w30213 <= w1685 and not w30083;
w30214 <= not w30212 and not w30213;
w30215 <= b(1) and not w30214;
w30216 <= not b(1) and not w30213;
w30217 <= not w30212 and w30216;
w30218 <= not w30215 and not w30217;
w30219 <= not w1902 and not w30218;
w30220 <= not b(1) and not w30214;
w30221 <= not w30219 and not w30220;
w30222 <= b(2) and not w30208;
w30223 <= not w30206 and w30222;
w30224 <= not w30210 and not w30223;
w30225 <= not w30221 and w30224;
w30226 <= not w30210 and not w30225;
w30227 <= b(3) and not w30200;
w30228 <= not w30198 and w30227;
w30229 <= not w30202 and not w30228;
w30230 <= not w30226 and w30229;
w30231 <= not w30202 and not w30230;
w30232 <= b(4) and not w30191;
w30233 <= not w30189 and w30232;
w30234 <= not w30193 and not w30233;
w30235 <= not w30231 and w30234;
w30236 <= not w30193 and not w30235;
w30237 <= b(5) and not w30182;
w30238 <= not w30180 and w30237;
w30239 <= not w30184 and not w30238;
w30240 <= not w30236 and w30239;
w30241 <= not w30184 and not w30240;
w30242 <= b(6) and not w30173;
w30243 <= not w30171 and w30242;
w30244 <= not w30175 and not w30243;
w30245 <= not w30241 and w30244;
w30246 <= not w30175 and not w30245;
w30247 <= b(7) and not w30164;
w30248 <= not w30162 and w30247;
w30249 <= not w30166 and not w30248;
w30250 <= not w30246 and w30249;
w30251 <= not w30166 and not w30250;
w30252 <= b(8) and not w30155;
w30253 <= not w30153 and w30252;
w30254 <= not w30157 and not w30253;
w30255 <= not w30251 and w30254;
w30256 <= not w30157 and not w30255;
w30257 <= b(9) and not w30146;
w30258 <= not w30144 and w30257;
w30259 <= not w30148 and not w30258;
w30260 <= not w30256 and w30259;
w30261 <= not w30148 and not w30260;
w30262 <= b(10) and not w30137;
w30263 <= not w30135 and w30262;
w30264 <= not w30139 and not w30263;
w30265 <= not w30261 and w30264;
w30266 <= not w30139 and not w30265;
w30267 <= b(11) and not w30128;
w30268 <= not w30126 and w30267;
w30269 <= not w30130 and not w30268;
w30270 <= not w30266 and w30269;
w30271 <= not w30130 and not w30270;
w30272 <= b(12) and not w30119;
w30273 <= not w30117 and w30272;
w30274 <= not w30121 and not w30273;
w30275 <= not w30271 and w30274;
w30276 <= not w30121 and not w30275;
w30277 <= b(13) and not w30110;
w30278 <= not w30108 and w30277;
w30279 <= not w30112 and not w30278;
w30280 <= not w30276 and w30279;
w30281 <= not w30112 and not w30280;
w30282 <= b(14) and not w30090;
w30283 <= not w30088 and w30282;
w30284 <= not w30103 and not w30283;
w30285 <= not w30281 and w30284;
w30286 <= not w30103 and not w30285;
w30287 <= b(15) and not w30100;
w30288 <= not w30098 and w30287;
w30289 <= not w30102 and not w30288;
w30290 <= not w30286 and w30289;
w30291 <= not w30102 and not w30290;
w30292 <= w89 and not w30291;
w30293 <= not w30091 and not w30292;
w30294 <= not w30112 and w30284;
w30295 <= not w30280 and w30294;
w30296 <= not w30281 and not w30284;
w30297 <= not w30295 and not w30296;
w30298 <= w89 and not w30297;
w30299 <= not w30291 and w30298;
w30300 <= not w30293 and not w30299;
w30301 <= not w30101 and not w30292;
w30302 <= not w30103 and w30289;
w30303 <= not w30285 and w30302;
w30304 <= not w30286 and not w30289;
w30305 <= not w30303 and not w30304;
w30306 <= w30292 and not w30305;
w30307 <= not w30301 and not w30306;
w30308 <= not b(16) and not w30307;
w30309 <= not b(15) and not w30300;
w30310 <= not w30111 and not w30292;
w30311 <= not w30121 and w30279;
w30312 <= not w30275 and w30311;
w30313 <= not w30276 and not w30279;
w30314 <= not w30312 and not w30313;
w30315 <= w89 and not w30314;
w30316 <= not w30291 and w30315;
w30317 <= not w30310 and not w30316;
w30318 <= not b(14) and not w30317;
w30319 <= not w30120 and not w30292;
w30320 <= not w30130 and w30274;
w30321 <= not w30270 and w30320;
w30322 <= not w30271 and not w30274;
w30323 <= not w30321 and not w30322;
w30324 <= w89 and not w30323;
w30325 <= not w30291 and w30324;
w30326 <= not w30319 and not w30325;
w30327 <= not b(13) and not w30326;
w30328 <= not w30129 and not w30292;
w30329 <= not w30139 and w30269;
w30330 <= not w30265 and w30329;
w30331 <= not w30266 and not w30269;
w30332 <= not w30330 and not w30331;
w30333 <= w89 and not w30332;
w30334 <= not w30291 and w30333;
w30335 <= not w30328 and not w30334;
w30336 <= not b(12) and not w30335;
w30337 <= not w30138 and not w30292;
w30338 <= not w30148 and w30264;
w30339 <= not w30260 and w30338;
w30340 <= not w30261 and not w30264;
w30341 <= not w30339 and not w30340;
w30342 <= w89 and not w30341;
w30343 <= not w30291 and w30342;
w30344 <= not w30337 and not w30343;
w30345 <= not b(11) and not w30344;
w30346 <= not w30147 and not w30292;
w30347 <= not w30157 and w30259;
w30348 <= not w30255 and w30347;
w30349 <= not w30256 and not w30259;
w30350 <= not w30348 and not w30349;
w30351 <= w89 and not w30350;
w30352 <= not w30291 and w30351;
w30353 <= not w30346 and not w30352;
w30354 <= not b(10) and not w30353;
w30355 <= not w30156 and not w30292;
w30356 <= not w30166 and w30254;
w30357 <= not w30250 and w30356;
w30358 <= not w30251 and not w30254;
w30359 <= not w30357 and not w30358;
w30360 <= w89 and not w30359;
w30361 <= not w30291 and w30360;
w30362 <= not w30355 and not w30361;
w30363 <= not b(9) and not w30362;
w30364 <= not w30165 and not w30292;
w30365 <= not w30175 and w30249;
w30366 <= not w30245 and w30365;
w30367 <= not w30246 and not w30249;
w30368 <= not w30366 and not w30367;
w30369 <= w89 and not w30368;
w30370 <= not w30291 and w30369;
w30371 <= not w30364 and not w30370;
w30372 <= not b(8) and not w30371;
w30373 <= not w30174 and not w30292;
w30374 <= not w30184 and w30244;
w30375 <= not w30240 and w30374;
w30376 <= not w30241 and not w30244;
w30377 <= not w30375 and not w30376;
w30378 <= w89 and not w30377;
w30379 <= not w30291 and w30378;
w30380 <= not w30373 and not w30379;
w30381 <= not b(7) and not w30380;
w30382 <= not w30183 and not w30292;
w30383 <= not w30193 and w30239;
w30384 <= not w30235 and w30383;
w30385 <= not w30236 and not w30239;
w30386 <= not w30384 and not w30385;
w30387 <= w89 and not w30386;
w30388 <= not w30291 and w30387;
w30389 <= not w30382 and not w30388;
w30390 <= not b(6) and not w30389;
w30391 <= not w30192 and not w30292;
w30392 <= not w30202 and w30234;
w30393 <= not w30230 and w30392;
w30394 <= not w30231 and not w30234;
w30395 <= not w30393 and not w30394;
w30396 <= w89 and not w30395;
w30397 <= not w30291 and w30396;
w30398 <= not w30391 and not w30397;
w30399 <= not b(5) and not w30398;
w30400 <= not w30201 and not w30292;
w30401 <= not w30210 and w30229;
w30402 <= not w30225 and w30401;
w30403 <= not w30226 and not w30229;
w30404 <= not w30402 and not w30403;
w30405 <= w89 and not w30404;
w30406 <= not w30291 and w30405;
w30407 <= not w30400 and not w30406;
w30408 <= not b(4) and not w30407;
w30409 <= not w30209 and not w30292;
w30410 <= not w30220 and w30224;
w30411 <= not w30219 and w30410;
w30412 <= not w30221 and not w30224;
w30413 <= not w30411 and not w30412;
w30414 <= w89 and not w30413;
w30415 <= not w30291 and w30414;
w30416 <= not w30409 and not w30415;
w30417 <= not b(3) and not w30416;
w30418 <= not w30214 and not w30292;
w30419 <= w1902 and not w30217;
w30420 <= not w30215 and w30419;
w30421 <= w89 and not w30420;
w30422 <= not w30219 and w30421;
w30423 <= not w30291 and w30422;
w30424 <= not w30418 and not w30423;
w30425 <= not b(2) and not w30424;
w30426 <= w2113 and not w30291;
w30427 <= a(48) and not w30426;
w30428 <= w2118 and not w30291;
w30429 <= not w30427 and not w30428;
w30430 <= b(1) and not w30429;
w30431 <= not b(1) and not w30428;
w30432 <= not w30427 and w30431;
w30433 <= not w30430 and not w30432;
w30434 <= not w2125 and not w30433;
w30435 <= not b(1) and not w30429;
w30436 <= not w30434 and not w30435;
w30437 <= b(2) and not w30423;
w30438 <= not w30418 and w30437;
w30439 <= not w30425 and not w30438;
w30440 <= not w30436 and w30439;
w30441 <= not w30425 and not w30440;
w30442 <= b(3) and not w30415;
w30443 <= not w30409 and w30442;
w30444 <= not w30417 and not w30443;
w30445 <= not w30441 and w30444;
w30446 <= not w30417 and not w30445;
w30447 <= b(4) and not w30406;
w30448 <= not w30400 and w30447;
w30449 <= not w30408 and not w30448;
w30450 <= not w30446 and w30449;
w30451 <= not w30408 and not w30450;
w30452 <= b(5) and not w30397;
w30453 <= not w30391 and w30452;
w30454 <= not w30399 and not w30453;
w30455 <= not w30451 and w30454;
w30456 <= not w30399 and not w30455;
w30457 <= b(6) and not w30388;
w30458 <= not w30382 and w30457;
w30459 <= not w30390 and not w30458;
w30460 <= not w30456 and w30459;
w30461 <= not w30390 and not w30460;
w30462 <= b(7) and not w30379;
w30463 <= not w30373 and w30462;
w30464 <= not w30381 and not w30463;
w30465 <= not w30461 and w30464;
w30466 <= not w30381 and not w30465;
w30467 <= b(8) and not w30370;
w30468 <= not w30364 and w30467;
w30469 <= not w30372 and not w30468;
w30470 <= not w30466 and w30469;
w30471 <= not w30372 and not w30470;
w30472 <= b(9) and not w30361;
w30473 <= not w30355 and w30472;
w30474 <= not w30363 and not w30473;
w30475 <= not w30471 and w30474;
w30476 <= not w30363 and not w30475;
w30477 <= b(10) and not w30352;
w30478 <= not w30346 and w30477;
w30479 <= not w30354 and not w30478;
w30480 <= not w30476 and w30479;
w30481 <= not w30354 and not w30480;
w30482 <= b(11) and not w30343;
w30483 <= not w30337 and w30482;
w30484 <= not w30345 and not w30483;
w30485 <= not w30481 and w30484;
w30486 <= not w30345 and not w30485;
w30487 <= b(12) and not w30334;
w30488 <= not w30328 and w30487;
w30489 <= not w30336 and not w30488;
w30490 <= not w30486 and w30489;
w30491 <= not w30336 and not w30490;
w30492 <= b(13) and not w30325;
w30493 <= not w30319 and w30492;
w30494 <= not w30327 and not w30493;
w30495 <= not w30491 and w30494;
w30496 <= not w30327 and not w30495;
w30497 <= b(14) and not w30316;
w30498 <= not w30310 and w30497;
w30499 <= not w30318 and not w30498;
w30500 <= not w30496 and w30499;
w30501 <= not w30318 and not w30500;
w30502 <= b(15) and not w30299;
w30503 <= not w30293 and w30502;
w30504 <= not w30309 and not w30503;
w30505 <= not w30501 and w30504;
w30506 <= not w30309 and not w30505;
w30507 <= b(16) and not w30301;
w30508 <= not w30306 and w30507;
w30509 <= not w30308 and not w30508;
w30510 <= not w30506 and w30509;
w30511 <= not w30308 and not w30510;
w30512 <= w218 and not w30511;
w30513 <= not w30300 and not w30512;
w30514 <= not w30318 and w30504;
w30515 <= not w30500 and w30514;
w30516 <= not w30501 and not w30504;
w30517 <= not w30515 and not w30516;
w30518 <= w218 and not w30517;
w30519 <= not w30511 and w30518;
w30520 <= not w30513 and not w30519;
w30521 <= not b(16) and not w30520;
w30522 <= not w30317 and not w30512;
w30523 <= not w30327 and w30499;
w30524 <= not w30495 and w30523;
w30525 <= not w30496 and not w30499;
w30526 <= not w30524 and not w30525;
w30527 <= w218 and not w30526;
w30528 <= not w30511 and w30527;
w30529 <= not w30522 and not w30528;
w30530 <= not b(15) and not w30529;
w30531 <= not w30326 and not w30512;
w30532 <= not w30336 and w30494;
w30533 <= not w30490 and w30532;
w30534 <= not w30491 and not w30494;
w30535 <= not w30533 and not w30534;
w30536 <= w218 and not w30535;
w30537 <= not w30511 and w30536;
w30538 <= not w30531 and not w30537;
w30539 <= not b(14) and not w30538;
w30540 <= not w30335 and not w30512;
w30541 <= not w30345 and w30489;
w30542 <= not w30485 and w30541;
w30543 <= not w30486 and not w30489;
w30544 <= not w30542 and not w30543;
w30545 <= w218 and not w30544;
w30546 <= not w30511 and w30545;
w30547 <= not w30540 and not w30546;
w30548 <= not b(13) and not w30547;
w30549 <= not w30344 and not w30512;
w30550 <= not w30354 and w30484;
w30551 <= not w30480 and w30550;
w30552 <= not w30481 and not w30484;
w30553 <= not w30551 and not w30552;
w30554 <= w218 and not w30553;
w30555 <= not w30511 and w30554;
w30556 <= not w30549 and not w30555;
w30557 <= not b(12) and not w30556;
w30558 <= not w30353 and not w30512;
w30559 <= not w30363 and w30479;
w30560 <= not w30475 and w30559;
w30561 <= not w30476 and not w30479;
w30562 <= not w30560 and not w30561;
w30563 <= w218 and not w30562;
w30564 <= not w30511 and w30563;
w30565 <= not w30558 and not w30564;
w30566 <= not b(11) and not w30565;
w30567 <= not w30362 and not w30512;
w30568 <= not w30372 and w30474;
w30569 <= not w30470 and w30568;
w30570 <= not w30471 and not w30474;
w30571 <= not w30569 and not w30570;
w30572 <= w218 and not w30571;
w30573 <= not w30511 and w30572;
w30574 <= not w30567 and not w30573;
w30575 <= not b(10) and not w30574;
w30576 <= not w30371 and not w30512;
w30577 <= not w30381 and w30469;
w30578 <= not w30465 and w30577;
w30579 <= not w30466 and not w30469;
w30580 <= not w30578 and not w30579;
w30581 <= w218 and not w30580;
w30582 <= not w30511 and w30581;
w30583 <= not w30576 and not w30582;
w30584 <= not b(9) and not w30583;
w30585 <= not w30380 and not w30512;
w30586 <= not w30390 and w30464;
w30587 <= not w30460 and w30586;
w30588 <= not w30461 and not w30464;
w30589 <= not w30587 and not w30588;
w30590 <= w218 and not w30589;
w30591 <= not w30511 and w30590;
w30592 <= not w30585 and not w30591;
w30593 <= not b(8) and not w30592;
w30594 <= not w30389 and not w30512;
w30595 <= not w30399 and w30459;
w30596 <= not w30455 and w30595;
w30597 <= not w30456 and not w30459;
w30598 <= not w30596 and not w30597;
w30599 <= w218 and not w30598;
w30600 <= not w30511 and w30599;
w30601 <= not w30594 and not w30600;
w30602 <= not b(7) and not w30601;
w30603 <= not w30398 and not w30512;
w30604 <= not w30408 and w30454;
w30605 <= not w30450 and w30604;
w30606 <= not w30451 and not w30454;
w30607 <= not w30605 and not w30606;
w30608 <= w218 and not w30607;
w30609 <= not w30511 and w30608;
w30610 <= not w30603 and not w30609;
w30611 <= not b(6) and not w30610;
w30612 <= not w30407 and not w30512;
w30613 <= not w30417 and w30449;
w30614 <= not w30445 and w30613;
w30615 <= not w30446 and not w30449;
w30616 <= not w30614 and not w30615;
w30617 <= w218 and not w30616;
w30618 <= not w30511 and w30617;
w30619 <= not w30612 and not w30618;
w30620 <= not b(5) and not w30619;
w30621 <= not w30416 and not w30512;
w30622 <= not w30425 and w30444;
w30623 <= not w30440 and w30622;
w30624 <= not w30441 and not w30444;
w30625 <= not w30623 and not w30624;
w30626 <= w218 and not w30625;
w30627 <= not w30511 and w30626;
w30628 <= not w30621 and not w30627;
w30629 <= not b(4) and not w30628;
w30630 <= not w30424 and not w30512;
w30631 <= not w30435 and w30439;
w30632 <= not w30434 and w30631;
w30633 <= not w30436 and not w30439;
w30634 <= not w30632 and not w30633;
w30635 <= w218 and not w30634;
w30636 <= not w30511 and w30635;
w30637 <= not w30630 and not w30636;
w30638 <= not b(3) and not w30637;
w30639 <= not w30429 and not w30512;
w30640 <= w2125 and not w30432;
w30641 <= not w30430 and w30640;
w30642 <= w218 and not w30641;
w30643 <= not w30434 and w30642;
w30644 <= not w30511 and w30643;
w30645 <= not w30639 and not w30644;
w30646 <= not b(2) and not w30645;
w30647 <= w2344 and not w30511;
w30648 <= a(47) and not w30647;
w30649 <= w2349 and not w30511;
w30650 <= not w30648 and not w30649;
w30651 <= b(1) and not w30650;
w30652 <= not b(1) and not w30649;
w30653 <= not w30648 and w30652;
w30654 <= not w30651 and not w30653;
w30655 <= not w2356 and not w30654;
w30656 <= not b(1) and not w30650;
w30657 <= not w30655 and not w30656;
w30658 <= b(2) and not w30644;
w30659 <= not w30639 and w30658;
w30660 <= not w30646 and not w30659;
w30661 <= not w30657 and w30660;
w30662 <= not w30646 and not w30661;
w30663 <= b(3) and not w30636;
w30664 <= not w30630 and w30663;
w30665 <= not w30638 and not w30664;
w30666 <= not w30662 and w30665;
w30667 <= not w30638 and not w30666;
w30668 <= b(4) and not w30627;
w30669 <= not w30621 and w30668;
w30670 <= not w30629 and not w30669;
w30671 <= not w30667 and w30670;
w30672 <= not w30629 and not w30671;
w30673 <= b(5) and not w30618;
w30674 <= not w30612 and w30673;
w30675 <= not w30620 and not w30674;
w30676 <= not w30672 and w30675;
w30677 <= not w30620 and not w30676;
w30678 <= b(6) and not w30609;
w30679 <= not w30603 and w30678;
w30680 <= not w30611 and not w30679;
w30681 <= not w30677 and w30680;
w30682 <= not w30611 and not w30681;
w30683 <= b(7) and not w30600;
w30684 <= not w30594 and w30683;
w30685 <= not w30602 and not w30684;
w30686 <= not w30682 and w30685;
w30687 <= not w30602 and not w30686;
w30688 <= b(8) and not w30591;
w30689 <= not w30585 and w30688;
w30690 <= not w30593 and not w30689;
w30691 <= not w30687 and w30690;
w30692 <= not w30593 and not w30691;
w30693 <= b(9) and not w30582;
w30694 <= not w30576 and w30693;
w30695 <= not w30584 and not w30694;
w30696 <= not w30692 and w30695;
w30697 <= not w30584 and not w30696;
w30698 <= b(10) and not w30573;
w30699 <= not w30567 and w30698;
w30700 <= not w30575 and not w30699;
w30701 <= not w30697 and w30700;
w30702 <= not w30575 and not w30701;
w30703 <= b(11) and not w30564;
w30704 <= not w30558 and w30703;
w30705 <= not w30566 and not w30704;
w30706 <= not w30702 and w30705;
w30707 <= not w30566 and not w30706;
w30708 <= b(12) and not w30555;
w30709 <= not w30549 and w30708;
w30710 <= not w30557 and not w30709;
w30711 <= not w30707 and w30710;
w30712 <= not w30557 and not w30711;
w30713 <= b(13) and not w30546;
w30714 <= not w30540 and w30713;
w30715 <= not w30548 and not w30714;
w30716 <= not w30712 and w30715;
w30717 <= not w30548 and not w30716;
w30718 <= b(14) and not w30537;
w30719 <= not w30531 and w30718;
w30720 <= not w30539 and not w30719;
w30721 <= not w30717 and w30720;
w30722 <= not w30539 and not w30721;
w30723 <= b(15) and not w30528;
w30724 <= not w30522 and w30723;
w30725 <= not w30530 and not w30724;
w30726 <= not w30722 and w30725;
w30727 <= not w30530 and not w30726;
w30728 <= b(16) and not w30519;
w30729 <= not w30513 and w30728;
w30730 <= not w30521 and not w30729;
w30731 <= not w30727 and w30730;
w30732 <= not w30521 and not w30731;
w30733 <= not w30307 and not w30512;
w30734 <= not w30309 and w30509;
w30735 <= not w30505 and w30734;
w30736 <= not w30506 and not w30509;
w30737 <= not w30735 and not w30736;
w30738 <= w30512 and not w30737;
w30739 <= not w30733 and not w30738;
w30740 <= not b(17) and not w30739;
w30741 <= b(17) and not w30733;
w30742 <= not w30738 and w30741;
w30743 <= w2448 and not w30742;
w30744 <= not w30740 and w30743;
w30745 <= not w30732 and w30744;
w30746 <= w218 and not w30739;
w30747 <= not w30745 and not w30746;
w30748 <= not w30530 and w30730;
w30749 <= not w30726 and w30748;
w30750 <= not w30727 and not w30730;
w30751 <= not w30749 and not w30750;
w30752 <= not w30747 and not w30751;
w30753 <= not w30520 and not w30746;
w30754 <= not w30745 and w30753;
w30755 <= not w30752 and not w30754;
w30756 <= not w30521 and not w30742;
w30757 <= not w30740 and w30756;
w30758 <= not w30731 and w30757;
w30759 <= not w30740 and not w30742;
w30760 <= not w30732 and not w30759;
w30761 <= not w30758 and not w30760;
w30762 <= not w30747 and not w30761;
w30763 <= not w30739 and not w30746;
w30764 <= not w30745 and w30763;
w30765 <= not w30762 and not w30764;
w30766 <= not b(18) and not w30765;
w30767 <= not b(17) and not w30755;
w30768 <= not w30539 and w30725;
w30769 <= not w30721 and w30768;
w30770 <= not w30722 and not w30725;
w30771 <= not w30769 and not w30770;
w30772 <= not w30747 and not w30771;
w30773 <= not w30529 and not w30746;
w30774 <= not w30745 and w30773;
w30775 <= not w30772 and not w30774;
w30776 <= not b(16) and not w30775;
w30777 <= not w30548 and w30720;
w30778 <= not w30716 and w30777;
w30779 <= not w30717 and not w30720;
w30780 <= not w30778 and not w30779;
w30781 <= not w30747 and not w30780;
w30782 <= not w30538 and not w30746;
w30783 <= not w30745 and w30782;
w30784 <= not w30781 and not w30783;
w30785 <= not b(15) and not w30784;
w30786 <= not w30557 and w30715;
w30787 <= not w30711 and w30786;
w30788 <= not w30712 and not w30715;
w30789 <= not w30787 and not w30788;
w30790 <= not w30747 and not w30789;
w30791 <= not w30547 and not w30746;
w30792 <= not w30745 and w30791;
w30793 <= not w30790 and not w30792;
w30794 <= not b(14) and not w30793;
w30795 <= not w30566 and w30710;
w30796 <= not w30706 and w30795;
w30797 <= not w30707 and not w30710;
w30798 <= not w30796 and not w30797;
w30799 <= not w30747 and not w30798;
w30800 <= not w30556 and not w30746;
w30801 <= not w30745 and w30800;
w30802 <= not w30799 and not w30801;
w30803 <= not b(13) and not w30802;
w30804 <= not w30575 and w30705;
w30805 <= not w30701 and w30804;
w30806 <= not w30702 and not w30705;
w30807 <= not w30805 and not w30806;
w30808 <= not w30747 and not w30807;
w30809 <= not w30565 and not w30746;
w30810 <= not w30745 and w30809;
w30811 <= not w30808 and not w30810;
w30812 <= not b(12) and not w30811;
w30813 <= not w30584 and w30700;
w30814 <= not w30696 and w30813;
w30815 <= not w30697 and not w30700;
w30816 <= not w30814 and not w30815;
w30817 <= not w30747 and not w30816;
w30818 <= not w30574 and not w30746;
w30819 <= not w30745 and w30818;
w30820 <= not w30817 and not w30819;
w30821 <= not b(11) and not w30820;
w30822 <= not w30593 and w30695;
w30823 <= not w30691 and w30822;
w30824 <= not w30692 and not w30695;
w30825 <= not w30823 and not w30824;
w30826 <= not w30747 and not w30825;
w30827 <= not w30583 and not w30746;
w30828 <= not w30745 and w30827;
w30829 <= not w30826 and not w30828;
w30830 <= not b(10) and not w30829;
w30831 <= not w30602 and w30690;
w30832 <= not w30686 and w30831;
w30833 <= not w30687 and not w30690;
w30834 <= not w30832 and not w30833;
w30835 <= not w30747 and not w30834;
w30836 <= not w30592 and not w30746;
w30837 <= not w30745 and w30836;
w30838 <= not w30835 and not w30837;
w30839 <= not b(9) and not w30838;
w30840 <= not w30611 and w30685;
w30841 <= not w30681 and w30840;
w30842 <= not w30682 and not w30685;
w30843 <= not w30841 and not w30842;
w30844 <= not w30747 and not w30843;
w30845 <= not w30601 and not w30746;
w30846 <= not w30745 and w30845;
w30847 <= not w30844 and not w30846;
w30848 <= not b(8) and not w30847;
w30849 <= not w30620 and w30680;
w30850 <= not w30676 and w30849;
w30851 <= not w30677 and not w30680;
w30852 <= not w30850 and not w30851;
w30853 <= not w30747 and not w30852;
w30854 <= not w30610 and not w30746;
w30855 <= not w30745 and w30854;
w30856 <= not w30853 and not w30855;
w30857 <= not b(7) and not w30856;
w30858 <= not w30629 and w30675;
w30859 <= not w30671 and w30858;
w30860 <= not w30672 and not w30675;
w30861 <= not w30859 and not w30860;
w30862 <= not w30747 and not w30861;
w30863 <= not w30619 and not w30746;
w30864 <= not w30745 and w30863;
w30865 <= not w30862 and not w30864;
w30866 <= not b(6) and not w30865;
w30867 <= not w30638 and w30670;
w30868 <= not w30666 and w30867;
w30869 <= not w30667 and not w30670;
w30870 <= not w30868 and not w30869;
w30871 <= not w30747 and not w30870;
w30872 <= not w30628 and not w30746;
w30873 <= not w30745 and w30872;
w30874 <= not w30871 and not w30873;
w30875 <= not b(5) and not w30874;
w30876 <= not w30646 and w30665;
w30877 <= not w30661 and w30876;
w30878 <= not w30662 and not w30665;
w30879 <= not w30877 and not w30878;
w30880 <= not w30747 and not w30879;
w30881 <= not w30637 and not w30746;
w30882 <= not w30745 and w30881;
w30883 <= not w30880 and not w30882;
w30884 <= not b(4) and not w30883;
w30885 <= not w30656 and w30660;
w30886 <= not w30655 and w30885;
w30887 <= not w30657 and not w30660;
w30888 <= not w30886 and not w30887;
w30889 <= not w30747 and not w30888;
w30890 <= not w30645 and not w30746;
w30891 <= not w30745 and w30890;
w30892 <= not w30889 and not w30891;
w30893 <= not b(3) and not w30892;
w30894 <= w2356 and not w30653;
w30895 <= not w30651 and w30894;
w30896 <= not w30655 and not w30895;
w30897 <= not w30747 and w30896;
w30898 <= not w30650 and not w30746;
w30899 <= not w30745 and w30898;
w30900 <= not w30897 and not w30899;
w30901 <= not b(2) and not w30900;
w30902 <= b(0) and not w30747;
w30903 <= a(46) and not w30902;
w30904 <= w2356 and not w30747;
w30905 <= not w30903 and not w30904;
w30906 <= b(1) and not w30905;
w30907 <= not b(1) and not w30904;
w30908 <= not w30903 and w30907;
w30909 <= not w30906 and not w30908;
w30910 <= not w2616 and not w30909;
w30911 <= not b(1) and not w30905;
w30912 <= not w30910 and not w30911;
w30913 <= b(2) and not w30899;
w30914 <= not w30897 and w30913;
w30915 <= not w30901 and not w30914;
w30916 <= not w30912 and w30915;
w30917 <= not w30901 and not w30916;
w30918 <= b(3) and not w30891;
w30919 <= not w30889 and w30918;
w30920 <= not w30893 and not w30919;
w30921 <= not w30917 and w30920;
w30922 <= not w30893 and not w30921;
w30923 <= b(4) and not w30882;
w30924 <= not w30880 and w30923;
w30925 <= not w30884 and not w30924;
w30926 <= not w30922 and w30925;
w30927 <= not w30884 and not w30926;
w30928 <= b(5) and not w30873;
w30929 <= not w30871 and w30928;
w30930 <= not w30875 and not w30929;
w30931 <= not w30927 and w30930;
w30932 <= not w30875 and not w30931;
w30933 <= b(6) and not w30864;
w30934 <= not w30862 and w30933;
w30935 <= not w30866 and not w30934;
w30936 <= not w30932 and w30935;
w30937 <= not w30866 and not w30936;
w30938 <= b(7) and not w30855;
w30939 <= not w30853 and w30938;
w30940 <= not w30857 and not w30939;
w30941 <= not w30937 and w30940;
w30942 <= not w30857 and not w30941;
w30943 <= b(8) and not w30846;
w30944 <= not w30844 and w30943;
w30945 <= not w30848 and not w30944;
w30946 <= not w30942 and w30945;
w30947 <= not w30848 and not w30946;
w30948 <= b(9) and not w30837;
w30949 <= not w30835 and w30948;
w30950 <= not w30839 and not w30949;
w30951 <= not w30947 and w30950;
w30952 <= not w30839 and not w30951;
w30953 <= b(10) and not w30828;
w30954 <= not w30826 and w30953;
w30955 <= not w30830 and not w30954;
w30956 <= not w30952 and w30955;
w30957 <= not w30830 and not w30956;
w30958 <= b(11) and not w30819;
w30959 <= not w30817 and w30958;
w30960 <= not w30821 and not w30959;
w30961 <= not w30957 and w30960;
w30962 <= not w30821 and not w30961;
w30963 <= b(12) and not w30810;
w30964 <= not w30808 and w30963;
w30965 <= not w30812 and not w30964;
w30966 <= not w30962 and w30965;
w30967 <= not w30812 and not w30966;
w30968 <= b(13) and not w30801;
w30969 <= not w30799 and w30968;
w30970 <= not w30803 and not w30969;
w30971 <= not w30967 and w30970;
w30972 <= not w30803 and not w30971;
w30973 <= b(14) and not w30792;
w30974 <= not w30790 and w30973;
w30975 <= not w30794 and not w30974;
w30976 <= not w30972 and w30975;
w30977 <= not w30794 and not w30976;
w30978 <= b(15) and not w30783;
w30979 <= not w30781 and w30978;
w30980 <= not w30785 and not w30979;
w30981 <= not w30977 and w30980;
w30982 <= not w30785 and not w30981;
w30983 <= b(16) and not w30774;
w30984 <= not w30772 and w30983;
w30985 <= not w30776 and not w30984;
w30986 <= not w30982 and w30985;
w30987 <= not w30776 and not w30986;
w30988 <= b(17) and not w30754;
w30989 <= not w30752 and w30988;
w30990 <= not w30767 and not w30989;
w30991 <= not w30987 and w30990;
w30992 <= not w30767 and not w30991;
w30993 <= b(18) and not w30764;
w30994 <= not w30762 and w30993;
w30995 <= not w30766 and not w30994;
w30996 <= not w30992 and w30995;
w30997 <= not w30766 and not w30996;
w30998 <= w2708 and not w30997;
w30999 <= not w30755 and not w30998;
w31000 <= not w30776 and w30990;
w31001 <= not w30986 and w31000;
w31002 <= not w30987 and not w30990;
w31003 <= not w31001 and not w31002;
w31004 <= w2708 and not w31003;
w31005 <= not w30997 and w31004;
w31006 <= not w30999 and not w31005;
w31007 <= not w30765 and not w30998;
w31008 <= not w30767 and w30995;
w31009 <= not w30991 and w31008;
w31010 <= not w30992 and not w30995;
w31011 <= not w31009 and not w31010;
w31012 <= w30998 and not w31011;
w31013 <= not w31007 and not w31012;
w31014 <= not b(19) and not w31013;
w31015 <= not b(18) and not w31006;
w31016 <= not w30775 and not w30998;
w31017 <= not w30785 and w30985;
w31018 <= not w30981 and w31017;
w31019 <= not w30982 and not w30985;
w31020 <= not w31018 and not w31019;
w31021 <= w2708 and not w31020;
w31022 <= not w30997 and w31021;
w31023 <= not w31016 and not w31022;
w31024 <= not b(17) and not w31023;
w31025 <= not w30784 and not w30998;
w31026 <= not w30794 and w30980;
w31027 <= not w30976 and w31026;
w31028 <= not w30977 and not w30980;
w31029 <= not w31027 and not w31028;
w31030 <= w2708 and not w31029;
w31031 <= not w30997 and w31030;
w31032 <= not w31025 and not w31031;
w31033 <= not b(16) and not w31032;
w31034 <= not w30793 and not w30998;
w31035 <= not w30803 and w30975;
w31036 <= not w30971 and w31035;
w31037 <= not w30972 and not w30975;
w31038 <= not w31036 and not w31037;
w31039 <= w2708 and not w31038;
w31040 <= not w30997 and w31039;
w31041 <= not w31034 and not w31040;
w31042 <= not b(15) and not w31041;
w31043 <= not w30802 and not w30998;
w31044 <= not w30812 and w30970;
w31045 <= not w30966 and w31044;
w31046 <= not w30967 and not w30970;
w31047 <= not w31045 and not w31046;
w31048 <= w2708 and not w31047;
w31049 <= not w30997 and w31048;
w31050 <= not w31043 and not w31049;
w31051 <= not b(14) and not w31050;
w31052 <= not w30811 and not w30998;
w31053 <= not w30821 and w30965;
w31054 <= not w30961 and w31053;
w31055 <= not w30962 and not w30965;
w31056 <= not w31054 and not w31055;
w31057 <= w2708 and not w31056;
w31058 <= not w30997 and w31057;
w31059 <= not w31052 and not w31058;
w31060 <= not b(13) and not w31059;
w31061 <= not w30820 and not w30998;
w31062 <= not w30830 and w30960;
w31063 <= not w30956 and w31062;
w31064 <= not w30957 and not w30960;
w31065 <= not w31063 and not w31064;
w31066 <= w2708 and not w31065;
w31067 <= not w30997 and w31066;
w31068 <= not w31061 and not w31067;
w31069 <= not b(12) and not w31068;
w31070 <= not w30829 and not w30998;
w31071 <= not w30839 and w30955;
w31072 <= not w30951 and w31071;
w31073 <= not w30952 and not w30955;
w31074 <= not w31072 and not w31073;
w31075 <= w2708 and not w31074;
w31076 <= not w30997 and w31075;
w31077 <= not w31070 and not w31076;
w31078 <= not b(11) and not w31077;
w31079 <= not w30838 and not w30998;
w31080 <= not w30848 and w30950;
w31081 <= not w30946 and w31080;
w31082 <= not w30947 and not w30950;
w31083 <= not w31081 and not w31082;
w31084 <= w2708 and not w31083;
w31085 <= not w30997 and w31084;
w31086 <= not w31079 and not w31085;
w31087 <= not b(10) and not w31086;
w31088 <= not w30847 and not w30998;
w31089 <= not w30857 and w30945;
w31090 <= not w30941 and w31089;
w31091 <= not w30942 and not w30945;
w31092 <= not w31090 and not w31091;
w31093 <= w2708 and not w31092;
w31094 <= not w30997 and w31093;
w31095 <= not w31088 and not w31094;
w31096 <= not b(9) and not w31095;
w31097 <= not w30856 and not w30998;
w31098 <= not w30866 and w30940;
w31099 <= not w30936 and w31098;
w31100 <= not w30937 and not w30940;
w31101 <= not w31099 and not w31100;
w31102 <= w2708 and not w31101;
w31103 <= not w30997 and w31102;
w31104 <= not w31097 and not w31103;
w31105 <= not b(8) and not w31104;
w31106 <= not w30865 and not w30998;
w31107 <= not w30875 and w30935;
w31108 <= not w30931 and w31107;
w31109 <= not w30932 and not w30935;
w31110 <= not w31108 and not w31109;
w31111 <= w2708 and not w31110;
w31112 <= not w30997 and w31111;
w31113 <= not w31106 and not w31112;
w31114 <= not b(7) and not w31113;
w31115 <= not w30874 and not w30998;
w31116 <= not w30884 and w30930;
w31117 <= not w30926 and w31116;
w31118 <= not w30927 and not w30930;
w31119 <= not w31117 and not w31118;
w31120 <= w2708 and not w31119;
w31121 <= not w30997 and w31120;
w31122 <= not w31115 and not w31121;
w31123 <= not b(6) and not w31122;
w31124 <= not w30883 and not w30998;
w31125 <= not w30893 and w30925;
w31126 <= not w30921 and w31125;
w31127 <= not w30922 and not w30925;
w31128 <= not w31126 and not w31127;
w31129 <= w2708 and not w31128;
w31130 <= not w30997 and w31129;
w31131 <= not w31124 and not w31130;
w31132 <= not b(5) and not w31131;
w31133 <= not w30892 and not w30998;
w31134 <= not w30901 and w30920;
w31135 <= not w30916 and w31134;
w31136 <= not w30917 and not w30920;
w31137 <= not w31135 and not w31136;
w31138 <= w2708 and not w31137;
w31139 <= not w30997 and w31138;
w31140 <= not w31133 and not w31139;
w31141 <= not b(4) and not w31140;
w31142 <= not w30900 and not w30998;
w31143 <= not w30911 and w30915;
w31144 <= not w30910 and w31143;
w31145 <= not w30912 and not w30915;
w31146 <= not w31144 and not w31145;
w31147 <= w2708 and not w31146;
w31148 <= not w30997 and w31147;
w31149 <= not w31142 and not w31148;
w31150 <= not b(3) and not w31149;
w31151 <= not w30905 and not w30998;
w31152 <= w2616 and not w30908;
w31153 <= not w30906 and w31152;
w31154 <= w2708 and not w31153;
w31155 <= not w30910 and w31154;
w31156 <= not w30997 and w31155;
w31157 <= not w31151 and not w31156;
w31158 <= not b(2) and not w31157;
w31159 <= w2874 and not w30997;
w31160 <= a(45) and not w31159;
w31161 <= w2881 and not w30997;
w31162 <= not w31160 and not w31161;
w31163 <= b(1) and not w31162;
w31164 <= not b(1) and not w31161;
w31165 <= not w31160 and w31164;
w31166 <= not w31163 and not w31165;
w31167 <= not w2888 and not w31166;
w31168 <= not b(1) and not w31162;
w31169 <= not w31167 and not w31168;
w31170 <= b(2) and not w31156;
w31171 <= not w31151 and w31170;
w31172 <= not w31158 and not w31171;
w31173 <= not w31169 and w31172;
w31174 <= not w31158 and not w31173;
w31175 <= b(3) and not w31148;
w31176 <= not w31142 and w31175;
w31177 <= not w31150 and not w31176;
w31178 <= not w31174 and w31177;
w31179 <= not w31150 and not w31178;
w31180 <= b(4) and not w31139;
w31181 <= not w31133 and w31180;
w31182 <= not w31141 and not w31181;
w31183 <= not w31179 and w31182;
w31184 <= not w31141 and not w31183;
w31185 <= b(5) and not w31130;
w31186 <= not w31124 and w31185;
w31187 <= not w31132 and not w31186;
w31188 <= not w31184 and w31187;
w31189 <= not w31132 and not w31188;
w31190 <= b(6) and not w31121;
w31191 <= not w31115 and w31190;
w31192 <= not w31123 and not w31191;
w31193 <= not w31189 and w31192;
w31194 <= not w31123 and not w31193;
w31195 <= b(7) and not w31112;
w31196 <= not w31106 and w31195;
w31197 <= not w31114 and not w31196;
w31198 <= not w31194 and w31197;
w31199 <= not w31114 and not w31198;
w31200 <= b(8) and not w31103;
w31201 <= not w31097 and w31200;
w31202 <= not w31105 and not w31201;
w31203 <= not w31199 and w31202;
w31204 <= not w31105 and not w31203;
w31205 <= b(9) and not w31094;
w31206 <= not w31088 and w31205;
w31207 <= not w31096 and not w31206;
w31208 <= not w31204 and w31207;
w31209 <= not w31096 and not w31208;
w31210 <= b(10) and not w31085;
w31211 <= not w31079 and w31210;
w31212 <= not w31087 and not w31211;
w31213 <= not w31209 and w31212;
w31214 <= not w31087 and not w31213;
w31215 <= b(11) and not w31076;
w31216 <= not w31070 and w31215;
w31217 <= not w31078 and not w31216;
w31218 <= not w31214 and w31217;
w31219 <= not w31078 and not w31218;
w31220 <= b(12) and not w31067;
w31221 <= not w31061 and w31220;
w31222 <= not w31069 and not w31221;
w31223 <= not w31219 and w31222;
w31224 <= not w31069 and not w31223;
w31225 <= b(13) and not w31058;
w31226 <= not w31052 and w31225;
w31227 <= not w31060 and not w31226;
w31228 <= not w31224 and w31227;
w31229 <= not w31060 and not w31228;
w31230 <= b(14) and not w31049;
w31231 <= not w31043 and w31230;
w31232 <= not w31051 and not w31231;
w31233 <= not w31229 and w31232;
w31234 <= not w31051 and not w31233;
w31235 <= b(15) and not w31040;
w31236 <= not w31034 and w31235;
w31237 <= not w31042 and not w31236;
w31238 <= not w31234 and w31237;
w31239 <= not w31042 and not w31238;
w31240 <= b(16) and not w31031;
w31241 <= not w31025 and w31240;
w31242 <= not w31033 and not w31241;
w31243 <= not w31239 and w31242;
w31244 <= not w31033 and not w31243;
w31245 <= b(17) and not w31022;
w31246 <= not w31016 and w31245;
w31247 <= not w31024 and not w31246;
w31248 <= not w31244 and w31247;
w31249 <= not w31024 and not w31248;
w31250 <= b(18) and not w31005;
w31251 <= not w30999 and w31250;
w31252 <= not w31015 and not w31251;
w31253 <= not w31249 and w31252;
w31254 <= not w31015 and not w31253;
w31255 <= b(19) and not w31007;
w31256 <= not w31012 and w31255;
w31257 <= not w31014 and not w31256;
w31258 <= not w31254 and w31257;
w31259 <= not w31014 and not w31258;
w31260 <= w63 and not w31259;
w31261 <= not w31006 and not w31260;
w31262 <= not w31024 and w31252;
w31263 <= not w31248 and w31262;
w31264 <= not w31249 and not w31252;
w31265 <= not w31263 and not w31264;
w31266 <= w63 and not w31265;
w31267 <= not w31259 and w31266;
w31268 <= not w31261 and not w31267;
w31269 <= not b(19) and not w31268;
w31270 <= not w31023 and not w31260;
w31271 <= not w31033 and w31247;
w31272 <= not w31243 and w31271;
w31273 <= not w31244 and not w31247;
w31274 <= not w31272 and not w31273;
w31275 <= w63 and not w31274;
w31276 <= not w31259 and w31275;
w31277 <= not w31270 and not w31276;
w31278 <= not b(18) and not w31277;
w31279 <= not w31032 and not w31260;
w31280 <= not w31042 and w31242;
w31281 <= not w31238 and w31280;
w31282 <= not w31239 and not w31242;
w31283 <= not w31281 and not w31282;
w31284 <= w63 and not w31283;
w31285 <= not w31259 and w31284;
w31286 <= not w31279 and not w31285;
w31287 <= not b(17) and not w31286;
w31288 <= not w31041 and not w31260;
w31289 <= not w31051 and w31237;
w31290 <= not w31233 and w31289;
w31291 <= not w31234 and not w31237;
w31292 <= not w31290 and not w31291;
w31293 <= w63 and not w31292;
w31294 <= not w31259 and w31293;
w31295 <= not w31288 and not w31294;
w31296 <= not b(16) and not w31295;
w31297 <= not w31050 and not w31260;
w31298 <= not w31060 and w31232;
w31299 <= not w31228 and w31298;
w31300 <= not w31229 and not w31232;
w31301 <= not w31299 and not w31300;
w31302 <= w63 and not w31301;
w31303 <= not w31259 and w31302;
w31304 <= not w31297 and not w31303;
w31305 <= not b(15) and not w31304;
w31306 <= not w31059 and not w31260;
w31307 <= not w31069 and w31227;
w31308 <= not w31223 and w31307;
w31309 <= not w31224 and not w31227;
w31310 <= not w31308 and not w31309;
w31311 <= w63 and not w31310;
w31312 <= not w31259 and w31311;
w31313 <= not w31306 and not w31312;
w31314 <= not b(14) and not w31313;
w31315 <= not w31068 and not w31260;
w31316 <= not w31078 and w31222;
w31317 <= not w31218 and w31316;
w31318 <= not w31219 and not w31222;
w31319 <= not w31317 and not w31318;
w31320 <= w63 and not w31319;
w31321 <= not w31259 and w31320;
w31322 <= not w31315 and not w31321;
w31323 <= not b(13) and not w31322;
w31324 <= not w31077 and not w31260;
w31325 <= not w31087 and w31217;
w31326 <= not w31213 and w31325;
w31327 <= not w31214 and not w31217;
w31328 <= not w31326 and not w31327;
w31329 <= w63 and not w31328;
w31330 <= not w31259 and w31329;
w31331 <= not w31324 and not w31330;
w31332 <= not b(12) and not w31331;
w31333 <= not w31086 and not w31260;
w31334 <= not w31096 and w31212;
w31335 <= not w31208 and w31334;
w31336 <= not w31209 and not w31212;
w31337 <= not w31335 and not w31336;
w31338 <= w63 and not w31337;
w31339 <= not w31259 and w31338;
w31340 <= not w31333 and not w31339;
w31341 <= not b(11) and not w31340;
w31342 <= not w31095 and not w31260;
w31343 <= not w31105 and w31207;
w31344 <= not w31203 and w31343;
w31345 <= not w31204 and not w31207;
w31346 <= not w31344 and not w31345;
w31347 <= w63 and not w31346;
w31348 <= not w31259 and w31347;
w31349 <= not w31342 and not w31348;
w31350 <= not b(10) and not w31349;
w31351 <= not w31104 and not w31260;
w31352 <= not w31114 and w31202;
w31353 <= not w31198 and w31352;
w31354 <= not w31199 and not w31202;
w31355 <= not w31353 and not w31354;
w31356 <= w63 and not w31355;
w31357 <= not w31259 and w31356;
w31358 <= not w31351 and not w31357;
w31359 <= not b(9) and not w31358;
w31360 <= not w31113 and not w31260;
w31361 <= not w31123 and w31197;
w31362 <= not w31193 and w31361;
w31363 <= not w31194 and not w31197;
w31364 <= not w31362 and not w31363;
w31365 <= w63 and not w31364;
w31366 <= not w31259 and w31365;
w31367 <= not w31360 and not w31366;
w31368 <= not b(8) and not w31367;
w31369 <= not w31122 and not w31260;
w31370 <= not w31132 and w31192;
w31371 <= not w31188 and w31370;
w31372 <= not w31189 and not w31192;
w31373 <= not w31371 and not w31372;
w31374 <= w63 and not w31373;
w31375 <= not w31259 and w31374;
w31376 <= not w31369 and not w31375;
w31377 <= not b(7) and not w31376;
w31378 <= not w31131 and not w31260;
w31379 <= not w31141 and w31187;
w31380 <= not w31183 and w31379;
w31381 <= not w31184 and not w31187;
w31382 <= not w31380 and not w31381;
w31383 <= w63 and not w31382;
w31384 <= not w31259 and w31383;
w31385 <= not w31378 and not w31384;
w31386 <= not b(6) and not w31385;
w31387 <= not w31140 and not w31260;
w31388 <= not w31150 and w31182;
w31389 <= not w31178 and w31388;
w31390 <= not w31179 and not w31182;
w31391 <= not w31389 and not w31390;
w31392 <= w63 and not w31391;
w31393 <= not w31259 and w31392;
w31394 <= not w31387 and not w31393;
w31395 <= not b(5) and not w31394;
w31396 <= not w31149 and not w31260;
w31397 <= not w31158 and w31177;
w31398 <= not w31173 and w31397;
w31399 <= not w31174 and not w31177;
w31400 <= not w31398 and not w31399;
w31401 <= w63 and not w31400;
w31402 <= not w31259 and w31401;
w31403 <= not w31396 and not w31402;
w31404 <= not b(4) and not w31403;
w31405 <= not w31157 and not w31260;
w31406 <= not w31168 and w31172;
w31407 <= not w31167 and w31406;
w31408 <= not w31169 and not w31172;
w31409 <= not w31407 and not w31408;
w31410 <= w63 and not w31409;
w31411 <= not w31259 and w31410;
w31412 <= not w31405 and not w31411;
w31413 <= not b(3) and not w31412;
w31414 <= not w31162 and not w31260;
w31415 <= w2888 and not w31165;
w31416 <= not w31163 and w31415;
w31417 <= w63 and not w31416;
w31418 <= not w31167 and w31417;
w31419 <= not w31259 and w31418;
w31420 <= not w31414 and not w31419;
w31421 <= not b(2) and not w31420;
w31422 <= w3148 and not w31259;
w31423 <= a(44) and not w31422;
w31424 <= w3154 and not w31259;
w31425 <= not w31423 and not w31424;
w31426 <= b(1) and not w31425;
w31427 <= not b(1) and not w31424;
w31428 <= not w31423 and w31427;
w31429 <= not w31426 and not w31428;
w31430 <= not w3161 and not w31429;
w31431 <= not b(1) and not w31425;
w31432 <= not w31430 and not w31431;
w31433 <= b(2) and not w31419;
w31434 <= not w31414 and w31433;
w31435 <= not w31421 and not w31434;
w31436 <= not w31432 and w31435;
w31437 <= not w31421 and not w31436;
w31438 <= b(3) and not w31411;
w31439 <= not w31405 and w31438;
w31440 <= not w31413 and not w31439;
w31441 <= not w31437 and w31440;
w31442 <= not w31413 and not w31441;
w31443 <= b(4) and not w31402;
w31444 <= not w31396 and w31443;
w31445 <= not w31404 and not w31444;
w31446 <= not w31442 and w31445;
w31447 <= not w31404 and not w31446;
w31448 <= b(5) and not w31393;
w31449 <= not w31387 and w31448;
w31450 <= not w31395 and not w31449;
w31451 <= not w31447 and w31450;
w31452 <= not w31395 and not w31451;
w31453 <= b(6) and not w31384;
w31454 <= not w31378 and w31453;
w31455 <= not w31386 and not w31454;
w31456 <= not w31452 and w31455;
w31457 <= not w31386 and not w31456;
w31458 <= b(7) and not w31375;
w31459 <= not w31369 and w31458;
w31460 <= not w31377 and not w31459;
w31461 <= not w31457 and w31460;
w31462 <= not w31377 and not w31461;
w31463 <= b(8) and not w31366;
w31464 <= not w31360 and w31463;
w31465 <= not w31368 and not w31464;
w31466 <= not w31462 and w31465;
w31467 <= not w31368 and not w31466;
w31468 <= b(9) and not w31357;
w31469 <= not w31351 and w31468;
w31470 <= not w31359 and not w31469;
w31471 <= not w31467 and w31470;
w31472 <= not w31359 and not w31471;
w31473 <= b(10) and not w31348;
w31474 <= not w31342 and w31473;
w31475 <= not w31350 and not w31474;
w31476 <= not w31472 and w31475;
w31477 <= not w31350 and not w31476;
w31478 <= b(11) and not w31339;
w31479 <= not w31333 and w31478;
w31480 <= not w31341 and not w31479;
w31481 <= not w31477 and w31480;
w31482 <= not w31341 and not w31481;
w31483 <= b(12) and not w31330;
w31484 <= not w31324 and w31483;
w31485 <= not w31332 and not w31484;
w31486 <= not w31482 and w31485;
w31487 <= not w31332 and not w31486;
w31488 <= b(13) and not w31321;
w31489 <= not w31315 and w31488;
w31490 <= not w31323 and not w31489;
w31491 <= not w31487 and w31490;
w31492 <= not w31323 and not w31491;
w31493 <= b(14) and not w31312;
w31494 <= not w31306 and w31493;
w31495 <= not w31314 and not w31494;
w31496 <= not w31492 and w31495;
w31497 <= not w31314 and not w31496;
w31498 <= b(15) and not w31303;
w31499 <= not w31297 and w31498;
w31500 <= not w31305 and not w31499;
w31501 <= not w31497 and w31500;
w31502 <= not w31305 and not w31501;
w31503 <= b(16) and not w31294;
w31504 <= not w31288 and w31503;
w31505 <= not w31296 and not w31504;
w31506 <= not w31502 and w31505;
w31507 <= not w31296 and not w31506;
w31508 <= b(17) and not w31285;
w31509 <= not w31279 and w31508;
w31510 <= not w31287 and not w31509;
w31511 <= not w31507 and w31510;
w31512 <= not w31287 and not w31511;
w31513 <= b(18) and not w31276;
w31514 <= not w31270 and w31513;
w31515 <= not w31278 and not w31514;
w31516 <= not w31512 and w31515;
w31517 <= not w31278 and not w31516;
w31518 <= b(19) and not w31267;
w31519 <= not w31261 and w31518;
w31520 <= not w31269 and not w31519;
w31521 <= not w31517 and w31520;
w31522 <= not w31269 and not w31521;
w31523 <= not w31013 and not w31260;
w31524 <= not w31015 and w31257;
w31525 <= not w31253 and w31524;
w31526 <= not w31254 and not w31257;
w31527 <= not w31525 and not w31526;
w31528 <= w31260 and not w31527;
w31529 <= not w31523 and not w31528;
w31530 <= not b(20) and not w31529;
w31531 <= b(20) and not w31523;
w31532 <= not w31528 and w31531;
w31533 <= w386 and not w31532;
w31534 <= not w31530 and w31533;
w31535 <= not w31522 and w31534;
w31536 <= w63 and not w31529;
w31537 <= not w31535 and not w31536;
w31538 <= not w31278 and w31520;
w31539 <= not w31516 and w31538;
w31540 <= not w31517 and not w31520;
w31541 <= not w31539 and not w31540;
w31542 <= not w31537 and not w31541;
w31543 <= not w31268 and not w31536;
w31544 <= not w31535 and w31543;
w31545 <= not w31542 and not w31544;
w31546 <= not w31269 and not w31532;
w31547 <= not w31530 and w31546;
w31548 <= not w31521 and w31547;
w31549 <= not w31530 and not w31532;
w31550 <= not w31522 and not w31549;
w31551 <= not w31548 and not w31550;
w31552 <= not w31537 and not w31551;
w31553 <= not w31529 and not w31536;
w31554 <= not w31535 and w31553;
w31555 <= not w31552 and not w31554;
w31556 <= not b(21) and not w31555;
w31557 <= not b(20) and not w31545;
w31558 <= not w31287 and w31515;
w31559 <= not w31511 and w31558;
w31560 <= not w31512 and not w31515;
w31561 <= not w31559 and not w31560;
w31562 <= not w31537 and not w31561;
w31563 <= not w31277 and not w31536;
w31564 <= not w31535 and w31563;
w31565 <= not w31562 and not w31564;
w31566 <= not b(19) and not w31565;
w31567 <= not w31296 and w31510;
w31568 <= not w31506 and w31567;
w31569 <= not w31507 and not w31510;
w31570 <= not w31568 and not w31569;
w31571 <= not w31537 and not w31570;
w31572 <= not w31286 and not w31536;
w31573 <= not w31535 and w31572;
w31574 <= not w31571 and not w31573;
w31575 <= not b(18) and not w31574;
w31576 <= not w31305 and w31505;
w31577 <= not w31501 and w31576;
w31578 <= not w31502 and not w31505;
w31579 <= not w31577 and not w31578;
w31580 <= not w31537 and not w31579;
w31581 <= not w31295 and not w31536;
w31582 <= not w31535 and w31581;
w31583 <= not w31580 and not w31582;
w31584 <= not b(17) and not w31583;
w31585 <= not w31314 and w31500;
w31586 <= not w31496 and w31585;
w31587 <= not w31497 and not w31500;
w31588 <= not w31586 and not w31587;
w31589 <= not w31537 and not w31588;
w31590 <= not w31304 and not w31536;
w31591 <= not w31535 and w31590;
w31592 <= not w31589 and not w31591;
w31593 <= not b(16) and not w31592;
w31594 <= not w31323 and w31495;
w31595 <= not w31491 and w31594;
w31596 <= not w31492 and not w31495;
w31597 <= not w31595 and not w31596;
w31598 <= not w31537 and not w31597;
w31599 <= not w31313 and not w31536;
w31600 <= not w31535 and w31599;
w31601 <= not w31598 and not w31600;
w31602 <= not b(15) and not w31601;
w31603 <= not w31332 and w31490;
w31604 <= not w31486 and w31603;
w31605 <= not w31487 and not w31490;
w31606 <= not w31604 and not w31605;
w31607 <= not w31537 and not w31606;
w31608 <= not w31322 and not w31536;
w31609 <= not w31535 and w31608;
w31610 <= not w31607 and not w31609;
w31611 <= not b(14) and not w31610;
w31612 <= not w31341 and w31485;
w31613 <= not w31481 and w31612;
w31614 <= not w31482 and not w31485;
w31615 <= not w31613 and not w31614;
w31616 <= not w31537 and not w31615;
w31617 <= not w31331 and not w31536;
w31618 <= not w31535 and w31617;
w31619 <= not w31616 and not w31618;
w31620 <= not b(13) and not w31619;
w31621 <= not w31350 and w31480;
w31622 <= not w31476 and w31621;
w31623 <= not w31477 and not w31480;
w31624 <= not w31622 and not w31623;
w31625 <= not w31537 and not w31624;
w31626 <= not w31340 and not w31536;
w31627 <= not w31535 and w31626;
w31628 <= not w31625 and not w31627;
w31629 <= not b(12) and not w31628;
w31630 <= not w31359 and w31475;
w31631 <= not w31471 and w31630;
w31632 <= not w31472 and not w31475;
w31633 <= not w31631 and not w31632;
w31634 <= not w31537 and not w31633;
w31635 <= not w31349 and not w31536;
w31636 <= not w31535 and w31635;
w31637 <= not w31634 and not w31636;
w31638 <= not b(11) and not w31637;
w31639 <= not w31368 and w31470;
w31640 <= not w31466 and w31639;
w31641 <= not w31467 and not w31470;
w31642 <= not w31640 and not w31641;
w31643 <= not w31537 and not w31642;
w31644 <= not w31358 and not w31536;
w31645 <= not w31535 and w31644;
w31646 <= not w31643 and not w31645;
w31647 <= not b(10) and not w31646;
w31648 <= not w31377 and w31465;
w31649 <= not w31461 and w31648;
w31650 <= not w31462 and not w31465;
w31651 <= not w31649 and not w31650;
w31652 <= not w31537 and not w31651;
w31653 <= not w31367 and not w31536;
w31654 <= not w31535 and w31653;
w31655 <= not w31652 and not w31654;
w31656 <= not b(9) and not w31655;
w31657 <= not w31386 and w31460;
w31658 <= not w31456 and w31657;
w31659 <= not w31457 and not w31460;
w31660 <= not w31658 and not w31659;
w31661 <= not w31537 and not w31660;
w31662 <= not w31376 and not w31536;
w31663 <= not w31535 and w31662;
w31664 <= not w31661 and not w31663;
w31665 <= not b(8) and not w31664;
w31666 <= not w31395 and w31455;
w31667 <= not w31451 and w31666;
w31668 <= not w31452 and not w31455;
w31669 <= not w31667 and not w31668;
w31670 <= not w31537 and not w31669;
w31671 <= not w31385 and not w31536;
w31672 <= not w31535 and w31671;
w31673 <= not w31670 and not w31672;
w31674 <= not b(7) and not w31673;
w31675 <= not w31404 and w31450;
w31676 <= not w31446 and w31675;
w31677 <= not w31447 and not w31450;
w31678 <= not w31676 and not w31677;
w31679 <= not w31537 and not w31678;
w31680 <= not w31394 and not w31536;
w31681 <= not w31535 and w31680;
w31682 <= not w31679 and not w31681;
w31683 <= not b(6) and not w31682;
w31684 <= not w31413 and w31445;
w31685 <= not w31441 and w31684;
w31686 <= not w31442 and not w31445;
w31687 <= not w31685 and not w31686;
w31688 <= not w31537 and not w31687;
w31689 <= not w31403 and not w31536;
w31690 <= not w31535 and w31689;
w31691 <= not w31688 and not w31690;
w31692 <= not b(5) and not w31691;
w31693 <= not w31421 and w31440;
w31694 <= not w31436 and w31693;
w31695 <= not w31437 and not w31440;
w31696 <= not w31694 and not w31695;
w31697 <= not w31537 and not w31696;
w31698 <= not w31412 and not w31536;
w31699 <= not w31535 and w31698;
w31700 <= not w31697 and not w31699;
w31701 <= not b(4) and not w31700;
w31702 <= not w31431 and w31435;
w31703 <= not w31430 and w31702;
w31704 <= not w31432 and not w31435;
w31705 <= not w31703 and not w31704;
w31706 <= not w31537 and not w31705;
w31707 <= not w31420 and not w31536;
w31708 <= not w31535 and w31707;
w31709 <= not w31706 and not w31708;
w31710 <= not b(3) and not w31709;
w31711 <= w3161 and not w31428;
w31712 <= not w31426 and w31711;
w31713 <= not w31430 and not w31712;
w31714 <= not w31537 and w31713;
w31715 <= not w31425 and not w31536;
w31716 <= not w31535 and w31715;
w31717 <= not w31714 and not w31716;
w31718 <= not b(2) and not w31717;
w31719 <= b(0) and not w31537;
w31720 <= a(43) and not w31719;
w31721 <= w3161 and not w31537;
w31722 <= not w31720 and not w31721;
w31723 <= b(1) and not w31722;
w31724 <= not b(1) and not w31721;
w31725 <= not w31720 and w31724;
w31726 <= not w31723 and not w31725;
w31727 <= not w3459 and not w31726;
w31728 <= not b(1) and not w31722;
w31729 <= not w31727 and not w31728;
w31730 <= b(2) and not w31716;
w31731 <= not w31714 and w31730;
w31732 <= not w31718 and not w31731;
w31733 <= not w31729 and w31732;
w31734 <= not w31718 and not w31733;
w31735 <= b(3) and not w31708;
w31736 <= not w31706 and w31735;
w31737 <= not w31710 and not w31736;
w31738 <= not w31734 and w31737;
w31739 <= not w31710 and not w31738;
w31740 <= b(4) and not w31699;
w31741 <= not w31697 and w31740;
w31742 <= not w31701 and not w31741;
w31743 <= not w31739 and w31742;
w31744 <= not w31701 and not w31743;
w31745 <= b(5) and not w31690;
w31746 <= not w31688 and w31745;
w31747 <= not w31692 and not w31746;
w31748 <= not w31744 and w31747;
w31749 <= not w31692 and not w31748;
w31750 <= b(6) and not w31681;
w31751 <= not w31679 and w31750;
w31752 <= not w31683 and not w31751;
w31753 <= not w31749 and w31752;
w31754 <= not w31683 and not w31753;
w31755 <= b(7) and not w31672;
w31756 <= not w31670 and w31755;
w31757 <= not w31674 and not w31756;
w31758 <= not w31754 and w31757;
w31759 <= not w31674 and not w31758;
w31760 <= b(8) and not w31663;
w31761 <= not w31661 and w31760;
w31762 <= not w31665 and not w31761;
w31763 <= not w31759 and w31762;
w31764 <= not w31665 and not w31763;
w31765 <= b(9) and not w31654;
w31766 <= not w31652 and w31765;
w31767 <= not w31656 and not w31766;
w31768 <= not w31764 and w31767;
w31769 <= not w31656 and not w31768;
w31770 <= b(10) and not w31645;
w31771 <= not w31643 and w31770;
w31772 <= not w31647 and not w31771;
w31773 <= not w31769 and w31772;
w31774 <= not w31647 and not w31773;
w31775 <= b(11) and not w31636;
w31776 <= not w31634 and w31775;
w31777 <= not w31638 and not w31776;
w31778 <= not w31774 and w31777;
w31779 <= not w31638 and not w31778;
w31780 <= b(12) and not w31627;
w31781 <= not w31625 and w31780;
w31782 <= not w31629 and not w31781;
w31783 <= not w31779 and w31782;
w31784 <= not w31629 and not w31783;
w31785 <= b(13) and not w31618;
w31786 <= not w31616 and w31785;
w31787 <= not w31620 and not w31786;
w31788 <= not w31784 and w31787;
w31789 <= not w31620 and not w31788;
w31790 <= b(14) and not w31609;
w31791 <= not w31607 and w31790;
w31792 <= not w31611 and not w31791;
w31793 <= not w31789 and w31792;
w31794 <= not w31611 and not w31793;
w31795 <= b(15) and not w31600;
w31796 <= not w31598 and w31795;
w31797 <= not w31602 and not w31796;
w31798 <= not w31794 and w31797;
w31799 <= not w31602 and not w31798;
w31800 <= b(16) and not w31591;
w31801 <= not w31589 and w31800;
w31802 <= not w31593 and not w31801;
w31803 <= not w31799 and w31802;
w31804 <= not w31593 and not w31803;
w31805 <= b(17) and not w31582;
w31806 <= not w31580 and w31805;
w31807 <= not w31584 and not w31806;
w31808 <= not w31804 and w31807;
w31809 <= not w31584 and not w31808;
w31810 <= b(18) and not w31573;
w31811 <= not w31571 and w31810;
w31812 <= not w31575 and not w31811;
w31813 <= not w31809 and w31812;
w31814 <= not w31575 and not w31813;
w31815 <= b(19) and not w31564;
w31816 <= not w31562 and w31815;
w31817 <= not w31566 and not w31816;
w31818 <= not w31814 and w31817;
w31819 <= not w31566 and not w31818;
w31820 <= b(20) and not w31544;
w31821 <= not w31542 and w31820;
w31822 <= not w31557 and not w31821;
w31823 <= not w31819 and w31822;
w31824 <= not w31557 and not w31823;
w31825 <= b(21) and not w31554;
w31826 <= not w31552 and w31825;
w31827 <= not w31556 and not w31826;
w31828 <= not w31824 and w31827;
w31829 <= not w31556 and not w31828;
w31830 <= w3566 and not w31829;
w31831 <= not w31545 and not w31830;
w31832 <= not w31566 and w31822;
w31833 <= not w31818 and w31832;
w31834 <= not w31819 and not w31822;
w31835 <= not w31833 and not w31834;
w31836 <= w3566 and not w31835;
w31837 <= not w31829 and w31836;
w31838 <= not w31831 and not w31837;
w31839 <= not w31555 and not w31830;
w31840 <= not w31557 and w31827;
w31841 <= not w31823 and w31840;
w31842 <= not w31824 and not w31827;
w31843 <= not w31841 and not w31842;
w31844 <= w31830 and not w31843;
w31845 <= not w31839 and not w31844;
w31846 <= not b(22) and not w31845;
w31847 <= not b(21) and not w31838;
w31848 <= not w31565 and not w31830;
w31849 <= not w31575 and w31817;
w31850 <= not w31813 and w31849;
w31851 <= not w31814 and not w31817;
w31852 <= not w31850 and not w31851;
w31853 <= w3566 and not w31852;
w31854 <= not w31829 and w31853;
w31855 <= not w31848 and not w31854;
w31856 <= not b(20) and not w31855;
w31857 <= not w31574 and not w31830;
w31858 <= not w31584 and w31812;
w31859 <= not w31808 and w31858;
w31860 <= not w31809 and not w31812;
w31861 <= not w31859 and not w31860;
w31862 <= w3566 and not w31861;
w31863 <= not w31829 and w31862;
w31864 <= not w31857 and not w31863;
w31865 <= not b(19) and not w31864;
w31866 <= not w31583 and not w31830;
w31867 <= not w31593 and w31807;
w31868 <= not w31803 and w31867;
w31869 <= not w31804 and not w31807;
w31870 <= not w31868 and not w31869;
w31871 <= w3566 and not w31870;
w31872 <= not w31829 and w31871;
w31873 <= not w31866 and not w31872;
w31874 <= not b(18) and not w31873;
w31875 <= not w31592 and not w31830;
w31876 <= not w31602 and w31802;
w31877 <= not w31798 and w31876;
w31878 <= not w31799 and not w31802;
w31879 <= not w31877 and not w31878;
w31880 <= w3566 and not w31879;
w31881 <= not w31829 and w31880;
w31882 <= not w31875 and not w31881;
w31883 <= not b(17) and not w31882;
w31884 <= not w31601 and not w31830;
w31885 <= not w31611 and w31797;
w31886 <= not w31793 and w31885;
w31887 <= not w31794 and not w31797;
w31888 <= not w31886 and not w31887;
w31889 <= w3566 and not w31888;
w31890 <= not w31829 and w31889;
w31891 <= not w31884 and not w31890;
w31892 <= not b(16) and not w31891;
w31893 <= not w31610 and not w31830;
w31894 <= not w31620 and w31792;
w31895 <= not w31788 and w31894;
w31896 <= not w31789 and not w31792;
w31897 <= not w31895 and not w31896;
w31898 <= w3566 and not w31897;
w31899 <= not w31829 and w31898;
w31900 <= not w31893 and not w31899;
w31901 <= not b(15) and not w31900;
w31902 <= not w31619 and not w31830;
w31903 <= not w31629 and w31787;
w31904 <= not w31783 and w31903;
w31905 <= not w31784 and not w31787;
w31906 <= not w31904 and not w31905;
w31907 <= w3566 and not w31906;
w31908 <= not w31829 and w31907;
w31909 <= not w31902 and not w31908;
w31910 <= not b(14) and not w31909;
w31911 <= not w31628 and not w31830;
w31912 <= not w31638 and w31782;
w31913 <= not w31778 and w31912;
w31914 <= not w31779 and not w31782;
w31915 <= not w31913 and not w31914;
w31916 <= w3566 and not w31915;
w31917 <= not w31829 and w31916;
w31918 <= not w31911 and not w31917;
w31919 <= not b(13) and not w31918;
w31920 <= not w31637 and not w31830;
w31921 <= not w31647 and w31777;
w31922 <= not w31773 and w31921;
w31923 <= not w31774 and not w31777;
w31924 <= not w31922 and not w31923;
w31925 <= w3566 and not w31924;
w31926 <= not w31829 and w31925;
w31927 <= not w31920 and not w31926;
w31928 <= not b(12) and not w31927;
w31929 <= not w31646 and not w31830;
w31930 <= not w31656 and w31772;
w31931 <= not w31768 and w31930;
w31932 <= not w31769 and not w31772;
w31933 <= not w31931 and not w31932;
w31934 <= w3566 and not w31933;
w31935 <= not w31829 and w31934;
w31936 <= not w31929 and not w31935;
w31937 <= not b(11) and not w31936;
w31938 <= not w31655 and not w31830;
w31939 <= not w31665 and w31767;
w31940 <= not w31763 and w31939;
w31941 <= not w31764 and not w31767;
w31942 <= not w31940 and not w31941;
w31943 <= w3566 and not w31942;
w31944 <= not w31829 and w31943;
w31945 <= not w31938 and not w31944;
w31946 <= not b(10) and not w31945;
w31947 <= not w31664 and not w31830;
w31948 <= not w31674 and w31762;
w31949 <= not w31758 and w31948;
w31950 <= not w31759 and not w31762;
w31951 <= not w31949 and not w31950;
w31952 <= w3566 and not w31951;
w31953 <= not w31829 and w31952;
w31954 <= not w31947 and not w31953;
w31955 <= not b(9) and not w31954;
w31956 <= not w31673 and not w31830;
w31957 <= not w31683 and w31757;
w31958 <= not w31753 and w31957;
w31959 <= not w31754 and not w31757;
w31960 <= not w31958 and not w31959;
w31961 <= w3566 and not w31960;
w31962 <= not w31829 and w31961;
w31963 <= not w31956 and not w31962;
w31964 <= not b(8) and not w31963;
w31965 <= not w31682 and not w31830;
w31966 <= not w31692 and w31752;
w31967 <= not w31748 and w31966;
w31968 <= not w31749 and not w31752;
w31969 <= not w31967 and not w31968;
w31970 <= w3566 and not w31969;
w31971 <= not w31829 and w31970;
w31972 <= not w31965 and not w31971;
w31973 <= not b(7) and not w31972;
w31974 <= not w31691 and not w31830;
w31975 <= not w31701 and w31747;
w31976 <= not w31743 and w31975;
w31977 <= not w31744 and not w31747;
w31978 <= not w31976 and not w31977;
w31979 <= w3566 and not w31978;
w31980 <= not w31829 and w31979;
w31981 <= not w31974 and not w31980;
w31982 <= not b(6) and not w31981;
w31983 <= not w31700 and not w31830;
w31984 <= not w31710 and w31742;
w31985 <= not w31738 and w31984;
w31986 <= not w31739 and not w31742;
w31987 <= not w31985 and not w31986;
w31988 <= w3566 and not w31987;
w31989 <= not w31829 and w31988;
w31990 <= not w31983 and not w31989;
w31991 <= not b(5) and not w31990;
w31992 <= not w31709 and not w31830;
w31993 <= not w31718 and w31737;
w31994 <= not w31733 and w31993;
w31995 <= not w31734 and not w31737;
w31996 <= not w31994 and not w31995;
w31997 <= w3566 and not w31996;
w31998 <= not w31829 and w31997;
w31999 <= not w31992 and not w31998;
w32000 <= not b(4) and not w31999;
w32001 <= not w31717 and not w31830;
w32002 <= not w31728 and w31732;
w32003 <= not w31727 and w32002;
w32004 <= not w31729 and not w31732;
w32005 <= not w32003 and not w32004;
w32006 <= w3566 and not w32005;
w32007 <= not w31829 and w32006;
w32008 <= not w32001 and not w32007;
w32009 <= not b(3) and not w32008;
w32010 <= not w31722 and not w31830;
w32011 <= w3459 and not w31725;
w32012 <= not w31723 and w32011;
w32013 <= w3566 and not w32012;
w32014 <= not w31727 and w32013;
w32015 <= not w31829 and w32014;
w32016 <= not w32010 and not w32015;
w32017 <= not b(2) and not w32016;
w32018 <= w3760 and not w31829;
w32019 <= a(42) and not w32018;
w32020 <= w3767 and not w31829;
w32021 <= not w32019 and not w32020;
w32022 <= b(1) and not w32021;
w32023 <= not b(1) and not w32020;
w32024 <= not w32019 and w32023;
w32025 <= not w32022 and not w32024;
w32026 <= not w3774 and not w32025;
w32027 <= not b(1) and not w32021;
w32028 <= not w32026 and not w32027;
w32029 <= b(2) and not w32015;
w32030 <= not w32010 and w32029;
w32031 <= not w32017 and not w32030;
w32032 <= not w32028 and w32031;
w32033 <= not w32017 and not w32032;
w32034 <= b(3) and not w32007;
w32035 <= not w32001 and w32034;
w32036 <= not w32009 and not w32035;
w32037 <= not w32033 and w32036;
w32038 <= not w32009 and not w32037;
w32039 <= b(4) and not w31998;
w32040 <= not w31992 and w32039;
w32041 <= not w32000 and not w32040;
w32042 <= not w32038 and w32041;
w32043 <= not w32000 and not w32042;
w32044 <= b(5) and not w31989;
w32045 <= not w31983 and w32044;
w32046 <= not w31991 and not w32045;
w32047 <= not w32043 and w32046;
w32048 <= not w31991 and not w32047;
w32049 <= b(6) and not w31980;
w32050 <= not w31974 and w32049;
w32051 <= not w31982 and not w32050;
w32052 <= not w32048 and w32051;
w32053 <= not w31982 and not w32052;
w32054 <= b(7) and not w31971;
w32055 <= not w31965 and w32054;
w32056 <= not w31973 and not w32055;
w32057 <= not w32053 and w32056;
w32058 <= not w31973 and not w32057;
w32059 <= b(8) and not w31962;
w32060 <= not w31956 and w32059;
w32061 <= not w31964 and not w32060;
w32062 <= not w32058 and w32061;
w32063 <= not w31964 and not w32062;
w32064 <= b(9) and not w31953;
w32065 <= not w31947 and w32064;
w32066 <= not w31955 and not w32065;
w32067 <= not w32063 and w32066;
w32068 <= not w31955 and not w32067;
w32069 <= b(10) and not w31944;
w32070 <= not w31938 and w32069;
w32071 <= not w31946 and not w32070;
w32072 <= not w32068 and w32071;
w32073 <= not w31946 and not w32072;
w32074 <= b(11) and not w31935;
w32075 <= not w31929 and w32074;
w32076 <= not w31937 and not w32075;
w32077 <= not w32073 and w32076;
w32078 <= not w31937 and not w32077;
w32079 <= b(12) and not w31926;
w32080 <= not w31920 and w32079;
w32081 <= not w31928 and not w32080;
w32082 <= not w32078 and w32081;
w32083 <= not w31928 and not w32082;
w32084 <= b(13) and not w31917;
w32085 <= not w31911 and w32084;
w32086 <= not w31919 and not w32085;
w32087 <= not w32083 and w32086;
w32088 <= not w31919 and not w32087;
w32089 <= b(14) and not w31908;
w32090 <= not w31902 and w32089;
w32091 <= not w31910 and not w32090;
w32092 <= not w32088 and w32091;
w32093 <= not w31910 and not w32092;
w32094 <= b(15) and not w31899;
w32095 <= not w31893 and w32094;
w32096 <= not w31901 and not w32095;
w32097 <= not w32093 and w32096;
w32098 <= not w31901 and not w32097;
w32099 <= b(16) and not w31890;
w32100 <= not w31884 and w32099;
w32101 <= not w31892 and not w32100;
w32102 <= not w32098 and w32101;
w32103 <= not w31892 and not w32102;
w32104 <= b(17) and not w31881;
w32105 <= not w31875 and w32104;
w32106 <= not w31883 and not w32105;
w32107 <= not w32103 and w32106;
w32108 <= not w31883 and not w32107;
w32109 <= b(18) and not w31872;
w32110 <= not w31866 and w32109;
w32111 <= not w31874 and not w32110;
w32112 <= not w32108 and w32111;
w32113 <= not w31874 and not w32112;
w32114 <= b(19) and not w31863;
w32115 <= not w31857 and w32114;
w32116 <= not w31865 and not w32115;
w32117 <= not w32113 and w32116;
w32118 <= not w31865 and not w32117;
w32119 <= b(20) and not w31854;
w32120 <= not w31848 and w32119;
w32121 <= not w31856 and not w32120;
w32122 <= not w32118 and w32121;
w32123 <= not w31856 and not w32122;
w32124 <= b(21) and not w31837;
w32125 <= not w31831 and w32124;
w32126 <= not w31847 and not w32125;
w32127 <= not w32123 and w32126;
w32128 <= not w31847 and not w32127;
w32129 <= b(22) and not w31839;
w32130 <= not w31844 and w32129;
w32131 <= not w31846 and not w32130;
w32132 <= not w32128 and w32131;
w32133 <= not w31846 and not w32132;
w32134 <= w3886 and not w32133;
w32135 <= not w31838 and not w32134;
w32136 <= not w31856 and w32126;
w32137 <= not w32122 and w32136;
w32138 <= not w32123 and not w32126;
w32139 <= not w32137 and not w32138;
w32140 <= w3886 and not w32139;
w32141 <= not w32133 and w32140;
w32142 <= not w32135 and not w32141;
w32143 <= not b(22) and not w32142;
w32144 <= not w31855 and not w32134;
w32145 <= not w31865 and w32121;
w32146 <= not w32117 and w32145;
w32147 <= not w32118 and not w32121;
w32148 <= not w32146 and not w32147;
w32149 <= w3886 and not w32148;
w32150 <= not w32133 and w32149;
w32151 <= not w32144 and not w32150;
w32152 <= not b(21) and not w32151;
w32153 <= not w31864 and not w32134;
w32154 <= not w31874 and w32116;
w32155 <= not w32112 and w32154;
w32156 <= not w32113 and not w32116;
w32157 <= not w32155 and not w32156;
w32158 <= w3886 and not w32157;
w32159 <= not w32133 and w32158;
w32160 <= not w32153 and not w32159;
w32161 <= not b(20) and not w32160;
w32162 <= not w31873 and not w32134;
w32163 <= not w31883 and w32111;
w32164 <= not w32107 and w32163;
w32165 <= not w32108 and not w32111;
w32166 <= not w32164 and not w32165;
w32167 <= w3886 and not w32166;
w32168 <= not w32133 and w32167;
w32169 <= not w32162 and not w32168;
w32170 <= not b(19) and not w32169;
w32171 <= not w31882 and not w32134;
w32172 <= not w31892 and w32106;
w32173 <= not w32102 and w32172;
w32174 <= not w32103 and not w32106;
w32175 <= not w32173 and not w32174;
w32176 <= w3886 and not w32175;
w32177 <= not w32133 and w32176;
w32178 <= not w32171 and not w32177;
w32179 <= not b(18) and not w32178;
w32180 <= not w31891 and not w32134;
w32181 <= not w31901 and w32101;
w32182 <= not w32097 and w32181;
w32183 <= not w32098 and not w32101;
w32184 <= not w32182 and not w32183;
w32185 <= w3886 and not w32184;
w32186 <= not w32133 and w32185;
w32187 <= not w32180 and not w32186;
w32188 <= not b(17) and not w32187;
w32189 <= not w31900 and not w32134;
w32190 <= not w31910 and w32096;
w32191 <= not w32092 and w32190;
w32192 <= not w32093 and not w32096;
w32193 <= not w32191 and not w32192;
w32194 <= w3886 and not w32193;
w32195 <= not w32133 and w32194;
w32196 <= not w32189 and not w32195;
w32197 <= not b(16) and not w32196;
w32198 <= not w31909 and not w32134;
w32199 <= not w31919 and w32091;
w32200 <= not w32087 and w32199;
w32201 <= not w32088 and not w32091;
w32202 <= not w32200 and not w32201;
w32203 <= w3886 and not w32202;
w32204 <= not w32133 and w32203;
w32205 <= not w32198 and not w32204;
w32206 <= not b(15) and not w32205;
w32207 <= not w31918 and not w32134;
w32208 <= not w31928 and w32086;
w32209 <= not w32082 and w32208;
w32210 <= not w32083 and not w32086;
w32211 <= not w32209 and not w32210;
w32212 <= w3886 and not w32211;
w32213 <= not w32133 and w32212;
w32214 <= not w32207 and not w32213;
w32215 <= not b(14) and not w32214;
w32216 <= not w31927 and not w32134;
w32217 <= not w31937 and w32081;
w32218 <= not w32077 and w32217;
w32219 <= not w32078 and not w32081;
w32220 <= not w32218 and not w32219;
w32221 <= w3886 and not w32220;
w32222 <= not w32133 and w32221;
w32223 <= not w32216 and not w32222;
w32224 <= not b(13) and not w32223;
w32225 <= not w31936 and not w32134;
w32226 <= not w31946 and w32076;
w32227 <= not w32072 and w32226;
w32228 <= not w32073 and not w32076;
w32229 <= not w32227 and not w32228;
w32230 <= w3886 and not w32229;
w32231 <= not w32133 and w32230;
w32232 <= not w32225 and not w32231;
w32233 <= not b(12) and not w32232;
w32234 <= not w31945 and not w32134;
w32235 <= not w31955 and w32071;
w32236 <= not w32067 and w32235;
w32237 <= not w32068 and not w32071;
w32238 <= not w32236 and not w32237;
w32239 <= w3886 and not w32238;
w32240 <= not w32133 and w32239;
w32241 <= not w32234 and not w32240;
w32242 <= not b(11) and not w32241;
w32243 <= not w31954 and not w32134;
w32244 <= not w31964 and w32066;
w32245 <= not w32062 and w32244;
w32246 <= not w32063 and not w32066;
w32247 <= not w32245 and not w32246;
w32248 <= w3886 and not w32247;
w32249 <= not w32133 and w32248;
w32250 <= not w32243 and not w32249;
w32251 <= not b(10) and not w32250;
w32252 <= not w31963 and not w32134;
w32253 <= not w31973 and w32061;
w32254 <= not w32057 and w32253;
w32255 <= not w32058 and not w32061;
w32256 <= not w32254 and not w32255;
w32257 <= w3886 and not w32256;
w32258 <= not w32133 and w32257;
w32259 <= not w32252 and not w32258;
w32260 <= not b(9) and not w32259;
w32261 <= not w31972 and not w32134;
w32262 <= not w31982 and w32056;
w32263 <= not w32052 and w32262;
w32264 <= not w32053 and not w32056;
w32265 <= not w32263 and not w32264;
w32266 <= w3886 and not w32265;
w32267 <= not w32133 and w32266;
w32268 <= not w32261 and not w32267;
w32269 <= not b(8) and not w32268;
w32270 <= not w31981 and not w32134;
w32271 <= not w31991 and w32051;
w32272 <= not w32047 and w32271;
w32273 <= not w32048 and not w32051;
w32274 <= not w32272 and not w32273;
w32275 <= w3886 and not w32274;
w32276 <= not w32133 and w32275;
w32277 <= not w32270 and not w32276;
w32278 <= not b(7) and not w32277;
w32279 <= not w31990 and not w32134;
w32280 <= not w32000 and w32046;
w32281 <= not w32042 and w32280;
w32282 <= not w32043 and not w32046;
w32283 <= not w32281 and not w32282;
w32284 <= w3886 and not w32283;
w32285 <= not w32133 and w32284;
w32286 <= not w32279 and not w32285;
w32287 <= not b(6) and not w32286;
w32288 <= not w31999 and not w32134;
w32289 <= not w32009 and w32041;
w32290 <= not w32037 and w32289;
w32291 <= not w32038 and not w32041;
w32292 <= not w32290 and not w32291;
w32293 <= w3886 and not w32292;
w32294 <= not w32133 and w32293;
w32295 <= not w32288 and not w32294;
w32296 <= not b(5) and not w32295;
w32297 <= not w32008 and not w32134;
w32298 <= not w32017 and w32036;
w32299 <= not w32032 and w32298;
w32300 <= not w32033 and not w32036;
w32301 <= not w32299 and not w32300;
w32302 <= w3886 and not w32301;
w32303 <= not w32133 and w32302;
w32304 <= not w32297 and not w32303;
w32305 <= not b(4) and not w32304;
w32306 <= not w32016 and not w32134;
w32307 <= not w32027 and w32031;
w32308 <= not w32026 and w32307;
w32309 <= not w32028 and not w32031;
w32310 <= not w32308 and not w32309;
w32311 <= w3886 and not w32310;
w32312 <= not w32133 and w32311;
w32313 <= not w32306 and not w32312;
w32314 <= not b(3) and not w32313;
w32315 <= not w32021 and not w32134;
w32316 <= w3774 and not w32024;
w32317 <= not w32022 and w32316;
w32318 <= w3886 and not w32317;
w32319 <= not w32026 and w32318;
w32320 <= not w32133 and w32319;
w32321 <= not w32315 and not w32320;
w32322 <= not b(2) and not w32321;
w32323 <= w4080 and not w32133;
w32324 <= a(41) and not w32323;
w32325 <= w4087 and not w32133;
w32326 <= not w32324 and not w32325;
w32327 <= b(1) and not w32326;
w32328 <= not b(1) and not w32325;
w32329 <= not w32324 and w32328;
w32330 <= not w32327 and not w32329;
w32331 <= not w4094 and not w32330;
w32332 <= not b(1) and not w32326;
w32333 <= not w32331 and not w32332;
w32334 <= b(2) and not w32320;
w32335 <= not w32315 and w32334;
w32336 <= not w32322 and not w32335;
w32337 <= not w32333 and w32336;
w32338 <= not w32322 and not w32337;
w32339 <= b(3) and not w32312;
w32340 <= not w32306 and w32339;
w32341 <= not w32314 and not w32340;
w32342 <= not w32338 and w32341;
w32343 <= not w32314 and not w32342;
w32344 <= b(4) and not w32303;
w32345 <= not w32297 and w32344;
w32346 <= not w32305 and not w32345;
w32347 <= not w32343 and w32346;
w32348 <= not w32305 and not w32347;
w32349 <= b(5) and not w32294;
w32350 <= not w32288 and w32349;
w32351 <= not w32296 and not w32350;
w32352 <= not w32348 and w32351;
w32353 <= not w32296 and not w32352;
w32354 <= b(6) and not w32285;
w32355 <= not w32279 and w32354;
w32356 <= not w32287 and not w32355;
w32357 <= not w32353 and w32356;
w32358 <= not w32287 and not w32357;
w32359 <= b(7) and not w32276;
w32360 <= not w32270 and w32359;
w32361 <= not w32278 and not w32360;
w32362 <= not w32358 and w32361;
w32363 <= not w32278 and not w32362;
w32364 <= b(8) and not w32267;
w32365 <= not w32261 and w32364;
w32366 <= not w32269 and not w32365;
w32367 <= not w32363 and w32366;
w32368 <= not w32269 and not w32367;
w32369 <= b(9) and not w32258;
w32370 <= not w32252 and w32369;
w32371 <= not w32260 and not w32370;
w32372 <= not w32368 and w32371;
w32373 <= not w32260 and not w32372;
w32374 <= b(10) and not w32249;
w32375 <= not w32243 and w32374;
w32376 <= not w32251 and not w32375;
w32377 <= not w32373 and w32376;
w32378 <= not w32251 and not w32377;
w32379 <= b(11) and not w32240;
w32380 <= not w32234 and w32379;
w32381 <= not w32242 and not w32380;
w32382 <= not w32378 and w32381;
w32383 <= not w32242 and not w32382;
w32384 <= b(12) and not w32231;
w32385 <= not w32225 and w32384;
w32386 <= not w32233 and not w32385;
w32387 <= not w32383 and w32386;
w32388 <= not w32233 and not w32387;
w32389 <= b(13) and not w32222;
w32390 <= not w32216 and w32389;
w32391 <= not w32224 and not w32390;
w32392 <= not w32388 and w32391;
w32393 <= not w32224 and not w32392;
w32394 <= b(14) and not w32213;
w32395 <= not w32207 and w32394;
w32396 <= not w32215 and not w32395;
w32397 <= not w32393 and w32396;
w32398 <= not w32215 and not w32397;
w32399 <= b(15) and not w32204;
w32400 <= not w32198 and w32399;
w32401 <= not w32206 and not w32400;
w32402 <= not w32398 and w32401;
w32403 <= not w32206 and not w32402;
w32404 <= b(16) and not w32195;
w32405 <= not w32189 and w32404;
w32406 <= not w32197 and not w32405;
w32407 <= not w32403 and w32406;
w32408 <= not w32197 and not w32407;
w32409 <= b(17) and not w32186;
w32410 <= not w32180 and w32409;
w32411 <= not w32188 and not w32410;
w32412 <= not w32408 and w32411;
w32413 <= not w32188 and not w32412;
w32414 <= b(18) and not w32177;
w32415 <= not w32171 and w32414;
w32416 <= not w32179 and not w32415;
w32417 <= not w32413 and w32416;
w32418 <= not w32179 and not w32417;
w32419 <= b(19) and not w32168;
w32420 <= not w32162 and w32419;
w32421 <= not w32170 and not w32420;
w32422 <= not w32418 and w32421;
w32423 <= not w32170 and not w32422;
w32424 <= b(20) and not w32159;
w32425 <= not w32153 and w32424;
w32426 <= not w32161 and not w32425;
w32427 <= not w32423 and w32426;
w32428 <= not w32161 and not w32427;
w32429 <= b(21) and not w32150;
w32430 <= not w32144 and w32429;
w32431 <= not w32152 and not w32430;
w32432 <= not w32428 and w32431;
w32433 <= not w32152 and not w32432;
w32434 <= b(22) and not w32141;
w32435 <= not w32135 and w32434;
w32436 <= not w32143 and not w32435;
w32437 <= not w32433 and w32436;
w32438 <= not w32143 and not w32437;
w32439 <= not w31845 and not w32134;
w32440 <= not w31847 and w32131;
w32441 <= not w32127 and w32440;
w32442 <= not w32128 and not w32131;
w32443 <= not w32441 and not w32442;
w32444 <= w32134 and not w32443;
w32445 <= not w32439 and not w32444;
w32446 <= not b(23) and not w32445;
w32447 <= b(23) and not w32439;
w32448 <= not w32444 and w32447;
w32449 <= w4214 and not w32448;
w32450 <= not w32446 and w32449;
w32451 <= not w32438 and w32450;
w32452 <= w3886 and not w32445;
w32453 <= not w32451 and not w32452;
w32454 <= not w32152 and w32436;
w32455 <= not w32432 and w32454;
w32456 <= not w32433 and not w32436;
w32457 <= not w32455 and not w32456;
w32458 <= not w32453 and not w32457;
w32459 <= not w32142 and not w32452;
w32460 <= not w32451 and w32459;
w32461 <= not w32458 and not w32460;
w32462 <= not w32143 and not w32448;
w32463 <= not w32446 and w32462;
w32464 <= not w32437 and w32463;
w32465 <= not w32446 and not w32448;
w32466 <= not w32438 and not w32465;
w32467 <= not w32464 and not w32466;
w32468 <= not w32453 and not w32467;
w32469 <= not w32445 and not w32452;
w32470 <= not w32451 and w32469;
w32471 <= not w32468 and not w32470;
w32472 <= not b(24) and not w32471;
w32473 <= not b(23) and not w32461;
w32474 <= not w32161 and w32431;
w32475 <= not w32427 and w32474;
w32476 <= not w32428 and not w32431;
w32477 <= not w32475 and not w32476;
w32478 <= not w32453 and not w32477;
w32479 <= not w32151 and not w32452;
w32480 <= not w32451 and w32479;
w32481 <= not w32478 and not w32480;
w32482 <= not b(22) and not w32481;
w32483 <= not w32170 and w32426;
w32484 <= not w32422 and w32483;
w32485 <= not w32423 and not w32426;
w32486 <= not w32484 and not w32485;
w32487 <= not w32453 and not w32486;
w32488 <= not w32160 and not w32452;
w32489 <= not w32451 and w32488;
w32490 <= not w32487 and not w32489;
w32491 <= not b(21) and not w32490;
w32492 <= not w32179 and w32421;
w32493 <= not w32417 and w32492;
w32494 <= not w32418 and not w32421;
w32495 <= not w32493 and not w32494;
w32496 <= not w32453 and not w32495;
w32497 <= not w32169 and not w32452;
w32498 <= not w32451 and w32497;
w32499 <= not w32496 and not w32498;
w32500 <= not b(20) and not w32499;
w32501 <= not w32188 and w32416;
w32502 <= not w32412 and w32501;
w32503 <= not w32413 and not w32416;
w32504 <= not w32502 and not w32503;
w32505 <= not w32453 and not w32504;
w32506 <= not w32178 and not w32452;
w32507 <= not w32451 and w32506;
w32508 <= not w32505 and not w32507;
w32509 <= not b(19) and not w32508;
w32510 <= not w32197 and w32411;
w32511 <= not w32407 and w32510;
w32512 <= not w32408 and not w32411;
w32513 <= not w32511 and not w32512;
w32514 <= not w32453 and not w32513;
w32515 <= not w32187 and not w32452;
w32516 <= not w32451 and w32515;
w32517 <= not w32514 and not w32516;
w32518 <= not b(18) and not w32517;
w32519 <= not w32206 and w32406;
w32520 <= not w32402 and w32519;
w32521 <= not w32403 and not w32406;
w32522 <= not w32520 and not w32521;
w32523 <= not w32453 and not w32522;
w32524 <= not w32196 and not w32452;
w32525 <= not w32451 and w32524;
w32526 <= not w32523 and not w32525;
w32527 <= not b(17) and not w32526;
w32528 <= not w32215 and w32401;
w32529 <= not w32397 and w32528;
w32530 <= not w32398 and not w32401;
w32531 <= not w32529 and not w32530;
w32532 <= not w32453 and not w32531;
w32533 <= not w32205 and not w32452;
w32534 <= not w32451 and w32533;
w32535 <= not w32532 and not w32534;
w32536 <= not b(16) and not w32535;
w32537 <= not w32224 and w32396;
w32538 <= not w32392 and w32537;
w32539 <= not w32393 and not w32396;
w32540 <= not w32538 and not w32539;
w32541 <= not w32453 and not w32540;
w32542 <= not w32214 and not w32452;
w32543 <= not w32451 and w32542;
w32544 <= not w32541 and not w32543;
w32545 <= not b(15) and not w32544;
w32546 <= not w32233 and w32391;
w32547 <= not w32387 and w32546;
w32548 <= not w32388 and not w32391;
w32549 <= not w32547 and not w32548;
w32550 <= not w32453 and not w32549;
w32551 <= not w32223 and not w32452;
w32552 <= not w32451 and w32551;
w32553 <= not w32550 and not w32552;
w32554 <= not b(14) and not w32553;
w32555 <= not w32242 and w32386;
w32556 <= not w32382 and w32555;
w32557 <= not w32383 and not w32386;
w32558 <= not w32556 and not w32557;
w32559 <= not w32453 and not w32558;
w32560 <= not w32232 and not w32452;
w32561 <= not w32451 and w32560;
w32562 <= not w32559 and not w32561;
w32563 <= not b(13) and not w32562;
w32564 <= not w32251 and w32381;
w32565 <= not w32377 and w32564;
w32566 <= not w32378 and not w32381;
w32567 <= not w32565 and not w32566;
w32568 <= not w32453 and not w32567;
w32569 <= not w32241 and not w32452;
w32570 <= not w32451 and w32569;
w32571 <= not w32568 and not w32570;
w32572 <= not b(12) and not w32571;
w32573 <= not w32260 and w32376;
w32574 <= not w32372 and w32573;
w32575 <= not w32373 and not w32376;
w32576 <= not w32574 and not w32575;
w32577 <= not w32453 and not w32576;
w32578 <= not w32250 and not w32452;
w32579 <= not w32451 and w32578;
w32580 <= not w32577 and not w32579;
w32581 <= not b(11) and not w32580;
w32582 <= not w32269 and w32371;
w32583 <= not w32367 and w32582;
w32584 <= not w32368 and not w32371;
w32585 <= not w32583 and not w32584;
w32586 <= not w32453 and not w32585;
w32587 <= not w32259 and not w32452;
w32588 <= not w32451 and w32587;
w32589 <= not w32586 and not w32588;
w32590 <= not b(10) and not w32589;
w32591 <= not w32278 and w32366;
w32592 <= not w32362 and w32591;
w32593 <= not w32363 and not w32366;
w32594 <= not w32592 and not w32593;
w32595 <= not w32453 and not w32594;
w32596 <= not w32268 and not w32452;
w32597 <= not w32451 and w32596;
w32598 <= not w32595 and not w32597;
w32599 <= not b(9) and not w32598;
w32600 <= not w32287 and w32361;
w32601 <= not w32357 and w32600;
w32602 <= not w32358 and not w32361;
w32603 <= not w32601 and not w32602;
w32604 <= not w32453 and not w32603;
w32605 <= not w32277 and not w32452;
w32606 <= not w32451 and w32605;
w32607 <= not w32604 and not w32606;
w32608 <= not b(8) and not w32607;
w32609 <= not w32296 and w32356;
w32610 <= not w32352 and w32609;
w32611 <= not w32353 and not w32356;
w32612 <= not w32610 and not w32611;
w32613 <= not w32453 and not w32612;
w32614 <= not w32286 and not w32452;
w32615 <= not w32451 and w32614;
w32616 <= not w32613 and not w32615;
w32617 <= not b(7) and not w32616;
w32618 <= not w32305 and w32351;
w32619 <= not w32347 and w32618;
w32620 <= not w32348 and not w32351;
w32621 <= not w32619 and not w32620;
w32622 <= not w32453 and not w32621;
w32623 <= not w32295 and not w32452;
w32624 <= not w32451 and w32623;
w32625 <= not w32622 and not w32624;
w32626 <= not b(6) and not w32625;
w32627 <= not w32314 and w32346;
w32628 <= not w32342 and w32627;
w32629 <= not w32343 and not w32346;
w32630 <= not w32628 and not w32629;
w32631 <= not w32453 and not w32630;
w32632 <= not w32304 and not w32452;
w32633 <= not w32451 and w32632;
w32634 <= not w32631 and not w32633;
w32635 <= not b(5) and not w32634;
w32636 <= not w32322 and w32341;
w32637 <= not w32337 and w32636;
w32638 <= not w32338 and not w32341;
w32639 <= not w32637 and not w32638;
w32640 <= not w32453 and not w32639;
w32641 <= not w32313 and not w32452;
w32642 <= not w32451 and w32641;
w32643 <= not w32640 and not w32642;
w32644 <= not b(4) and not w32643;
w32645 <= not w32332 and w32336;
w32646 <= not w32331 and w32645;
w32647 <= not w32333 and not w32336;
w32648 <= not w32646 and not w32647;
w32649 <= not w32453 and not w32648;
w32650 <= not w32321 and not w32452;
w32651 <= not w32451 and w32650;
w32652 <= not w32649 and not w32651;
w32653 <= not b(3) and not w32652;
w32654 <= w4094 and not w32329;
w32655 <= not w32327 and w32654;
w32656 <= not w32331 and not w32655;
w32657 <= not w32453 and w32656;
w32658 <= not w32326 and not w32452;
w32659 <= not w32451 and w32658;
w32660 <= not w32657 and not w32659;
w32661 <= not b(2) and not w32660;
w32662 <= b(0) and not w32453;
w32663 <= a(40) and not w32662;
w32664 <= w4094 and not w32453;
w32665 <= not w32663 and not w32664;
w32666 <= b(1) and not w32665;
w32667 <= not b(1) and not w32664;
w32668 <= not w32663 and w32667;
w32669 <= not w32666 and not w32668;
w32670 <= not w4436 and not w32669;
w32671 <= not b(1) and not w32665;
w32672 <= not w32670 and not w32671;
w32673 <= b(2) and not w32659;
w32674 <= not w32657 and w32673;
w32675 <= not w32661 and not w32674;
w32676 <= not w32672 and w32675;
w32677 <= not w32661 and not w32676;
w32678 <= b(3) and not w32651;
w32679 <= not w32649 and w32678;
w32680 <= not w32653 and not w32679;
w32681 <= not w32677 and w32680;
w32682 <= not w32653 and not w32681;
w32683 <= b(4) and not w32642;
w32684 <= not w32640 and w32683;
w32685 <= not w32644 and not w32684;
w32686 <= not w32682 and w32685;
w32687 <= not w32644 and not w32686;
w32688 <= b(5) and not w32633;
w32689 <= not w32631 and w32688;
w32690 <= not w32635 and not w32689;
w32691 <= not w32687 and w32690;
w32692 <= not w32635 and not w32691;
w32693 <= b(6) and not w32624;
w32694 <= not w32622 and w32693;
w32695 <= not w32626 and not w32694;
w32696 <= not w32692 and w32695;
w32697 <= not w32626 and not w32696;
w32698 <= b(7) and not w32615;
w32699 <= not w32613 and w32698;
w32700 <= not w32617 and not w32699;
w32701 <= not w32697 and w32700;
w32702 <= not w32617 and not w32701;
w32703 <= b(8) and not w32606;
w32704 <= not w32604 and w32703;
w32705 <= not w32608 and not w32704;
w32706 <= not w32702 and w32705;
w32707 <= not w32608 and not w32706;
w32708 <= b(9) and not w32597;
w32709 <= not w32595 and w32708;
w32710 <= not w32599 and not w32709;
w32711 <= not w32707 and w32710;
w32712 <= not w32599 and not w32711;
w32713 <= b(10) and not w32588;
w32714 <= not w32586 and w32713;
w32715 <= not w32590 and not w32714;
w32716 <= not w32712 and w32715;
w32717 <= not w32590 and not w32716;
w32718 <= b(11) and not w32579;
w32719 <= not w32577 and w32718;
w32720 <= not w32581 and not w32719;
w32721 <= not w32717 and w32720;
w32722 <= not w32581 and not w32721;
w32723 <= b(12) and not w32570;
w32724 <= not w32568 and w32723;
w32725 <= not w32572 and not w32724;
w32726 <= not w32722 and w32725;
w32727 <= not w32572 and not w32726;
w32728 <= b(13) and not w32561;
w32729 <= not w32559 and w32728;
w32730 <= not w32563 and not w32729;
w32731 <= not w32727 and w32730;
w32732 <= not w32563 and not w32731;
w32733 <= b(14) and not w32552;
w32734 <= not w32550 and w32733;
w32735 <= not w32554 and not w32734;
w32736 <= not w32732 and w32735;
w32737 <= not w32554 and not w32736;
w32738 <= b(15) and not w32543;
w32739 <= not w32541 and w32738;
w32740 <= not w32545 and not w32739;
w32741 <= not w32737 and w32740;
w32742 <= not w32545 and not w32741;
w32743 <= b(16) and not w32534;
w32744 <= not w32532 and w32743;
w32745 <= not w32536 and not w32744;
w32746 <= not w32742 and w32745;
w32747 <= not w32536 and not w32746;
w32748 <= b(17) and not w32525;
w32749 <= not w32523 and w32748;
w32750 <= not w32527 and not w32749;
w32751 <= not w32747 and w32750;
w32752 <= not w32527 and not w32751;
w32753 <= b(18) and not w32516;
w32754 <= not w32514 and w32753;
w32755 <= not w32518 and not w32754;
w32756 <= not w32752 and w32755;
w32757 <= not w32518 and not w32756;
w32758 <= b(19) and not w32507;
w32759 <= not w32505 and w32758;
w32760 <= not w32509 and not w32759;
w32761 <= not w32757 and w32760;
w32762 <= not w32509 and not w32761;
w32763 <= b(20) and not w32498;
w32764 <= not w32496 and w32763;
w32765 <= not w32500 and not w32764;
w32766 <= not w32762 and w32765;
w32767 <= not w32500 and not w32766;
w32768 <= b(21) and not w32489;
w32769 <= not w32487 and w32768;
w32770 <= not w32491 and not w32769;
w32771 <= not w32767 and w32770;
w32772 <= not w32491 and not w32771;
w32773 <= b(22) and not w32480;
w32774 <= not w32478 and w32773;
w32775 <= not w32482 and not w32774;
w32776 <= not w32772 and w32775;
w32777 <= not w32482 and not w32776;
w32778 <= b(23) and not w32460;
w32779 <= not w32458 and w32778;
w32780 <= not w32473 and not w32779;
w32781 <= not w32777 and w32780;
w32782 <= not w32473 and not w32781;
w32783 <= b(24) and not w32470;
w32784 <= not w32468 and w32783;
w32785 <= not w32472 and not w32784;
w32786 <= not w32782 and w32785;
w32787 <= not w32472 and not w32786;
w32788 <= w4556 and not w32787;
w32789 <= not w32461 and not w32788;
w32790 <= not w32482 and w32780;
w32791 <= not w32776 and w32790;
w32792 <= not w32777 and not w32780;
w32793 <= not w32791 and not w32792;
w32794 <= w4556 and not w32793;
w32795 <= not w32787 and w32794;
w32796 <= not w32789 and not w32795;
w32797 <= not w32471 and not w32788;
w32798 <= not w32473 and w32785;
w32799 <= not w32781 and w32798;
w32800 <= not w32782 and not w32785;
w32801 <= not w32799 and not w32800;
w32802 <= w32788 and not w32801;
w32803 <= not w32797 and not w32802;
w32804 <= not b(25) and not w32803;
w32805 <= not b(24) and not w32796;
w32806 <= not w32481 and not w32788;
w32807 <= not w32491 and w32775;
w32808 <= not w32771 and w32807;
w32809 <= not w32772 and not w32775;
w32810 <= not w32808 and not w32809;
w32811 <= w4556 and not w32810;
w32812 <= not w32787 and w32811;
w32813 <= not w32806 and not w32812;
w32814 <= not b(23) and not w32813;
w32815 <= not w32490 and not w32788;
w32816 <= not w32500 and w32770;
w32817 <= not w32766 and w32816;
w32818 <= not w32767 and not w32770;
w32819 <= not w32817 and not w32818;
w32820 <= w4556 and not w32819;
w32821 <= not w32787 and w32820;
w32822 <= not w32815 and not w32821;
w32823 <= not b(22) and not w32822;
w32824 <= not w32499 and not w32788;
w32825 <= not w32509 and w32765;
w32826 <= not w32761 and w32825;
w32827 <= not w32762 and not w32765;
w32828 <= not w32826 and not w32827;
w32829 <= w4556 and not w32828;
w32830 <= not w32787 and w32829;
w32831 <= not w32824 and not w32830;
w32832 <= not b(21) and not w32831;
w32833 <= not w32508 and not w32788;
w32834 <= not w32518 and w32760;
w32835 <= not w32756 and w32834;
w32836 <= not w32757 and not w32760;
w32837 <= not w32835 and not w32836;
w32838 <= w4556 and not w32837;
w32839 <= not w32787 and w32838;
w32840 <= not w32833 and not w32839;
w32841 <= not b(20) and not w32840;
w32842 <= not w32517 and not w32788;
w32843 <= not w32527 and w32755;
w32844 <= not w32751 and w32843;
w32845 <= not w32752 and not w32755;
w32846 <= not w32844 and not w32845;
w32847 <= w4556 and not w32846;
w32848 <= not w32787 and w32847;
w32849 <= not w32842 and not w32848;
w32850 <= not b(19) and not w32849;
w32851 <= not w32526 and not w32788;
w32852 <= not w32536 and w32750;
w32853 <= not w32746 and w32852;
w32854 <= not w32747 and not w32750;
w32855 <= not w32853 and not w32854;
w32856 <= w4556 and not w32855;
w32857 <= not w32787 and w32856;
w32858 <= not w32851 and not w32857;
w32859 <= not b(18) and not w32858;
w32860 <= not w32535 and not w32788;
w32861 <= not w32545 and w32745;
w32862 <= not w32741 and w32861;
w32863 <= not w32742 and not w32745;
w32864 <= not w32862 and not w32863;
w32865 <= w4556 and not w32864;
w32866 <= not w32787 and w32865;
w32867 <= not w32860 and not w32866;
w32868 <= not b(17) and not w32867;
w32869 <= not w32544 and not w32788;
w32870 <= not w32554 and w32740;
w32871 <= not w32736 and w32870;
w32872 <= not w32737 and not w32740;
w32873 <= not w32871 and not w32872;
w32874 <= w4556 and not w32873;
w32875 <= not w32787 and w32874;
w32876 <= not w32869 and not w32875;
w32877 <= not b(16) and not w32876;
w32878 <= not w32553 and not w32788;
w32879 <= not w32563 and w32735;
w32880 <= not w32731 and w32879;
w32881 <= not w32732 and not w32735;
w32882 <= not w32880 and not w32881;
w32883 <= w4556 and not w32882;
w32884 <= not w32787 and w32883;
w32885 <= not w32878 and not w32884;
w32886 <= not b(15) and not w32885;
w32887 <= not w32562 and not w32788;
w32888 <= not w32572 and w32730;
w32889 <= not w32726 and w32888;
w32890 <= not w32727 and not w32730;
w32891 <= not w32889 and not w32890;
w32892 <= w4556 and not w32891;
w32893 <= not w32787 and w32892;
w32894 <= not w32887 and not w32893;
w32895 <= not b(14) and not w32894;
w32896 <= not w32571 and not w32788;
w32897 <= not w32581 and w32725;
w32898 <= not w32721 and w32897;
w32899 <= not w32722 and not w32725;
w32900 <= not w32898 and not w32899;
w32901 <= w4556 and not w32900;
w32902 <= not w32787 and w32901;
w32903 <= not w32896 and not w32902;
w32904 <= not b(13) and not w32903;
w32905 <= not w32580 and not w32788;
w32906 <= not w32590 and w32720;
w32907 <= not w32716 and w32906;
w32908 <= not w32717 and not w32720;
w32909 <= not w32907 and not w32908;
w32910 <= w4556 and not w32909;
w32911 <= not w32787 and w32910;
w32912 <= not w32905 and not w32911;
w32913 <= not b(12) and not w32912;
w32914 <= not w32589 and not w32788;
w32915 <= not w32599 and w32715;
w32916 <= not w32711 and w32915;
w32917 <= not w32712 and not w32715;
w32918 <= not w32916 and not w32917;
w32919 <= w4556 and not w32918;
w32920 <= not w32787 and w32919;
w32921 <= not w32914 and not w32920;
w32922 <= not b(11) and not w32921;
w32923 <= not w32598 and not w32788;
w32924 <= not w32608 and w32710;
w32925 <= not w32706 and w32924;
w32926 <= not w32707 and not w32710;
w32927 <= not w32925 and not w32926;
w32928 <= w4556 and not w32927;
w32929 <= not w32787 and w32928;
w32930 <= not w32923 and not w32929;
w32931 <= not b(10) and not w32930;
w32932 <= not w32607 and not w32788;
w32933 <= not w32617 and w32705;
w32934 <= not w32701 and w32933;
w32935 <= not w32702 and not w32705;
w32936 <= not w32934 and not w32935;
w32937 <= w4556 and not w32936;
w32938 <= not w32787 and w32937;
w32939 <= not w32932 and not w32938;
w32940 <= not b(9) and not w32939;
w32941 <= not w32616 and not w32788;
w32942 <= not w32626 and w32700;
w32943 <= not w32696 and w32942;
w32944 <= not w32697 and not w32700;
w32945 <= not w32943 and not w32944;
w32946 <= w4556 and not w32945;
w32947 <= not w32787 and w32946;
w32948 <= not w32941 and not w32947;
w32949 <= not b(8) and not w32948;
w32950 <= not w32625 and not w32788;
w32951 <= not w32635 and w32695;
w32952 <= not w32691 and w32951;
w32953 <= not w32692 and not w32695;
w32954 <= not w32952 and not w32953;
w32955 <= w4556 and not w32954;
w32956 <= not w32787 and w32955;
w32957 <= not w32950 and not w32956;
w32958 <= not b(7) and not w32957;
w32959 <= not w32634 and not w32788;
w32960 <= not w32644 and w32690;
w32961 <= not w32686 and w32960;
w32962 <= not w32687 and not w32690;
w32963 <= not w32961 and not w32962;
w32964 <= w4556 and not w32963;
w32965 <= not w32787 and w32964;
w32966 <= not w32959 and not w32965;
w32967 <= not b(6) and not w32966;
w32968 <= not w32643 and not w32788;
w32969 <= not w32653 and w32685;
w32970 <= not w32681 and w32969;
w32971 <= not w32682 and not w32685;
w32972 <= not w32970 and not w32971;
w32973 <= w4556 and not w32972;
w32974 <= not w32787 and w32973;
w32975 <= not w32968 and not w32974;
w32976 <= not b(5) and not w32975;
w32977 <= not w32652 and not w32788;
w32978 <= not w32661 and w32680;
w32979 <= not w32676 and w32978;
w32980 <= not w32677 and not w32680;
w32981 <= not w32979 and not w32980;
w32982 <= w4556 and not w32981;
w32983 <= not w32787 and w32982;
w32984 <= not w32977 and not w32983;
w32985 <= not b(4) and not w32984;
w32986 <= not w32660 and not w32788;
w32987 <= not w32671 and w32675;
w32988 <= not w32670 and w32987;
w32989 <= not w32672 and not w32675;
w32990 <= not w32988 and not w32989;
w32991 <= w4556 and not w32990;
w32992 <= not w32787 and w32991;
w32993 <= not w32986 and not w32992;
w32994 <= not b(3) and not w32993;
w32995 <= not w32665 and not w32788;
w32996 <= w4436 and not w32668;
w32997 <= not w32666 and w32996;
w32998 <= w4556 and not w32997;
w32999 <= not w32670 and w32998;
w33000 <= not w32787 and w32999;
w33001 <= not w32995 and not w33000;
w33002 <= not b(2) and not w33001;
w33003 <= w4776 and not w32787;
w33004 <= a(39) and not w33003;
w33005 <= w4782 and not w32787;
w33006 <= not w33004 and not w33005;
w33007 <= b(1) and not w33006;
w33008 <= not b(1) and not w33005;
w33009 <= not w33004 and w33008;
w33010 <= not w33007 and not w33009;
w33011 <= not w4789 and not w33010;
w33012 <= not b(1) and not w33006;
w33013 <= not w33011 and not w33012;
w33014 <= b(2) and not w33000;
w33015 <= not w32995 and w33014;
w33016 <= not w33002 and not w33015;
w33017 <= not w33013 and w33016;
w33018 <= not w33002 and not w33017;
w33019 <= b(3) and not w32992;
w33020 <= not w32986 and w33019;
w33021 <= not w32994 and not w33020;
w33022 <= not w33018 and w33021;
w33023 <= not w32994 and not w33022;
w33024 <= b(4) and not w32983;
w33025 <= not w32977 and w33024;
w33026 <= not w32985 and not w33025;
w33027 <= not w33023 and w33026;
w33028 <= not w32985 and not w33027;
w33029 <= b(5) and not w32974;
w33030 <= not w32968 and w33029;
w33031 <= not w32976 and not w33030;
w33032 <= not w33028 and w33031;
w33033 <= not w32976 and not w33032;
w33034 <= b(6) and not w32965;
w33035 <= not w32959 and w33034;
w33036 <= not w32967 and not w33035;
w33037 <= not w33033 and w33036;
w33038 <= not w32967 and not w33037;
w33039 <= b(7) and not w32956;
w33040 <= not w32950 and w33039;
w33041 <= not w32958 and not w33040;
w33042 <= not w33038 and w33041;
w33043 <= not w32958 and not w33042;
w33044 <= b(8) and not w32947;
w33045 <= not w32941 and w33044;
w33046 <= not w32949 and not w33045;
w33047 <= not w33043 and w33046;
w33048 <= not w32949 and not w33047;
w33049 <= b(9) and not w32938;
w33050 <= not w32932 and w33049;
w33051 <= not w32940 and not w33050;
w33052 <= not w33048 and w33051;
w33053 <= not w32940 and not w33052;
w33054 <= b(10) and not w32929;
w33055 <= not w32923 and w33054;
w33056 <= not w32931 and not w33055;
w33057 <= not w33053 and w33056;
w33058 <= not w32931 and not w33057;
w33059 <= b(11) and not w32920;
w33060 <= not w32914 and w33059;
w33061 <= not w32922 and not w33060;
w33062 <= not w33058 and w33061;
w33063 <= not w32922 and not w33062;
w33064 <= b(12) and not w32911;
w33065 <= not w32905 and w33064;
w33066 <= not w32913 and not w33065;
w33067 <= not w33063 and w33066;
w33068 <= not w32913 and not w33067;
w33069 <= b(13) and not w32902;
w33070 <= not w32896 and w33069;
w33071 <= not w32904 and not w33070;
w33072 <= not w33068 and w33071;
w33073 <= not w32904 and not w33072;
w33074 <= b(14) and not w32893;
w33075 <= not w32887 and w33074;
w33076 <= not w32895 and not w33075;
w33077 <= not w33073 and w33076;
w33078 <= not w32895 and not w33077;
w33079 <= b(15) and not w32884;
w33080 <= not w32878 and w33079;
w33081 <= not w32886 and not w33080;
w33082 <= not w33078 and w33081;
w33083 <= not w32886 and not w33082;
w33084 <= b(16) and not w32875;
w33085 <= not w32869 and w33084;
w33086 <= not w32877 and not w33085;
w33087 <= not w33083 and w33086;
w33088 <= not w32877 and not w33087;
w33089 <= b(17) and not w32866;
w33090 <= not w32860 and w33089;
w33091 <= not w32868 and not w33090;
w33092 <= not w33088 and w33091;
w33093 <= not w32868 and not w33092;
w33094 <= b(18) and not w32857;
w33095 <= not w32851 and w33094;
w33096 <= not w32859 and not w33095;
w33097 <= not w33093 and w33096;
w33098 <= not w32859 and not w33097;
w33099 <= b(19) and not w32848;
w33100 <= not w32842 and w33099;
w33101 <= not w32850 and not w33100;
w33102 <= not w33098 and w33101;
w33103 <= not w32850 and not w33102;
w33104 <= b(20) and not w32839;
w33105 <= not w32833 and w33104;
w33106 <= not w32841 and not w33105;
w33107 <= not w33103 and w33106;
w33108 <= not w32841 and not w33107;
w33109 <= b(21) and not w32830;
w33110 <= not w32824 and w33109;
w33111 <= not w32832 and not w33110;
w33112 <= not w33108 and w33111;
w33113 <= not w32832 and not w33112;
w33114 <= b(22) and not w32821;
w33115 <= not w32815 and w33114;
w33116 <= not w32823 and not w33115;
w33117 <= not w33113 and w33116;
w33118 <= not w32823 and not w33117;
w33119 <= b(23) and not w32812;
w33120 <= not w32806 and w33119;
w33121 <= not w32814 and not w33120;
w33122 <= not w33118 and w33121;
w33123 <= not w32814 and not w33122;
w33124 <= b(24) and not w32795;
w33125 <= not w32789 and w33124;
w33126 <= not w32805 and not w33125;
w33127 <= not w33123 and w33126;
w33128 <= not w32805 and not w33127;
w33129 <= b(25) and not w32797;
w33130 <= not w32802 and w33129;
w33131 <= not w32804 and not w33130;
w33132 <= not w33128 and w33131;
w33133 <= not w32804 and not w33132;
w33134 <= w4915 and not w33133;
w33135 <= not w32796 and not w33134;
w33136 <= not w32814 and w33126;
w33137 <= not w33122 and w33136;
w33138 <= not w33123 and not w33126;
w33139 <= not w33137 and not w33138;
w33140 <= w4915 and not w33139;
w33141 <= not w33133 and w33140;
w33142 <= not w33135 and not w33141;
w33143 <= not b(25) and not w33142;
w33144 <= not w32813 and not w33134;
w33145 <= not w32823 and w33121;
w33146 <= not w33117 and w33145;
w33147 <= not w33118 and not w33121;
w33148 <= not w33146 and not w33147;
w33149 <= w4915 and not w33148;
w33150 <= not w33133 and w33149;
w33151 <= not w33144 and not w33150;
w33152 <= not b(24) and not w33151;
w33153 <= not w32822 and not w33134;
w33154 <= not w32832 and w33116;
w33155 <= not w33112 and w33154;
w33156 <= not w33113 and not w33116;
w33157 <= not w33155 and not w33156;
w33158 <= w4915 and not w33157;
w33159 <= not w33133 and w33158;
w33160 <= not w33153 and not w33159;
w33161 <= not b(23) and not w33160;
w33162 <= not w32831 and not w33134;
w33163 <= not w32841 and w33111;
w33164 <= not w33107 and w33163;
w33165 <= not w33108 and not w33111;
w33166 <= not w33164 and not w33165;
w33167 <= w4915 and not w33166;
w33168 <= not w33133 and w33167;
w33169 <= not w33162 and not w33168;
w33170 <= not b(22) and not w33169;
w33171 <= not w32840 and not w33134;
w33172 <= not w32850 and w33106;
w33173 <= not w33102 and w33172;
w33174 <= not w33103 and not w33106;
w33175 <= not w33173 and not w33174;
w33176 <= w4915 and not w33175;
w33177 <= not w33133 and w33176;
w33178 <= not w33171 and not w33177;
w33179 <= not b(21) and not w33178;
w33180 <= not w32849 and not w33134;
w33181 <= not w32859 and w33101;
w33182 <= not w33097 and w33181;
w33183 <= not w33098 and not w33101;
w33184 <= not w33182 and not w33183;
w33185 <= w4915 and not w33184;
w33186 <= not w33133 and w33185;
w33187 <= not w33180 and not w33186;
w33188 <= not b(20) and not w33187;
w33189 <= not w32858 and not w33134;
w33190 <= not w32868 and w33096;
w33191 <= not w33092 and w33190;
w33192 <= not w33093 and not w33096;
w33193 <= not w33191 and not w33192;
w33194 <= w4915 and not w33193;
w33195 <= not w33133 and w33194;
w33196 <= not w33189 and not w33195;
w33197 <= not b(19) and not w33196;
w33198 <= not w32867 and not w33134;
w33199 <= not w32877 and w33091;
w33200 <= not w33087 and w33199;
w33201 <= not w33088 and not w33091;
w33202 <= not w33200 and not w33201;
w33203 <= w4915 and not w33202;
w33204 <= not w33133 and w33203;
w33205 <= not w33198 and not w33204;
w33206 <= not b(18) and not w33205;
w33207 <= not w32876 and not w33134;
w33208 <= not w32886 and w33086;
w33209 <= not w33082 and w33208;
w33210 <= not w33083 and not w33086;
w33211 <= not w33209 and not w33210;
w33212 <= w4915 and not w33211;
w33213 <= not w33133 and w33212;
w33214 <= not w33207 and not w33213;
w33215 <= not b(17) and not w33214;
w33216 <= not w32885 and not w33134;
w33217 <= not w32895 and w33081;
w33218 <= not w33077 and w33217;
w33219 <= not w33078 and not w33081;
w33220 <= not w33218 and not w33219;
w33221 <= w4915 and not w33220;
w33222 <= not w33133 and w33221;
w33223 <= not w33216 and not w33222;
w33224 <= not b(16) and not w33223;
w33225 <= not w32894 and not w33134;
w33226 <= not w32904 and w33076;
w33227 <= not w33072 and w33226;
w33228 <= not w33073 and not w33076;
w33229 <= not w33227 and not w33228;
w33230 <= w4915 and not w33229;
w33231 <= not w33133 and w33230;
w33232 <= not w33225 and not w33231;
w33233 <= not b(15) and not w33232;
w33234 <= not w32903 and not w33134;
w33235 <= not w32913 and w33071;
w33236 <= not w33067 and w33235;
w33237 <= not w33068 and not w33071;
w33238 <= not w33236 and not w33237;
w33239 <= w4915 and not w33238;
w33240 <= not w33133 and w33239;
w33241 <= not w33234 and not w33240;
w33242 <= not b(14) and not w33241;
w33243 <= not w32912 and not w33134;
w33244 <= not w32922 and w33066;
w33245 <= not w33062 and w33244;
w33246 <= not w33063 and not w33066;
w33247 <= not w33245 and not w33246;
w33248 <= w4915 and not w33247;
w33249 <= not w33133 and w33248;
w33250 <= not w33243 and not w33249;
w33251 <= not b(13) and not w33250;
w33252 <= not w32921 and not w33134;
w33253 <= not w32931 and w33061;
w33254 <= not w33057 and w33253;
w33255 <= not w33058 and not w33061;
w33256 <= not w33254 and not w33255;
w33257 <= w4915 and not w33256;
w33258 <= not w33133 and w33257;
w33259 <= not w33252 and not w33258;
w33260 <= not b(12) and not w33259;
w33261 <= not w32930 and not w33134;
w33262 <= not w32940 and w33056;
w33263 <= not w33052 and w33262;
w33264 <= not w33053 and not w33056;
w33265 <= not w33263 and not w33264;
w33266 <= w4915 and not w33265;
w33267 <= not w33133 and w33266;
w33268 <= not w33261 and not w33267;
w33269 <= not b(11) and not w33268;
w33270 <= not w32939 and not w33134;
w33271 <= not w32949 and w33051;
w33272 <= not w33047 and w33271;
w33273 <= not w33048 and not w33051;
w33274 <= not w33272 and not w33273;
w33275 <= w4915 and not w33274;
w33276 <= not w33133 and w33275;
w33277 <= not w33270 and not w33276;
w33278 <= not b(10) and not w33277;
w33279 <= not w32948 and not w33134;
w33280 <= not w32958 and w33046;
w33281 <= not w33042 and w33280;
w33282 <= not w33043 and not w33046;
w33283 <= not w33281 and not w33282;
w33284 <= w4915 and not w33283;
w33285 <= not w33133 and w33284;
w33286 <= not w33279 and not w33285;
w33287 <= not b(9) and not w33286;
w33288 <= not w32957 and not w33134;
w33289 <= not w32967 and w33041;
w33290 <= not w33037 and w33289;
w33291 <= not w33038 and not w33041;
w33292 <= not w33290 and not w33291;
w33293 <= w4915 and not w33292;
w33294 <= not w33133 and w33293;
w33295 <= not w33288 and not w33294;
w33296 <= not b(8) and not w33295;
w33297 <= not w32966 and not w33134;
w33298 <= not w32976 and w33036;
w33299 <= not w33032 and w33298;
w33300 <= not w33033 and not w33036;
w33301 <= not w33299 and not w33300;
w33302 <= w4915 and not w33301;
w33303 <= not w33133 and w33302;
w33304 <= not w33297 and not w33303;
w33305 <= not b(7) and not w33304;
w33306 <= not w32975 and not w33134;
w33307 <= not w32985 and w33031;
w33308 <= not w33027 and w33307;
w33309 <= not w33028 and not w33031;
w33310 <= not w33308 and not w33309;
w33311 <= w4915 and not w33310;
w33312 <= not w33133 and w33311;
w33313 <= not w33306 and not w33312;
w33314 <= not b(6) and not w33313;
w33315 <= not w32984 and not w33134;
w33316 <= not w32994 and w33026;
w33317 <= not w33022 and w33316;
w33318 <= not w33023 and not w33026;
w33319 <= not w33317 and not w33318;
w33320 <= w4915 and not w33319;
w33321 <= not w33133 and w33320;
w33322 <= not w33315 and not w33321;
w33323 <= not b(5) and not w33322;
w33324 <= not w32993 and not w33134;
w33325 <= not w33002 and w33021;
w33326 <= not w33017 and w33325;
w33327 <= not w33018 and not w33021;
w33328 <= not w33326 and not w33327;
w33329 <= w4915 and not w33328;
w33330 <= not w33133 and w33329;
w33331 <= not w33324 and not w33330;
w33332 <= not b(4) and not w33331;
w33333 <= not w33001 and not w33134;
w33334 <= not w33012 and w33016;
w33335 <= not w33011 and w33334;
w33336 <= not w33013 and not w33016;
w33337 <= not w33335 and not w33336;
w33338 <= w4915 and not w33337;
w33339 <= not w33133 and w33338;
w33340 <= not w33333 and not w33339;
w33341 <= not b(3) and not w33340;
w33342 <= not w33006 and not w33134;
w33343 <= w4789 and not w33009;
w33344 <= not w33007 and w33343;
w33345 <= w4915 and not w33344;
w33346 <= not w33011 and w33345;
w33347 <= not w33133 and w33346;
w33348 <= not w33342 and not w33347;
w33349 <= not b(2) and not w33348;
w33350 <= w5136 and not w33133;
w33351 <= a(38) and not w33350;
w33352 <= w5142 and not w33133;
w33353 <= not w33351 and not w33352;
w33354 <= b(1) and not w33353;
w33355 <= not b(1) and not w33352;
w33356 <= not w33351 and w33355;
w33357 <= not w33354 and not w33356;
w33358 <= not w5149 and not w33357;
w33359 <= not b(1) and not w33353;
w33360 <= not w33358 and not w33359;
w33361 <= b(2) and not w33347;
w33362 <= not w33342 and w33361;
w33363 <= not w33349 and not w33362;
w33364 <= not w33360 and w33363;
w33365 <= not w33349 and not w33364;
w33366 <= b(3) and not w33339;
w33367 <= not w33333 and w33366;
w33368 <= not w33341 and not w33367;
w33369 <= not w33365 and w33368;
w33370 <= not w33341 and not w33369;
w33371 <= b(4) and not w33330;
w33372 <= not w33324 and w33371;
w33373 <= not w33332 and not w33372;
w33374 <= not w33370 and w33373;
w33375 <= not w33332 and not w33374;
w33376 <= b(5) and not w33321;
w33377 <= not w33315 and w33376;
w33378 <= not w33323 and not w33377;
w33379 <= not w33375 and w33378;
w33380 <= not w33323 and not w33379;
w33381 <= b(6) and not w33312;
w33382 <= not w33306 and w33381;
w33383 <= not w33314 and not w33382;
w33384 <= not w33380 and w33383;
w33385 <= not w33314 and not w33384;
w33386 <= b(7) and not w33303;
w33387 <= not w33297 and w33386;
w33388 <= not w33305 and not w33387;
w33389 <= not w33385 and w33388;
w33390 <= not w33305 and not w33389;
w33391 <= b(8) and not w33294;
w33392 <= not w33288 and w33391;
w33393 <= not w33296 and not w33392;
w33394 <= not w33390 and w33393;
w33395 <= not w33296 and not w33394;
w33396 <= b(9) and not w33285;
w33397 <= not w33279 and w33396;
w33398 <= not w33287 and not w33397;
w33399 <= not w33395 and w33398;
w33400 <= not w33287 and not w33399;
w33401 <= b(10) and not w33276;
w33402 <= not w33270 and w33401;
w33403 <= not w33278 and not w33402;
w33404 <= not w33400 and w33403;
w33405 <= not w33278 and not w33404;
w33406 <= b(11) and not w33267;
w33407 <= not w33261 and w33406;
w33408 <= not w33269 and not w33407;
w33409 <= not w33405 and w33408;
w33410 <= not w33269 and not w33409;
w33411 <= b(12) and not w33258;
w33412 <= not w33252 and w33411;
w33413 <= not w33260 and not w33412;
w33414 <= not w33410 and w33413;
w33415 <= not w33260 and not w33414;
w33416 <= b(13) and not w33249;
w33417 <= not w33243 and w33416;
w33418 <= not w33251 and not w33417;
w33419 <= not w33415 and w33418;
w33420 <= not w33251 and not w33419;
w33421 <= b(14) and not w33240;
w33422 <= not w33234 and w33421;
w33423 <= not w33242 and not w33422;
w33424 <= not w33420 and w33423;
w33425 <= not w33242 and not w33424;
w33426 <= b(15) and not w33231;
w33427 <= not w33225 and w33426;
w33428 <= not w33233 and not w33427;
w33429 <= not w33425 and w33428;
w33430 <= not w33233 and not w33429;
w33431 <= b(16) and not w33222;
w33432 <= not w33216 and w33431;
w33433 <= not w33224 and not w33432;
w33434 <= not w33430 and w33433;
w33435 <= not w33224 and not w33434;
w33436 <= b(17) and not w33213;
w33437 <= not w33207 and w33436;
w33438 <= not w33215 and not w33437;
w33439 <= not w33435 and w33438;
w33440 <= not w33215 and not w33439;
w33441 <= b(18) and not w33204;
w33442 <= not w33198 and w33441;
w33443 <= not w33206 and not w33442;
w33444 <= not w33440 and w33443;
w33445 <= not w33206 and not w33444;
w33446 <= b(19) and not w33195;
w33447 <= not w33189 and w33446;
w33448 <= not w33197 and not w33447;
w33449 <= not w33445 and w33448;
w33450 <= not w33197 and not w33449;
w33451 <= b(20) and not w33186;
w33452 <= not w33180 and w33451;
w33453 <= not w33188 and not w33452;
w33454 <= not w33450 and w33453;
w33455 <= not w33188 and not w33454;
w33456 <= b(21) and not w33177;
w33457 <= not w33171 and w33456;
w33458 <= not w33179 and not w33457;
w33459 <= not w33455 and w33458;
w33460 <= not w33179 and not w33459;
w33461 <= b(22) and not w33168;
w33462 <= not w33162 and w33461;
w33463 <= not w33170 and not w33462;
w33464 <= not w33460 and w33463;
w33465 <= not w33170 and not w33464;
w33466 <= b(23) and not w33159;
w33467 <= not w33153 and w33466;
w33468 <= not w33161 and not w33467;
w33469 <= not w33465 and w33468;
w33470 <= not w33161 and not w33469;
w33471 <= b(24) and not w33150;
w33472 <= not w33144 and w33471;
w33473 <= not w33152 and not w33472;
w33474 <= not w33470 and w33473;
w33475 <= not w33152 and not w33474;
w33476 <= b(25) and not w33141;
w33477 <= not w33135 and w33476;
w33478 <= not w33143 and not w33477;
w33479 <= not w33475 and w33478;
w33480 <= not w33143 and not w33479;
w33481 <= not w32803 and not w33134;
w33482 <= not w32805 and w33131;
w33483 <= not w33127 and w33482;
w33484 <= not w33128 and not w33131;
w33485 <= not w33483 and not w33484;
w33486 <= w33134 and not w33485;
w33487 <= not w33481 and not w33486;
w33488 <= not b(26) and not w33487;
w33489 <= b(26) and not w33481;
w33490 <= not w33486 and w33489;
w33491 <= w5285 and not w33490;
w33492 <= not w33488 and w33491;
w33493 <= not w33480 and w33492;
w33494 <= w4915 and not w33487;
w33495 <= not w33493 and not w33494;
w33496 <= not w33152 and w33478;
w33497 <= not w33474 and w33496;
w33498 <= not w33475 and not w33478;
w33499 <= not w33497 and not w33498;
w33500 <= not w33495 and not w33499;
w33501 <= not w33142 and not w33494;
w33502 <= not w33493 and w33501;
w33503 <= not w33500 and not w33502;
w33504 <= not w33143 and not w33490;
w33505 <= not w33488 and w33504;
w33506 <= not w33479 and w33505;
w33507 <= not w33488 and not w33490;
w33508 <= not w33480 and not w33507;
w33509 <= not w33506 and not w33508;
w33510 <= not w33495 and not w33509;
w33511 <= not w33487 and not w33494;
w33512 <= not w33493 and w33511;
w33513 <= not w33510 and not w33512;
w33514 <= not b(27) and not w33513;
w33515 <= not b(26) and not w33503;
w33516 <= not w33161 and w33473;
w33517 <= not w33469 and w33516;
w33518 <= not w33470 and not w33473;
w33519 <= not w33517 and not w33518;
w33520 <= not w33495 and not w33519;
w33521 <= not w33151 and not w33494;
w33522 <= not w33493 and w33521;
w33523 <= not w33520 and not w33522;
w33524 <= not b(25) and not w33523;
w33525 <= not w33170 and w33468;
w33526 <= not w33464 and w33525;
w33527 <= not w33465 and not w33468;
w33528 <= not w33526 and not w33527;
w33529 <= not w33495 and not w33528;
w33530 <= not w33160 and not w33494;
w33531 <= not w33493 and w33530;
w33532 <= not w33529 and not w33531;
w33533 <= not b(24) and not w33532;
w33534 <= not w33179 and w33463;
w33535 <= not w33459 and w33534;
w33536 <= not w33460 and not w33463;
w33537 <= not w33535 and not w33536;
w33538 <= not w33495 and not w33537;
w33539 <= not w33169 and not w33494;
w33540 <= not w33493 and w33539;
w33541 <= not w33538 and not w33540;
w33542 <= not b(23) and not w33541;
w33543 <= not w33188 and w33458;
w33544 <= not w33454 and w33543;
w33545 <= not w33455 and not w33458;
w33546 <= not w33544 and not w33545;
w33547 <= not w33495 and not w33546;
w33548 <= not w33178 and not w33494;
w33549 <= not w33493 and w33548;
w33550 <= not w33547 and not w33549;
w33551 <= not b(22) and not w33550;
w33552 <= not w33197 and w33453;
w33553 <= not w33449 and w33552;
w33554 <= not w33450 and not w33453;
w33555 <= not w33553 and not w33554;
w33556 <= not w33495 and not w33555;
w33557 <= not w33187 and not w33494;
w33558 <= not w33493 and w33557;
w33559 <= not w33556 and not w33558;
w33560 <= not b(21) and not w33559;
w33561 <= not w33206 and w33448;
w33562 <= not w33444 and w33561;
w33563 <= not w33445 and not w33448;
w33564 <= not w33562 and not w33563;
w33565 <= not w33495 and not w33564;
w33566 <= not w33196 and not w33494;
w33567 <= not w33493 and w33566;
w33568 <= not w33565 and not w33567;
w33569 <= not b(20) and not w33568;
w33570 <= not w33215 and w33443;
w33571 <= not w33439 and w33570;
w33572 <= not w33440 and not w33443;
w33573 <= not w33571 and not w33572;
w33574 <= not w33495 and not w33573;
w33575 <= not w33205 and not w33494;
w33576 <= not w33493 and w33575;
w33577 <= not w33574 and not w33576;
w33578 <= not b(19) and not w33577;
w33579 <= not w33224 and w33438;
w33580 <= not w33434 and w33579;
w33581 <= not w33435 and not w33438;
w33582 <= not w33580 and not w33581;
w33583 <= not w33495 and not w33582;
w33584 <= not w33214 and not w33494;
w33585 <= not w33493 and w33584;
w33586 <= not w33583 and not w33585;
w33587 <= not b(18) and not w33586;
w33588 <= not w33233 and w33433;
w33589 <= not w33429 and w33588;
w33590 <= not w33430 and not w33433;
w33591 <= not w33589 and not w33590;
w33592 <= not w33495 and not w33591;
w33593 <= not w33223 and not w33494;
w33594 <= not w33493 and w33593;
w33595 <= not w33592 and not w33594;
w33596 <= not b(17) and not w33595;
w33597 <= not w33242 and w33428;
w33598 <= not w33424 and w33597;
w33599 <= not w33425 and not w33428;
w33600 <= not w33598 and not w33599;
w33601 <= not w33495 and not w33600;
w33602 <= not w33232 and not w33494;
w33603 <= not w33493 and w33602;
w33604 <= not w33601 and not w33603;
w33605 <= not b(16) and not w33604;
w33606 <= not w33251 and w33423;
w33607 <= not w33419 and w33606;
w33608 <= not w33420 and not w33423;
w33609 <= not w33607 and not w33608;
w33610 <= not w33495 and not w33609;
w33611 <= not w33241 and not w33494;
w33612 <= not w33493 and w33611;
w33613 <= not w33610 and not w33612;
w33614 <= not b(15) and not w33613;
w33615 <= not w33260 and w33418;
w33616 <= not w33414 and w33615;
w33617 <= not w33415 and not w33418;
w33618 <= not w33616 and not w33617;
w33619 <= not w33495 and not w33618;
w33620 <= not w33250 and not w33494;
w33621 <= not w33493 and w33620;
w33622 <= not w33619 and not w33621;
w33623 <= not b(14) and not w33622;
w33624 <= not w33269 and w33413;
w33625 <= not w33409 and w33624;
w33626 <= not w33410 and not w33413;
w33627 <= not w33625 and not w33626;
w33628 <= not w33495 and not w33627;
w33629 <= not w33259 and not w33494;
w33630 <= not w33493 and w33629;
w33631 <= not w33628 and not w33630;
w33632 <= not b(13) and not w33631;
w33633 <= not w33278 and w33408;
w33634 <= not w33404 and w33633;
w33635 <= not w33405 and not w33408;
w33636 <= not w33634 and not w33635;
w33637 <= not w33495 and not w33636;
w33638 <= not w33268 and not w33494;
w33639 <= not w33493 and w33638;
w33640 <= not w33637 and not w33639;
w33641 <= not b(12) and not w33640;
w33642 <= not w33287 and w33403;
w33643 <= not w33399 and w33642;
w33644 <= not w33400 and not w33403;
w33645 <= not w33643 and not w33644;
w33646 <= not w33495 and not w33645;
w33647 <= not w33277 and not w33494;
w33648 <= not w33493 and w33647;
w33649 <= not w33646 and not w33648;
w33650 <= not b(11) and not w33649;
w33651 <= not w33296 and w33398;
w33652 <= not w33394 and w33651;
w33653 <= not w33395 and not w33398;
w33654 <= not w33652 and not w33653;
w33655 <= not w33495 and not w33654;
w33656 <= not w33286 and not w33494;
w33657 <= not w33493 and w33656;
w33658 <= not w33655 and not w33657;
w33659 <= not b(10) and not w33658;
w33660 <= not w33305 and w33393;
w33661 <= not w33389 and w33660;
w33662 <= not w33390 and not w33393;
w33663 <= not w33661 and not w33662;
w33664 <= not w33495 and not w33663;
w33665 <= not w33295 and not w33494;
w33666 <= not w33493 and w33665;
w33667 <= not w33664 and not w33666;
w33668 <= not b(9) and not w33667;
w33669 <= not w33314 and w33388;
w33670 <= not w33384 and w33669;
w33671 <= not w33385 and not w33388;
w33672 <= not w33670 and not w33671;
w33673 <= not w33495 and not w33672;
w33674 <= not w33304 and not w33494;
w33675 <= not w33493 and w33674;
w33676 <= not w33673 and not w33675;
w33677 <= not b(8) and not w33676;
w33678 <= not w33323 and w33383;
w33679 <= not w33379 and w33678;
w33680 <= not w33380 and not w33383;
w33681 <= not w33679 and not w33680;
w33682 <= not w33495 and not w33681;
w33683 <= not w33313 and not w33494;
w33684 <= not w33493 and w33683;
w33685 <= not w33682 and not w33684;
w33686 <= not b(7) and not w33685;
w33687 <= not w33332 and w33378;
w33688 <= not w33374 and w33687;
w33689 <= not w33375 and not w33378;
w33690 <= not w33688 and not w33689;
w33691 <= not w33495 and not w33690;
w33692 <= not w33322 and not w33494;
w33693 <= not w33493 and w33692;
w33694 <= not w33691 and not w33693;
w33695 <= not b(6) and not w33694;
w33696 <= not w33341 and w33373;
w33697 <= not w33369 and w33696;
w33698 <= not w33370 and not w33373;
w33699 <= not w33697 and not w33698;
w33700 <= not w33495 and not w33699;
w33701 <= not w33331 and not w33494;
w33702 <= not w33493 and w33701;
w33703 <= not w33700 and not w33702;
w33704 <= not b(5) and not w33703;
w33705 <= not w33349 and w33368;
w33706 <= not w33364 and w33705;
w33707 <= not w33365 and not w33368;
w33708 <= not w33706 and not w33707;
w33709 <= not w33495 and not w33708;
w33710 <= not w33340 and not w33494;
w33711 <= not w33493 and w33710;
w33712 <= not w33709 and not w33711;
w33713 <= not b(4) and not w33712;
w33714 <= not w33359 and w33363;
w33715 <= not w33358 and w33714;
w33716 <= not w33360 and not w33363;
w33717 <= not w33715 and not w33716;
w33718 <= not w33495 and not w33717;
w33719 <= not w33348 and not w33494;
w33720 <= not w33493 and w33719;
w33721 <= not w33718 and not w33720;
w33722 <= not b(3) and not w33721;
w33723 <= w5149 and not w33356;
w33724 <= not w33354 and w33723;
w33725 <= not w33358 and not w33724;
w33726 <= not w33495 and w33725;
w33727 <= not w33353 and not w33494;
w33728 <= not w33493 and w33727;
w33729 <= not w33726 and not w33728;
w33730 <= not b(2) and not w33729;
w33731 <= b(0) and not w33495;
w33732 <= a(37) and not w33731;
w33733 <= w5149 and not w33495;
w33734 <= not w33732 and not w33733;
w33735 <= b(1) and not w33734;
w33736 <= not b(1) and not w33733;
w33737 <= not w33732 and w33736;
w33738 <= not w33735 and not w33737;
w33739 <= not w5534 and not w33738;
w33740 <= not b(1) and not w33734;
w33741 <= not w33739 and not w33740;
w33742 <= b(2) and not w33728;
w33743 <= not w33726 and w33742;
w33744 <= not w33730 and not w33743;
w33745 <= not w33741 and w33744;
w33746 <= not w33730 and not w33745;
w33747 <= b(3) and not w33720;
w33748 <= not w33718 and w33747;
w33749 <= not w33722 and not w33748;
w33750 <= not w33746 and w33749;
w33751 <= not w33722 and not w33750;
w33752 <= b(4) and not w33711;
w33753 <= not w33709 and w33752;
w33754 <= not w33713 and not w33753;
w33755 <= not w33751 and w33754;
w33756 <= not w33713 and not w33755;
w33757 <= b(5) and not w33702;
w33758 <= not w33700 and w33757;
w33759 <= not w33704 and not w33758;
w33760 <= not w33756 and w33759;
w33761 <= not w33704 and not w33760;
w33762 <= b(6) and not w33693;
w33763 <= not w33691 and w33762;
w33764 <= not w33695 and not w33763;
w33765 <= not w33761 and w33764;
w33766 <= not w33695 and not w33765;
w33767 <= b(7) and not w33684;
w33768 <= not w33682 and w33767;
w33769 <= not w33686 and not w33768;
w33770 <= not w33766 and w33769;
w33771 <= not w33686 and not w33770;
w33772 <= b(8) and not w33675;
w33773 <= not w33673 and w33772;
w33774 <= not w33677 and not w33773;
w33775 <= not w33771 and w33774;
w33776 <= not w33677 and not w33775;
w33777 <= b(9) and not w33666;
w33778 <= not w33664 and w33777;
w33779 <= not w33668 and not w33778;
w33780 <= not w33776 and w33779;
w33781 <= not w33668 and not w33780;
w33782 <= b(10) and not w33657;
w33783 <= not w33655 and w33782;
w33784 <= not w33659 and not w33783;
w33785 <= not w33781 and w33784;
w33786 <= not w33659 and not w33785;
w33787 <= b(11) and not w33648;
w33788 <= not w33646 and w33787;
w33789 <= not w33650 and not w33788;
w33790 <= not w33786 and w33789;
w33791 <= not w33650 and not w33790;
w33792 <= b(12) and not w33639;
w33793 <= not w33637 and w33792;
w33794 <= not w33641 and not w33793;
w33795 <= not w33791 and w33794;
w33796 <= not w33641 and not w33795;
w33797 <= b(13) and not w33630;
w33798 <= not w33628 and w33797;
w33799 <= not w33632 and not w33798;
w33800 <= not w33796 and w33799;
w33801 <= not w33632 and not w33800;
w33802 <= b(14) and not w33621;
w33803 <= not w33619 and w33802;
w33804 <= not w33623 and not w33803;
w33805 <= not w33801 and w33804;
w33806 <= not w33623 and not w33805;
w33807 <= b(15) and not w33612;
w33808 <= not w33610 and w33807;
w33809 <= not w33614 and not w33808;
w33810 <= not w33806 and w33809;
w33811 <= not w33614 and not w33810;
w33812 <= b(16) and not w33603;
w33813 <= not w33601 and w33812;
w33814 <= not w33605 and not w33813;
w33815 <= not w33811 and w33814;
w33816 <= not w33605 and not w33815;
w33817 <= b(17) and not w33594;
w33818 <= not w33592 and w33817;
w33819 <= not w33596 and not w33818;
w33820 <= not w33816 and w33819;
w33821 <= not w33596 and not w33820;
w33822 <= b(18) and not w33585;
w33823 <= not w33583 and w33822;
w33824 <= not w33587 and not w33823;
w33825 <= not w33821 and w33824;
w33826 <= not w33587 and not w33825;
w33827 <= b(19) and not w33576;
w33828 <= not w33574 and w33827;
w33829 <= not w33578 and not w33828;
w33830 <= not w33826 and w33829;
w33831 <= not w33578 and not w33830;
w33832 <= b(20) and not w33567;
w33833 <= not w33565 and w33832;
w33834 <= not w33569 and not w33833;
w33835 <= not w33831 and w33834;
w33836 <= not w33569 and not w33835;
w33837 <= b(21) and not w33558;
w33838 <= not w33556 and w33837;
w33839 <= not w33560 and not w33838;
w33840 <= not w33836 and w33839;
w33841 <= not w33560 and not w33840;
w33842 <= b(22) and not w33549;
w33843 <= not w33547 and w33842;
w33844 <= not w33551 and not w33843;
w33845 <= not w33841 and w33844;
w33846 <= not w33551 and not w33845;
w33847 <= b(23) and not w33540;
w33848 <= not w33538 and w33847;
w33849 <= not w33542 and not w33848;
w33850 <= not w33846 and w33849;
w33851 <= not w33542 and not w33850;
w33852 <= b(24) and not w33531;
w33853 <= not w33529 and w33852;
w33854 <= not w33533 and not w33853;
w33855 <= not w33851 and w33854;
w33856 <= not w33533 and not w33855;
w33857 <= b(25) and not w33522;
w33858 <= not w33520 and w33857;
w33859 <= not w33524 and not w33858;
w33860 <= not w33856 and w33859;
w33861 <= not w33524 and not w33860;
w33862 <= b(26) and not w33502;
w33863 <= not w33500 and w33862;
w33864 <= not w33515 and not w33863;
w33865 <= not w33861 and w33864;
w33866 <= not w33515 and not w33865;
w33867 <= b(27) and not w33512;
w33868 <= not w33510 and w33867;
w33869 <= not w33514 and not w33868;
w33870 <= not w33866 and w33869;
w33871 <= not w33514 and not w33870;
w33872 <= w5669 and not w33871;
w33873 <= not w33503 and not w33872;
w33874 <= not w33524 and w33864;
w33875 <= not w33860 and w33874;
w33876 <= not w33861 and not w33864;
w33877 <= not w33875 and not w33876;
w33878 <= w5669 and not w33877;
w33879 <= not w33871 and w33878;
w33880 <= not w33873 and not w33879;
w33881 <= not w33513 and not w33872;
w33882 <= not w33515 and w33869;
w33883 <= not w33865 and w33882;
w33884 <= not w33866 and not w33869;
w33885 <= not w33883 and not w33884;
w33886 <= w33872 and not w33885;
w33887 <= not w33881 and not w33886;
w33888 <= not b(28) and not w33887;
w33889 <= not b(27) and not w33880;
w33890 <= not w33523 and not w33872;
w33891 <= not w33533 and w33859;
w33892 <= not w33855 and w33891;
w33893 <= not w33856 and not w33859;
w33894 <= not w33892 and not w33893;
w33895 <= w5669 and not w33894;
w33896 <= not w33871 and w33895;
w33897 <= not w33890 and not w33896;
w33898 <= not b(26) and not w33897;
w33899 <= not w33532 and not w33872;
w33900 <= not w33542 and w33854;
w33901 <= not w33850 and w33900;
w33902 <= not w33851 and not w33854;
w33903 <= not w33901 and not w33902;
w33904 <= w5669 and not w33903;
w33905 <= not w33871 and w33904;
w33906 <= not w33899 and not w33905;
w33907 <= not b(25) and not w33906;
w33908 <= not w33541 and not w33872;
w33909 <= not w33551 and w33849;
w33910 <= not w33845 and w33909;
w33911 <= not w33846 and not w33849;
w33912 <= not w33910 and not w33911;
w33913 <= w5669 and not w33912;
w33914 <= not w33871 and w33913;
w33915 <= not w33908 and not w33914;
w33916 <= not b(24) and not w33915;
w33917 <= not w33550 and not w33872;
w33918 <= not w33560 and w33844;
w33919 <= not w33840 and w33918;
w33920 <= not w33841 and not w33844;
w33921 <= not w33919 and not w33920;
w33922 <= w5669 and not w33921;
w33923 <= not w33871 and w33922;
w33924 <= not w33917 and not w33923;
w33925 <= not b(23) and not w33924;
w33926 <= not w33559 and not w33872;
w33927 <= not w33569 and w33839;
w33928 <= not w33835 and w33927;
w33929 <= not w33836 and not w33839;
w33930 <= not w33928 and not w33929;
w33931 <= w5669 and not w33930;
w33932 <= not w33871 and w33931;
w33933 <= not w33926 and not w33932;
w33934 <= not b(22) and not w33933;
w33935 <= not w33568 and not w33872;
w33936 <= not w33578 and w33834;
w33937 <= not w33830 and w33936;
w33938 <= not w33831 and not w33834;
w33939 <= not w33937 and not w33938;
w33940 <= w5669 and not w33939;
w33941 <= not w33871 and w33940;
w33942 <= not w33935 and not w33941;
w33943 <= not b(21) and not w33942;
w33944 <= not w33577 and not w33872;
w33945 <= not w33587 and w33829;
w33946 <= not w33825 and w33945;
w33947 <= not w33826 and not w33829;
w33948 <= not w33946 and not w33947;
w33949 <= w5669 and not w33948;
w33950 <= not w33871 and w33949;
w33951 <= not w33944 and not w33950;
w33952 <= not b(20) and not w33951;
w33953 <= not w33586 and not w33872;
w33954 <= not w33596 and w33824;
w33955 <= not w33820 and w33954;
w33956 <= not w33821 and not w33824;
w33957 <= not w33955 and not w33956;
w33958 <= w5669 and not w33957;
w33959 <= not w33871 and w33958;
w33960 <= not w33953 and not w33959;
w33961 <= not b(19) and not w33960;
w33962 <= not w33595 and not w33872;
w33963 <= not w33605 and w33819;
w33964 <= not w33815 and w33963;
w33965 <= not w33816 and not w33819;
w33966 <= not w33964 and not w33965;
w33967 <= w5669 and not w33966;
w33968 <= not w33871 and w33967;
w33969 <= not w33962 and not w33968;
w33970 <= not b(18) and not w33969;
w33971 <= not w33604 and not w33872;
w33972 <= not w33614 and w33814;
w33973 <= not w33810 and w33972;
w33974 <= not w33811 and not w33814;
w33975 <= not w33973 and not w33974;
w33976 <= w5669 and not w33975;
w33977 <= not w33871 and w33976;
w33978 <= not w33971 and not w33977;
w33979 <= not b(17) and not w33978;
w33980 <= not w33613 and not w33872;
w33981 <= not w33623 and w33809;
w33982 <= not w33805 and w33981;
w33983 <= not w33806 and not w33809;
w33984 <= not w33982 and not w33983;
w33985 <= w5669 and not w33984;
w33986 <= not w33871 and w33985;
w33987 <= not w33980 and not w33986;
w33988 <= not b(16) and not w33987;
w33989 <= not w33622 and not w33872;
w33990 <= not w33632 and w33804;
w33991 <= not w33800 and w33990;
w33992 <= not w33801 and not w33804;
w33993 <= not w33991 and not w33992;
w33994 <= w5669 and not w33993;
w33995 <= not w33871 and w33994;
w33996 <= not w33989 and not w33995;
w33997 <= not b(15) and not w33996;
w33998 <= not w33631 and not w33872;
w33999 <= not w33641 and w33799;
w34000 <= not w33795 and w33999;
w34001 <= not w33796 and not w33799;
w34002 <= not w34000 and not w34001;
w34003 <= w5669 and not w34002;
w34004 <= not w33871 and w34003;
w34005 <= not w33998 and not w34004;
w34006 <= not b(14) and not w34005;
w34007 <= not w33640 and not w33872;
w34008 <= not w33650 and w33794;
w34009 <= not w33790 and w34008;
w34010 <= not w33791 and not w33794;
w34011 <= not w34009 and not w34010;
w34012 <= w5669 and not w34011;
w34013 <= not w33871 and w34012;
w34014 <= not w34007 and not w34013;
w34015 <= not b(13) and not w34014;
w34016 <= not w33649 and not w33872;
w34017 <= not w33659 and w33789;
w34018 <= not w33785 and w34017;
w34019 <= not w33786 and not w33789;
w34020 <= not w34018 and not w34019;
w34021 <= w5669 and not w34020;
w34022 <= not w33871 and w34021;
w34023 <= not w34016 and not w34022;
w34024 <= not b(12) and not w34023;
w34025 <= not w33658 and not w33872;
w34026 <= not w33668 and w33784;
w34027 <= not w33780 and w34026;
w34028 <= not w33781 and not w33784;
w34029 <= not w34027 and not w34028;
w34030 <= w5669 and not w34029;
w34031 <= not w33871 and w34030;
w34032 <= not w34025 and not w34031;
w34033 <= not b(11) and not w34032;
w34034 <= not w33667 and not w33872;
w34035 <= not w33677 and w33779;
w34036 <= not w33775 and w34035;
w34037 <= not w33776 and not w33779;
w34038 <= not w34036 and not w34037;
w34039 <= w5669 and not w34038;
w34040 <= not w33871 and w34039;
w34041 <= not w34034 and not w34040;
w34042 <= not b(10) and not w34041;
w34043 <= not w33676 and not w33872;
w34044 <= not w33686 and w33774;
w34045 <= not w33770 and w34044;
w34046 <= not w33771 and not w33774;
w34047 <= not w34045 and not w34046;
w34048 <= w5669 and not w34047;
w34049 <= not w33871 and w34048;
w34050 <= not w34043 and not w34049;
w34051 <= not b(9) and not w34050;
w34052 <= not w33685 and not w33872;
w34053 <= not w33695 and w33769;
w34054 <= not w33765 and w34053;
w34055 <= not w33766 and not w33769;
w34056 <= not w34054 and not w34055;
w34057 <= w5669 and not w34056;
w34058 <= not w33871 and w34057;
w34059 <= not w34052 and not w34058;
w34060 <= not b(8) and not w34059;
w34061 <= not w33694 and not w33872;
w34062 <= not w33704 and w33764;
w34063 <= not w33760 and w34062;
w34064 <= not w33761 and not w33764;
w34065 <= not w34063 and not w34064;
w34066 <= w5669 and not w34065;
w34067 <= not w33871 and w34066;
w34068 <= not w34061 and not w34067;
w34069 <= not b(7) and not w34068;
w34070 <= not w33703 and not w33872;
w34071 <= not w33713 and w33759;
w34072 <= not w33755 and w34071;
w34073 <= not w33756 and not w33759;
w34074 <= not w34072 and not w34073;
w34075 <= w5669 and not w34074;
w34076 <= not w33871 and w34075;
w34077 <= not w34070 and not w34076;
w34078 <= not b(6) and not w34077;
w34079 <= not w33712 and not w33872;
w34080 <= not w33722 and w33754;
w34081 <= not w33750 and w34080;
w34082 <= not w33751 and not w33754;
w34083 <= not w34081 and not w34082;
w34084 <= w5669 and not w34083;
w34085 <= not w33871 and w34084;
w34086 <= not w34079 and not w34085;
w34087 <= not b(5) and not w34086;
w34088 <= not w33721 and not w33872;
w34089 <= not w33730 and w33749;
w34090 <= not w33745 and w34089;
w34091 <= not w33746 and not w33749;
w34092 <= not w34090 and not w34091;
w34093 <= w5669 and not w34092;
w34094 <= not w33871 and w34093;
w34095 <= not w34088 and not w34094;
w34096 <= not b(4) and not w34095;
w34097 <= not w33729 and not w33872;
w34098 <= not w33740 and w33744;
w34099 <= not w33739 and w34098;
w34100 <= not w33741 and not w33744;
w34101 <= not w34099 and not w34100;
w34102 <= w5669 and not w34101;
w34103 <= not w33871 and w34102;
w34104 <= not w34097 and not w34103;
w34105 <= not b(3) and not w34104;
w34106 <= not w33734 and not w33872;
w34107 <= w5534 and not w33737;
w34108 <= not w33735 and w34107;
w34109 <= w5669 and not w34108;
w34110 <= not w33739 and w34109;
w34111 <= not w33871 and w34110;
w34112 <= not w34106 and not w34111;
w34113 <= not b(2) and not w34112;
w34114 <= w5915 and not w33871;
w34115 <= a(36) and not w34114;
w34116 <= w5920 and not w33871;
w34117 <= not w34115 and not w34116;
w34118 <= b(1) and not w34117;
w34119 <= not b(1) and not w34116;
w34120 <= not w34115 and w34119;
w34121 <= not w34118 and not w34120;
w34122 <= not w5927 and not w34121;
w34123 <= not b(1) and not w34117;
w34124 <= not w34122 and not w34123;
w34125 <= b(2) and not w34111;
w34126 <= not w34106 and w34125;
w34127 <= not w34113 and not w34126;
w34128 <= not w34124 and w34127;
w34129 <= not w34113 and not w34128;
w34130 <= b(3) and not w34103;
w34131 <= not w34097 and w34130;
w34132 <= not w34105 and not w34131;
w34133 <= not w34129 and w34132;
w34134 <= not w34105 and not w34133;
w34135 <= b(4) and not w34094;
w34136 <= not w34088 and w34135;
w34137 <= not w34096 and not w34136;
w34138 <= not w34134 and w34137;
w34139 <= not w34096 and not w34138;
w34140 <= b(5) and not w34085;
w34141 <= not w34079 and w34140;
w34142 <= not w34087 and not w34141;
w34143 <= not w34139 and w34142;
w34144 <= not w34087 and not w34143;
w34145 <= b(6) and not w34076;
w34146 <= not w34070 and w34145;
w34147 <= not w34078 and not w34146;
w34148 <= not w34144 and w34147;
w34149 <= not w34078 and not w34148;
w34150 <= b(7) and not w34067;
w34151 <= not w34061 and w34150;
w34152 <= not w34069 and not w34151;
w34153 <= not w34149 and w34152;
w34154 <= not w34069 and not w34153;
w34155 <= b(8) and not w34058;
w34156 <= not w34052 and w34155;
w34157 <= not w34060 and not w34156;
w34158 <= not w34154 and w34157;
w34159 <= not w34060 and not w34158;
w34160 <= b(9) and not w34049;
w34161 <= not w34043 and w34160;
w34162 <= not w34051 and not w34161;
w34163 <= not w34159 and w34162;
w34164 <= not w34051 and not w34163;
w34165 <= b(10) and not w34040;
w34166 <= not w34034 and w34165;
w34167 <= not w34042 and not w34166;
w34168 <= not w34164 and w34167;
w34169 <= not w34042 and not w34168;
w34170 <= b(11) and not w34031;
w34171 <= not w34025 and w34170;
w34172 <= not w34033 and not w34171;
w34173 <= not w34169 and w34172;
w34174 <= not w34033 and not w34173;
w34175 <= b(12) and not w34022;
w34176 <= not w34016 and w34175;
w34177 <= not w34024 and not w34176;
w34178 <= not w34174 and w34177;
w34179 <= not w34024 and not w34178;
w34180 <= b(13) and not w34013;
w34181 <= not w34007 and w34180;
w34182 <= not w34015 and not w34181;
w34183 <= not w34179 and w34182;
w34184 <= not w34015 and not w34183;
w34185 <= b(14) and not w34004;
w34186 <= not w33998 and w34185;
w34187 <= not w34006 and not w34186;
w34188 <= not w34184 and w34187;
w34189 <= not w34006 and not w34188;
w34190 <= b(15) and not w33995;
w34191 <= not w33989 and w34190;
w34192 <= not w33997 and not w34191;
w34193 <= not w34189 and w34192;
w34194 <= not w33997 and not w34193;
w34195 <= b(16) and not w33986;
w34196 <= not w33980 and w34195;
w34197 <= not w33988 and not w34196;
w34198 <= not w34194 and w34197;
w34199 <= not w33988 and not w34198;
w34200 <= b(17) and not w33977;
w34201 <= not w33971 and w34200;
w34202 <= not w33979 and not w34201;
w34203 <= not w34199 and w34202;
w34204 <= not w33979 and not w34203;
w34205 <= b(18) and not w33968;
w34206 <= not w33962 and w34205;
w34207 <= not w33970 and not w34206;
w34208 <= not w34204 and w34207;
w34209 <= not w33970 and not w34208;
w34210 <= b(19) and not w33959;
w34211 <= not w33953 and w34210;
w34212 <= not w33961 and not w34211;
w34213 <= not w34209 and w34212;
w34214 <= not w33961 and not w34213;
w34215 <= b(20) and not w33950;
w34216 <= not w33944 and w34215;
w34217 <= not w33952 and not w34216;
w34218 <= not w34214 and w34217;
w34219 <= not w33952 and not w34218;
w34220 <= b(21) and not w33941;
w34221 <= not w33935 and w34220;
w34222 <= not w33943 and not w34221;
w34223 <= not w34219 and w34222;
w34224 <= not w33943 and not w34223;
w34225 <= b(22) and not w33932;
w34226 <= not w33926 and w34225;
w34227 <= not w33934 and not w34226;
w34228 <= not w34224 and w34227;
w34229 <= not w33934 and not w34228;
w34230 <= b(23) and not w33923;
w34231 <= not w33917 and w34230;
w34232 <= not w33925 and not w34231;
w34233 <= not w34229 and w34232;
w34234 <= not w33925 and not w34233;
w34235 <= b(24) and not w33914;
w34236 <= not w33908 and w34235;
w34237 <= not w33916 and not w34236;
w34238 <= not w34234 and w34237;
w34239 <= not w33916 and not w34238;
w34240 <= b(25) and not w33905;
w34241 <= not w33899 and w34240;
w34242 <= not w33907 and not w34241;
w34243 <= not w34239 and w34242;
w34244 <= not w33907 and not w34243;
w34245 <= b(26) and not w33896;
w34246 <= not w33890 and w34245;
w34247 <= not w33898 and not w34246;
w34248 <= not w34244 and w34247;
w34249 <= not w33898 and not w34248;
w34250 <= b(27) and not w33879;
w34251 <= not w33873 and w34250;
w34252 <= not w33889 and not w34251;
w34253 <= not w34249 and w34252;
w34254 <= not w33889 and not w34253;
w34255 <= b(28) and not w33881;
w34256 <= not w33886 and w34255;
w34257 <= not w33888 and not w34256;
w34258 <= not w34254 and w34257;
w34259 <= not w33888 and not w34258;
w34260 <= w6067 and not w34259;
w34261 <= not w33880 and not w34260;
w34262 <= not w33898 and w34252;
w34263 <= not w34248 and w34262;
w34264 <= not w34249 and not w34252;
w34265 <= not w34263 and not w34264;
w34266 <= w6067 and not w34265;
w34267 <= not w34259 and w34266;
w34268 <= not w34261 and not w34267;
w34269 <= not b(28) and not w34268;
w34270 <= not w33897 and not w34260;
w34271 <= not w33907 and w34247;
w34272 <= not w34243 and w34271;
w34273 <= not w34244 and not w34247;
w34274 <= not w34272 and not w34273;
w34275 <= w6067 and not w34274;
w34276 <= not w34259 and w34275;
w34277 <= not w34270 and not w34276;
w34278 <= not b(27) and not w34277;
w34279 <= not w33906 and not w34260;
w34280 <= not w33916 and w34242;
w34281 <= not w34238 and w34280;
w34282 <= not w34239 and not w34242;
w34283 <= not w34281 and not w34282;
w34284 <= w6067 and not w34283;
w34285 <= not w34259 and w34284;
w34286 <= not w34279 and not w34285;
w34287 <= not b(26) and not w34286;
w34288 <= not w33915 and not w34260;
w34289 <= not w33925 and w34237;
w34290 <= not w34233 and w34289;
w34291 <= not w34234 and not w34237;
w34292 <= not w34290 and not w34291;
w34293 <= w6067 and not w34292;
w34294 <= not w34259 and w34293;
w34295 <= not w34288 and not w34294;
w34296 <= not b(25) and not w34295;
w34297 <= not w33924 and not w34260;
w34298 <= not w33934 and w34232;
w34299 <= not w34228 and w34298;
w34300 <= not w34229 and not w34232;
w34301 <= not w34299 and not w34300;
w34302 <= w6067 and not w34301;
w34303 <= not w34259 and w34302;
w34304 <= not w34297 and not w34303;
w34305 <= not b(24) and not w34304;
w34306 <= not w33933 and not w34260;
w34307 <= not w33943 and w34227;
w34308 <= not w34223 and w34307;
w34309 <= not w34224 and not w34227;
w34310 <= not w34308 and not w34309;
w34311 <= w6067 and not w34310;
w34312 <= not w34259 and w34311;
w34313 <= not w34306 and not w34312;
w34314 <= not b(23) and not w34313;
w34315 <= not w33942 and not w34260;
w34316 <= not w33952 and w34222;
w34317 <= not w34218 and w34316;
w34318 <= not w34219 and not w34222;
w34319 <= not w34317 and not w34318;
w34320 <= w6067 and not w34319;
w34321 <= not w34259 and w34320;
w34322 <= not w34315 and not w34321;
w34323 <= not b(22) and not w34322;
w34324 <= not w33951 and not w34260;
w34325 <= not w33961 and w34217;
w34326 <= not w34213 and w34325;
w34327 <= not w34214 and not w34217;
w34328 <= not w34326 and not w34327;
w34329 <= w6067 and not w34328;
w34330 <= not w34259 and w34329;
w34331 <= not w34324 and not w34330;
w34332 <= not b(21) and not w34331;
w34333 <= not w33960 and not w34260;
w34334 <= not w33970 and w34212;
w34335 <= not w34208 and w34334;
w34336 <= not w34209 and not w34212;
w34337 <= not w34335 and not w34336;
w34338 <= w6067 and not w34337;
w34339 <= not w34259 and w34338;
w34340 <= not w34333 and not w34339;
w34341 <= not b(20) and not w34340;
w34342 <= not w33969 and not w34260;
w34343 <= not w33979 and w34207;
w34344 <= not w34203 and w34343;
w34345 <= not w34204 and not w34207;
w34346 <= not w34344 and not w34345;
w34347 <= w6067 and not w34346;
w34348 <= not w34259 and w34347;
w34349 <= not w34342 and not w34348;
w34350 <= not b(19) and not w34349;
w34351 <= not w33978 and not w34260;
w34352 <= not w33988 and w34202;
w34353 <= not w34198 and w34352;
w34354 <= not w34199 and not w34202;
w34355 <= not w34353 and not w34354;
w34356 <= w6067 and not w34355;
w34357 <= not w34259 and w34356;
w34358 <= not w34351 and not w34357;
w34359 <= not b(18) and not w34358;
w34360 <= not w33987 and not w34260;
w34361 <= not w33997 and w34197;
w34362 <= not w34193 and w34361;
w34363 <= not w34194 and not w34197;
w34364 <= not w34362 and not w34363;
w34365 <= w6067 and not w34364;
w34366 <= not w34259 and w34365;
w34367 <= not w34360 and not w34366;
w34368 <= not b(17) and not w34367;
w34369 <= not w33996 and not w34260;
w34370 <= not w34006 and w34192;
w34371 <= not w34188 and w34370;
w34372 <= not w34189 and not w34192;
w34373 <= not w34371 and not w34372;
w34374 <= w6067 and not w34373;
w34375 <= not w34259 and w34374;
w34376 <= not w34369 and not w34375;
w34377 <= not b(16) and not w34376;
w34378 <= not w34005 and not w34260;
w34379 <= not w34015 and w34187;
w34380 <= not w34183 and w34379;
w34381 <= not w34184 and not w34187;
w34382 <= not w34380 and not w34381;
w34383 <= w6067 and not w34382;
w34384 <= not w34259 and w34383;
w34385 <= not w34378 and not w34384;
w34386 <= not b(15) and not w34385;
w34387 <= not w34014 and not w34260;
w34388 <= not w34024 and w34182;
w34389 <= not w34178 and w34388;
w34390 <= not w34179 and not w34182;
w34391 <= not w34389 and not w34390;
w34392 <= w6067 and not w34391;
w34393 <= not w34259 and w34392;
w34394 <= not w34387 and not w34393;
w34395 <= not b(14) and not w34394;
w34396 <= not w34023 and not w34260;
w34397 <= not w34033 and w34177;
w34398 <= not w34173 and w34397;
w34399 <= not w34174 and not w34177;
w34400 <= not w34398 and not w34399;
w34401 <= w6067 and not w34400;
w34402 <= not w34259 and w34401;
w34403 <= not w34396 and not w34402;
w34404 <= not b(13) and not w34403;
w34405 <= not w34032 and not w34260;
w34406 <= not w34042 and w34172;
w34407 <= not w34168 and w34406;
w34408 <= not w34169 and not w34172;
w34409 <= not w34407 and not w34408;
w34410 <= w6067 and not w34409;
w34411 <= not w34259 and w34410;
w34412 <= not w34405 and not w34411;
w34413 <= not b(12) and not w34412;
w34414 <= not w34041 and not w34260;
w34415 <= not w34051 and w34167;
w34416 <= not w34163 and w34415;
w34417 <= not w34164 and not w34167;
w34418 <= not w34416 and not w34417;
w34419 <= w6067 and not w34418;
w34420 <= not w34259 and w34419;
w34421 <= not w34414 and not w34420;
w34422 <= not b(11) and not w34421;
w34423 <= not w34050 and not w34260;
w34424 <= not w34060 and w34162;
w34425 <= not w34158 and w34424;
w34426 <= not w34159 and not w34162;
w34427 <= not w34425 and not w34426;
w34428 <= w6067 and not w34427;
w34429 <= not w34259 and w34428;
w34430 <= not w34423 and not w34429;
w34431 <= not b(10) and not w34430;
w34432 <= not w34059 and not w34260;
w34433 <= not w34069 and w34157;
w34434 <= not w34153 and w34433;
w34435 <= not w34154 and not w34157;
w34436 <= not w34434 and not w34435;
w34437 <= w6067 and not w34436;
w34438 <= not w34259 and w34437;
w34439 <= not w34432 and not w34438;
w34440 <= not b(9) and not w34439;
w34441 <= not w34068 and not w34260;
w34442 <= not w34078 and w34152;
w34443 <= not w34148 and w34442;
w34444 <= not w34149 and not w34152;
w34445 <= not w34443 and not w34444;
w34446 <= w6067 and not w34445;
w34447 <= not w34259 and w34446;
w34448 <= not w34441 and not w34447;
w34449 <= not b(8) and not w34448;
w34450 <= not w34077 and not w34260;
w34451 <= not w34087 and w34147;
w34452 <= not w34143 and w34451;
w34453 <= not w34144 and not w34147;
w34454 <= not w34452 and not w34453;
w34455 <= w6067 and not w34454;
w34456 <= not w34259 and w34455;
w34457 <= not w34450 and not w34456;
w34458 <= not b(7) and not w34457;
w34459 <= not w34086 and not w34260;
w34460 <= not w34096 and w34142;
w34461 <= not w34138 and w34460;
w34462 <= not w34139 and not w34142;
w34463 <= not w34461 and not w34462;
w34464 <= w6067 and not w34463;
w34465 <= not w34259 and w34464;
w34466 <= not w34459 and not w34465;
w34467 <= not b(6) and not w34466;
w34468 <= not w34095 and not w34260;
w34469 <= not w34105 and w34137;
w34470 <= not w34133 and w34469;
w34471 <= not w34134 and not w34137;
w34472 <= not w34470 and not w34471;
w34473 <= w6067 and not w34472;
w34474 <= not w34259 and w34473;
w34475 <= not w34468 and not w34474;
w34476 <= not b(5) and not w34475;
w34477 <= not w34104 and not w34260;
w34478 <= not w34113 and w34132;
w34479 <= not w34128 and w34478;
w34480 <= not w34129 and not w34132;
w34481 <= not w34479 and not w34480;
w34482 <= w6067 and not w34481;
w34483 <= not w34259 and w34482;
w34484 <= not w34477 and not w34483;
w34485 <= not b(4) and not w34484;
w34486 <= not w34112 and not w34260;
w34487 <= not w34123 and w34127;
w34488 <= not w34122 and w34487;
w34489 <= not w34124 and not w34127;
w34490 <= not w34488 and not w34489;
w34491 <= w6067 and not w34490;
w34492 <= not w34259 and w34491;
w34493 <= not w34486 and not w34492;
w34494 <= not b(3) and not w34493;
w34495 <= not w34117 and not w34260;
w34496 <= w5927 and not w34120;
w34497 <= not w34118 and w34496;
w34498 <= w6067 and not w34497;
w34499 <= not w34122 and w34498;
w34500 <= not w34259 and w34499;
w34501 <= not w34495 and not w34500;
w34502 <= not b(2) and not w34501;
w34503 <= w6315 and not w34259;
w34504 <= a(35) and not w34503;
w34505 <= w6320 and not w34259;
w34506 <= not w34504 and not w34505;
w34507 <= b(1) and not w34506;
w34508 <= not b(1) and not w34505;
w34509 <= not w34504 and w34508;
w34510 <= not w34507 and not w34509;
w34511 <= not w6327 and not w34510;
w34512 <= not b(1) and not w34506;
w34513 <= not w34511 and not w34512;
w34514 <= b(2) and not w34500;
w34515 <= not w34495 and w34514;
w34516 <= not w34502 and not w34515;
w34517 <= not w34513 and w34516;
w34518 <= not w34502 and not w34517;
w34519 <= b(3) and not w34492;
w34520 <= not w34486 and w34519;
w34521 <= not w34494 and not w34520;
w34522 <= not w34518 and w34521;
w34523 <= not w34494 and not w34522;
w34524 <= b(4) and not w34483;
w34525 <= not w34477 and w34524;
w34526 <= not w34485 and not w34525;
w34527 <= not w34523 and w34526;
w34528 <= not w34485 and not w34527;
w34529 <= b(5) and not w34474;
w34530 <= not w34468 and w34529;
w34531 <= not w34476 and not w34530;
w34532 <= not w34528 and w34531;
w34533 <= not w34476 and not w34532;
w34534 <= b(6) and not w34465;
w34535 <= not w34459 and w34534;
w34536 <= not w34467 and not w34535;
w34537 <= not w34533 and w34536;
w34538 <= not w34467 and not w34537;
w34539 <= b(7) and not w34456;
w34540 <= not w34450 and w34539;
w34541 <= not w34458 and not w34540;
w34542 <= not w34538 and w34541;
w34543 <= not w34458 and not w34542;
w34544 <= b(8) and not w34447;
w34545 <= not w34441 and w34544;
w34546 <= not w34449 and not w34545;
w34547 <= not w34543 and w34546;
w34548 <= not w34449 and not w34547;
w34549 <= b(9) and not w34438;
w34550 <= not w34432 and w34549;
w34551 <= not w34440 and not w34550;
w34552 <= not w34548 and w34551;
w34553 <= not w34440 and not w34552;
w34554 <= b(10) and not w34429;
w34555 <= not w34423 and w34554;
w34556 <= not w34431 and not w34555;
w34557 <= not w34553 and w34556;
w34558 <= not w34431 and not w34557;
w34559 <= b(11) and not w34420;
w34560 <= not w34414 and w34559;
w34561 <= not w34422 and not w34560;
w34562 <= not w34558 and w34561;
w34563 <= not w34422 and not w34562;
w34564 <= b(12) and not w34411;
w34565 <= not w34405 and w34564;
w34566 <= not w34413 and not w34565;
w34567 <= not w34563 and w34566;
w34568 <= not w34413 and not w34567;
w34569 <= b(13) and not w34402;
w34570 <= not w34396 and w34569;
w34571 <= not w34404 and not w34570;
w34572 <= not w34568 and w34571;
w34573 <= not w34404 and not w34572;
w34574 <= b(14) and not w34393;
w34575 <= not w34387 and w34574;
w34576 <= not w34395 and not w34575;
w34577 <= not w34573 and w34576;
w34578 <= not w34395 and not w34577;
w34579 <= b(15) and not w34384;
w34580 <= not w34378 and w34579;
w34581 <= not w34386 and not w34580;
w34582 <= not w34578 and w34581;
w34583 <= not w34386 and not w34582;
w34584 <= b(16) and not w34375;
w34585 <= not w34369 and w34584;
w34586 <= not w34377 and not w34585;
w34587 <= not w34583 and w34586;
w34588 <= not w34377 and not w34587;
w34589 <= b(17) and not w34366;
w34590 <= not w34360 and w34589;
w34591 <= not w34368 and not w34590;
w34592 <= not w34588 and w34591;
w34593 <= not w34368 and not w34592;
w34594 <= b(18) and not w34357;
w34595 <= not w34351 and w34594;
w34596 <= not w34359 and not w34595;
w34597 <= not w34593 and w34596;
w34598 <= not w34359 and not w34597;
w34599 <= b(19) and not w34348;
w34600 <= not w34342 and w34599;
w34601 <= not w34350 and not w34600;
w34602 <= not w34598 and w34601;
w34603 <= not w34350 and not w34602;
w34604 <= b(20) and not w34339;
w34605 <= not w34333 and w34604;
w34606 <= not w34341 and not w34605;
w34607 <= not w34603 and w34606;
w34608 <= not w34341 and not w34607;
w34609 <= b(21) and not w34330;
w34610 <= not w34324 and w34609;
w34611 <= not w34332 and not w34610;
w34612 <= not w34608 and w34611;
w34613 <= not w34332 and not w34612;
w34614 <= b(22) and not w34321;
w34615 <= not w34315 and w34614;
w34616 <= not w34323 and not w34615;
w34617 <= not w34613 and w34616;
w34618 <= not w34323 and not w34617;
w34619 <= b(23) and not w34312;
w34620 <= not w34306 and w34619;
w34621 <= not w34314 and not w34620;
w34622 <= not w34618 and w34621;
w34623 <= not w34314 and not w34622;
w34624 <= b(24) and not w34303;
w34625 <= not w34297 and w34624;
w34626 <= not w34305 and not w34625;
w34627 <= not w34623 and w34626;
w34628 <= not w34305 and not w34627;
w34629 <= b(25) and not w34294;
w34630 <= not w34288 and w34629;
w34631 <= not w34296 and not w34630;
w34632 <= not w34628 and w34631;
w34633 <= not w34296 and not w34632;
w34634 <= b(26) and not w34285;
w34635 <= not w34279 and w34634;
w34636 <= not w34287 and not w34635;
w34637 <= not w34633 and w34636;
w34638 <= not w34287 and not w34637;
w34639 <= b(27) and not w34276;
w34640 <= not w34270 and w34639;
w34641 <= not w34278 and not w34640;
w34642 <= not w34638 and w34641;
w34643 <= not w34278 and not w34642;
w34644 <= b(28) and not w34267;
w34645 <= not w34261 and w34644;
w34646 <= not w34269 and not w34645;
w34647 <= not w34643 and w34646;
w34648 <= not w34269 and not w34647;
w34649 <= not w33887 and not w34260;
w34650 <= not w33889 and w34257;
w34651 <= not w34253 and w34650;
w34652 <= not w34254 and not w34257;
w34653 <= not w34651 and not w34652;
w34654 <= w34260 and not w34653;
w34655 <= not w34649 and not w34654;
w34656 <= not b(29) and not w34655;
w34657 <= b(29) and not w34649;
w34658 <= not w34654 and w34657;
w34659 <= w6478 and not w34658;
w34660 <= not w34656 and w34659;
w34661 <= not w34648 and w34660;
w34662 <= w6067 and not w34655;
w34663 <= not w34661 and not w34662;
w34664 <= not w34278 and w34646;
w34665 <= not w34642 and w34664;
w34666 <= not w34643 and not w34646;
w34667 <= not w34665 and not w34666;
w34668 <= not w34663 and not w34667;
w34669 <= not w34268 and not w34662;
w34670 <= not w34661 and w34669;
w34671 <= not w34668 and not w34670;
w34672 <= not w34269 and not w34658;
w34673 <= not w34656 and w34672;
w34674 <= not w34647 and w34673;
w34675 <= not w34656 and not w34658;
w34676 <= not w34648 and not w34675;
w34677 <= not w34674 and not w34676;
w34678 <= not w34663 and not w34677;
w34679 <= not w34655 and not w34662;
w34680 <= not w34661 and w34679;
w34681 <= not w34678 and not w34680;
w34682 <= not b(30) and not w34681;
w34683 <= not b(29) and not w34671;
w34684 <= not w34287 and w34641;
w34685 <= not w34637 and w34684;
w34686 <= not w34638 and not w34641;
w34687 <= not w34685 and not w34686;
w34688 <= not w34663 and not w34687;
w34689 <= not w34277 and not w34662;
w34690 <= not w34661 and w34689;
w34691 <= not w34688 and not w34690;
w34692 <= not b(28) and not w34691;
w34693 <= not w34296 and w34636;
w34694 <= not w34632 and w34693;
w34695 <= not w34633 and not w34636;
w34696 <= not w34694 and not w34695;
w34697 <= not w34663 and not w34696;
w34698 <= not w34286 and not w34662;
w34699 <= not w34661 and w34698;
w34700 <= not w34697 and not w34699;
w34701 <= not b(27) and not w34700;
w34702 <= not w34305 and w34631;
w34703 <= not w34627 and w34702;
w34704 <= not w34628 and not w34631;
w34705 <= not w34703 and not w34704;
w34706 <= not w34663 and not w34705;
w34707 <= not w34295 and not w34662;
w34708 <= not w34661 and w34707;
w34709 <= not w34706 and not w34708;
w34710 <= not b(26) and not w34709;
w34711 <= not w34314 and w34626;
w34712 <= not w34622 and w34711;
w34713 <= not w34623 and not w34626;
w34714 <= not w34712 and not w34713;
w34715 <= not w34663 and not w34714;
w34716 <= not w34304 and not w34662;
w34717 <= not w34661 and w34716;
w34718 <= not w34715 and not w34717;
w34719 <= not b(25) and not w34718;
w34720 <= not w34323 and w34621;
w34721 <= not w34617 and w34720;
w34722 <= not w34618 and not w34621;
w34723 <= not w34721 and not w34722;
w34724 <= not w34663 and not w34723;
w34725 <= not w34313 and not w34662;
w34726 <= not w34661 and w34725;
w34727 <= not w34724 and not w34726;
w34728 <= not b(24) and not w34727;
w34729 <= not w34332 and w34616;
w34730 <= not w34612 and w34729;
w34731 <= not w34613 and not w34616;
w34732 <= not w34730 and not w34731;
w34733 <= not w34663 and not w34732;
w34734 <= not w34322 and not w34662;
w34735 <= not w34661 and w34734;
w34736 <= not w34733 and not w34735;
w34737 <= not b(23) and not w34736;
w34738 <= not w34341 and w34611;
w34739 <= not w34607 and w34738;
w34740 <= not w34608 and not w34611;
w34741 <= not w34739 and not w34740;
w34742 <= not w34663 and not w34741;
w34743 <= not w34331 and not w34662;
w34744 <= not w34661 and w34743;
w34745 <= not w34742 and not w34744;
w34746 <= not b(22) and not w34745;
w34747 <= not w34350 and w34606;
w34748 <= not w34602 and w34747;
w34749 <= not w34603 and not w34606;
w34750 <= not w34748 and not w34749;
w34751 <= not w34663 and not w34750;
w34752 <= not w34340 and not w34662;
w34753 <= not w34661 and w34752;
w34754 <= not w34751 and not w34753;
w34755 <= not b(21) and not w34754;
w34756 <= not w34359 and w34601;
w34757 <= not w34597 and w34756;
w34758 <= not w34598 and not w34601;
w34759 <= not w34757 and not w34758;
w34760 <= not w34663 and not w34759;
w34761 <= not w34349 and not w34662;
w34762 <= not w34661 and w34761;
w34763 <= not w34760 and not w34762;
w34764 <= not b(20) and not w34763;
w34765 <= not w34368 and w34596;
w34766 <= not w34592 and w34765;
w34767 <= not w34593 and not w34596;
w34768 <= not w34766 and not w34767;
w34769 <= not w34663 and not w34768;
w34770 <= not w34358 and not w34662;
w34771 <= not w34661 and w34770;
w34772 <= not w34769 and not w34771;
w34773 <= not b(19) and not w34772;
w34774 <= not w34377 and w34591;
w34775 <= not w34587 and w34774;
w34776 <= not w34588 and not w34591;
w34777 <= not w34775 and not w34776;
w34778 <= not w34663 and not w34777;
w34779 <= not w34367 and not w34662;
w34780 <= not w34661 and w34779;
w34781 <= not w34778 and not w34780;
w34782 <= not b(18) and not w34781;
w34783 <= not w34386 and w34586;
w34784 <= not w34582 and w34783;
w34785 <= not w34583 and not w34586;
w34786 <= not w34784 and not w34785;
w34787 <= not w34663 and not w34786;
w34788 <= not w34376 and not w34662;
w34789 <= not w34661 and w34788;
w34790 <= not w34787 and not w34789;
w34791 <= not b(17) and not w34790;
w34792 <= not w34395 and w34581;
w34793 <= not w34577 and w34792;
w34794 <= not w34578 and not w34581;
w34795 <= not w34793 and not w34794;
w34796 <= not w34663 and not w34795;
w34797 <= not w34385 and not w34662;
w34798 <= not w34661 and w34797;
w34799 <= not w34796 and not w34798;
w34800 <= not b(16) and not w34799;
w34801 <= not w34404 and w34576;
w34802 <= not w34572 and w34801;
w34803 <= not w34573 and not w34576;
w34804 <= not w34802 and not w34803;
w34805 <= not w34663 and not w34804;
w34806 <= not w34394 and not w34662;
w34807 <= not w34661 and w34806;
w34808 <= not w34805 and not w34807;
w34809 <= not b(15) and not w34808;
w34810 <= not w34413 and w34571;
w34811 <= not w34567 and w34810;
w34812 <= not w34568 and not w34571;
w34813 <= not w34811 and not w34812;
w34814 <= not w34663 and not w34813;
w34815 <= not w34403 and not w34662;
w34816 <= not w34661 and w34815;
w34817 <= not w34814 and not w34816;
w34818 <= not b(14) and not w34817;
w34819 <= not w34422 and w34566;
w34820 <= not w34562 and w34819;
w34821 <= not w34563 and not w34566;
w34822 <= not w34820 and not w34821;
w34823 <= not w34663 and not w34822;
w34824 <= not w34412 and not w34662;
w34825 <= not w34661 and w34824;
w34826 <= not w34823 and not w34825;
w34827 <= not b(13) and not w34826;
w34828 <= not w34431 and w34561;
w34829 <= not w34557 and w34828;
w34830 <= not w34558 and not w34561;
w34831 <= not w34829 and not w34830;
w34832 <= not w34663 and not w34831;
w34833 <= not w34421 and not w34662;
w34834 <= not w34661 and w34833;
w34835 <= not w34832 and not w34834;
w34836 <= not b(12) and not w34835;
w34837 <= not w34440 and w34556;
w34838 <= not w34552 and w34837;
w34839 <= not w34553 and not w34556;
w34840 <= not w34838 and not w34839;
w34841 <= not w34663 and not w34840;
w34842 <= not w34430 and not w34662;
w34843 <= not w34661 and w34842;
w34844 <= not w34841 and not w34843;
w34845 <= not b(11) and not w34844;
w34846 <= not w34449 and w34551;
w34847 <= not w34547 and w34846;
w34848 <= not w34548 and not w34551;
w34849 <= not w34847 and not w34848;
w34850 <= not w34663 and not w34849;
w34851 <= not w34439 and not w34662;
w34852 <= not w34661 and w34851;
w34853 <= not w34850 and not w34852;
w34854 <= not b(10) and not w34853;
w34855 <= not w34458 and w34546;
w34856 <= not w34542 and w34855;
w34857 <= not w34543 and not w34546;
w34858 <= not w34856 and not w34857;
w34859 <= not w34663 and not w34858;
w34860 <= not w34448 and not w34662;
w34861 <= not w34661 and w34860;
w34862 <= not w34859 and not w34861;
w34863 <= not b(9) and not w34862;
w34864 <= not w34467 and w34541;
w34865 <= not w34537 and w34864;
w34866 <= not w34538 and not w34541;
w34867 <= not w34865 and not w34866;
w34868 <= not w34663 and not w34867;
w34869 <= not w34457 and not w34662;
w34870 <= not w34661 and w34869;
w34871 <= not w34868 and not w34870;
w34872 <= not b(8) and not w34871;
w34873 <= not w34476 and w34536;
w34874 <= not w34532 and w34873;
w34875 <= not w34533 and not w34536;
w34876 <= not w34874 and not w34875;
w34877 <= not w34663 and not w34876;
w34878 <= not w34466 and not w34662;
w34879 <= not w34661 and w34878;
w34880 <= not w34877 and not w34879;
w34881 <= not b(7) and not w34880;
w34882 <= not w34485 and w34531;
w34883 <= not w34527 and w34882;
w34884 <= not w34528 and not w34531;
w34885 <= not w34883 and not w34884;
w34886 <= not w34663 and not w34885;
w34887 <= not w34475 and not w34662;
w34888 <= not w34661 and w34887;
w34889 <= not w34886 and not w34888;
w34890 <= not b(6) and not w34889;
w34891 <= not w34494 and w34526;
w34892 <= not w34522 and w34891;
w34893 <= not w34523 and not w34526;
w34894 <= not w34892 and not w34893;
w34895 <= not w34663 and not w34894;
w34896 <= not w34484 and not w34662;
w34897 <= not w34661 and w34896;
w34898 <= not w34895 and not w34897;
w34899 <= not b(5) and not w34898;
w34900 <= not w34502 and w34521;
w34901 <= not w34517 and w34900;
w34902 <= not w34518 and not w34521;
w34903 <= not w34901 and not w34902;
w34904 <= not w34663 and not w34903;
w34905 <= not w34493 and not w34662;
w34906 <= not w34661 and w34905;
w34907 <= not w34904 and not w34906;
w34908 <= not b(4) and not w34907;
w34909 <= not w34512 and w34516;
w34910 <= not w34511 and w34909;
w34911 <= not w34513 and not w34516;
w34912 <= not w34910 and not w34911;
w34913 <= not w34663 and not w34912;
w34914 <= not w34501 and not w34662;
w34915 <= not w34661 and w34914;
w34916 <= not w34913 and not w34915;
w34917 <= not b(3) and not w34916;
w34918 <= w6327 and not w34509;
w34919 <= not w34507 and w34918;
w34920 <= not w34511 and not w34919;
w34921 <= not w34663 and w34920;
w34922 <= not w34506 and not w34662;
w34923 <= not w34661 and w34922;
w34924 <= not w34921 and not w34923;
w34925 <= not b(2) and not w34924;
w34926 <= b(0) and not w34663;
w34927 <= a(34) and not w34926;
w34928 <= w6327 and not w34663;
w34929 <= not w34927 and not w34928;
w34930 <= b(1) and not w34929;
w34931 <= not b(1) and not w34928;
w34932 <= not w34927 and w34931;
w34933 <= not w34930 and not w34932;
w34934 <= not w6754 and not w34933;
w34935 <= not b(1) and not w34929;
w34936 <= not w34934 and not w34935;
w34937 <= b(2) and not w34923;
w34938 <= not w34921 and w34937;
w34939 <= not w34925 and not w34938;
w34940 <= not w34936 and w34939;
w34941 <= not w34925 and not w34940;
w34942 <= b(3) and not w34915;
w34943 <= not w34913 and w34942;
w34944 <= not w34917 and not w34943;
w34945 <= not w34941 and w34944;
w34946 <= not w34917 and not w34945;
w34947 <= b(4) and not w34906;
w34948 <= not w34904 and w34947;
w34949 <= not w34908 and not w34948;
w34950 <= not w34946 and w34949;
w34951 <= not w34908 and not w34950;
w34952 <= b(5) and not w34897;
w34953 <= not w34895 and w34952;
w34954 <= not w34899 and not w34953;
w34955 <= not w34951 and w34954;
w34956 <= not w34899 and not w34955;
w34957 <= b(6) and not w34888;
w34958 <= not w34886 and w34957;
w34959 <= not w34890 and not w34958;
w34960 <= not w34956 and w34959;
w34961 <= not w34890 and not w34960;
w34962 <= b(7) and not w34879;
w34963 <= not w34877 and w34962;
w34964 <= not w34881 and not w34963;
w34965 <= not w34961 and w34964;
w34966 <= not w34881 and not w34965;
w34967 <= b(8) and not w34870;
w34968 <= not w34868 and w34967;
w34969 <= not w34872 and not w34968;
w34970 <= not w34966 and w34969;
w34971 <= not w34872 and not w34970;
w34972 <= b(9) and not w34861;
w34973 <= not w34859 and w34972;
w34974 <= not w34863 and not w34973;
w34975 <= not w34971 and w34974;
w34976 <= not w34863 and not w34975;
w34977 <= b(10) and not w34852;
w34978 <= not w34850 and w34977;
w34979 <= not w34854 and not w34978;
w34980 <= not w34976 and w34979;
w34981 <= not w34854 and not w34980;
w34982 <= b(11) and not w34843;
w34983 <= not w34841 and w34982;
w34984 <= not w34845 and not w34983;
w34985 <= not w34981 and w34984;
w34986 <= not w34845 and not w34985;
w34987 <= b(12) and not w34834;
w34988 <= not w34832 and w34987;
w34989 <= not w34836 and not w34988;
w34990 <= not w34986 and w34989;
w34991 <= not w34836 and not w34990;
w34992 <= b(13) and not w34825;
w34993 <= not w34823 and w34992;
w34994 <= not w34827 and not w34993;
w34995 <= not w34991 and w34994;
w34996 <= not w34827 and not w34995;
w34997 <= b(14) and not w34816;
w34998 <= not w34814 and w34997;
w34999 <= not w34818 and not w34998;
w35000 <= not w34996 and w34999;
w35001 <= not w34818 and not w35000;
w35002 <= b(15) and not w34807;
w35003 <= not w34805 and w35002;
w35004 <= not w34809 and not w35003;
w35005 <= not w35001 and w35004;
w35006 <= not w34809 and not w35005;
w35007 <= b(16) and not w34798;
w35008 <= not w34796 and w35007;
w35009 <= not w34800 and not w35008;
w35010 <= not w35006 and w35009;
w35011 <= not w34800 and not w35010;
w35012 <= b(17) and not w34789;
w35013 <= not w34787 and w35012;
w35014 <= not w34791 and not w35013;
w35015 <= not w35011 and w35014;
w35016 <= not w34791 and not w35015;
w35017 <= b(18) and not w34780;
w35018 <= not w34778 and w35017;
w35019 <= not w34782 and not w35018;
w35020 <= not w35016 and w35019;
w35021 <= not w34782 and not w35020;
w35022 <= b(19) and not w34771;
w35023 <= not w34769 and w35022;
w35024 <= not w34773 and not w35023;
w35025 <= not w35021 and w35024;
w35026 <= not w34773 and not w35025;
w35027 <= b(20) and not w34762;
w35028 <= not w34760 and w35027;
w35029 <= not w34764 and not w35028;
w35030 <= not w35026 and w35029;
w35031 <= not w34764 and not w35030;
w35032 <= b(21) and not w34753;
w35033 <= not w34751 and w35032;
w35034 <= not w34755 and not w35033;
w35035 <= not w35031 and w35034;
w35036 <= not w34755 and not w35035;
w35037 <= b(22) and not w34744;
w35038 <= not w34742 and w35037;
w35039 <= not w34746 and not w35038;
w35040 <= not w35036 and w35039;
w35041 <= not w34746 and not w35040;
w35042 <= b(23) and not w34735;
w35043 <= not w34733 and w35042;
w35044 <= not w34737 and not w35043;
w35045 <= not w35041 and w35044;
w35046 <= not w34737 and not w35045;
w35047 <= b(24) and not w34726;
w35048 <= not w34724 and w35047;
w35049 <= not w34728 and not w35048;
w35050 <= not w35046 and w35049;
w35051 <= not w34728 and not w35050;
w35052 <= b(25) and not w34717;
w35053 <= not w34715 and w35052;
w35054 <= not w34719 and not w35053;
w35055 <= not w35051 and w35054;
w35056 <= not w34719 and not w35055;
w35057 <= b(26) and not w34708;
w35058 <= not w34706 and w35057;
w35059 <= not w34710 and not w35058;
w35060 <= not w35056 and w35059;
w35061 <= not w34710 and not w35060;
w35062 <= b(27) and not w34699;
w35063 <= not w34697 and w35062;
w35064 <= not w34701 and not w35063;
w35065 <= not w35061 and w35064;
w35066 <= not w34701 and not w35065;
w35067 <= b(28) and not w34690;
w35068 <= not w34688 and w35067;
w35069 <= not w34692 and not w35068;
w35070 <= not w35066 and w35069;
w35071 <= not w34692 and not w35070;
w35072 <= b(29) and not w34670;
w35073 <= not w34668 and w35072;
w35074 <= not w34683 and not w35073;
w35075 <= not w35071 and w35074;
w35076 <= not w34683 and not w35075;
w35077 <= b(30) and not w34680;
w35078 <= not w34678 and w35077;
w35079 <= not w34682 and not w35078;
w35080 <= not w35076 and w35079;
w35081 <= not w34682 and not w35080;
w35082 <= w6905 and not w35081;
w35083 <= not w34671 and not w35082;
w35084 <= not w34692 and w35074;
w35085 <= not w35070 and w35084;
w35086 <= not w35071 and not w35074;
w35087 <= not w35085 and not w35086;
w35088 <= w6905 and not w35087;
w35089 <= not w35081 and w35088;
w35090 <= not w35083 and not w35089;
w35091 <= not w34681 and not w35082;
w35092 <= not w34683 and w35079;
w35093 <= not w35075 and w35092;
w35094 <= not w35076 and not w35079;
w35095 <= not w35093 and not w35094;
w35096 <= w35082 and not w35095;
w35097 <= not w35091 and not w35096;
w35098 <= not b(31) and not w35097;
w35099 <= not b(30) and not w35090;
w35100 <= not w34691 and not w35082;
w35101 <= not w34701 and w35069;
w35102 <= not w35065 and w35101;
w35103 <= not w35066 and not w35069;
w35104 <= not w35102 and not w35103;
w35105 <= w6905 and not w35104;
w35106 <= not w35081 and w35105;
w35107 <= not w35100 and not w35106;
w35108 <= not b(29) and not w35107;
w35109 <= not w34700 and not w35082;
w35110 <= not w34710 and w35064;
w35111 <= not w35060 and w35110;
w35112 <= not w35061 and not w35064;
w35113 <= not w35111 and not w35112;
w35114 <= w6905 and not w35113;
w35115 <= not w35081 and w35114;
w35116 <= not w35109 and not w35115;
w35117 <= not b(28) and not w35116;
w35118 <= not w34709 and not w35082;
w35119 <= not w34719 and w35059;
w35120 <= not w35055 and w35119;
w35121 <= not w35056 and not w35059;
w35122 <= not w35120 and not w35121;
w35123 <= w6905 and not w35122;
w35124 <= not w35081 and w35123;
w35125 <= not w35118 and not w35124;
w35126 <= not b(27) and not w35125;
w35127 <= not w34718 and not w35082;
w35128 <= not w34728 and w35054;
w35129 <= not w35050 and w35128;
w35130 <= not w35051 and not w35054;
w35131 <= not w35129 and not w35130;
w35132 <= w6905 and not w35131;
w35133 <= not w35081 and w35132;
w35134 <= not w35127 and not w35133;
w35135 <= not b(26) and not w35134;
w35136 <= not w34727 and not w35082;
w35137 <= not w34737 and w35049;
w35138 <= not w35045 and w35137;
w35139 <= not w35046 and not w35049;
w35140 <= not w35138 and not w35139;
w35141 <= w6905 and not w35140;
w35142 <= not w35081 and w35141;
w35143 <= not w35136 and not w35142;
w35144 <= not b(25) and not w35143;
w35145 <= not w34736 and not w35082;
w35146 <= not w34746 and w35044;
w35147 <= not w35040 and w35146;
w35148 <= not w35041 and not w35044;
w35149 <= not w35147 and not w35148;
w35150 <= w6905 and not w35149;
w35151 <= not w35081 and w35150;
w35152 <= not w35145 and not w35151;
w35153 <= not b(24) and not w35152;
w35154 <= not w34745 and not w35082;
w35155 <= not w34755 and w35039;
w35156 <= not w35035 and w35155;
w35157 <= not w35036 and not w35039;
w35158 <= not w35156 and not w35157;
w35159 <= w6905 and not w35158;
w35160 <= not w35081 and w35159;
w35161 <= not w35154 and not w35160;
w35162 <= not b(23) and not w35161;
w35163 <= not w34754 and not w35082;
w35164 <= not w34764 and w35034;
w35165 <= not w35030 and w35164;
w35166 <= not w35031 and not w35034;
w35167 <= not w35165 and not w35166;
w35168 <= w6905 and not w35167;
w35169 <= not w35081 and w35168;
w35170 <= not w35163 and not w35169;
w35171 <= not b(22) and not w35170;
w35172 <= not w34763 and not w35082;
w35173 <= not w34773 and w35029;
w35174 <= not w35025 and w35173;
w35175 <= not w35026 and not w35029;
w35176 <= not w35174 and not w35175;
w35177 <= w6905 and not w35176;
w35178 <= not w35081 and w35177;
w35179 <= not w35172 and not w35178;
w35180 <= not b(21) and not w35179;
w35181 <= not w34772 and not w35082;
w35182 <= not w34782 and w35024;
w35183 <= not w35020 and w35182;
w35184 <= not w35021 and not w35024;
w35185 <= not w35183 and not w35184;
w35186 <= w6905 and not w35185;
w35187 <= not w35081 and w35186;
w35188 <= not w35181 and not w35187;
w35189 <= not b(20) and not w35188;
w35190 <= not w34781 and not w35082;
w35191 <= not w34791 and w35019;
w35192 <= not w35015 and w35191;
w35193 <= not w35016 and not w35019;
w35194 <= not w35192 and not w35193;
w35195 <= w6905 and not w35194;
w35196 <= not w35081 and w35195;
w35197 <= not w35190 and not w35196;
w35198 <= not b(19) and not w35197;
w35199 <= not w34790 and not w35082;
w35200 <= not w34800 and w35014;
w35201 <= not w35010 and w35200;
w35202 <= not w35011 and not w35014;
w35203 <= not w35201 and not w35202;
w35204 <= w6905 and not w35203;
w35205 <= not w35081 and w35204;
w35206 <= not w35199 and not w35205;
w35207 <= not b(18) and not w35206;
w35208 <= not w34799 and not w35082;
w35209 <= not w34809 and w35009;
w35210 <= not w35005 and w35209;
w35211 <= not w35006 and not w35009;
w35212 <= not w35210 and not w35211;
w35213 <= w6905 and not w35212;
w35214 <= not w35081 and w35213;
w35215 <= not w35208 and not w35214;
w35216 <= not b(17) and not w35215;
w35217 <= not w34808 and not w35082;
w35218 <= not w34818 and w35004;
w35219 <= not w35000 and w35218;
w35220 <= not w35001 and not w35004;
w35221 <= not w35219 and not w35220;
w35222 <= w6905 and not w35221;
w35223 <= not w35081 and w35222;
w35224 <= not w35217 and not w35223;
w35225 <= not b(16) and not w35224;
w35226 <= not w34817 and not w35082;
w35227 <= not w34827 and w34999;
w35228 <= not w34995 and w35227;
w35229 <= not w34996 and not w34999;
w35230 <= not w35228 and not w35229;
w35231 <= w6905 and not w35230;
w35232 <= not w35081 and w35231;
w35233 <= not w35226 and not w35232;
w35234 <= not b(15) and not w35233;
w35235 <= not w34826 and not w35082;
w35236 <= not w34836 and w34994;
w35237 <= not w34990 and w35236;
w35238 <= not w34991 and not w34994;
w35239 <= not w35237 and not w35238;
w35240 <= w6905 and not w35239;
w35241 <= not w35081 and w35240;
w35242 <= not w35235 and not w35241;
w35243 <= not b(14) and not w35242;
w35244 <= not w34835 and not w35082;
w35245 <= not w34845 and w34989;
w35246 <= not w34985 and w35245;
w35247 <= not w34986 and not w34989;
w35248 <= not w35246 and not w35247;
w35249 <= w6905 and not w35248;
w35250 <= not w35081 and w35249;
w35251 <= not w35244 and not w35250;
w35252 <= not b(13) and not w35251;
w35253 <= not w34844 and not w35082;
w35254 <= not w34854 and w34984;
w35255 <= not w34980 and w35254;
w35256 <= not w34981 and not w34984;
w35257 <= not w35255 and not w35256;
w35258 <= w6905 and not w35257;
w35259 <= not w35081 and w35258;
w35260 <= not w35253 and not w35259;
w35261 <= not b(12) and not w35260;
w35262 <= not w34853 and not w35082;
w35263 <= not w34863 and w34979;
w35264 <= not w34975 and w35263;
w35265 <= not w34976 and not w34979;
w35266 <= not w35264 and not w35265;
w35267 <= w6905 and not w35266;
w35268 <= not w35081 and w35267;
w35269 <= not w35262 and not w35268;
w35270 <= not b(11) and not w35269;
w35271 <= not w34862 and not w35082;
w35272 <= not w34872 and w34974;
w35273 <= not w34970 and w35272;
w35274 <= not w34971 and not w34974;
w35275 <= not w35273 and not w35274;
w35276 <= w6905 and not w35275;
w35277 <= not w35081 and w35276;
w35278 <= not w35271 and not w35277;
w35279 <= not b(10) and not w35278;
w35280 <= not w34871 and not w35082;
w35281 <= not w34881 and w34969;
w35282 <= not w34965 and w35281;
w35283 <= not w34966 and not w34969;
w35284 <= not w35282 and not w35283;
w35285 <= w6905 and not w35284;
w35286 <= not w35081 and w35285;
w35287 <= not w35280 and not w35286;
w35288 <= not b(9) and not w35287;
w35289 <= not w34880 and not w35082;
w35290 <= not w34890 and w34964;
w35291 <= not w34960 and w35290;
w35292 <= not w34961 and not w34964;
w35293 <= not w35291 and not w35292;
w35294 <= w6905 and not w35293;
w35295 <= not w35081 and w35294;
w35296 <= not w35289 and not w35295;
w35297 <= not b(8) and not w35296;
w35298 <= not w34889 and not w35082;
w35299 <= not w34899 and w34959;
w35300 <= not w34955 and w35299;
w35301 <= not w34956 and not w34959;
w35302 <= not w35300 and not w35301;
w35303 <= w6905 and not w35302;
w35304 <= not w35081 and w35303;
w35305 <= not w35298 and not w35304;
w35306 <= not b(7) and not w35305;
w35307 <= not w34898 and not w35082;
w35308 <= not w34908 and w34954;
w35309 <= not w34950 and w35308;
w35310 <= not w34951 and not w34954;
w35311 <= not w35309 and not w35310;
w35312 <= w6905 and not w35311;
w35313 <= not w35081 and w35312;
w35314 <= not w35307 and not w35313;
w35315 <= not b(6) and not w35314;
w35316 <= not w34907 and not w35082;
w35317 <= not w34917 and w34949;
w35318 <= not w34945 and w35317;
w35319 <= not w34946 and not w34949;
w35320 <= not w35318 and not w35319;
w35321 <= w6905 and not w35320;
w35322 <= not w35081 and w35321;
w35323 <= not w35316 and not w35322;
w35324 <= not b(5) and not w35323;
w35325 <= not w34916 and not w35082;
w35326 <= not w34925 and w34944;
w35327 <= not w34940 and w35326;
w35328 <= not w34941 and not w34944;
w35329 <= not w35327 and not w35328;
w35330 <= w6905 and not w35329;
w35331 <= not w35081 and w35330;
w35332 <= not w35325 and not w35331;
w35333 <= not b(4) and not w35332;
w35334 <= not w34924 and not w35082;
w35335 <= not w34935 and w34939;
w35336 <= not w34934 and w35335;
w35337 <= not w34936 and not w34939;
w35338 <= not w35336 and not w35337;
w35339 <= w6905 and not w35338;
w35340 <= not w35081 and w35339;
w35341 <= not w35334 and not w35340;
w35342 <= not b(3) and not w35341;
w35343 <= not w34929 and not w35082;
w35344 <= w6754 and not w34932;
w35345 <= not w34930 and w35344;
w35346 <= w6905 and not w35345;
w35347 <= not w34934 and w35346;
w35348 <= not w35081 and w35347;
w35349 <= not w35343 and not w35348;
w35350 <= not b(2) and not w35349;
w35351 <= w7178 and not w35081;
w35352 <= a(33) and not w35351;
w35353 <= w7184 and not w35081;
w35354 <= not w35352 and not w35353;
w35355 <= b(1) and not w35354;
w35356 <= not b(1) and not w35353;
w35357 <= not w35352 and w35356;
w35358 <= not w35355 and not w35357;
w35359 <= not w7191 and not w35358;
w35360 <= not b(1) and not w35354;
w35361 <= not w35359 and not w35360;
w35362 <= b(2) and not w35348;
w35363 <= not w35343 and w35362;
w35364 <= not w35350 and not w35363;
w35365 <= not w35361 and w35364;
w35366 <= not w35350 and not w35365;
w35367 <= b(3) and not w35340;
w35368 <= not w35334 and w35367;
w35369 <= not w35342 and not w35368;
w35370 <= not w35366 and w35369;
w35371 <= not w35342 and not w35370;
w35372 <= b(4) and not w35331;
w35373 <= not w35325 and w35372;
w35374 <= not w35333 and not w35373;
w35375 <= not w35371 and w35374;
w35376 <= not w35333 and not w35375;
w35377 <= b(5) and not w35322;
w35378 <= not w35316 and w35377;
w35379 <= not w35324 and not w35378;
w35380 <= not w35376 and w35379;
w35381 <= not w35324 and not w35380;
w35382 <= b(6) and not w35313;
w35383 <= not w35307 and w35382;
w35384 <= not w35315 and not w35383;
w35385 <= not w35381 and w35384;
w35386 <= not w35315 and not w35385;
w35387 <= b(7) and not w35304;
w35388 <= not w35298 and w35387;
w35389 <= not w35306 and not w35388;
w35390 <= not w35386 and w35389;
w35391 <= not w35306 and not w35390;
w35392 <= b(8) and not w35295;
w35393 <= not w35289 and w35392;
w35394 <= not w35297 and not w35393;
w35395 <= not w35391 and w35394;
w35396 <= not w35297 and not w35395;
w35397 <= b(9) and not w35286;
w35398 <= not w35280 and w35397;
w35399 <= not w35288 and not w35398;
w35400 <= not w35396 and w35399;
w35401 <= not w35288 and not w35400;
w35402 <= b(10) and not w35277;
w35403 <= not w35271 and w35402;
w35404 <= not w35279 and not w35403;
w35405 <= not w35401 and w35404;
w35406 <= not w35279 and not w35405;
w35407 <= b(11) and not w35268;
w35408 <= not w35262 and w35407;
w35409 <= not w35270 and not w35408;
w35410 <= not w35406 and w35409;
w35411 <= not w35270 and not w35410;
w35412 <= b(12) and not w35259;
w35413 <= not w35253 and w35412;
w35414 <= not w35261 and not w35413;
w35415 <= not w35411 and w35414;
w35416 <= not w35261 and not w35415;
w35417 <= b(13) and not w35250;
w35418 <= not w35244 and w35417;
w35419 <= not w35252 and not w35418;
w35420 <= not w35416 and w35419;
w35421 <= not w35252 and not w35420;
w35422 <= b(14) and not w35241;
w35423 <= not w35235 and w35422;
w35424 <= not w35243 and not w35423;
w35425 <= not w35421 and w35424;
w35426 <= not w35243 and not w35425;
w35427 <= b(15) and not w35232;
w35428 <= not w35226 and w35427;
w35429 <= not w35234 and not w35428;
w35430 <= not w35426 and w35429;
w35431 <= not w35234 and not w35430;
w35432 <= b(16) and not w35223;
w35433 <= not w35217 and w35432;
w35434 <= not w35225 and not w35433;
w35435 <= not w35431 and w35434;
w35436 <= not w35225 and not w35435;
w35437 <= b(17) and not w35214;
w35438 <= not w35208 and w35437;
w35439 <= not w35216 and not w35438;
w35440 <= not w35436 and w35439;
w35441 <= not w35216 and not w35440;
w35442 <= b(18) and not w35205;
w35443 <= not w35199 and w35442;
w35444 <= not w35207 and not w35443;
w35445 <= not w35441 and w35444;
w35446 <= not w35207 and not w35445;
w35447 <= b(19) and not w35196;
w35448 <= not w35190 and w35447;
w35449 <= not w35198 and not w35448;
w35450 <= not w35446 and w35449;
w35451 <= not w35198 and not w35450;
w35452 <= b(20) and not w35187;
w35453 <= not w35181 and w35452;
w35454 <= not w35189 and not w35453;
w35455 <= not w35451 and w35454;
w35456 <= not w35189 and not w35455;
w35457 <= b(21) and not w35178;
w35458 <= not w35172 and w35457;
w35459 <= not w35180 and not w35458;
w35460 <= not w35456 and w35459;
w35461 <= not w35180 and not w35460;
w35462 <= b(22) and not w35169;
w35463 <= not w35163 and w35462;
w35464 <= not w35171 and not w35463;
w35465 <= not w35461 and w35464;
w35466 <= not w35171 and not w35465;
w35467 <= b(23) and not w35160;
w35468 <= not w35154 and w35467;
w35469 <= not w35162 and not w35468;
w35470 <= not w35466 and w35469;
w35471 <= not w35162 and not w35470;
w35472 <= b(24) and not w35151;
w35473 <= not w35145 and w35472;
w35474 <= not w35153 and not w35473;
w35475 <= not w35471 and w35474;
w35476 <= not w35153 and not w35475;
w35477 <= b(25) and not w35142;
w35478 <= not w35136 and w35477;
w35479 <= not w35144 and not w35478;
w35480 <= not w35476 and w35479;
w35481 <= not w35144 and not w35480;
w35482 <= b(26) and not w35133;
w35483 <= not w35127 and w35482;
w35484 <= not w35135 and not w35483;
w35485 <= not w35481 and w35484;
w35486 <= not w35135 and not w35485;
w35487 <= b(27) and not w35124;
w35488 <= not w35118 and w35487;
w35489 <= not w35126 and not w35488;
w35490 <= not w35486 and w35489;
w35491 <= not w35126 and not w35490;
w35492 <= b(28) and not w35115;
w35493 <= not w35109 and w35492;
w35494 <= not w35117 and not w35493;
w35495 <= not w35491 and w35494;
w35496 <= not w35117 and not w35495;
w35497 <= b(29) and not w35106;
w35498 <= not w35100 and w35497;
w35499 <= not w35108 and not w35498;
w35500 <= not w35496 and w35499;
w35501 <= not w35108 and not w35500;
w35502 <= b(30) and not w35089;
w35503 <= not w35083 and w35502;
w35504 <= not w35099 and not w35503;
w35505 <= not w35501 and w35504;
w35506 <= not w35099 and not w35505;
w35507 <= b(31) and not w35091;
w35508 <= not w35096 and w35507;
w35509 <= not w35098 and not w35508;
w35510 <= not w35506 and w35509;
w35511 <= not w35098 and not w35510;
w35512 <= w175 and not w35511;
w35513 <= not w35090 and not w35512;
w35514 <= not w35108 and w35504;
w35515 <= not w35500 and w35514;
w35516 <= not w35501 and not w35504;
w35517 <= not w35515 and not w35516;
w35518 <= w175 and not w35517;
w35519 <= not w35511 and w35518;
w35520 <= not w35513 and not w35519;
w35521 <= not b(31) and not w35520;
w35522 <= not w35107 and not w35512;
w35523 <= not w35117 and w35499;
w35524 <= not w35495 and w35523;
w35525 <= not w35496 and not w35499;
w35526 <= not w35524 and not w35525;
w35527 <= w175 and not w35526;
w35528 <= not w35511 and w35527;
w35529 <= not w35522 and not w35528;
w35530 <= not b(30) and not w35529;
w35531 <= not w35116 and not w35512;
w35532 <= not w35126 and w35494;
w35533 <= not w35490 and w35532;
w35534 <= not w35491 and not w35494;
w35535 <= not w35533 and not w35534;
w35536 <= w175 and not w35535;
w35537 <= not w35511 and w35536;
w35538 <= not w35531 and not w35537;
w35539 <= not b(29) and not w35538;
w35540 <= not w35125 and not w35512;
w35541 <= not w35135 and w35489;
w35542 <= not w35485 and w35541;
w35543 <= not w35486 and not w35489;
w35544 <= not w35542 and not w35543;
w35545 <= w175 and not w35544;
w35546 <= not w35511 and w35545;
w35547 <= not w35540 and not w35546;
w35548 <= not b(28) and not w35547;
w35549 <= not w35134 and not w35512;
w35550 <= not w35144 and w35484;
w35551 <= not w35480 and w35550;
w35552 <= not w35481 and not w35484;
w35553 <= not w35551 and not w35552;
w35554 <= w175 and not w35553;
w35555 <= not w35511 and w35554;
w35556 <= not w35549 and not w35555;
w35557 <= not b(27) and not w35556;
w35558 <= not w35143 and not w35512;
w35559 <= not w35153 and w35479;
w35560 <= not w35475 and w35559;
w35561 <= not w35476 and not w35479;
w35562 <= not w35560 and not w35561;
w35563 <= w175 and not w35562;
w35564 <= not w35511 and w35563;
w35565 <= not w35558 and not w35564;
w35566 <= not b(26) and not w35565;
w35567 <= not w35152 and not w35512;
w35568 <= not w35162 and w35474;
w35569 <= not w35470 and w35568;
w35570 <= not w35471 and not w35474;
w35571 <= not w35569 and not w35570;
w35572 <= w175 and not w35571;
w35573 <= not w35511 and w35572;
w35574 <= not w35567 and not w35573;
w35575 <= not b(25) and not w35574;
w35576 <= not w35161 and not w35512;
w35577 <= not w35171 and w35469;
w35578 <= not w35465 and w35577;
w35579 <= not w35466 and not w35469;
w35580 <= not w35578 and not w35579;
w35581 <= w175 and not w35580;
w35582 <= not w35511 and w35581;
w35583 <= not w35576 and not w35582;
w35584 <= not b(24) and not w35583;
w35585 <= not w35170 and not w35512;
w35586 <= not w35180 and w35464;
w35587 <= not w35460 and w35586;
w35588 <= not w35461 and not w35464;
w35589 <= not w35587 and not w35588;
w35590 <= w175 and not w35589;
w35591 <= not w35511 and w35590;
w35592 <= not w35585 and not w35591;
w35593 <= not b(23) and not w35592;
w35594 <= not w35179 and not w35512;
w35595 <= not w35189 and w35459;
w35596 <= not w35455 and w35595;
w35597 <= not w35456 and not w35459;
w35598 <= not w35596 and not w35597;
w35599 <= w175 and not w35598;
w35600 <= not w35511 and w35599;
w35601 <= not w35594 and not w35600;
w35602 <= not b(22) and not w35601;
w35603 <= not w35188 and not w35512;
w35604 <= not w35198 and w35454;
w35605 <= not w35450 and w35604;
w35606 <= not w35451 and not w35454;
w35607 <= not w35605 and not w35606;
w35608 <= w175 and not w35607;
w35609 <= not w35511 and w35608;
w35610 <= not w35603 and not w35609;
w35611 <= not b(21) and not w35610;
w35612 <= not w35197 and not w35512;
w35613 <= not w35207 and w35449;
w35614 <= not w35445 and w35613;
w35615 <= not w35446 and not w35449;
w35616 <= not w35614 and not w35615;
w35617 <= w175 and not w35616;
w35618 <= not w35511 and w35617;
w35619 <= not w35612 and not w35618;
w35620 <= not b(20) and not w35619;
w35621 <= not w35206 and not w35512;
w35622 <= not w35216 and w35444;
w35623 <= not w35440 and w35622;
w35624 <= not w35441 and not w35444;
w35625 <= not w35623 and not w35624;
w35626 <= w175 and not w35625;
w35627 <= not w35511 and w35626;
w35628 <= not w35621 and not w35627;
w35629 <= not b(19) and not w35628;
w35630 <= not w35215 and not w35512;
w35631 <= not w35225 and w35439;
w35632 <= not w35435 and w35631;
w35633 <= not w35436 and not w35439;
w35634 <= not w35632 and not w35633;
w35635 <= w175 and not w35634;
w35636 <= not w35511 and w35635;
w35637 <= not w35630 and not w35636;
w35638 <= not b(18) and not w35637;
w35639 <= not w35224 and not w35512;
w35640 <= not w35234 and w35434;
w35641 <= not w35430 and w35640;
w35642 <= not w35431 and not w35434;
w35643 <= not w35641 and not w35642;
w35644 <= w175 and not w35643;
w35645 <= not w35511 and w35644;
w35646 <= not w35639 and not w35645;
w35647 <= not b(17) and not w35646;
w35648 <= not w35233 and not w35512;
w35649 <= not w35243 and w35429;
w35650 <= not w35425 and w35649;
w35651 <= not w35426 and not w35429;
w35652 <= not w35650 and not w35651;
w35653 <= w175 and not w35652;
w35654 <= not w35511 and w35653;
w35655 <= not w35648 and not w35654;
w35656 <= not b(16) and not w35655;
w35657 <= not w35242 and not w35512;
w35658 <= not w35252 and w35424;
w35659 <= not w35420 and w35658;
w35660 <= not w35421 and not w35424;
w35661 <= not w35659 and not w35660;
w35662 <= w175 and not w35661;
w35663 <= not w35511 and w35662;
w35664 <= not w35657 and not w35663;
w35665 <= not b(15) and not w35664;
w35666 <= not w35251 and not w35512;
w35667 <= not w35261 and w35419;
w35668 <= not w35415 and w35667;
w35669 <= not w35416 and not w35419;
w35670 <= not w35668 and not w35669;
w35671 <= w175 and not w35670;
w35672 <= not w35511 and w35671;
w35673 <= not w35666 and not w35672;
w35674 <= not b(14) and not w35673;
w35675 <= not w35260 and not w35512;
w35676 <= not w35270 and w35414;
w35677 <= not w35410 and w35676;
w35678 <= not w35411 and not w35414;
w35679 <= not w35677 and not w35678;
w35680 <= w175 and not w35679;
w35681 <= not w35511 and w35680;
w35682 <= not w35675 and not w35681;
w35683 <= not b(13) and not w35682;
w35684 <= not w35269 and not w35512;
w35685 <= not w35279 and w35409;
w35686 <= not w35405 and w35685;
w35687 <= not w35406 and not w35409;
w35688 <= not w35686 and not w35687;
w35689 <= w175 and not w35688;
w35690 <= not w35511 and w35689;
w35691 <= not w35684 and not w35690;
w35692 <= not b(12) and not w35691;
w35693 <= not w35278 and not w35512;
w35694 <= not w35288 and w35404;
w35695 <= not w35400 and w35694;
w35696 <= not w35401 and not w35404;
w35697 <= not w35695 and not w35696;
w35698 <= w175 and not w35697;
w35699 <= not w35511 and w35698;
w35700 <= not w35693 and not w35699;
w35701 <= not b(11) and not w35700;
w35702 <= not w35287 and not w35512;
w35703 <= not w35297 and w35399;
w35704 <= not w35395 and w35703;
w35705 <= not w35396 and not w35399;
w35706 <= not w35704 and not w35705;
w35707 <= w175 and not w35706;
w35708 <= not w35511 and w35707;
w35709 <= not w35702 and not w35708;
w35710 <= not b(10) and not w35709;
w35711 <= not w35296 and not w35512;
w35712 <= not w35306 and w35394;
w35713 <= not w35390 and w35712;
w35714 <= not w35391 and not w35394;
w35715 <= not w35713 and not w35714;
w35716 <= w175 and not w35715;
w35717 <= not w35511 and w35716;
w35718 <= not w35711 and not w35717;
w35719 <= not b(9) and not w35718;
w35720 <= not w35305 and not w35512;
w35721 <= not w35315 and w35389;
w35722 <= not w35385 and w35721;
w35723 <= not w35386 and not w35389;
w35724 <= not w35722 and not w35723;
w35725 <= w175 and not w35724;
w35726 <= not w35511 and w35725;
w35727 <= not w35720 and not w35726;
w35728 <= not b(8) and not w35727;
w35729 <= not w35314 and not w35512;
w35730 <= not w35324 and w35384;
w35731 <= not w35380 and w35730;
w35732 <= not w35381 and not w35384;
w35733 <= not w35731 and not w35732;
w35734 <= w175 and not w35733;
w35735 <= not w35511 and w35734;
w35736 <= not w35729 and not w35735;
w35737 <= not b(7) and not w35736;
w35738 <= not w35323 and not w35512;
w35739 <= not w35333 and w35379;
w35740 <= not w35375 and w35739;
w35741 <= not w35376 and not w35379;
w35742 <= not w35740 and not w35741;
w35743 <= w175 and not w35742;
w35744 <= not w35511 and w35743;
w35745 <= not w35738 and not w35744;
w35746 <= not b(6) and not w35745;
w35747 <= not w35332 and not w35512;
w35748 <= not w35342 and w35374;
w35749 <= not w35370 and w35748;
w35750 <= not w35371 and not w35374;
w35751 <= not w35749 and not w35750;
w35752 <= w175 and not w35751;
w35753 <= not w35511 and w35752;
w35754 <= not w35747 and not w35753;
w35755 <= not b(5) and not w35754;
w35756 <= not w35341 and not w35512;
w35757 <= not w35350 and w35369;
w35758 <= not w35365 and w35757;
w35759 <= not w35366 and not w35369;
w35760 <= not w35758 and not w35759;
w35761 <= w175 and not w35760;
w35762 <= not w35511 and w35761;
w35763 <= not w35756 and not w35762;
w35764 <= not b(4) and not w35763;
w35765 <= not w35349 and not w35512;
w35766 <= not w35360 and w35364;
w35767 <= not w35359 and w35766;
w35768 <= not w35361 and not w35364;
w35769 <= not w35767 and not w35768;
w35770 <= w175 and not w35769;
w35771 <= not w35511 and w35770;
w35772 <= not w35765 and not w35771;
w35773 <= not b(3) and not w35772;
w35774 <= not w35354 and not w35512;
w35775 <= w7191 and not w35357;
w35776 <= not w35355 and w35775;
w35777 <= w175 and not w35776;
w35778 <= not w35359 and w35777;
w35779 <= not w35511 and w35778;
w35780 <= not w35774 and not w35779;
w35781 <= not b(2) and not w35780;
w35782 <= w7618 and not w35511;
w35783 <= a(32) and not w35782;
w35784 <= w7623 and not w35511;
w35785 <= not w35783 and not w35784;
w35786 <= b(1) and not w35785;
w35787 <= not b(1) and not w35784;
w35788 <= not w35783 and w35787;
w35789 <= not w35786 and not w35788;
w35790 <= not w7630 and not w35789;
w35791 <= not b(1) and not w35785;
w35792 <= not w35790 and not w35791;
w35793 <= b(2) and not w35779;
w35794 <= not w35774 and w35793;
w35795 <= not w35781 and not w35794;
w35796 <= not w35792 and w35795;
w35797 <= not w35781 and not w35796;
w35798 <= b(3) and not w35771;
w35799 <= not w35765 and w35798;
w35800 <= not w35773 and not w35799;
w35801 <= not w35797 and w35800;
w35802 <= not w35773 and not w35801;
w35803 <= b(4) and not w35762;
w35804 <= not w35756 and w35803;
w35805 <= not w35764 and not w35804;
w35806 <= not w35802 and w35805;
w35807 <= not w35764 and not w35806;
w35808 <= b(5) and not w35753;
w35809 <= not w35747 and w35808;
w35810 <= not w35755 and not w35809;
w35811 <= not w35807 and w35810;
w35812 <= not w35755 and not w35811;
w35813 <= b(6) and not w35744;
w35814 <= not w35738 and w35813;
w35815 <= not w35746 and not w35814;
w35816 <= not w35812 and w35815;
w35817 <= not w35746 and not w35816;
w35818 <= b(7) and not w35735;
w35819 <= not w35729 and w35818;
w35820 <= not w35737 and not w35819;
w35821 <= not w35817 and w35820;
w35822 <= not w35737 and not w35821;
w35823 <= b(8) and not w35726;
w35824 <= not w35720 and w35823;
w35825 <= not w35728 and not w35824;
w35826 <= not w35822 and w35825;
w35827 <= not w35728 and not w35826;
w35828 <= b(9) and not w35717;
w35829 <= not w35711 and w35828;
w35830 <= not w35719 and not w35829;
w35831 <= not w35827 and w35830;
w35832 <= not w35719 and not w35831;
w35833 <= b(10) and not w35708;
w35834 <= not w35702 and w35833;
w35835 <= not w35710 and not w35834;
w35836 <= not w35832 and w35835;
w35837 <= not w35710 and not w35836;
w35838 <= b(11) and not w35699;
w35839 <= not w35693 and w35838;
w35840 <= not w35701 and not w35839;
w35841 <= not w35837 and w35840;
w35842 <= not w35701 and not w35841;
w35843 <= b(12) and not w35690;
w35844 <= not w35684 and w35843;
w35845 <= not w35692 and not w35844;
w35846 <= not w35842 and w35845;
w35847 <= not w35692 and not w35846;
w35848 <= b(13) and not w35681;
w35849 <= not w35675 and w35848;
w35850 <= not w35683 and not w35849;
w35851 <= not w35847 and w35850;
w35852 <= not w35683 and not w35851;
w35853 <= b(14) and not w35672;
w35854 <= not w35666 and w35853;
w35855 <= not w35674 and not w35854;
w35856 <= not w35852 and w35855;
w35857 <= not w35674 and not w35856;
w35858 <= b(15) and not w35663;
w35859 <= not w35657 and w35858;
w35860 <= not w35665 and not w35859;
w35861 <= not w35857 and w35860;
w35862 <= not w35665 and not w35861;
w35863 <= b(16) and not w35654;
w35864 <= not w35648 and w35863;
w35865 <= not w35656 and not w35864;
w35866 <= not w35862 and w35865;
w35867 <= not w35656 and not w35866;
w35868 <= b(17) and not w35645;
w35869 <= not w35639 and w35868;
w35870 <= not w35647 and not w35869;
w35871 <= not w35867 and w35870;
w35872 <= not w35647 and not w35871;
w35873 <= b(18) and not w35636;
w35874 <= not w35630 and w35873;
w35875 <= not w35638 and not w35874;
w35876 <= not w35872 and w35875;
w35877 <= not w35638 and not w35876;
w35878 <= b(19) and not w35627;
w35879 <= not w35621 and w35878;
w35880 <= not w35629 and not w35879;
w35881 <= not w35877 and w35880;
w35882 <= not w35629 and not w35881;
w35883 <= b(20) and not w35618;
w35884 <= not w35612 and w35883;
w35885 <= not w35620 and not w35884;
w35886 <= not w35882 and w35885;
w35887 <= not w35620 and not w35886;
w35888 <= b(21) and not w35609;
w35889 <= not w35603 and w35888;
w35890 <= not w35611 and not w35889;
w35891 <= not w35887 and w35890;
w35892 <= not w35611 and not w35891;
w35893 <= b(22) and not w35600;
w35894 <= not w35594 and w35893;
w35895 <= not w35602 and not w35894;
w35896 <= not w35892 and w35895;
w35897 <= not w35602 and not w35896;
w35898 <= b(23) and not w35591;
w35899 <= not w35585 and w35898;
w35900 <= not w35593 and not w35899;
w35901 <= not w35897 and w35900;
w35902 <= not w35593 and not w35901;
w35903 <= b(24) and not w35582;
w35904 <= not w35576 and w35903;
w35905 <= not w35584 and not w35904;
w35906 <= not w35902 and w35905;
w35907 <= not w35584 and not w35906;
w35908 <= b(25) and not w35573;
w35909 <= not w35567 and w35908;
w35910 <= not w35575 and not w35909;
w35911 <= not w35907 and w35910;
w35912 <= not w35575 and not w35911;
w35913 <= b(26) and not w35564;
w35914 <= not w35558 and w35913;
w35915 <= not w35566 and not w35914;
w35916 <= not w35912 and w35915;
w35917 <= not w35566 and not w35916;
w35918 <= b(27) and not w35555;
w35919 <= not w35549 and w35918;
w35920 <= not w35557 and not w35919;
w35921 <= not w35917 and w35920;
w35922 <= not w35557 and not w35921;
w35923 <= b(28) and not w35546;
w35924 <= not w35540 and w35923;
w35925 <= not w35548 and not w35924;
w35926 <= not w35922 and w35925;
w35927 <= not w35548 and not w35926;
w35928 <= b(29) and not w35537;
w35929 <= not w35531 and w35928;
w35930 <= not w35539 and not w35929;
w35931 <= not w35927 and w35930;
w35932 <= not w35539 and not w35931;
w35933 <= b(30) and not w35528;
w35934 <= not w35522 and w35933;
w35935 <= not w35530 and not w35934;
w35936 <= not w35932 and w35935;
w35937 <= not w35530 and not w35936;
w35938 <= b(31) and not w35519;
w35939 <= not w35513 and w35938;
w35940 <= not w35521 and not w35939;
w35941 <= not w35937 and w35940;
w35942 <= not w35521 and not w35941;
w35943 <= not w35097 and not w35512;
w35944 <= not w35099 and w35509;
w35945 <= not w35505 and w35944;
w35946 <= not w35506 and not w35509;
w35947 <= not w35945 and not w35946;
w35948 <= w35512 and not w35947;
w35949 <= not w35943 and not w35948;
w35950 <= not b(32) and not w35949;
w35951 <= b(32) and not w35943;
w35952 <= not w35948 and w35951;
w35953 <= w167 and not w35952;
w35954 <= not w35950 and w35953;
w35955 <= not w35942 and w35954;
w35956 <= w175 and not w35949;
w35957 <= not w35955 and not w35956;
w35958 <= not w35530 and w35940;
w35959 <= not w35936 and w35958;
w35960 <= not w35937 and not w35940;
w35961 <= not w35959 and not w35960;
w35962 <= not w35957 and not w35961;
w35963 <= not w35520 and not w35956;
w35964 <= not w35955 and w35963;
w35965 <= not w35962 and not w35964;
w35966 <= not w35521 and not w35952;
w35967 <= not w35950 and w35966;
w35968 <= not w35941 and w35967;
w35969 <= not w35950 and not w35952;
w35970 <= not w35942 and not w35969;
w35971 <= not w35968 and not w35970;
w35972 <= not w35957 and not w35971;
w35973 <= not w35949 and not w35956;
w35974 <= not w35955 and w35973;
w35975 <= not w35972 and not w35974;
w35976 <= not b(33) and not w35975;
w35977 <= not b(32) and not w35965;
w35978 <= not w35539 and w35935;
w35979 <= not w35931 and w35978;
w35980 <= not w35932 and not w35935;
w35981 <= not w35979 and not w35980;
w35982 <= not w35957 and not w35981;
w35983 <= not w35529 and not w35956;
w35984 <= not w35955 and w35983;
w35985 <= not w35982 and not w35984;
w35986 <= not b(31) and not w35985;
w35987 <= not w35548 and w35930;
w35988 <= not w35926 and w35987;
w35989 <= not w35927 and not w35930;
w35990 <= not w35988 and not w35989;
w35991 <= not w35957 and not w35990;
w35992 <= not w35538 and not w35956;
w35993 <= not w35955 and w35992;
w35994 <= not w35991 and not w35993;
w35995 <= not b(30) and not w35994;
w35996 <= not w35557 and w35925;
w35997 <= not w35921 and w35996;
w35998 <= not w35922 and not w35925;
w35999 <= not w35997 and not w35998;
w36000 <= not w35957 and not w35999;
w36001 <= not w35547 and not w35956;
w36002 <= not w35955 and w36001;
w36003 <= not w36000 and not w36002;
w36004 <= not b(29) and not w36003;
w36005 <= not w35566 and w35920;
w36006 <= not w35916 and w36005;
w36007 <= not w35917 and not w35920;
w36008 <= not w36006 and not w36007;
w36009 <= not w35957 and not w36008;
w36010 <= not w35556 and not w35956;
w36011 <= not w35955 and w36010;
w36012 <= not w36009 and not w36011;
w36013 <= not b(28) and not w36012;
w36014 <= not w35575 and w35915;
w36015 <= not w35911 and w36014;
w36016 <= not w35912 and not w35915;
w36017 <= not w36015 and not w36016;
w36018 <= not w35957 and not w36017;
w36019 <= not w35565 and not w35956;
w36020 <= not w35955 and w36019;
w36021 <= not w36018 and not w36020;
w36022 <= not b(27) and not w36021;
w36023 <= not w35584 and w35910;
w36024 <= not w35906 and w36023;
w36025 <= not w35907 and not w35910;
w36026 <= not w36024 and not w36025;
w36027 <= not w35957 and not w36026;
w36028 <= not w35574 and not w35956;
w36029 <= not w35955 and w36028;
w36030 <= not w36027 and not w36029;
w36031 <= not b(26) and not w36030;
w36032 <= not w35593 and w35905;
w36033 <= not w35901 and w36032;
w36034 <= not w35902 and not w35905;
w36035 <= not w36033 and not w36034;
w36036 <= not w35957 and not w36035;
w36037 <= not w35583 and not w35956;
w36038 <= not w35955 and w36037;
w36039 <= not w36036 and not w36038;
w36040 <= not b(25) and not w36039;
w36041 <= not w35602 and w35900;
w36042 <= not w35896 and w36041;
w36043 <= not w35897 and not w35900;
w36044 <= not w36042 and not w36043;
w36045 <= not w35957 and not w36044;
w36046 <= not w35592 and not w35956;
w36047 <= not w35955 and w36046;
w36048 <= not w36045 and not w36047;
w36049 <= not b(24) and not w36048;
w36050 <= not w35611 and w35895;
w36051 <= not w35891 and w36050;
w36052 <= not w35892 and not w35895;
w36053 <= not w36051 and not w36052;
w36054 <= not w35957 and not w36053;
w36055 <= not w35601 and not w35956;
w36056 <= not w35955 and w36055;
w36057 <= not w36054 and not w36056;
w36058 <= not b(23) and not w36057;
w36059 <= not w35620 and w35890;
w36060 <= not w35886 and w36059;
w36061 <= not w35887 and not w35890;
w36062 <= not w36060 and not w36061;
w36063 <= not w35957 and not w36062;
w36064 <= not w35610 and not w35956;
w36065 <= not w35955 and w36064;
w36066 <= not w36063 and not w36065;
w36067 <= not b(22) and not w36066;
w36068 <= not w35629 and w35885;
w36069 <= not w35881 and w36068;
w36070 <= not w35882 and not w35885;
w36071 <= not w36069 and not w36070;
w36072 <= not w35957 and not w36071;
w36073 <= not w35619 and not w35956;
w36074 <= not w35955 and w36073;
w36075 <= not w36072 and not w36074;
w36076 <= not b(21) and not w36075;
w36077 <= not w35638 and w35880;
w36078 <= not w35876 and w36077;
w36079 <= not w35877 and not w35880;
w36080 <= not w36078 and not w36079;
w36081 <= not w35957 and not w36080;
w36082 <= not w35628 and not w35956;
w36083 <= not w35955 and w36082;
w36084 <= not w36081 and not w36083;
w36085 <= not b(20) and not w36084;
w36086 <= not w35647 and w35875;
w36087 <= not w35871 and w36086;
w36088 <= not w35872 and not w35875;
w36089 <= not w36087 and not w36088;
w36090 <= not w35957 and not w36089;
w36091 <= not w35637 and not w35956;
w36092 <= not w35955 and w36091;
w36093 <= not w36090 and not w36092;
w36094 <= not b(19) and not w36093;
w36095 <= not w35656 and w35870;
w36096 <= not w35866 and w36095;
w36097 <= not w35867 and not w35870;
w36098 <= not w36096 and not w36097;
w36099 <= not w35957 and not w36098;
w36100 <= not w35646 and not w35956;
w36101 <= not w35955 and w36100;
w36102 <= not w36099 and not w36101;
w36103 <= not b(18) and not w36102;
w36104 <= not w35665 and w35865;
w36105 <= not w35861 and w36104;
w36106 <= not w35862 and not w35865;
w36107 <= not w36105 and not w36106;
w36108 <= not w35957 and not w36107;
w36109 <= not w35655 and not w35956;
w36110 <= not w35955 and w36109;
w36111 <= not w36108 and not w36110;
w36112 <= not b(17) and not w36111;
w36113 <= not w35674 and w35860;
w36114 <= not w35856 and w36113;
w36115 <= not w35857 and not w35860;
w36116 <= not w36114 and not w36115;
w36117 <= not w35957 and not w36116;
w36118 <= not w35664 and not w35956;
w36119 <= not w35955 and w36118;
w36120 <= not w36117 and not w36119;
w36121 <= not b(16) and not w36120;
w36122 <= not w35683 and w35855;
w36123 <= not w35851 and w36122;
w36124 <= not w35852 and not w35855;
w36125 <= not w36123 and not w36124;
w36126 <= not w35957 and not w36125;
w36127 <= not w35673 and not w35956;
w36128 <= not w35955 and w36127;
w36129 <= not w36126 and not w36128;
w36130 <= not b(15) and not w36129;
w36131 <= not w35692 and w35850;
w36132 <= not w35846 and w36131;
w36133 <= not w35847 and not w35850;
w36134 <= not w36132 and not w36133;
w36135 <= not w35957 and not w36134;
w36136 <= not w35682 and not w35956;
w36137 <= not w35955 and w36136;
w36138 <= not w36135 and not w36137;
w36139 <= not b(14) and not w36138;
w36140 <= not w35701 and w35845;
w36141 <= not w35841 and w36140;
w36142 <= not w35842 and not w35845;
w36143 <= not w36141 and not w36142;
w36144 <= not w35957 and not w36143;
w36145 <= not w35691 and not w35956;
w36146 <= not w35955 and w36145;
w36147 <= not w36144 and not w36146;
w36148 <= not b(13) and not w36147;
w36149 <= not w35710 and w35840;
w36150 <= not w35836 and w36149;
w36151 <= not w35837 and not w35840;
w36152 <= not w36150 and not w36151;
w36153 <= not w35957 and not w36152;
w36154 <= not w35700 and not w35956;
w36155 <= not w35955 and w36154;
w36156 <= not w36153 and not w36155;
w36157 <= not b(12) and not w36156;
w36158 <= not w35719 and w35835;
w36159 <= not w35831 and w36158;
w36160 <= not w35832 and not w35835;
w36161 <= not w36159 and not w36160;
w36162 <= not w35957 and not w36161;
w36163 <= not w35709 and not w35956;
w36164 <= not w35955 and w36163;
w36165 <= not w36162 and not w36164;
w36166 <= not b(11) and not w36165;
w36167 <= not w35728 and w35830;
w36168 <= not w35826 and w36167;
w36169 <= not w35827 and not w35830;
w36170 <= not w36168 and not w36169;
w36171 <= not w35957 and not w36170;
w36172 <= not w35718 and not w35956;
w36173 <= not w35955 and w36172;
w36174 <= not w36171 and not w36173;
w36175 <= not b(10) and not w36174;
w36176 <= not w35737 and w35825;
w36177 <= not w35821 and w36176;
w36178 <= not w35822 and not w35825;
w36179 <= not w36177 and not w36178;
w36180 <= not w35957 and not w36179;
w36181 <= not w35727 and not w35956;
w36182 <= not w35955 and w36181;
w36183 <= not w36180 and not w36182;
w36184 <= not b(9) and not w36183;
w36185 <= not w35746 and w35820;
w36186 <= not w35816 and w36185;
w36187 <= not w35817 and not w35820;
w36188 <= not w36186 and not w36187;
w36189 <= not w35957 and not w36188;
w36190 <= not w35736 and not w35956;
w36191 <= not w35955 and w36190;
w36192 <= not w36189 and not w36191;
w36193 <= not b(8) and not w36192;
w36194 <= not w35755 and w35815;
w36195 <= not w35811 and w36194;
w36196 <= not w35812 and not w35815;
w36197 <= not w36195 and not w36196;
w36198 <= not w35957 and not w36197;
w36199 <= not w35745 and not w35956;
w36200 <= not w35955 and w36199;
w36201 <= not w36198 and not w36200;
w36202 <= not b(7) and not w36201;
w36203 <= not w35764 and w35810;
w36204 <= not w35806 and w36203;
w36205 <= not w35807 and not w35810;
w36206 <= not w36204 and not w36205;
w36207 <= not w35957 and not w36206;
w36208 <= not w35754 and not w35956;
w36209 <= not w35955 and w36208;
w36210 <= not w36207 and not w36209;
w36211 <= not b(6) and not w36210;
w36212 <= not w35773 and w35805;
w36213 <= not w35801 and w36212;
w36214 <= not w35802 and not w35805;
w36215 <= not w36213 and not w36214;
w36216 <= not w35957 and not w36215;
w36217 <= not w35763 and not w35956;
w36218 <= not w35955 and w36217;
w36219 <= not w36216 and not w36218;
w36220 <= not b(5) and not w36219;
w36221 <= not w35781 and w35800;
w36222 <= not w35796 and w36221;
w36223 <= not w35797 and not w35800;
w36224 <= not w36222 and not w36223;
w36225 <= not w35957 and not w36224;
w36226 <= not w35772 and not w35956;
w36227 <= not w35955 and w36226;
w36228 <= not w36225 and not w36227;
w36229 <= not b(4) and not w36228;
w36230 <= not w35791 and w35795;
w36231 <= not w35790 and w36230;
w36232 <= not w35792 and not w35795;
w36233 <= not w36231 and not w36232;
w36234 <= not w35957 and not w36233;
w36235 <= not w35780 and not w35956;
w36236 <= not w35955 and w36235;
w36237 <= not w36234 and not w36236;
w36238 <= not b(3) and not w36237;
w36239 <= w7630 and not w35788;
w36240 <= not w35786 and w36239;
w36241 <= not w35790 and not w36240;
w36242 <= not w35957 and w36241;
w36243 <= not w35785 and not w35956;
w36244 <= not w35955 and w36243;
w36245 <= not w36242 and not w36244;
w36246 <= not b(2) and not w36245;
w36247 <= b(0) and not w35957;
w36248 <= a(31) and not w36247;
w36249 <= w7630 and not w35957;
w36250 <= not w36248 and not w36249;
w36251 <= b(1) and not w36250;
w36252 <= not b(1) and not w36249;
w36253 <= not w36248 and w36252;
w36254 <= not w36251 and not w36253;
w36255 <= not w8096 and not w36254;
w36256 <= not b(1) and not w36250;
w36257 <= not w36255 and not w36256;
w36258 <= b(2) and not w36244;
w36259 <= not w36242 and w36258;
w36260 <= not w36246 and not w36259;
w36261 <= not w36257 and w36260;
w36262 <= not w36246 and not w36261;
w36263 <= b(3) and not w36236;
w36264 <= not w36234 and w36263;
w36265 <= not w36238 and not w36264;
w36266 <= not w36262 and w36265;
w36267 <= not w36238 and not w36266;
w36268 <= b(4) and not w36227;
w36269 <= not w36225 and w36268;
w36270 <= not w36229 and not w36269;
w36271 <= not w36267 and w36270;
w36272 <= not w36229 and not w36271;
w36273 <= b(5) and not w36218;
w36274 <= not w36216 and w36273;
w36275 <= not w36220 and not w36274;
w36276 <= not w36272 and w36275;
w36277 <= not w36220 and not w36276;
w36278 <= b(6) and not w36209;
w36279 <= not w36207 and w36278;
w36280 <= not w36211 and not w36279;
w36281 <= not w36277 and w36280;
w36282 <= not w36211 and not w36281;
w36283 <= b(7) and not w36200;
w36284 <= not w36198 and w36283;
w36285 <= not w36202 and not w36284;
w36286 <= not w36282 and w36285;
w36287 <= not w36202 and not w36286;
w36288 <= b(8) and not w36191;
w36289 <= not w36189 and w36288;
w36290 <= not w36193 and not w36289;
w36291 <= not w36287 and w36290;
w36292 <= not w36193 and not w36291;
w36293 <= b(9) and not w36182;
w36294 <= not w36180 and w36293;
w36295 <= not w36184 and not w36294;
w36296 <= not w36292 and w36295;
w36297 <= not w36184 and not w36296;
w36298 <= b(10) and not w36173;
w36299 <= not w36171 and w36298;
w36300 <= not w36175 and not w36299;
w36301 <= not w36297 and w36300;
w36302 <= not w36175 and not w36301;
w36303 <= b(11) and not w36164;
w36304 <= not w36162 and w36303;
w36305 <= not w36166 and not w36304;
w36306 <= not w36302 and w36305;
w36307 <= not w36166 and not w36306;
w36308 <= b(12) and not w36155;
w36309 <= not w36153 and w36308;
w36310 <= not w36157 and not w36309;
w36311 <= not w36307 and w36310;
w36312 <= not w36157 and not w36311;
w36313 <= b(13) and not w36146;
w36314 <= not w36144 and w36313;
w36315 <= not w36148 and not w36314;
w36316 <= not w36312 and w36315;
w36317 <= not w36148 and not w36316;
w36318 <= b(14) and not w36137;
w36319 <= not w36135 and w36318;
w36320 <= not w36139 and not w36319;
w36321 <= not w36317 and w36320;
w36322 <= not w36139 and not w36321;
w36323 <= b(15) and not w36128;
w36324 <= not w36126 and w36323;
w36325 <= not w36130 and not w36324;
w36326 <= not w36322 and w36325;
w36327 <= not w36130 and not w36326;
w36328 <= b(16) and not w36119;
w36329 <= not w36117 and w36328;
w36330 <= not w36121 and not w36329;
w36331 <= not w36327 and w36330;
w36332 <= not w36121 and not w36331;
w36333 <= b(17) and not w36110;
w36334 <= not w36108 and w36333;
w36335 <= not w36112 and not w36334;
w36336 <= not w36332 and w36335;
w36337 <= not w36112 and not w36336;
w36338 <= b(18) and not w36101;
w36339 <= not w36099 and w36338;
w36340 <= not w36103 and not w36339;
w36341 <= not w36337 and w36340;
w36342 <= not w36103 and not w36341;
w36343 <= b(19) and not w36092;
w36344 <= not w36090 and w36343;
w36345 <= not w36094 and not w36344;
w36346 <= not w36342 and w36345;
w36347 <= not w36094 and not w36346;
w36348 <= b(20) and not w36083;
w36349 <= not w36081 and w36348;
w36350 <= not w36085 and not w36349;
w36351 <= not w36347 and w36350;
w36352 <= not w36085 and not w36351;
w36353 <= b(21) and not w36074;
w36354 <= not w36072 and w36353;
w36355 <= not w36076 and not w36354;
w36356 <= not w36352 and w36355;
w36357 <= not w36076 and not w36356;
w36358 <= b(22) and not w36065;
w36359 <= not w36063 and w36358;
w36360 <= not w36067 and not w36359;
w36361 <= not w36357 and w36360;
w36362 <= not w36067 and not w36361;
w36363 <= b(23) and not w36056;
w36364 <= not w36054 and w36363;
w36365 <= not w36058 and not w36364;
w36366 <= not w36362 and w36365;
w36367 <= not w36058 and not w36366;
w36368 <= b(24) and not w36047;
w36369 <= not w36045 and w36368;
w36370 <= not w36049 and not w36369;
w36371 <= not w36367 and w36370;
w36372 <= not w36049 and not w36371;
w36373 <= b(25) and not w36038;
w36374 <= not w36036 and w36373;
w36375 <= not w36040 and not w36374;
w36376 <= not w36372 and w36375;
w36377 <= not w36040 and not w36376;
w36378 <= b(26) and not w36029;
w36379 <= not w36027 and w36378;
w36380 <= not w36031 and not w36379;
w36381 <= not w36377 and w36380;
w36382 <= not w36031 and not w36381;
w36383 <= b(27) and not w36020;
w36384 <= not w36018 and w36383;
w36385 <= not w36022 and not w36384;
w36386 <= not w36382 and w36385;
w36387 <= not w36022 and not w36386;
w36388 <= b(28) and not w36011;
w36389 <= not w36009 and w36388;
w36390 <= not w36013 and not w36389;
w36391 <= not w36387 and w36390;
w36392 <= not w36013 and not w36391;
w36393 <= b(29) and not w36002;
w36394 <= not w36000 and w36393;
w36395 <= not w36004 and not w36394;
w36396 <= not w36392 and w36395;
w36397 <= not w36004 and not w36396;
w36398 <= b(30) and not w35993;
w36399 <= not w35991 and w36398;
w36400 <= not w35995 and not w36399;
w36401 <= not w36397 and w36400;
w36402 <= not w35995 and not w36401;
w36403 <= b(31) and not w35984;
w36404 <= not w35982 and w36403;
w36405 <= not w35986 and not w36404;
w36406 <= not w36402 and w36405;
w36407 <= not w35986 and not w36406;
w36408 <= b(32) and not w35964;
w36409 <= not w35962 and w36408;
w36410 <= not w35977 and not w36409;
w36411 <= not w36407 and w36410;
w36412 <= not w35977 and not w36411;
w36413 <= b(33) and not w35974;
w36414 <= not w35972 and w36413;
w36415 <= not w35976 and not w36414;
w36416 <= not w36412 and w36415;
w36417 <= not w35976 and not w36416;
w36418 <= w8262 and not w36417;
w36419 <= not w35965 and not w36418;
w36420 <= not w35986 and w36410;
w36421 <= not w36406 and w36420;
w36422 <= not w36407 and not w36410;
w36423 <= not w36421 and not w36422;
w36424 <= w8262 and not w36423;
w36425 <= not w36417 and w36424;
w36426 <= not w36419 and not w36425;
w36427 <= not w35975 and not w36418;
w36428 <= not w35977 and w36415;
w36429 <= not w36411 and w36428;
w36430 <= not w36412 and not w36415;
w36431 <= not w36429 and not w36430;
w36432 <= w36418 and not w36431;
w36433 <= not w36427 and not w36432;
w36434 <= not b(34) and not w36433;
w36435 <= not b(33) and not w36426;
w36436 <= not w35985 and not w36418;
w36437 <= not w35995 and w36405;
w36438 <= not w36401 and w36437;
w36439 <= not w36402 and not w36405;
w36440 <= not w36438 and not w36439;
w36441 <= w8262 and not w36440;
w36442 <= not w36417 and w36441;
w36443 <= not w36436 and not w36442;
w36444 <= not b(32) and not w36443;
w36445 <= not w35994 and not w36418;
w36446 <= not w36004 and w36400;
w36447 <= not w36396 and w36446;
w36448 <= not w36397 and not w36400;
w36449 <= not w36447 and not w36448;
w36450 <= w8262 and not w36449;
w36451 <= not w36417 and w36450;
w36452 <= not w36445 and not w36451;
w36453 <= not b(31) and not w36452;
w36454 <= not w36003 and not w36418;
w36455 <= not w36013 and w36395;
w36456 <= not w36391 and w36455;
w36457 <= not w36392 and not w36395;
w36458 <= not w36456 and not w36457;
w36459 <= w8262 and not w36458;
w36460 <= not w36417 and w36459;
w36461 <= not w36454 and not w36460;
w36462 <= not b(30) and not w36461;
w36463 <= not w36012 and not w36418;
w36464 <= not w36022 and w36390;
w36465 <= not w36386 and w36464;
w36466 <= not w36387 and not w36390;
w36467 <= not w36465 and not w36466;
w36468 <= w8262 and not w36467;
w36469 <= not w36417 and w36468;
w36470 <= not w36463 and not w36469;
w36471 <= not b(29) and not w36470;
w36472 <= not w36021 and not w36418;
w36473 <= not w36031 and w36385;
w36474 <= not w36381 and w36473;
w36475 <= not w36382 and not w36385;
w36476 <= not w36474 and not w36475;
w36477 <= w8262 and not w36476;
w36478 <= not w36417 and w36477;
w36479 <= not w36472 and not w36478;
w36480 <= not b(28) and not w36479;
w36481 <= not w36030 and not w36418;
w36482 <= not w36040 and w36380;
w36483 <= not w36376 and w36482;
w36484 <= not w36377 and not w36380;
w36485 <= not w36483 and not w36484;
w36486 <= w8262 and not w36485;
w36487 <= not w36417 and w36486;
w36488 <= not w36481 and not w36487;
w36489 <= not b(27) and not w36488;
w36490 <= not w36039 and not w36418;
w36491 <= not w36049 and w36375;
w36492 <= not w36371 and w36491;
w36493 <= not w36372 and not w36375;
w36494 <= not w36492 and not w36493;
w36495 <= w8262 and not w36494;
w36496 <= not w36417 and w36495;
w36497 <= not w36490 and not w36496;
w36498 <= not b(26) and not w36497;
w36499 <= not w36048 and not w36418;
w36500 <= not w36058 and w36370;
w36501 <= not w36366 and w36500;
w36502 <= not w36367 and not w36370;
w36503 <= not w36501 and not w36502;
w36504 <= w8262 and not w36503;
w36505 <= not w36417 and w36504;
w36506 <= not w36499 and not w36505;
w36507 <= not b(25) and not w36506;
w36508 <= not w36057 and not w36418;
w36509 <= not w36067 and w36365;
w36510 <= not w36361 and w36509;
w36511 <= not w36362 and not w36365;
w36512 <= not w36510 and not w36511;
w36513 <= w8262 and not w36512;
w36514 <= not w36417 and w36513;
w36515 <= not w36508 and not w36514;
w36516 <= not b(24) and not w36515;
w36517 <= not w36066 and not w36418;
w36518 <= not w36076 and w36360;
w36519 <= not w36356 and w36518;
w36520 <= not w36357 and not w36360;
w36521 <= not w36519 and not w36520;
w36522 <= w8262 and not w36521;
w36523 <= not w36417 and w36522;
w36524 <= not w36517 and not w36523;
w36525 <= not b(23) and not w36524;
w36526 <= not w36075 and not w36418;
w36527 <= not w36085 and w36355;
w36528 <= not w36351 and w36527;
w36529 <= not w36352 and not w36355;
w36530 <= not w36528 and not w36529;
w36531 <= w8262 and not w36530;
w36532 <= not w36417 and w36531;
w36533 <= not w36526 and not w36532;
w36534 <= not b(22) and not w36533;
w36535 <= not w36084 and not w36418;
w36536 <= not w36094 and w36350;
w36537 <= not w36346 and w36536;
w36538 <= not w36347 and not w36350;
w36539 <= not w36537 and not w36538;
w36540 <= w8262 and not w36539;
w36541 <= not w36417 and w36540;
w36542 <= not w36535 and not w36541;
w36543 <= not b(21) and not w36542;
w36544 <= not w36093 and not w36418;
w36545 <= not w36103 and w36345;
w36546 <= not w36341 and w36545;
w36547 <= not w36342 and not w36345;
w36548 <= not w36546 and not w36547;
w36549 <= w8262 and not w36548;
w36550 <= not w36417 and w36549;
w36551 <= not w36544 and not w36550;
w36552 <= not b(20) and not w36551;
w36553 <= not w36102 and not w36418;
w36554 <= not w36112 and w36340;
w36555 <= not w36336 and w36554;
w36556 <= not w36337 and not w36340;
w36557 <= not w36555 and not w36556;
w36558 <= w8262 and not w36557;
w36559 <= not w36417 and w36558;
w36560 <= not w36553 and not w36559;
w36561 <= not b(19) and not w36560;
w36562 <= not w36111 and not w36418;
w36563 <= not w36121 and w36335;
w36564 <= not w36331 and w36563;
w36565 <= not w36332 and not w36335;
w36566 <= not w36564 and not w36565;
w36567 <= w8262 and not w36566;
w36568 <= not w36417 and w36567;
w36569 <= not w36562 and not w36568;
w36570 <= not b(18) and not w36569;
w36571 <= not w36120 and not w36418;
w36572 <= not w36130 and w36330;
w36573 <= not w36326 and w36572;
w36574 <= not w36327 and not w36330;
w36575 <= not w36573 and not w36574;
w36576 <= w8262 and not w36575;
w36577 <= not w36417 and w36576;
w36578 <= not w36571 and not w36577;
w36579 <= not b(17) and not w36578;
w36580 <= not w36129 and not w36418;
w36581 <= not w36139 and w36325;
w36582 <= not w36321 and w36581;
w36583 <= not w36322 and not w36325;
w36584 <= not w36582 and not w36583;
w36585 <= w8262 and not w36584;
w36586 <= not w36417 and w36585;
w36587 <= not w36580 and not w36586;
w36588 <= not b(16) and not w36587;
w36589 <= not w36138 and not w36418;
w36590 <= not w36148 and w36320;
w36591 <= not w36316 and w36590;
w36592 <= not w36317 and not w36320;
w36593 <= not w36591 and not w36592;
w36594 <= w8262 and not w36593;
w36595 <= not w36417 and w36594;
w36596 <= not w36589 and not w36595;
w36597 <= not b(15) and not w36596;
w36598 <= not w36147 and not w36418;
w36599 <= not w36157 and w36315;
w36600 <= not w36311 and w36599;
w36601 <= not w36312 and not w36315;
w36602 <= not w36600 and not w36601;
w36603 <= w8262 and not w36602;
w36604 <= not w36417 and w36603;
w36605 <= not w36598 and not w36604;
w36606 <= not b(14) and not w36605;
w36607 <= not w36156 and not w36418;
w36608 <= not w36166 and w36310;
w36609 <= not w36306 and w36608;
w36610 <= not w36307 and not w36310;
w36611 <= not w36609 and not w36610;
w36612 <= w8262 and not w36611;
w36613 <= not w36417 and w36612;
w36614 <= not w36607 and not w36613;
w36615 <= not b(13) and not w36614;
w36616 <= not w36165 and not w36418;
w36617 <= not w36175 and w36305;
w36618 <= not w36301 and w36617;
w36619 <= not w36302 and not w36305;
w36620 <= not w36618 and not w36619;
w36621 <= w8262 and not w36620;
w36622 <= not w36417 and w36621;
w36623 <= not w36616 and not w36622;
w36624 <= not b(12) and not w36623;
w36625 <= not w36174 and not w36418;
w36626 <= not w36184 and w36300;
w36627 <= not w36296 and w36626;
w36628 <= not w36297 and not w36300;
w36629 <= not w36627 and not w36628;
w36630 <= w8262 and not w36629;
w36631 <= not w36417 and w36630;
w36632 <= not w36625 and not w36631;
w36633 <= not b(11) and not w36632;
w36634 <= not w36183 and not w36418;
w36635 <= not w36193 and w36295;
w36636 <= not w36291 and w36635;
w36637 <= not w36292 and not w36295;
w36638 <= not w36636 and not w36637;
w36639 <= w8262 and not w36638;
w36640 <= not w36417 and w36639;
w36641 <= not w36634 and not w36640;
w36642 <= not b(10) and not w36641;
w36643 <= not w36192 and not w36418;
w36644 <= not w36202 and w36290;
w36645 <= not w36286 and w36644;
w36646 <= not w36287 and not w36290;
w36647 <= not w36645 and not w36646;
w36648 <= w8262 and not w36647;
w36649 <= not w36417 and w36648;
w36650 <= not w36643 and not w36649;
w36651 <= not b(9) and not w36650;
w36652 <= not w36201 and not w36418;
w36653 <= not w36211 and w36285;
w36654 <= not w36281 and w36653;
w36655 <= not w36282 and not w36285;
w36656 <= not w36654 and not w36655;
w36657 <= w8262 and not w36656;
w36658 <= not w36417 and w36657;
w36659 <= not w36652 and not w36658;
w36660 <= not b(8) and not w36659;
w36661 <= not w36210 and not w36418;
w36662 <= not w36220 and w36280;
w36663 <= not w36276 and w36662;
w36664 <= not w36277 and not w36280;
w36665 <= not w36663 and not w36664;
w36666 <= w8262 and not w36665;
w36667 <= not w36417 and w36666;
w36668 <= not w36661 and not w36667;
w36669 <= not b(7) and not w36668;
w36670 <= not w36219 and not w36418;
w36671 <= not w36229 and w36275;
w36672 <= not w36271 and w36671;
w36673 <= not w36272 and not w36275;
w36674 <= not w36672 and not w36673;
w36675 <= w8262 and not w36674;
w36676 <= not w36417 and w36675;
w36677 <= not w36670 and not w36676;
w36678 <= not b(6) and not w36677;
w36679 <= not w36228 and not w36418;
w36680 <= not w36238 and w36270;
w36681 <= not w36266 and w36680;
w36682 <= not w36267 and not w36270;
w36683 <= not w36681 and not w36682;
w36684 <= w8262 and not w36683;
w36685 <= not w36417 and w36684;
w36686 <= not w36679 and not w36685;
w36687 <= not b(5) and not w36686;
w36688 <= not w36237 and not w36418;
w36689 <= not w36246 and w36265;
w36690 <= not w36261 and w36689;
w36691 <= not w36262 and not w36265;
w36692 <= not w36690 and not w36691;
w36693 <= w8262 and not w36692;
w36694 <= not w36417 and w36693;
w36695 <= not w36688 and not w36694;
w36696 <= not b(4) and not w36695;
w36697 <= not w36245 and not w36418;
w36698 <= not w36256 and w36260;
w36699 <= not w36255 and w36698;
w36700 <= not w36257 and not w36260;
w36701 <= not w36699 and not w36700;
w36702 <= w8262 and not w36701;
w36703 <= not w36417 and w36702;
w36704 <= not w36697 and not w36703;
w36705 <= not b(3) and not w36704;
w36706 <= not w36250 and not w36418;
w36707 <= w8096 and not w36253;
w36708 <= not w36251 and w36707;
w36709 <= w8262 and not w36708;
w36710 <= not w36255 and w36709;
w36711 <= not w36417 and w36710;
w36712 <= not w36706 and not w36711;
w36713 <= not b(2) and not w36712;
w36714 <= w8563 and not w36417;
w36715 <= a(30) and not w36714;
w36716 <= w8569 and not w36417;
w36717 <= not w36715 and not w36716;
w36718 <= b(1) and not w36717;
w36719 <= not b(1) and not w36716;
w36720 <= not w36715 and w36719;
w36721 <= not w36718 and not w36720;
w36722 <= not w8576 and not w36721;
w36723 <= not b(1) and not w36717;
w36724 <= not w36722 and not w36723;
w36725 <= b(2) and not w36711;
w36726 <= not w36706 and w36725;
w36727 <= not w36713 and not w36726;
w36728 <= not w36724 and w36727;
w36729 <= not w36713 and not w36728;
w36730 <= b(3) and not w36703;
w36731 <= not w36697 and w36730;
w36732 <= not w36705 and not w36731;
w36733 <= not w36729 and w36732;
w36734 <= not w36705 and not w36733;
w36735 <= b(4) and not w36694;
w36736 <= not w36688 and w36735;
w36737 <= not w36696 and not w36736;
w36738 <= not w36734 and w36737;
w36739 <= not w36696 and not w36738;
w36740 <= b(5) and not w36685;
w36741 <= not w36679 and w36740;
w36742 <= not w36687 and not w36741;
w36743 <= not w36739 and w36742;
w36744 <= not w36687 and not w36743;
w36745 <= b(6) and not w36676;
w36746 <= not w36670 and w36745;
w36747 <= not w36678 and not w36746;
w36748 <= not w36744 and w36747;
w36749 <= not w36678 and not w36748;
w36750 <= b(7) and not w36667;
w36751 <= not w36661 and w36750;
w36752 <= not w36669 and not w36751;
w36753 <= not w36749 and w36752;
w36754 <= not w36669 and not w36753;
w36755 <= b(8) and not w36658;
w36756 <= not w36652 and w36755;
w36757 <= not w36660 and not w36756;
w36758 <= not w36754 and w36757;
w36759 <= not w36660 and not w36758;
w36760 <= b(9) and not w36649;
w36761 <= not w36643 and w36760;
w36762 <= not w36651 and not w36761;
w36763 <= not w36759 and w36762;
w36764 <= not w36651 and not w36763;
w36765 <= b(10) and not w36640;
w36766 <= not w36634 and w36765;
w36767 <= not w36642 and not w36766;
w36768 <= not w36764 and w36767;
w36769 <= not w36642 and not w36768;
w36770 <= b(11) and not w36631;
w36771 <= not w36625 and w36770;
w36772 <= not w36633 and not w36771;
w36773 <= not w36769 and w36772;
w36774 <= not w36633 and not w36773;
w36775 <= b(12) and not w36622;
w36776 <= not w36616 and w36775;
w36777 <= not w36624 and not w36776;
w36778 <= not w36774 and w36777;
w36779 <= not w36624 and not w36778;
w36780 <= b(13) and not w36613;
w36781 <= not w36607 and w36780;
w36782 <= not w36615 and not w36781;
w36783 <= not w36779 and w36782;
w36784 <= not w36615 and not w36783;
w36785 <= b(14) and not w36604;
w36786 <= not w36598 and w36785;
w36787 <= not w36606 and not w36786;
w36788 <= not w36784 and w36787;
w36789 <= not w36606 and not w36788;
w36790 <= b(15) and not w36595;
w36791 <= not w36589 and w36790;
w36792 <= not w36597 and not w36791;
w36793 <= not w36789 and w36792;
w36794 <= not w36597 and not w36793;
w36795 <= b(16) and not w36586;
w36796 <= not w36580 and w36795;
w36797 <= not w36588 and not w36796;
w36798 <= not w36794 and w36797;
w36799 <= not w36588 and not w36798;
w36800 <= b(17) and not w36577;
w36801 <= not w36571 and w36800;
w36802 <= not w36579 and not w36801;
w36803 <= not w36799 and w36802;
w36804 <= not w36579 and not w36803;
w36805 <= b(18) and not w36568;
w36806 <= not w36562 and w36805;
w36807 <= not w36570 and not w36806;
w36808 <= not w36804 and w36807;
w36809 <= not w36570 and not w36808;
w36810 <= b(19) and not w36559;
w36811 <= not w36553 and w36810;
w36812 <= not w36561 and not w36811;
w36813 <= not w36809 and w36812;
w36814 <= not w36561 and not w36813;
w36815 <= b(20) and not w36550;
w36816 <= not w36544 and w36815;
w36817 <= not w36552 and not w36816;
w36818 <= not w36814 and w36817;
w36819 <= not w36552 and not w36818;
w36820 <= b(21) and not w36541;
w36821 <= not w36535 and w36820;
w36822 <= not w36543 and not w36821;
w36823 <= not w36819 and w36822;
w36824 <= not w36543 and not w36823;
w36825 <= b(22) and not w36532;
w36826 <= not w36526 and w36825;
w36827 <= not w36534 and not w36826;
w36828 <= not w36824 and w36827;
w36829 <= not w36534 and not w36828;
w36830 <= b(23) and not w36523;
w36831 <= not w36517 and w36830;
w36832 <= not w36525 and not w36831;
w36833 <= not w36829 and w36832;
w36834 <= not w36525 and not w36833;
w36835 <= b(24) and not w36514;
w36836 <= not w36508 and w36835;
w36837 <= not w36516 and not w36836;
w36838 <= not w36834 and w36837;
w36839 <= not w36516 and not w36838;
w36840 <= b(25) and not w36505;
w36841 <= not w36499 and w36840;
w36842 <= not w36507 and not w36841;
w36843 <= not w36839 and w36842;
w36844 <= not w36507 and not w36843;
w36845 <= b(26) and not w36496;
w36846 <= not w36490 and w36845;
w36847 <= not w36498 and not w36846;
w36848 <= not w36844 and w36847;
w36849 <= not w36498 and not w36848;
w36850 <= b(27) and not w36487;
w36851 <= not w36481 and w36850;
w36852 <= not w36489 and not w36851;
w36853 <= not w36849 and w36852;
w36854 <= not w36489 and not w36853;
w36855 <= b(28) and not w36478;
w36856 <= not w36472 and w36855;
w36857 <= not w36480 and not w36856;
w36858 <= not w36854 and w36857;
w36859 <= not w36480 and not w36858;
w36860 <= b(29) and not w36469;
w36861 <= not w36463 and w36860;
w36862 <= not w36471 and not w36861;
w36863 <= not w36859 and w36862;
w36864 <= not w36471 and not w36863;
w36865 <= b(30) and not w36460;
w36866 <= not w36454 and w36865;
w36867 <= not w36462 and not w36866;
w36868 <= not w36864 and w36867;
w36869 <= not w36462 and not w36868;
w36870 <= b(31) and not w36451;
w36871 <= not w36445 and w36870;
w36872 <= not w36453 and not w36871;
w36873 <= not w36869 and w36872;
w36874 <= not w36453 and not w36873;
w36875 <= b(32) and not w36442;
w36876 <= not w36436 and w36875;
w36877 <= not w36444 and not w36876;
w36878 <= not w36874 and w36877;
w36879 <= not w36444 and not w36878;
w36880 <= b(33) and not w36425;
w36881 <= not w36419 and w36880;
w36882 <= not w36435 and not w36881;
w36883 <= not w36879 and w36882;
w36884 <= not w36435 and not w36883;
w36885 <= b(34) and not w36427;
w36886 <= not w36432 and w36885;
w36887 <= not w36434 and not w36886;
w36888 <= not w36884 and w36887;
w36889 <= not w36434 and not w36888;
w36890 <= w8747 and not w36889;
w36891 <= not w36426 and not w36890;
w36892 <= not w36444 and w36882;
w36893 <= not w36878 and w36892;
w36894 <= not w36879 and not w36882;
w36895 <= not w36893 and not w36894;
w36896 <= w8747 and not w36895;
w36897 <= not w36889 and w36896;
w36898 <= not w36891 and not w36897;
w36899 <= not b(34) and not w36898;
w36900 <= not w36443 and not w36890;
w36901 <= not w36453 and w36877;
w36902 <= not w36873 and w36901;
w36903 <= not w36874 and not w36877;
w36904 <= not w36902 and not w36903;
w36905 <= w8747 and not w36904;
w36906 <= not w36889 and w36905;
w36907 <= not w36900 and not w36906;
w36908 <= not b(33) and not w36907;
w36909 <= not w36452 and not w36890;
w36910 <= not w36462 and w36872;
w36911 <= not w36868 and w36910;
w36912 <= not w36869 and not w36872;
w36913 <= not w36911 and not w36912;
w36914 <= w8747 and not w36913;
w36915 <= not w36889 and w36914;
w36916 <= not w36909 and not w36915;
w36917 <= not b(32) and not w36916;
w36918 <= not w36461 and not w36890;
w36919 <= not w36471 and w36867;
w36920 <= not w36863 and w36919;
w36921 <= not w36864 and not w36867;
w36922 <= not w36920 and not w36921;
w36923 <= w8747 and not w36922;
w36924 <= not w36889 and w36923;
w36925 <= not w36918 and not w36924;
w36926 <= not b(31) and not w36925;
w36927 <= not w36470 and not w36890;
w36928 <= not w36480 and w36862;
w36929 <= not w36858 and w36928;
w36930 <= not w36859 and not w36862;
w36931 <= not w36929 and not w36930;
w36932 <= w8747 and not w36931;
w36933 <= not w36889 and w36932;
w36934 <= not w36927 and not w36933;
w36935 <= not b(30) and not w36934;
w36936 <= not w36479 and not w36890;
w36937 <= not w36489 and w36857;
w36938 <= not w36853 and w36937;
w36939 <= not w36854 and not w36857;
w36940 <= not w36938 and not w36939;
w36941 <= w8747 and not w36940;
w36942 <= not w36889 and w36941;
w36943 <= not w36936 and not w36942;
w36944 <= not b(29) and not w36943;
w36945 <= not w36488 and not w36890;
w36946 <= not w36498 and w36852;
w36947 <= not w36848 and w36946;
w36948 <= not w36849 and not w36852;
w36949 <= not w36947 and not w36948;
w36950 <= w8747 and not w36949;
w36951 <= not w36889 and w36950;
w36952 <= not w36945 and not w36951;
w36953 <= not b(28) and not w36952;
w36954 <= not w36497 and not w36890;
w36955 <= not w36507 and w36847;
w36956 <= not w36843 and w36955;
w36957 <= not w36844 and not w36847;
w36958 <= not w36956 and not w36957;
w36959 <= w8747 and not w36958;
w36960 <= not w36889 and w36959;
w36961 <= not w36954 and not w36960;
w36962 <= not b(27) and not w36961;
w36963 <= not w36506 and not w36890;
w36964 <= not w36516 and w36842;
w36965 <= not w36838 and w36964;
w36966 <= not w36839 and not w36842;
w36967 <= not w36965 and not w36966;
w36968 <= w8747 and not w36967;
w36969 <= not w36889 and w36968;
w36970 <= not w36963 and not w36969;
w36971 <= not b(26) and not w36970;
w36972 <= not w36515 and not w36890;
w36973 <= not w36525 and w36837;
w36974 <= not w36833 and w36973;
w36975 <= not w36834 and not w36837;
w36976 <= not w36974 and not w36975;
w36977 <= w8747 and not w36976;
w36978 <= not w36889 and w36977;
w36979 <= not w36972 and not w36978;
w36980 <= not b(25) and not w36979;
w36981 <= not w36524 and not w36890;
w36982 <= not w36534 and w36832;
w36983 <= not w36828 and w36982;
w36984 <= not w36829 and not w36832;
w36985 <= not w36983 and not w36984;
w36986 <= w8747 and not w36985;
w36987 <= not w36889 and w36986;
w36988 <= not w36981 and not w36987;
w36989 <= not b(24) and not w36988;
w36990 <= not w36533 and not w36890;
w36991 <= not w36543 and w36827;
w36992 <= not w36823 and w36991;
w36993 <= not w36824 and not w36827;
w36994 <= not w36992 and not w36993;
w36995 <= w8747 and not w36994;
w36996 <= not w36889 and w36995;
w36997 <= not w36990 and not w36996;
w36998 <= not b(23) and not w36997;
w36999 <= not w36542 and not w36890;
w37000 <= not w36552 and w36822;
w37001 <= not w36818 and w37000;
w37002 <= not w36819 and not w36822;
w37003 <= not w37001 and not w37002;
w37004 <= w8747 and not w37003;
w37005 <= not w36889 and w37004;
w37006 <= not w36999 and not w37005;
w37007 <= not b(22) and not w37006;
w37008 <= not w36551 and not w36890;
w37009 <= not w36561 and w36817;
w37010 <= not w36813 and w37009;
w37011 <= not w36814 and not w36817;
w37012 <= not w37010 and not w37011;
w37013 <= w8747 and not w37012;
w37014 <= not w36889 and w37013;
w37015 <= not w37008 and not w37014;
w37016 <= not b(21) and not w37015;
w37017 <= not w36560 and not w36890;
w37018 <= not w36570 and w36812;
w37019 <= not w36808 and w37018;
w37020 <= not w36809 and not w36812;
w37021 <= not w37019 and not w37020;
w37022 <= w8747 and not w37021;
w37023 <= not w36889 and w37022;
w37024 <= not w37017 and not w37023;
w37025 <= not b(20) and not w37024;
w37026 <= not w36569 and not w36890;
w37027 <= not w36579 and w36807;
w37028 <= not w36803 and w37027;
w37029 <= not w36804 and not w36807;
w37030 <= not w37028 and not w37029;
w37031 <= w8747 and not w37030;
w37032 <= not w36889 and w37031;
w37033 <= not w37026 and not w37032;
w37034 <= not b(19) and not w37033;
w37035 <= not w36578 and not w36890;
w37036 <= not w36588 and w36802;
w37037 <= not w36798 and w37036;
w37038 <= not w36799 and not w36802;
w37039 <= not w37037 and not w37038;
w37040 <= w8747 and not w37039;
w37041 <= not w36889 and w37040;
w37042 <= not w37035 and not w37041;
w37043 <= not b(18) and not w37042;
w37044 <= not w36587 and not w36890;
w37045 <= not w36597 and w36797;
w37046 <= not w36793 and w37045;
w37047 <= not w36794 and not w36797;
w37048 <= not w37046 and not w37047;
w37049 <= w8747 and not w37048;
w37050 <= not w36889 and w37049;
w37051 <= not w37044 and not w37050;
w37052 <= not b(17) and not w37051;
w37053 <= not w36596 and not w36890;
w37054 <= not w36606 and w36792;
w37055 <= not w36788 and w37054;
w37056 <= not w36789 and not w36792;
w37057 <= not w37055 and not w37056;
w37058 <= w8747 and not w37057;
w37059 <= not w36889 and w37058;
w37060 <= not w37053 and not w37059;
w37061 <= not b(16) and not w37060;
w37062 <= not w36605 and not w36890;
w37063 <= not w36615 and w36787;
w37064 <= not w36783 and w37063;
w37065 <= not w36784 and not w36787;
w37066 <= not w37064 and not w37065;
w37067 <= w8747 and not w37066;
w37068 <= not w36889 and w37067;
w37069 <= not w37062 and not w37068;
w37070 <= not b(15) and not w37069;
w37071 <= not w36614 and not w36890;
w37072 <= not w36624 and w36782;
w37073 <= not w36778 and w37072;
w37074 <= not w36779 and not w36782;
w37075 <= not w37073 and not w37074;
w37076 <= w8747 and not w37075;
w37077 <= not w36889 and w37076;
w37078 <= not w37071 and not w37077;
w37079 <= not b(14) and not w37078;
w37080 <= not w36623 and not w36890;
w37081 <= not w36633 and w36777;
w37082 <= not w36773 and w37081;
w37083 <= not w36774 and not w36777;
w37084 <= not w37082 and not w37083;
w37085 <= w8747 and not w37084;
w37086 <= not w36889 and w37085;
w37087 <= not w37080 and not w37086;
w37088 <= not b(13) and not w37087;
w37089 <= not w36632 and not w36890;
w37090 <= not w36642 and w36772;
w37091 <= not w36768 and w37090;
w37092 <= not w36769 and not w36772;
w37093 <= not w37091 and not w37092;
w37094 <= w8747 and not w37093;
w37095 <= not w36889 and w37094;
w37096 <= not w37089 and not w37095;
w37097 <= not b(12) and not w37096;
w37098 <= not w36641 and not w36890;
w37099 <= not w36651 and w36767;
w37100 <= not w36763 and w37099;
w37101 <= not w36764 and not w36767;
w37102 <= not w37100 and not w37101;
w37103 <= w8747 and not w37102;
w37104 <= not w36889 and w37103;
w37105 <= not w37098 and not w37104;
w37106 <= not b(11) and not w37105;
w37107 <= not w36650 and not w36890;
w37108 <= not w36660 and w36762;
w37109 <= not w36758 and w37108;
w37110 <= not w36759 and not w36762;
w37111 <= not w37109 and not w37110;
w37112 <= w8747 and not w37111;
w37113 <= not w36889 and w37112;
w37114 <= not w37107 and not w37113;
w37115 <= not b(10) and not w37114;
w37116 <= not w36659 and not w36890;
w37117 <= not w36669 and w36757;
w37118 <= not w36753 and w37117;
w37119 <= not w36754 and not w36757;
w37120 <= not w37118 and not w37119;
w37121 <= w8747 and not w37120;
w37122 <= not w36889 and w37121;
w37123 <= not w37116 and not w37122;
w37124 <= not b(9) and not w37123;
w37125 <= not w36668 and not w36890;
w37126 <= not w36678 and w36752;
w37127 <= not w36748 and w37126;
w37128 <= not w36749 and not w36752;
w37129 <= not w37127 and not w37128;
w37130 <= w8747 and not w37129;
w37131 <= not w36889 and w37130;
w37132 <= not w37125 and not w37131;
w37133 <= not b(8) and not w37132;
w37134 <= not w36677 and not w36890;
w37135 <= not w36687 and w36747;
w37136 <= not w36743 and w37135;
w37137 <= not w36744 and not w36747;
w37138 <= not w37136 and not w37137;
w37139 <= w8747 and not w37138;
w37140 <= not w36889 and w37139;
w37141 <= not w37134 and not w37140;
w37142 <= not b(7) and not w37141;
w37143 <= not w36686 and not w36890;
w37144 <= not w36696 and w36742;
w37145 <= not w36738 and w37144;
w37146 <= not w36739 and not w36742;
w37147 <= not w37145 and not w37146;
w37148 <= w8747 and not w37147;
w37149 <= not w36889 and w37148;
w37150 <= not w37143 and not w37149;
w37151 <= not b(6) and not w37150;
w37152 <= not w36695 and not w36890;
w37153 <= not w36705 and w36737;
w37154 <= not w36733 and w37153;
w37155 <= not w36734 and not w36737;
w37156 <= not w37154 and not w37155;
w37157 <= w8747 and not w37156;
w37158 <= not w36889 and w37157;
w37159 <= not w37152 and not w37158;
w37160 <= not b(5) and not w37159;
w37161 <= not w36704 and not w36890;
w37162 <= not w36713 and w36732;
w37163 <= not w36728 and w37162;
w37164 <= not w36729 and not w36732;
w37165 <= not w37163 and not w37164;
w37166 <= w8747 and not w37165;
w37167 <= not w36889 and w37166;
w37168 <= not w37161 and not w37167;
w37169 <= not b(4) and not w37168;
w37170 <= not w36712 and not w36890;
w37171 <= not w36723 and w36727;
w37172 <= not w36722 and w37171;
w37173 <= not w36724 and not w36727;
w37174 <= not w37172 and not w37173;
w37175 <= w8747 and not w37174;
w37176 <= not w36889 and w37175;
w37177 <= not w37170 and not w37176;
w37178 <= not b(3) and not w37177;
w37179 <= not w36717 and not w36890;
w37180 <= w8576 and not w36720;
w37181 <= not w36718 and w37180;
w37182 <= w8747 and not w37181;
w37183 <= not w36722 and w37182;
w37184 <= not w36889 and w37183;
w37185 <= not w37179 and not w37184;
w37186 <= not b(2) and not w37185;
w37187 <= w9048 and not w36889;
w37188 <= a(29) and not w37187;
w37189 <= w9054 and not w36889;
w37190 <= not w37188 and not w37189;
w37191 <= b(1) and not w37190;
w37192 <= not b(1) and not w37189;
w37193 <= not w37188 and w37192;
w37194 <= not w37191 and not w37193;
w37195 <= not w9061 and not w37194;
w37196 <= not b(1) and not w37190;
w37197 <= not w37195 and not w37196;
w37198 <= b(2) and not w37184;
w37199 <= not w37179 and w37198;
w37200 <= not w37186 and not w37199;
w37201 <= not w37197 and w37200;
w37202 <= not w37186 and not w37201;
w37203 <= b(3) and not w37176;
w37204 <= not w37170 and w37203;
w37205 <= not w37178 and not w37204;
w37206 <= not w37202 and w37205;
w37207 <= not w37178 and not w37206;
w37208 <= b(4) and not w37167;
w37209 <= not w37161 and w37208;
w37210 <= not w37169 and not w37209;
w37211 <= not w37207 and w37210;
w37212 <= not w37169 and not w37211;
w37213 <= b(5) and not w37158;
w37214 <= not w37152 and w37213;
w37215 <= not w37160 and not w37214;
w37216 <= not w37212 and w37215;
w37217 <= not w37160 and not w37216;
w37218 <= b(6) and not w37149;
w37219 <= not w37143 and w37218;
w37220 <= not w37151 and not w37219;
w37221 <= not w37217 and w37220;
w37222 <= not w37151 and not w37221;
w37223 <= b(7) and not w37140;
w37224 <= not w37134 and w37223;
w37225 <= not w37142 and not w37224;
w37226 <= not w37222 and w37225;
w37227 <= not w37142 and not w37226;
w37228 <= b(8) and not w37131;
w37229 <= not w37125 and w37228;
w37230 <= not w37133 and not w37229;
w37231 <= not w37227 and w37230;
w37232 <= not w37133 and not w37231;
w37233 <= b(9) and not w37122;
w37234 <= not w37116 and w37233;
w37235 <= not w37124 and not w37234;
w37236 <= not w37232 and w37235;
w37237 <= not w37124 and not w37236;
w37238 <= b(10) and not w37113;
w37239 <= not w37107 and w37238;
w37240 <= not w37115 and not w37239;
w37241 <= not w37237 and w37240;
w37242 <= not w37115 and not w37241;
w37243 <= b(11) and not w37104;
w37244 <= not w37098 and w37243;
w37245 <= not w37106 and not w37244;
w37246 <= not w37242 and w37245;
w37247 <= not w37106 and not w37246;
w37248 <= b(12) and not w37095;
w37249 <= not w37089 and w37248;
w37250 <= not w37097 and not w37249;
w37251 <= not w37247 and w37250;
w37252 <= not w37097 and not w37251;
w37253 <= b(13) and not w37086;
w37254 <= not w37080 and w37253;
w37255 <= not w37088 and not w37254;
w37256 <= not w37252 and w37255;
w37257 <= not w37088 and not w37256;
w37258 <= b(14) and not w37077;
w37259 <= not w37071 and w37258;
w37260 <= not w37079 and not w37259;
w37261 <= not w37257 and w37260;
w37262 <= not w37079 and not w37261;
w37263 <= b(15) and not w37068;
w37264 <= not w37062 and w37263;
w37265 <= not w37070 and not w37264;
w37266 <= not w37262 and w37265;
w37267 <= not w37070 and not w37266;
w37268 <= b(16) and not w37059;
w37269 <= not w37053 and w37268;
w37270 <= not w37061 and not w37269;
w37271 <= not w37267 and w37270;
w37272 <= not w37061 and not w37271;
w37273 <= b(17) and not w37050;
w37274 <= not w37044 and w37273;
w37275 <= not w37052 and not w37274;
w37276 <= not w37272 and w37275;
w37277 <= not w37052 and not w37276;
w37278 <= b(18) and not w37041;
w37279 <= not w37035 and w37278;
w37280 <= not w37043 and not w37279;
w37281 <= not w37277 and w37280;
w37282 <= not w37043 and not w37281;
w37283 <= b(19) and not w37032;
w37284 <= not w37026 and w37283;
w37285 <= not w37034 and not w37284;
w37286 <= not w37282 and w37285;
w37287 <= not w37034 and not w37286;
w37288 <= b(20) and not w37023;
w37289 <= not w37017 and w37288;
w37290 <= not w37025 and not w37289;
w37291 <= not w37287 and w37290;
w37292 <= not w37025 and not w37291;
w37293 <= b(21) and not w37014;
w37294 <= not w37008 and w37293;
w37295 <= not w37016 and not w37294;
w37296 <= not w37292 and w37295;
w37297 <= not w37016 and not w37296;
w37298 <= b(22) and not w37005;
w37299 <= not w36999 and w37298;
w37300 <= not w37007 and not w37299;
w37301 <= not w37297 and w37300;
w37302 <= not w37007 and not w37301;
w37303 <= b(23) and not w36996;
w37304 <= not w36990 and w37303;
w37305 <= not w36998 and not w37304;
w37306 <= not w37302 and w37305;
w37307 <= not w36998 and not w37306;
w37308 <= b(24) and not w36987;
w37309 <= not w36981 and w37308;
w37310 <= not w36989 and not w37309;
w37311 <= not w37307 and w37310;
w37312 <= not w36989 and not w37311;
w37313 <= b(25) and not w36978;
w37314 <= not w36972 and w37313;
w37315 <= not w36980 and not w37314;
w37316 <= not w37312 and w37315;
w37317 <= not w36980 and not w37316;
w37318 <= b(26) and not w36969;
w37319 <= not w36963 and w37318;
w37320 <= not w36971 and not w37319;
w37321 <= not w37317 and w37320;
w37322 <= not w36971 and not w37321;
w37323 <= b(27) and not w36960;
w37324 <= not w36954 and w37323;
w37325 <= not w36962 and not w37324;
w37326 <= not w37322 and w37325;
w37327 <= not w36962 and not w37326;
w37328 <= b(28) and not w36951;
w37329 <= not w36945 and w37328;
w37330 <= not w36953 and not w37329;
w37331 <= not w37327 and w37330;
w37332 <= not w36953 and not w37331;
w37333 <= b(29) and not w36942;
w37334 <= not w36936 and w37333;
w37335 <= not w36944 and not w37334;
w37336 <= not w37332 and w37335;
w37337 <= not w36944 and not w37336;
w37338 <= b(30) and not w36933;
w37339 <= not w36927 and w37338;
w37340 <= not w36935 and not w37339;
w37341 <= not w37337 and w37340;
w37342 <= not w36935 and not w37341;
w37343 <= b(31) and not w36924;
w37344 <= not w36918 and w37343;
w37345 <= not w36926 and not w37344;
w37346 <= not w37342 and w37345;
w37347 <= not w36926 and not w37346;
w37348 <= b(32) and not w36915;
w37349 <= not w36909 and w37348;
w37350 <= not w36917 and not w37349;
w37351 <= not w37347 and w37350;
w37352 <= not w36917 and not w37351;
w37353 <= b(33) and not w36906;
w37354 <= not w36900 and w37353;
w37355 <= not w36908 and not w37354;
w37356 <= not w37352 and w37355;
w37357 <= not w36908 and not w37356;
w37358 <= b(34) and not w36897;
w37359 <= not w36891 and w37358;
w37360 <= not w36899 and not w37359;
w37361 <= not w37357 and w37360;
w37362 <= not w36899 and not w37361;
w37363 <= not w36433 and not w36890;
w37364 <= not w36435 and w36887;
w37365 <= not w36883 and w37364;
w37366 <= not w36884 and not w36887;
w37367 <= not w37365 and not w37366;
w37368 <= w36890 and not w37367;
w37369 <= not w37363 and not w37368;
w37370 <= not b(35) and not w37369;
w37371 <= b(35) and not w37363;
w37372 <= not w37368 and w37371;
w37373 <= w255 and not w37372;
w37374 <= not w37370 and w37373;
w37375 <= not w37362 and w37374;
w37376 <= w8747 and not w37369;
w37377 <= not w37375 and not w37376;
w37378 <= not w36908 and w37360;
w37379 <= not w37356 and w37378;
w37380 <= not w37357 and not w37360;
w37381 <= not w37379 and not w37380;
w37382 <= not w37377 and not w37381;
w37383 <= not w36898 and not w37376;
w37384 <= not w37375 and w37383;
w37385 <= not w37382 and not w37384;
w37386 <= not w36899 and not w37372;
w37387 <= not w37370 and w37386;
w37388 <= not w37361 and w37387;
w37389 <= not w37370 and not w37372;
w37390 <= not w37362 and not w37389;
w37391 <= not w37388 and not w37390;
w37392 <= not w37377 and not w37391;
w37393 <= not w37369 and not w37376;
w37394 <= not w37375 and w37393;
w37395 <= not w37392 and not w37394;
w37396 <= not b(36) and not w37395;
w37397 <= not b(35) and not w37385;
w37398 <= not w36917 and w37355;
w37399 <= not w37351 and w37398;
w37400 <= not w37352 and not w37355;
w37401 <= not w37399 and not w37400;
w37402 <= not w37377 and not w37401;
w37403 <= not w36907 and not w37376;
w37404 <= not w37375 and w37403;
w37405 <= not w37402 and not w37404;
w37406 <= not b(34) and not w37405;
w37407 <= not w36926 and w37350;
w37408 <= not w37346 and w37407;
w37409 <= not w37347 and not w37350;
w37410 <= not w37408 and not w37409;
w37411 <= not w37377 and not w37410;
w37412 <= not w36916 and not w37376;
w37413 <= not w37375 and w37412;
w37414 <= not w37411 and not w37413;
w37415 <= not b(33) and not w37414;
w37416 <= not w36935 and w37345;
w37417 <= not w37341 and w37416;
w37418 <= not w37342 and not w37345;
w37419 <= not w37417 and not w37418;
w37420 <= not w37377 and not w37419;
w37421 <= not w36925 and not w37376;
w37422 <= not w37375 and w37421;
w37423 <= not w37420 and not w37422;
w37424 <= not b(32) and not w37423;
w37425 <= not w36944 and w37340;
w37426 <= not w37336 and w37425;
w37427 <= not w37337 and not w37340;
w37428 <= not w37426 and not w37427;
w37429 <= not w37377 and not w37428;
w37430 <= not w36934 and not w37376;
w37431 <= not w37375 and w37430;
w37432 <= not w37429 and not w37431;
w37433 <= not b(31) and not w37432;
w37434 <= not w36953 and w37335;
w37435 <= not w37331 and w37434;
w37436 <= not w37332 and not w37335;
w37437 <= not w37435 and not w37436;
w37438 <= not w37377 and not w37437;
w37439 <= not w36943 and not w37376;
w37440 <= not w37375 and w37439;
w37441 <= not w37438 and not w37440;
w37442 <= not b(30) and not w37441;
w37443 <= not w36962 and w37330;
w37444 <= not w37326 and w37443;
w37445 <= not w37327 and not w37330;
w37446 <= not w37444 and not w37445;
w37447 <= not w37377 and not w37446;
w37448 <= not w36952 and not w37376;
w37449 <= not w37375 and w37448;
w37450 <= not w37447 and not w37449;
w37451 <= not b(29) and not w37450;
w37452 <= not w36971 and w37325;
w37453 <= not w37321 and w37452;
w37454 <= not w37322 and not w37325;
w37455 <= not w37453 and not w37454;
w37456 <= not w37377 and not w37455;
w37457 <= not w36961 and not w37376;
w37458 <= not w37375 and w37457;
w37459 <= not w37456 and not w37458;
w37460 <= not b(28) and not w37459;
w37461 <= not w36980 and w37320;
w37462 <= not w37316 and w37461;
w37463 <= not w37317 and not w37320;
w37464 <= not w37462 and not w37463;
w37465 <= not w37377 and not w37464;
w37466 <= not w36970 and not w37376;
w37467 <= not w37375 and w37466;
w37468 <= not w37465 and not w37467;
w37469 <= not b(27) and not w37468;
w37470 <= not w36989 and w37315;
w37471 <= not w37311 and w37470;
w37472 <= not w37312 and not w37315;
w37473 <= not w37471 and not w37472;
w37474 <= not w37377 and not w37473;
w37475 <= not w36979 and not w37376;
w37476 <= not w37375 and w37475;
w37477 <= not w37474 and not w37476;
w37478 <= not b(26) and not w37477;
w37479 <= not w36998 and w37310;
w37480 <= not w37306 and w37479;
w37481 <= not w37307 and not w37310;
w37482 <= not w37480 and not w37481;
w37483 <= not w37377 and not w37482;
w37484 <= not w36988 and not w37376;
w37485 <= not w37375 and w37484;
w37486 <= not w37483 and not w37485;
w37487 <= not b(25) and not w37486;
w37488 <= not w37007 and w37305;
w37489 <= not w37301 and w37488;
w37490 <= not w37302 and not w37305;
w37491 <= not w37489 and not w37490;
w37492 <= not w37377 and not w37491;
w37493 <= not w36997 and not w37376;
w37494 <= not w37375 and w37493;
w37495 <= not w37492 and not w37494;
w37496 <= not b(24) and not w37495;
w37497 <= not w37016 and w37300;
w37498 <= not w37296 and w37497;
w37499 <= not w37297 and not w37300;
w37500 <= not w37498 and not w37499;
w37501 <= not w37377 and not w37500;
w37502 <= not w37006 and not w37376;
w37503 <= not w37375 and w37502;
w37504 <= not w37501 and not w37503;
w37505 <= not b(23) and not w37504;
w37506 <= not w37025 and w37295;
w37507 <= not w37291 and w37506;
w37508 <= not w37292 and not w37295;
w37509 <= not w37507 and not w37508;
w37510 <= not w37377 and not w37509;
w37511 <= not w37015 and not w37376;
w37512 <= not w37375 and w37511;
w37513 <= not w37510 and not w37512;
w37514 <= not b(22) and not w37513;
w37515 <= not w37034 and w37290;
w37516 <= not w37286 and w37515;
w37517 <= not w37287 and not w37290;
w37518 <= not w37516 and not w37517;
w37519 <= not w37377 and not w37518;
w37520 <= not w37024 and not w37376;
w37521 <= not w37375 and w37520;
w37522 <= not w37519 and not w37521;
w37523 <= not b(21) and not w37522;
w37524 <= not w37043 and w37285;
w37525 <= not w37281 and w37524;
w37526 <= not w37282 and not w37285;
w37527 <= not w37525 and not w37526;
w37528 <= not w37377 and not w37527;
w37529 <= not w37033 and not w37376;
w37530 <= not w37375 and w37529;
w37531 <= not w37528 and not w37530;
w37532 <= not b(20) and not w37531;
w37533 <= not w37052 and w37280;
w37534 <= not w37276 and w37533;
w37535 <= not w37277 and not w37280;
w37536 <= not w37534 and not w37535;
w37537 <= not w37377 and not w37536;
w37538 <= not w37042 and not w37376;
w37539 <= not w37375 and w37538;
w37540 <= not w37537 and not w37539;
w37541 <= not b(19) and not w37540;
w37542 <= not w37061 and w37275;
w37543 <= not w37271 and w37542;
w37544 <= not w37272 and not w37275;
w37545 <= not w37543 and not w37544;
w37546 <= not w37377 and not w37545;
w37547 <= not w37051 and not w37376;
w37548 <= not w37375 and w37547;
w37549 <= not w37546 and not w37548;
w37550 <= not b(18) and not w37549;
w37551 <= not w37070 and w37270;
w37552 <= not w37266 and w37551;
w37553 <= not w37267 and not w37270;
w37554 <= not w37552 and not w37553;
w37555 <= not w37377 and not w37554;
w37556 <= not w37060 and not w37376;
w37557 <= not w37375 and w37556;
w37558 <= not w37555 and not w37557;
w37559 <= not b(17) and not w37558;
w37560 <= not w37079 and w37265;
w37561 <= not w37261 and w37560;
w37562 <= not w37262 and not w37265;
w37563 <= not w37561 and not w37562;
w37564 <= not w37377 and not w37563;
w37565 <= not w37069 and not w37376;
w37566 <= not w37375 and w37565;
w37567 <= not w37564 and not w37566;
w37568 <= not b(16) and not w37567;
w37569 <= not w37088 and w37260;
w37570 <= not w37256 and w37569;
w37571 <= not w37257 and not w37260;
w37572 <= not w37570 and not w37571;
w37573 <= not w37377 and not w37572;
w37574 <= not w37078 and not w37376;
w37575 <= not w37375 and w37574;
w37576 <= not w37573 and not w37575;
w37577 <= not b(15) and not w37576;
w37578 <= not w37097 and w37255;
w37579 <= not w37251 and w37578;
w37580 <= not w37252 and not w37255;
w37581 <= not w37579 and not w37580;
w37582 <= not w37377 and not w37581;
w37583 <= not w37087 and not w37376;
w37584 <= not w37375 and w37583;
w37585 <= not w37582 and not w37584;
w37586 <= not b(14) and not w37585;
w37587 <= not w37106 and w37250;
w37588 <= not w37246 and w37587;
w37589 <= not w37247 and not w37250;
w37590 <= not w37588 and not w37589;
w37591 <= not w37377 and not w37590;
w37592 <= not w37096 and not w37376;
w37593 <= not w37375 and w37592;
w37594 <= not w37591 and not w37593;
w37595 <= not b(13) and not w37594;
w37596 <= not w37115 and w37245;
w37597 <= not w37241 and w37596;
w37598 <= not w37242 and not w37245;
w37599 <= not w37597 and not w37598;
w37600 <= not w37377 and not w37599;
w37601 <= not w37105 and not w37376;
w37602 <= not w37375 and w37601;
w37603 <= not w37600 and not w37602;
w37604 <= not b(12) and not w37603;
w37605 <= not w37124 and w37240;
w37606 <= not w37236 and w37605;
w37607 <= not w37237 and not w37240;
w37608 <= not w37606 and not w37607;
w37609 <= not w37377 and not w37608;
w37610 <= not w37114 and not w37376;
w37611 <= not w37375 and w37610;
w37612 <= not w37609 and not w37611;
w37613 <= not b(11) and not w37612;
w37614 <= not w37133 and w37235;
w37615 <= not w37231 and w37614;
w37616 <= not w37232 and not w37235;
w37617 <= not w37615 and not w37616;
w37618 <= not w37377 and not w37617;
w37619 <= not w37123 and not w37376;
w37620 <= not w37375 and w37619;
w37621 <= not w37618 and not w37620;
w37622 <= not b(10) and not w37621;
w37623 <= not w37142 and w37230;
w37624 <= not w37226 and w37623;
w37625 <= not w37227 and not w37230;
w37626 <= not w37624 and not w37625;
w37627 <= not w37377 and not w37626;
w37628 <= not w37132 and not w37376;
w37629 <= not w37375 and w37628;
w37630 <= not w37627 and not w37629;
w37631 <= not b(9) and not w37630;
w37632 <= not w37151 and w37225;
w37633 <= not w37221 and w37632;
w37634 <= not w37222 and not w37225;
w37635 <= not w37633 and not w37634;
w37636 <= not w37377 and not w37635;
w37637 <= not w37141 and not w37376;
w37638 <= not w37375 and w37637;
w37639 <= not w37636 and not w37638;
w37640 <= not b(8) and not w37639;
w37641 <= not w37160 and w37220;
w37642 <= not w37216 and w37641;
w37643 <= not w37217 and not w37220;
w37644 <= not w37642 and not w37643;
w37645 <= not w37377 and not w37644;
w37646 <= not w37150 and not w37376;
w37647 <= not w37375 and w37646;
w37648 <= not w37645 and not w37647;
w37649 <= not b(7) and not w37648;
w37650 <= not w37169 and w37215;
w37651 <= not w37211 and w37650;
w37652 <= not w37212 and not w37215;
w37653 <= not w37651 and not w37652;
w37654 <= not w37377 and not w37653;
w37655 <= not w37159 and not w37376;
w37656 <= not w37375 and w37655;
w37657 <= not w37654 and not w37656;
w37658 <= not b(6) and not w37657;
w37659 <= not w37178 and w37210;
w37660 <= not w37206 and w37659;
w37661 <= not w37207 and not w37210;
w37662 <= not w37660 and not w37661;
w37663 <= not w37377 and not w37662;
w37664 <= not w37168 and not w37376;
w37665 <= not w37375 and w37664;
w37666 <= not w37663 and not w37665;
w37667 <= not b(5) and not w37666;
w37668 <= not w37186 and w37205;
w37669 <= not w37201 and w37668;
w37670 <= not w37202 and not w37205;
w37671 <= not w37669 and not w37670;
w37672 <= not w37377 and not w37671;
w37673 <= not w37177 and not w37376;
w37674 <= not w37375 and w37673;
w37675 <= not w37672 and not w37674;
w37676 <= not b(4) and not w37675;
w37677 <= not w37196 and w37200;
w37678 <= not w37195 and w37677;
w37679 <= not w37197 and not w37200;
w37680 <= not w37678 and not w37679;
w37681 <= not w37377 and not w37680;
w37682 <= not w37185 and not w37376;
w37683 <= not w37375 and w37682;
w37684 <= not w37681 and not w37683;
w37685 <= not b(3) and not w37684;
w37686 <= w9061 and not w37193;
w37687 <= not w37191 and w37686;
w37688 <= not w37195 and not w37687;
w37689 <= not w37377 and w37688;
w37690 <= not w37190 and not w37376;
w37691 <= not w37375 and w37690;
w37692 <= not w37689 and not w37691;
w37693 <= not b(2) and not w37692;
w37694 <= b(0) and not w37377;
w37695 <= a(28) and not w37694;
w37696 <= w9061 and not w37377;
w37697 <= not w37695 and not w37696;
w37698 <= b(1) and not w37697;
w37699 <= not b(1) and not w37696;
w37700 <= not w37695 and w37699;
w37701 <= not w37698 and not w37700;
w37702 <= not w9569 and not w37701;
w37703 <= not b(1) and not w37697;
w37704 <= not w37702 and not w37703;
w37705 <= b(2) and not w37691;
w37706 <= not w37689 and w37705;
w37707 <= not w37693 and not w37706;
w37708 <= not w37704 and w37707;
w37709 <= not w37693 and not w37708;
w37710 <= b(3) and not w37683;
w37711 <= not w37681 and w37710;
w37712 <= not w37685 and not w37711;
w37713 <= not w37709 and w37712;
w37714 <= not w37685 and not w37713;
w37715 <= b(4) and not w37674;
w37716 <= not w37672 and w37715;
w37717 <= not w37676 and not w37716;
w37718 <= not w37714 and w37717;
w37719 <= not w37676 and not w37718;
w37720 <= b(5) and not w37665;
w37721 <= not w37663 and w37720;
w37722 <= not w37667 and not w37721;
w37723 <= not w37719 and w37722;
w37724 <= not w37667 and not w37723;
w37725 <= b(6) and not w37656;
w37726 <= not w37654 and w37725;
w37727 <= not w37658 and not w37726;
w37728 <= not w37724 and w37727;
w37729 <= not w37658 and not w37728;
w37730 <= b(7) and not w37647;
w37731 <= not w37645 and w37730;
w37732 <= not w37649 and not w37731;
w37733 <= not w37729 and w37732;
w37734 <= not w37649 and not w37733;
w37735 <= b(8) and not w37638;
w37736 <= not w37636 and w37735;
w37737 <= not w37640 and not w37736;
w37738 <= not w37734 and w37737;
w37739 <= not w37640 and not w37738;
w37740 <= b(9) and not w37629;
w37741 <= not w37627 and w37740;
w37742 <= not w37631 and not w37741;
w37743 <= not w37739 and w37742;
w37744 <= not w37631 and not w37743;
w37745 <= b(10) and not w37620;
w37746 <= not w37618 and w37745;
w37747 <= not w37622 and not w37746;
w37748 <= not w37744 and w37747;
w37749 <= not w37622 and not w37748;
w37750 <= b(11) and not w37611;
w37751 <= not w37609 and w37750;
w37752 <= not w37613 and not w37751;
w37753 <= not w37749 and w37752;
w37754 <= not w37613 and not w37753;
w37755 <= b(12) and not w37602;
w37756 <= not w37600 and w37755;
w37757 <= not w37604 and not w37756;
w37758 <= not w37754 and w37757;
w37759 <= not w37604 and not w37758;
w37760 <= b(13) and not w37593;
w37761 <= not w37591 and w37760;
w37762 <= not w37595 and not w37761;
w37763 <= not w37759 and w37762;
w37764 <= not w37595 and not w37763;
w37765 <= b(14) and not w37584;
w37766 <= not w37582 and w37765;
w37767 <= not w37586 and not w37766;
w37768 <= not w37764 and w37767;
w37769 <= not w37586 and not w37768;
w37770 <= b(15) and not w37575;
w37771 <= not w37573 and w37770;
w37772 <= not w37577 and not w37771;
w37773 <= not w37769 and w37772;
w37774 <= not w37577 and not w37773;
w37775 <= b(16) and not w37566;
w37776 <= not w37564 and w37775;
w37777 <= not w37568 and not w37776;
w37778 <= not w37774 and w37777;
w37779 <= not w37568 and not w37778;
w37780 <= b(17) and not w37557;
w37781 <= not w37555 and w37780;
w37782 <= not w37559 and not w37781;
w37783 <= not w37779 and w37782;
w37784 <= not w37559 and not w37783;
w37785 <= b(18) and not w37548;
w37786 <= not w37546 and w37785;
w37787 <= not w37550 and not w37786;
w37788 <= not w37784 and w37787;
w37789 <= not w37550 and not w37788;
w37790 <= b(19) and not w37539;
w37791 <= not w37537 and w37790;
w37792 <= not w37541 and not w37791;
w37793 <= not w37789 and w37792;
w37794 <= not w37541 and not w37793;
w37795 <= b(20) and not w37530;
w37796 <= not w37528 and w37795;
w37797 <= not w37532 and not w37796;
w37798 <= not w37794 and w37797;
w37799 <= not w37532 and not w37798;
w37800 <= b(21) and not w37521;
w37801 <= not w37519 and w37800;
w37802 <= not w37523 and not w37801;
w37803 <= not w37799 and w37802;
w37804 <= not w37523 and not w37803;
w37805 <= b(22) and not w37512;
w37806 <= not w37510 and w37805;
w37807 <= not w37514 and not w37806;
w37808 <= not w37804 and w37807;
w37809 <= not w37514 and not w37808;
w37810 <= b(23) and not w37503;
w37811 <= not w37501 and w37810;
w37812 <= not w37505 and not w37811;
w37813 <= not w37809 and w37812;
w37814 <= not w37505 and not w37813;
w37815 <= b(24) and not w37494;
w37816 <= not w37492 and w37815;
w37817 <= not w37496 and not w37816;
w37818 <= not w37814 and w37817;
w37819 <= not w37496 and not w37818;
w37820 <= b(25) and not w37485;
w37821 <= not w37483 and w37820;
w37822 <= not w37487 and not w37821;
w37823 <= not w37819 and w37822;
w37824 <= not w37487 and not w37823;
w37825 <= b(26) and not w37476;
w37826 <= not w37474 and w37825;
w37827 <= not w37478 and not w37826;
w37828 <= not w37824 and w37827;
w37829 <= not w37478 and not w37828;
w37830 <= b(27) and not w37467;
w37831 <= not w37465 and w37830;
w37832 <= not w37469 and not w37831;
w37833 <= not w37829 and w37832;
w37834 <= not w37469 and not w37833;
w37835 <= b(28) and not w37458;
w37836 <= not w37456 and w37835;
w37837 <= not w37460 and not w37836;
w37838 <= not w37834 and w37837;
w37839 <= not w37460 and not w37838;
w37840 <= b(29) and not w37449;
w37841 <= not w37447 and w37840;
w37842 <= not w37451 and not w37841;
w37843 <= not w37839 and w37842;
w37844 <= not w37451 and not w37843;
w37845 <= b(30) and not w37440;
w37846 <= not w37438 and w37845;
w37847 <= not w37442 and not w37846;
w37848 <= not w37844 and w37847;
w37849 <= not w37442 and not w37848;
w37850 <= b(31) and not w37431;
w37851 <= not w37429 and w37850;
w37852 <= not w37433 and not w37851;
w37853 <= not w37849 and w37852;
w37854 <= not w37433 and not w37853;
w37855 <= b(32) and not w37422;
w37856 <= not w37420 and w37855;
w37857 <= not w37424 and not w37856;
w37858 <= not w37854 and w37857;
w37859 <= not w37424 and not w37858;
w37860 <= b(33) and not w37413;
w37861 <= not w37411 and w37860;
w37862 <= not w37415 and not w37861;
w37863 <= not w37859 and w37862;
w37864 <= not w37415 and not w37863;
w37865 <= b(34) and not w37404;
w37866 <= not w37402 and w37865;
w37867 <= not w37406 and not w37866;
w37868 <= not w37864 and w37867;
w37869 <= not w37406 and not w37868;
w37870 <= b(35) and not w37384;
w37871 <= not w37382 and w37870;
w37872 <= not w37397 and not w37871;
w37873 <= not w37869 and w37872;
w37874 <= not w37397 and not w37873;
w37875 <= b(36) and not w37394;
w37876 <= not w37392 and w37875;
w37877 <= not w37396 and not w37876;
w37878 <= not w37874 and w37877;
w37879 <= not w37396 and not w37878;
w37880 <= w342 and not w37879;
w37881 <= not w37385 and not w37880;
w37882 <= not w37406 and w37872;
w37883 <= not w37868 and w37882;
w37884 <= not w37869 and not w37872;
w37885 <= not w37883 and not w37884;
w37886 <= w342 and not w37885;
w37887 <= not w37879 and w37886;
w37888 <= not w37881 and not w37887;
w37889 <= not w37395 and not w37880;
w37890 <= not w37397 and w37877;
w37891 <= not w37873 and w37890;
w37892 <= not w37874 and not w37877;
w37893 <= not w37891 and not w37892;
w37894 <= w37880 and not w37893;
w37895 <= not w37889 and not w37894;
w37896 <= not b(37) and not w37895;
w37897 <= not b(36) and not w37888;
w37898 <= not w37405 and not w37880;
w37899 <= not w37415 and w37867;
w37900 <= not w37863 and w37899;
w37901 <= not w37864 and not w37867;
w37902 <= not w37900 and not w37901;
w37903 <= w342 and not w37902;
w37904 <= not w37879 and w37903;
w37905 <= not w37898 and not w37904;
w37906 <= not b(35) and not w37905;
w37907 <= not w37414 and not w37880;
w37908 <= not w37424 and w37862;
w37909 <= not w37858 and w37908;
w37910 <= not w37859 and not w37862;
w37911 <= not w37909 and not w37910;
w37912 <= w342 and not w37911;
w37913 <= not w37879 and w37912;
w37914 <= not w37907 and not w37913;
w37915 <= not b(34) and not w37914;
w37916 <= not w37423 and not w37880;
w37917 <= not w37433 and w37857;
w37918 <= not w37853 and w37917;
w37919 <= not w37854 and not w37857;
w37920 <= not w37918 and not w37919;
w37921 <= w342 and not w37920;
w37922 <= not w37879 and w37921;
w37923 <= not w37916 and not w37922;
w37924 <= not b(33) and not w37923;
w37925 <= not w37432 and not w37880;
w37926 <= not w37442 and w37852;
w37927 <= not w37848 and w37926;
w37928 <= not w37849 and not w37852;
w37929 <= not w37927 and not w37928;
w37930 <= w342 and not w37929;
w37931 <= not w37879 and w37930;
w37932 <= not w37925 and not w37931;
w37933 <= not b(32) and not w37932;
w37934 <= not w37441 and not w37880;
w37935 <= not w37451 and w37847;
w37936 <= not w37843 and w37935;
w37937 <= not w37844 and not w37847;
w37938 <= not w37936 and not w37937;
w37939 <= w342 and not w37938;
w37940 <= not w37879 and w37939;
w37941 <= not w37934 and not w37940;
w37942 <= not b(31) and not w37941;
w37943 <= not w37450 and not w37880;
w37944 <= not w37460 and w37842;
w37945 <= not w37838 and w37944;
w37946 <= not w37839 and not w37842;
w37947 <= not w37945 and not w37946;
w37948 <= w342 and not w37947;
w37949 <= not w37879 and w37948;
w37950 <= not w37943 and not w37949;
w37951 <= not b(30) and not w37950;
w37952 <= not w37459 and not w37880;
w37953 <= not w37469 and w37837;
w37954 <= not w37833 and w37953;
w37955 <= not w37834 and not w37837;
w37956 <= not w37954 and not w37955;
w37957 <= w342 and not w37956;
w37958 <= not w37879 and w37957;
w37959 <= not w37952 and not w37958;
w37960 <= not b(29) and not w37959;
w37961 <= not w37468 and not w37880;
w37962 <= not w37478 and w37832;
w37963 <= not w37828 and w37962;
w37964 <= not w37829 and not w37832;
w37965 <= not w37963 and not w37964;
w37966 <= w342 and not w37965;
w37967 <= not w37879 and w37966;
w37968 <= not w37961 and not w37967;
w37969 <= not b(28) and not w37968;
w37970 <= not w37477 and not w37880;
w37971 <= not w37487 and w37827;
w37972 <= not w37823 and w37971;
w37973 <= not w37824 and not w37827;
w37974 <= not w37972 and not w37973;
w37975 <= w342 and not w37974;
w37976 <= not w37879 and w37975;
w37977 <= not w37970 and not w37976;
w37978 <= not b(27) and not w37977;
w37979 <= not w37486 and not w37880;
w37980 <= not w37496 and w37822;
w37981 <= not w37818 and w37980;
w37982 <= not w37819 and not w37822;
w37983 <= not w37981 and not w37982;
w37984 <= w342 and not w37983;
w37985 <= not w37879 and w37984;
w37986 <= not w37979 and not w37985;
w37987 <= not b(26) and not w37986;
w37988 <= not w37495 and not w37880;
w37989 <= not w37505 and w37817;
w37990 <= not w37813 and w37989;
w37991 <= not w37814 and not w37817;
w37992 <= not w37990 and not w37991;
w37993 <= w342 and not w37992;
w37994 <= not w37879 and w37993;
w37995 <= not w37988 and not w37994;
w37996 <= not b(25) and not w37995;
w37997 <= not w37504 and not w37880;
w37998 <= not w37514 and w37812;
w37999 <= not w37808 and w37998;
w38000 <= not w37809 and not w37812;
w38001 <= not w37999 and not w38000;
w38002 <= w342 and not w38001;
w38003 <= not w37879 and w38002;
w38004 <= not w37997 and not w38003;
w38005 <= not b(24) and not w38004;
w38006 <= not w37513 and not w37880;
w38007 <= not w37523 and w37807;
w38008 <= not w37803 and w38007;
w38009 <= not w37804 and not w37807;
w38010 <= not w38008 and not w38009;
w38011 <= w342 and not w38010;
w38012 <= not w37879 and w38011;
w38013 <= not w38006 and not w38012;
w38014 <= not b(23) and not w38013;
w38015 <= not w37522 and not w37880;
w38016 <= not w37532 and w37802;
w38017 <= not w37798 and w38016;
w38018 <= not w37799 and not w37802;
w38019 <= not w38017 and not w38018;
w38020 <= w342 and not w38019;
w38021 <= not w37879 and w38020;
w38022 <= not w38015 and not w38021;
w38023 <= not b(22) and not w38022;
w38024 <= not w37531 and not w37880;
w38025 <= not w37541 and w37797;
w38026 <= not w37793 and w38025;
w38027 <= not w37794 and not w37797;
w38028 <= not w38026 and not w38027;
w38029 <= w342 and not w38028;
w38030 <= not w37879 and w38029;
w38031 <= not w38024 and not w38030;
w38032 <= not b(21) and not w38031;
w38033 <= not w37540 and not w37880;
w38034 <= not w37550 and w37792;
w38035 <= not w37788 and w38034;
w38036 <= not w37789 and not w37792;
w38037 <= not w38035 and not w38036;
w38038 <= w342 and not w38037;
w38039 <= not w37879 and w38038;
w38040 <= not w38033 and not w38039;
w38041 <= not b(20) and not w38040;
w38042 <= not w37549 and not w37880;
w38043 <= not w37559 and w37787;
w38044 <= not w37783 and w38043;
w38045 <= not w37784 and not w37787;
w38046 <= not w38044 and not w38045;
w38047 <= w342 and not w38046;
w38048 <= not w37879 and w38047;
w38049 <= not w38042 and not w38048;
w38050 <= not b(19) and not w38049;
w38051 <= not w37558 and not w37880;
w38052 <= not w37568 and w37782;
w38053 <= not w37778 and w38052;
w38054 <= not w37779 and not w37782;
w38055 <= not w38053 and not w38054;
w38056 <= w342 and not w38055;
w38057 <= not w37879 and w38056;
w38058 <= not w38051 and not w38057;
w38059 <= not b(18) and not w38058;
w38060 <= not w37567 and not w37880;
w38061 <= not w37577 and w37777;
w38062 <= not w37773 and w38061;
w38063 <= not w37774 and not w37777;
w38064 <= not w38062 and not w38063;
w38065 <= w342 and not w38064;
w38066 <= not w37879 and w38065;
w38067 <= not w38060 and not w38066;
w38068 <= not b(17) and not w38067;
w38069 <= not w37576 and not w37880;
w38070 <= not w37586 and w37772;
w38071 <= not w37768 and w38070;
w38072 <= not w37769 and not w37772;
w38073 <= not w38071 and not w38072;
w38074 <= w342 and not w38073;
w38075 <= not w37879 and w38074;
w38076 <= not w38069 and not w38075;
w38077 <= not b(16) and not w38076;
w38078 <= not w37585 and not w37880;
w38079 <= not w37595 and w37767;
w38080 <= not w37763 and w38079;
w38081 <= not w37764 and not w37767;
w38082 <= not w38080 and not w38081;
w38083 <= w342 and not w38082;
w38084 <= not w37879 and w38083;
w38085 <= not w38078 and not w38084;
w38086 <= not b(15) and not w38085;
w38087 <= not w37594 and not w37880;
w38088 <= not w37604 and w37762;
w38089 <= not w37758 and w38088;
w38090 <= not w37759 and not w37762;
w38091 <= not w38089 and not w38090;
w38092 <= w342 and not w38091;
w38093 <= not w37879 and w38092;
w38094 <= not w38087 and not w38093;
w38095 <= not b(14) and not w38094;
w38096 <= not w37603 and not w37880;
w38097 <= not w37613 and w37757;
w38098 <= not w37753 and w38097;
w38099 <= not w37754 and not w37757;
w38100 <= not w38098 and not w38099;
w38101 <= w342 and not w38100;
w38102 <= not w37879 and w38101;
w38103 <= not w38096 and not w38102;
w38104 <= not b(13) and not w38103;
w38105 <= not w37612 and not w37880;
w38106 <= not w37622 and w37752;
w38107 <= not w37748 and w38106;
w38108 <= not w37749 and not w37752;
w38109 <= not w38107 and not w38108;
w38110 <= w342 and not w38109;
w38111 <= not w37879 and w38110;
w38112 <= not w38105 and not w38111;
w38113 <= not b(12) and not w38112;
w38114 <= not w37621 and not w37880;
w38115 <= not w37631 and w37747;
w38116 <= not w37743 and w38115;
w38117 <= not w37744 and not w37747;
w38118 <= not w38116 and not w38117;
w38119 <= w342 and not w38118;
w38120 <= not w37879 and w38119;
w38121 <= not w38114 and not w38120;
w38122 <= not b(11) and not w38121;
w38123 <= not w37630 and not w37880;
w38124 <= not w37640 and w37742;
w38125 <= not w37738 and w38124;
w38126 <= not w37739 and not w37742;
w38127 <= not w38125 and not w38126;
w38128 <= w342 and not w38127;
w38129 <= not w37879 and w38128;
w38130 <= not w38123 and not w38129;
w38131 <= not b(10) and not w38130;
w38132 <= not w37639 and not w37880;
w38133 <= not w37649 and w37737;
w38134 <= not w37733 and w38133;
w38135 <= not w37734 and not w37737;
w38136 <= not w38134 and not w38135;
w38137 <= w342 and not w38136;
w38138 <= not w37879 and w38137;
w38139 <= not w38132 and not w38138;
w38140 <= not b(9) and not w38139;
w38141 <= not w37648 and not w37880;
w38142 <= not w37658 and w37732;
w38143 <= not w37728 and w38142;
w38144 <= not w37729 and not w37732;
w38145 <= not w38143 and not w38144;
w38146 <= w342 and not w38145;
w38147 <= not w37879 and w38146;
w38148 <= not w38141 and not w38147;
w38149 <= not b(8) and not w38148;
w38150 <= not w37657 and not w37880;
w38151 <= not w37667 and w37727;
w38152 <= not w37723 and w38151;
w38153 <= not w37724 and not w37727;
w38154 <= not w38152 and not w38153;
w38155 <= w342 and not w38154;
w38156 <= not w37879 and w38155;
w38157 <= not w38150 and not w38156;
w38158 <= not b(7) and not w38157;
w38159 <= not w37666 and not w37880;
w38160 <= not w37676 and w37722;
w38161 <= not w37718 and w38160;
w38162 <= not w37719 and not w37722;
w38163 <= not w38161 and not w38162;
w38164 <= w342 and not w38163;
w38165 <= not w37879 and w38164;
w38166 <= not w38159 and not w38165;
w38167 <= not b(6) and not w38166;
w38168 <= not w37675 and not w37880;
w38169 <= not w37685 and w37717;
w38170 <= not w37713 and w38169;
w38171 <= not w37714 and not w37717;
w38172 <= not w38170 and not w38171;
w38173 <= w342 and not w38172;
w38174 <= not w37879 and w38173;
w38175 <= not w38168 and not w38174;
w38176 <= not b(5) and not w38175;
w38177 <= not w37684 and not w37880;
w38178 <= not w37693 and w37712;
w38179 <= not w37708 and w38178;
w38180 <= not w37709 and not w37712;
w38181 <= not w38179 and not w38180;
w38182 <= w342 and not w38181;
w38183 <= not w37879 and w38182;
w38184 <= not w38177 and not w38183;
w38185 <= not b(4) and not w38184;
w38186 <= not w37692 and not w37880;
w38187 <= not w37703 and w37707;
w38188 <= not w37702 and w38187;
w38189 <= not w37704 and not w37707;
w38190 <= not w38188 and not w38189;
w38191 <= w342 and not w38190;
w38192 <= not w37879 and w38191;
w38193 <= not w38186 and not w38192;
w38194 <= not b(3) and not w38193;
w38195 <= not w37697 and not w37880;
w38196 <= w9569 and not w37700;
w38197 <= not w37698 and w38196;
w38198 <= w342 and not w38197;
w38199 <= not w37702 and w38198;
w38200 <= not w37879 and w38199;
w38201 <= not w38195 and not w38200;
w38202 <= not b(2) and not w38201;
w38203 <= w10075 and not w37879;
w38204 <= a(27) and not w38203;
w38205 <= w10080 and not w37879;
w38206 <= not w38204 and not w38205;
w38207 <= b(1) and not w38206;
w38208 <= not b(1) and not w38205;
w38209 <= not w38204 and w38208;
w38210 <= not w38207 and not w38209;
w38211 <= not w10087 and not w38210;
w38212 <= not b(1) and not w38206;
w38213 <= not w38211 and not w38212;
w38214 <= b(2) and not w38200;
w38215 <= not w38195 and w38214;
w38216 <= not w38202 and not w38215;
w38217 <= not w38213 and w38216;
w38218 <= not w38202 and not w38217;
w38219 <= b(3) and not w38192;
w38220 <= not w38186 and w38219;
w38221 <= not w38194 and not w38220;
w38222 <= not w38218 and w38221;
w38223 <= not w38194 and not w38222;
w38224 <= b(4) and not w38183;
w38225 <= not w38177 and w38224;
w38226 <= not w38185 and not w38225;
w38227 <= not w38223 and w38226;
w38228 <= not w38185 and not w38227;
w38229 <= b(5) and not w38174;
w38230 <= not w38168 and w38229;
w38231 <= not w38176 and not w38230;
w38232 <= not w38228 and w38231;
w38233 <= not w38176 and not w38232;
w38234 <= b(6) and not w38165;
w38235 <= not w38159 and w38234;
w38236 <= not w38167 and not w38235;
w38237 <= not w38233 and w38236;
w38238 <= not w38167 and not w38237;
w38239 <= b(7) and not w38156;
w38240 <= not w38150 and w38239;
w38241 <= not w38158 and not w38240;
w38242 <= not w38238 and w38241;
w38243 <= not w38158 and not w38242;
w38244 <= b(8) and not w38147;
w38245 <= not w38141 and w38244;
w38246 <= not w38149 and not w38245;
w38247 <= not w38243 and w38246;
w38248 <= not w38149 and not w38247;
w38249 <= b(9) and not w38138;
w38250 <= not w38132 and w38249;
w38251 <= not w38140 and not w38250;
w38252 <= not w38248 and w38251;
w38253 <= not w38140 and not w38252;
w38254 <= b(10) and not w38129;
w38255 <= not w38123 and w38254;
w38256 <= not w38131 and not w38255;
w38257 <= not w38253 and w38256;
w38258 <= not w38131 and not w38257;
w38259 <= b(11) and not w38120;
w38260 <= not w38114 and w38259;
w38261 <= not w38122 and not w38260;
w38262 <= not w38258 and w38261;
w38263 <= not w38122 and not w38262;
w38264 <= b(12) and not w38111;
w38265 <= not w38105 and w38264;
w38266 <= not w38113 and not w38265;
w38267 <= not w38263 and w38266;
w38268 <= not w38113 and not w38267;
w38269 <= b(13) and not w38102;
w38270 <= not w38096 and w38269;
w38271 <= not w38104 and not w38270;
w38272 <= not w38268 and w38271;
w38273 <= not w38104 and not w38272;
w38274 <= b(14) and not w38093;
w38275 <= not w38087 and w38274;
w38276 <= not w38095 and not w38275;
w38277 <= not w38273 and w38276;
w38278 <= not w38095 and not w38277;
w38279 <= b(15) and not w38084;
w38280 <= not w38078 and w38279;
w38281 <= not w38086 and not w38280;
w38282 <= not w38278 and w38281;
w38283 <= not w38086 and not w38282;
w38284 <= b(16) and not w38075;
w38285 <= not w38069 and w38284;
w38286 <= not w38077 and not w38285;
w38287 <= not w38283 and w38286;
w38288 <= not w38077 and not w38287;
w38289 <= b(17) and not w38066;
w38290 <= not w38060 and w38289;
w38291 <= not w38068 and not w38290;
w38292 <= not w38288 and w38291;
w38293 <= not w38068 and not w38292;
w38294 <= b(18) and not w38057;
w38295 <= not w38051 and w38294;
w38296 <= not w38059 and not w38295;
w38297 <= not w38293 and w38296;
w38298 <= not w38059 and not w38297;
w38299 <= b(19) and not w38048;
w38300 <= not w38042 and w38299;
w38301 <= not w38050 and not w38300;
w38302 <= not w38298 and w38301;
w38303 <= not w38050 and not w38302;
w38304 <= b(20) and not w38039;
w38305 <= not w38033 and w38304;
w38306 <= not w38041 and not w38305;
w38307 <= not w38303 and w38306;
w38308 <= not w38041 and not w38307;
w38309 <= b(21) and not w38030;
w38310 <= not w38024 and w38309;
w38311 <= not w38032 and not w38310;
w38312 <= not w38308 and w38311;
w38313 <= not w38032 and not w38312;
w38314 <= b(22) and not w38021;
w38315 <= not w38015 and w38314;
w38316 <= not w38023 and not w38315;
w38317 <= not w38313 and w38316;
w38318 <= not w38023 and not w38317;
w38319 <= b(23) and not w38012;
w38320 <= not w38006 and w38319;
w38321 <= not w38014 and not w38320;
w38322 <= not w38318 and w38321;
w38323 <= not w38014 and not w38322;
w38324 <= b(24) and not w38003;
w38325 <= not w37997 and w38324;
w38326 <= not w38005 and not w38325;
w38327 <= not w38323 and w38326;
w38328 <= not w38005 and not w38327;
w38329 <= b(25) and not w37994;
w38330 <= not w37988 and w38329;
w38331 <= not w37996 and not w38330;
w38332 <= not w38328 and w38331;
w38333 <= not w37996 and not w38332;
w38334 <= b(26) and not w37985;
w38335 <= not w37979 and w38334;
w38336 <= not w37987 and not w38335;
w38337 <= not w38333 and w38336;
w38338 <= not w37987 and not w38337;
w38339 <= b(27) and not w37976;
w38340 <= not w37970 and w38339;
w38341 <= not w37978 and not w38340;
w38342 <= not w38338 and w38341;
w38343 <= not w37978 and not w38342;
w38344 <= b(28) and not w37967;
w38345 <= not w37961 and w38344;
w38346 <= not w37969 and not w38345;
w38347 <= not w38343 and w38346;
w38348 <= not w37969 and not w38347;
w38349 <= b(29) and not w37958;
w38350 <= not w37952 and w38349;
w38351 <= not w37960 and not w38350;
w38352 <= not w38348 and w38351;
w38353 <= not w37960 and not w38352;
w38354 <= b(30) and not w37949;
w38355 <= not w37943 and w38354;
w38356 <= not w37951 and not w38355;
w38357 <= not w38353 and w38356;
w38358 <= not w37951 and not w38357;
w38359 <= b(31) and not w37940;
w38360 <= not w37934 and w38359;
w38361 <= not w37942 and not w38360;
w38362 <= not w38358 and w38361;
w38363 <= not w37942 and not w38362;
w38364 <= b(32) and not w37931;
w38365 <= not w37925 and w38364;
w38366 <= not w37933 and not w38365;
w38367 <= not w38363 and w38366;
w38368 <= not w37933 and not w38367;
w38369 <= b(33) and not w37922;
w38370 <= not w37916 and w38369;
w38371 <= not w37924 and not w38370;
w38372 <= not w38368 and w38371;
w38373 <= not w37924 and not w38372;
w38374 <= b(34) and not w37913;
w38375 <= not w37907 and w38374;
w38376 <= not w37915 and not w38375;
w38377 <= not w38373 and w38376;
w38378 <= not w37915 and not w38377;
w38379 <= b(35) and not w37904;
w38380 <= not w37898 and w38379;
w38381 <= not w37906 and not w38380;
w38382 <= not w38378 and w38381;
w38383 <= not w37906 and not w38382;
w38384 <= b(36) and not w37887;
w38385 <= not w37881 and w38384;
w38386 <= not w37897 and not w38385;
w38387 <= not w38383 and w38386;
w38388 <= not w37897 and not w38387;
w38389 <= b(37) and not w37889;
w38390 <= not w37894 and w38389;
w38391 <= not w37896 and not w38390;
w38392 <= not w38388 and w38391;
w38393 <= not w37896 and not w38392;
w38394 <= w10273 and not w38393;
w38395 <= not w37888 and not w38394;
w38396 <= not w37906 and w38386;
w38397 <= not w38382 and w38396;
w38398 <= not w38383 and not w38386;
w38399 <= not w38397 and not w38398;
w38400 <= w10273 and not w38399;
w38401 <= not w38393 and w38400;
w38402 <= not w38395 and not w38401;
w38403 <= not b(37) and not w38402;
w38404 <= not w37905 and not w38394;
w38405 <= not w37915 and w38381;
w38406 <= not w38377 and w38405;
w38407 <= not w38378 and not w38381;
w38408 <= not w38406 and not w38407;
w38409 <= w10273 and not w38408;
w38410 <= not w38393 and w38409;
w38411 <= not w38404 and not w38410;
w38412 <= not b(36) and not w38411;
w38413 <= not w37914 and not w38394;
w38414 <= not w37924 and w38376;
w38415 <= not w38372 and w38414;
w38416 <= not w38373 and not w38376;
w38417 <= not w38415 and not w38416;
w38418 <= w10273 and not w38417;
w38419 <= not w38393 and w38418;
w38420 <= not w38413 and not w38419;
w38421 <= not b(35) and not w38420;
w38422 <= not w37923 and not w38394;
w38423 <= not w37933 and w38371;
w38424 <= not w38367 and w38423;
w38425 <= not w38368 and not w38371;
w38426 <= not w38424 and not w38425;
w38427 <= w10273 and not w38426;
w38428 <= not w38393 and w38427;
w38429 <= not w38422 and not w38428;
w38430 <= not b(34) and not w38429;
w38431 <= not w37932 and not w38394;
w38432 <= not w37942 and w38366;
w38433 <= not w38362 and w38432;
w38434 <= not w38363 and not w38366;
w38435 <= not w38433 and not w38434;
w38436 <= w10273 and not w38435;
w38437 <= not w38393 and w38436;
w38438 <= not w38431 and not w38437;
w38439 <= not b(33) and not w38438;
w38440 <= not w37941 and not w38394;
w38441 <= not w37951 and w38361;
w38442 <= not w38357 and w38441;
w38443 <= not w38358 and not w38361;
w38444 <= not w38442 and not w38443;
w38445 <= w10273 and not w38444;
w38446 <= not w38393 and w38445;
w38447 <= not w38440 and not w38446;
w38448 <= not b(32) and not w38447;
w38449 <= not w37950 and not w38394;
w38450 <= not w37960 and w38356;
w38451 <= not w38352 and w38450;
w38452 <= not w38353 and not w38356;
w38453 <= not w38451 and not w38452;
w38454 <= w10273 and not w38453;
w38455 <= not w38393 and w38454;
w38456 <= not w38449 and not w38455;
w38457 <= not b(31) and not w38456;
w38458 <= not w37959 and not w38394;
w38459 <= not w37969 and w38351;
w38460 <= not w38347 and w38459;
w38461 <= not w38348 and not w38351;
w38462 <= not w38460 and not w38461;
w38463 <= w10273 and not w38462;
w38464 <= not w38393 and w38463;
w38465 <= not w38458 and not w38464;
w38466 <= not b(30) and not w38465;
w38467 <= not w37968 and not w38394;
w38468 <= not w37978 and w38346;
w38469 <= not w38342 and w38468;
w38470 <= not w38343 and not w38346;
w38471 <= not w38469 and not w38470;
w38472 <= w10273 and not w38471;
w38473 <= not w38393 and w38472;
w38474 <= not w38467 and not w38473;
w38475 <= not b(29) and not w38474;
w38476 <= not w37977 and not w38394;
w38477 <= not w37987 and w38341;
w38478 <= not w38337 and w38477;
w38479 <= not w38338 and not w38341;
w38480 <= not w38478 and not w38479;
w38481 <= w10273 and not w38480;
w38482 <= not w38393 and w38481;
w38483 <= not w38476 and not w38482;
w38484 <= not b(28) and not w38483;
w38485 <= not w37986 and not w38394;
w38486 <= not w37996 and w38336;
w38487 <= not w38332 and w38486;
w38488 <= not w38333 and not w38336;
w38489 <= not w38487 and not w38488;
w38490 <= w10273 and not w38489;
w38491 <= not w38393 and w38490;
w38492 <= not w38485 and not w38491;
w38493 <= not b(27) and not w38492;
w38494 <= not w37995 and not w38394;
w38495 <= not w38005 and w38331;
w38496 <= not w38327 and w38495;
w38497 <= not w38328 and not w38331;
w38498 <= not w38496 and not w38497;
w38499 <= w10273 and not w38498;
w38500 <= not w38393 and w38499;
w38501 <= not w38494 and not w38500;
w38502 <= not b(26) and not w38501;
w38503 <= not w38004 and not w38394;
w38504 <= not w38014 and w38326;
w38505 <= not w38322 and w38504;
w38506 <= not w38323 and not w38326;
w38507 <= not w38505 and not w38506;
w38508 <= w10273 and not w38507;
w38509 <= not w38393 and w38508;
w38510 <= not w38503 and not w38509;
w38511 <= not b(25) and not w38510;
w38512 <= not w38013 and not w38394;
w38513 <= not w38023 and w38321;
w38514 <= not w38317 and w38513;
w38515 <= not w38318 and not w38321;
w38516 <= not w38514 and not w38515;
w38517 <= w10273 and not w38516;
w38518 <= not w38393 and w38517;
w38519 <= not w38512 and not w38518;
w38520 <= not b(24) and not w38519;
w38521 <= not w38022 and not w38394;
w38522 <= not w38032 and w38316;
w38523 <= not w38312 and w38522;
w38524 <= not w38313 and not w38316;
w38525 <= not w38523 and not w38524;
w38526 <= w10273 and not w38525;
w38527 <= not w38393 and w38526;
w38528 <= not w38521 and not w38527;
w38529 <= not b(23) and not w38528;
w38530 <= not w38031 and not w38394;
w38531 <= not w38041 and w38311;
w38532 <= not w38307 and w38531;
w38533 <= not w38308 and not w38311;
w38534 <= not w38532 and not w38533;
w38535 <= w10273 and not w38534;
w38536 <= not w38393 and w38535;
w38537 <= not w38530 and not w38536;
w38538 <= not b(22) and not w38537;
w38539 <= not w38040 and not w38394;
w38540 <= not w38050 and w38306;
w38541 <= not w38302 and w38540;
w38542 <= not w38303 and not w38306;
w38543 <= not w38541 and not w38542;
w38544 <= w10273 and not w38543;
w38545 <= not w38393 and w38544;
w38546 <= not w38539 and not w38545;
w38547 <= not b(21) and not w38546;
w38548 <= not w38049 and not w38394;
w38549 <= not w38059 and w38301;
w38550 <= not w38297 and w38549;
w38551 <= not w38298 and not w38301;
w38552 <= not w38550 and not w38551;
w38553 <= w10273 and not w38552;
w38554 <= not w38393 and w38553;
w38555 <= not w38548 and not w38554;
w38556 <= not b(20) and not w38555;
w38557 <= not w38058 and not w38394;
w38558 <= not w38068 and w38296;
w38559 <= not w38292 and w38558;
w38560 <= not w38293 and not w38296;
w38561 <= not w38559 and not w38560;
w38562 <= w10273 and not w38561;
w38563 <= not w38393 and w38562;
w38564 <= not w38557 and not w38563;
w38565 <= not b(19) and not w38564;
w38566 <= not w38067 and not w38394;
w38567 <= not w38077 and w38291;
w38568 <= not w38287 and w38567;
w38569 <= not w38288 and not w38291;
w38570 <= not w38568 and not w38569;
w38571 <= w10273 and not w38570;
w38572 <= not w38393 and w38571;
w38573 <= not w38566 and not w38572;
w38574 <= not b(18) and not w38573;
w38575 <= not w38076 and not w38394;
w38576 <= not w38086 and w38286;
w38577 <= not w38282 and w38576;
w38578 <= not w38283 and not w38286;
w38579 <= not w38577 and not w38578;
w38580 <= w10273 and not w38579;
w38581 <= not w38393 and w38580;
w38582 <= not w38575 and not w38581;
w38583 <= not b(17) and not w38582;
w38584 <= not w38085 and not w38394;
w38585 <= not w38095 and w38281;
w38586 <= not w38277 and w38585;
w38587 <= not w38278 and not w38281;
w38588 <= not w38586 and not w38587;
w38589 <= w10273 and not w38588;
w38590 <= not w38393 and w38589;
w38591 <= not w38584 and not w38590;
w38592 <= not b(16) and not w38591;
w38593 <= not w38094 and not w38394;
w38594 <= not w38104 and w38276;
w38595 <= not w38272 and w38594;
w38596 <= not w38273 and not w38276;
w38597 <= not w38595 and not w38596;
w38598 <= w10273 and not w38597;
w38599 <= not w38393 and w38598;
w38600 <= not w38593 and not w38599;
w38601 <= not b(15) and not w38600;
w38602 <= not w38103 and not w38394;
w38603 <= not w38113 and w38271;
w38604 <= not w38267 and w38603;
w38605 <= not w38268 and not w38271;
w38606 <= not w38604 and not w38605;
w38607 <= w10273 and not w38606;
w38608 <= not w38393 and w38607;
w38609 <= not w38602 and not w38608;
w38610 <= not b(14) and not w38609;
w38611 <= not w38112 and not w38394;
w38612 <= not w38122 and w38266;
w38613 <= not w38262 and w38612;
w38614 <= not w38263 and not w38266;
w38615 <= not w38613 and not w38614;
w38616 <= w10273 and not w38615;
w38617 <= not w38393 and w38616;
w38618 <= not w38611 and not w38617;
w38619 <= not b(13) and not w38618;
w38620 <= not w38121 and not w38394;
w38621 <= not w38131 and w38261;
w38622 <= not w38257 and w38621;
w38623 <= not w38258 and not w38261;
w38624 <= not w38622 and not w38623;
w38625 <= w10273 and not w38624;
w38626 <= not w38393 and w38625;
w38627 <= not w38620 and not w38626;
w38628 <= not b(12) and not w38627;
w38629 <= not w38130 and not w38394;
w38630 <= not w38140 and w38256;
w38631 <= not w38252 and w38630;
w38632 <= not w38253 and not w38256;
w38633 <= not w38631 and not w38632;
w38634 <= w10273 and not w38633;
w38635 <= not w38393 and w38634;
w38636 <= not w38629 and not w38635;
w38637 <= not b(11) and not w38636;
w38638 <= not w38139 and not w38394;
w38639 <= not w38149 and w38251;
w38640 <= not w38247 and w38639;
w38641 <= not w38248 and not w38251;
w38642 <= not w38640 and not w38641;
w38643 <= w10273 and not w38642;
w38644 <= not w38393 and w38643;
w38645 <= not w38638 and not w38644;
w38646 <= not b(10) and not w38645;
w38647 <= not w38148 and not w38394;
w38648 <= not w38158 and w38246;
w38649 <= not w38242 and w38648;
w38650 <= not w38243 and not w38246;
w38651 <= not w38649 and not w38650;
w38652 <= w10273 and not w38651;
w38653 <= not w38393 and w38652;
w38654 <= not w38647 and not w38653;
w38655 <= not b(9) and not w38654;
w38656 <= not w38157 and not w38394;
w38657 <= not w38167 and w38241;
w38658 <= not w38237 and w38657;
w38659 <= not w38238 and not w38241;
w38660 <= not w38658 and not w38659;
w38661 <= w10273 and not w38660;
w38662 <= not w38393 and w38661;
w38663 <= not w38656 and not w38662;
w38664 <= not b(8) and not w38663;
w38665 <= not w38166 and not w38394;
w38666 <= not w38176 and w38236;
w38667 <= not w38232 and w38666;
w38668 <= not w38233 and not w38236;
w38669 <= not w38667 and not w38668;
w38670 <= w10273 and not w38669;
w38671 <= not w38393 and w38670;
w38672 <= not w38665 and not w38671;
w38673 <= not b(7) and not w38672;
w38674 <= not w38175 and not w38394;
w38675 <= not w38185 and w38231;
w38676 <= not w38227 and w38675;
w38677 <= not w38228 and not w38231;
w38678 <= not w38676 and not w38677;
w38679 <= w10273 and not w38678;
w38680 <= not w38393 and w38679;
w38681 <= not w38674 and not w38680;
w38682 <= not b(6) and not w38681;
w38683 <= not w38184 and not w38394;
w38684 <= not w38194 and w38226;
w38685 <= not w38222 and w38684;
w38686 <= not w38223 and not w38226;
w38687 <= not w38685 and not w38686;
w38688 <= w10273 and not w38687;
w38689 <= not w38393 and w38688;
w38690 <= not w38683 and not w38689;
w38691 <= not b(5) and not w38690;
w38692 <= not w38193 and not w38394;
w38693 <= not w38202 and w38221;
w38694 <= not w38217 and w38693;
w38695 <= not w38218 and not w38221;
w38696 <= not w38694 and not w38695;
w38697 <= w10273 and not w38696;
w38698 <= not w38393 and w38697;
w38699 <= not w38692 and not w38698;
w38700 <= not b(4) and not w38699;
w38701 <= not w38201 and not w38394;
w38702 <= not w38212 and w38216;
w38703 <= not w38211 and w38702;
w38704 <= not w38213 and not w38216;
w38705 <= not w38703 and not w38704;
w38706 <= w10273 and not w38705;
w38707 <= not w38393 and w38706;
w38708 <= not w38701 and not w38707;
w38709 <= not b(3) and not w38708;
w38710 <= not w38206 and not w38394;
w38711 <= w10087 and not w38209;
w38712 <= not w38207 and w38711;
w38713 <= w10273 and not w38712;
w38714 <= not w38211 and w38713;
w38715 <= not w38393 and w38714;
w38716 <= not w38710 and not w38715;
w38717 <= not b(2) and not w38716;
w38718 <= w10602 and not w38393;
w38719 <= a(26) and not w38718;
w38720 <= w10608 and not w38393;
w38721 <= not w38719 and not w38720;
w38722 <= b(1) and not w38721;
w38723 <= not b(1) and not w38720;
w38724 <= not w38719 and w38723;
w38725 <= not w38722 and not w38724;
w38726 <= not w10615 and not w38725;
w38727 <= not b(1) and not w38721;
w38728 <= not w38726 and not w38727;
w38729 <= b(2) and not w38715;
w38730 <= not w38710 and w38729;
w38731 <= not w38717 and not w38730;
w38732 <= not w38728 and w38731;
w38733 <= not w38717 and not w38732;
w38734 <= b(3) and not w38707;
w38735 <= not w38701 and w38734;
w38736 <= not w38709 and not w38735;
w38737 <= not w38733 and w38736;
w38738 <= not w38709 and not w38737;
w38739 <= b(4) and not w38698;
w38740 <= not w38692 and w38739;
w38741 <= not w38700 and not w38740;
w38742 <= not w38738 and w38741;
w38743 <= not w38700 and not w38742;
w38744 <= b(5) and not w38689;
w38745 <= not w38683 and w38744;
w38746 <= not w38691 and not w38745;
w38747 <= not w38743 and w38746;
w38748 <= not w38691 and not w38747;
w38749 <= b(6) and not w38680;
w38750 <= not w38674 and w38749;
w38751 <= not w38682 and not w38750;
w38752 <= not w38748 and w38751;
w38753 <= not w38682 and not w38752;
w38754 <= b(7) and not w38671;
w38755 <= not w38665 and w38754;
w38756 <= not w38673 and not w38755;
w38757 <= not w38753 and w38756;
w38758 <= not w38673 and not w38757;
w38759 <= b(8) and not w38662;
w38760 <= not w38656 and w38759;
w38761 <= not w38664 and not w38760;
w38762 <= not w38758 and w38761;
w38763 <= not w38664 and not w38762;
w38764 <= b(9) and not w38653;
w38765 <= not w38647 and w38764;
w38766 <= not w38655 and not w38765;
w38767 <= not w38763 and w38766;
w38768 <= not w38655 and not w38767;
w38769 <= b(10) and not w38644;
w38770 <= not w38638 and w38769;
w38771 <= not w38646 and not w38770;
w38772 <= not w38768 and w38771;
w38773 <= not w38646 and not w38772;
w38774 <= b(11) and not w38635;
w38775 <= not w38629 and w38774;
w38776 <= not w38637 and not w38775;
w38777 <= not w38773 and w38776;
w38778 <= not w38637 and not w38777;
w38779 <= b(12) and not w38626;
w38780 <= not w38620 and w38779;
w38781 <= not w38628 and not w38780;
w38782 <= not w38778 and w38781;
w38783 <= not w38628 and not w38782;
w38784 <= b(13) and not w38617;
w38785 <= not w38611 and w38784;
w38786 <= not w38619 and not w38785;
w38787 <= not w38783 and w38786;
w38788 <= not w38619 and not w38787;
w38789 <= b(14) and not w38608;
w38790 <= not w38602 and w38789;
w38791 <= not w38610 and not w38790;
w38792 <= not w38788 and w38791;
w38793 <= not w38610 and not w38792;
w38794 <= b(15) and not w38599;
w38795 <= not w38593 and w38794;
w38796 <= not w38601 and not w38795;
w38797 <= not w38793 and w38796;
w38798 <= not w38601 and not w38797;
w38799 <= b(16) and not w38590;
w38800 <= not w38584 and w38799;
w38801 <= not w38592 and not w38800;
w38802 <= not w38798 and w38801;
w38803 <= not w38592 and not w38802;
w38804 <= b(17) and not w38581;
w38805 <= not w38575 and w38804;
w38806 <= not w38583 and not w38805;
w38807 <= not w38803 and w38806;
w38808 <= not w38583 and not w38807;
w38809 <= b(18) and not w38572;
w38810 <= not w38566 and w38809;
w38811 <= not w38574 and not w38810;
w38812 <= not w38808 and w38811;
w38813 <= not w38574 and not w38812;
w38814 <= b(19) and not w38563;
w38815 <= not w38557 and w38814;
w38816 <= not w38565 and not w38815;
w38817 <= not w38813 and w38816;
w38818 <= not w38565 and not w38817;
w38819 <= b(20) and not w38554;
w38820 <= not w38548 and w38819;
w38821 <= not w38556 and not w38820;
w38822 <= not w38818 and w38821;
w38823 <= not w38556 and not w38822;
w38824 <= b(21) and not w38545;
w38825 <= not w38539 and w38824;
w38826 <= not w38547 and not w38825;
w38827 <= not w38823 and w38826;
w38828 <= not w38547 and not w38827;
w38829 <= b(22) and not w38536;
w38830 <= not w38530 and w38829;
w38831 <= not w38538 and not w38830;
w38832 <= not w38828 and w38831;
w38833 <= not w38538 and not w38832;
w38834 <= b(23) and not w38527;
w38835 <= not w38521 and w38834;
w38836 <= not w38529 and not w38835;
w38837 <= not w38833 and w38836;
w38838 <= not w38529 and not w38837;
w38839 <= b(24) and not w38518;
w38840 <= not w38512 and w38839;
w38841 <= not w38520 and not w38840;
w38842 <= not w38838 and w38841;
w38843 <= not w38520 and not w38842;
w38844 <= b(25) and not w38509;
w38845 <= not w38503 and w38844;
w38846 <= not w38511 and not w38845;
w38847 <= not w38843 and w38846;
w38848 <= not w38511 and not w38847;
w38849 <= b(26) and not w38500;
w38850 <= not w38494 and w38849;
w38851 <= not w38502 and not w38850;
w38852 <= not w38848 and w38851;
w38853 <= not w38502 and not w38852;
w38854 <= b(27) and not w38491;
w38855 <= not w38485 and w38854;
w38856 <= not w38493 and not w38855;
w38857 <= not w38853 and w38856;
w38858 <= not w38493 and not w38857;
w38859 <= b(28) and not w38482;
w38860 <= not w38476 and w38859;
w38861 <= not w38484 and not w38860;
w38862 <= not w38858 and w38861;
w38863 <= not w38484 and not w38862;
w38864 <= b(29) and not w38473;
w38865 <= not w38467 and w38864;
w38866 <= not w38475 and not w38865;
w38867 <= not w38863 and w38866;
w38868 <= not w38475 and not w38867;
w38869 <= b(30) and not w38464;
w38870 <= not w38458 and w38869;
w38871 <= not w38466 and not w38870;
w38872 <= not w38868 and w38871;
w38873 <= not w38466 and not w38872;
w38874 <= b(31) and not w38455;
w38875 <= not w38449 and w38874;
w38876 <= not w38457 and not w38875;
w38877 <= not w38873 and w38876;
w38878 <= not w38457 and not w38877;
w38879 <= b(32) and not w38446;
w38880 <= not w38440 and w38879;
w38881 <= not w38448 and not w38880;
w38882 <= not w38878 and w38881;
w38883 <= not w38448 and not w38882;
w38884 <= b(33) and not w38437;
w38885 <= not w38431 and w38884;
w38886 <= not w38439 and not w38885;
w38887 <= not w38883 and w38886;
w38888 <= not w38439 and not w38887;
w38889 <= b(34) and not w38428;
w38890 <= not w38422 and w38889;
w38891 <= not w38430 and not w38890;
w38892 <= not w38888 and w38891;
w38893 <= not w38430 and not w38892;
w38894 <= b(35) and not w38419;
w38895 <= not w38413 and w38894;
w38896 <= not w38421 and not w38895;
w38897 <= not w38893 and w38896;
w38898 <= not w38421 and not w38897;
w38899 <= b(36) and not w38410;
w38900 <= not w38404 and w38899;
w38901 <= not w38412 and not w38900;
w38902 <= not w38898 and w38901;
w38903 <= not w38412 and not w38902;
w38904 <= b(37) and not w38401;
w38905 <= not w38395 and w38904;
w38906 <= not w38403 and not w38905;
w38907 <= not w38903 and w38906;
w38908 <= not w38403 and not w38907;
w38909 <= not w37895 and not w38394;
w38910 <= not w37897 and w38391;
w38911 <= not w38387 and w38910;
w38912 <= not w38388 and not w38391;
w38913 <= not w38911 and not w38912;
w38914 <= w38394 and not w38913;
w38915 <= not w38909 and not w38914;
w38916 <= not b(38) and not w38915;
w38917 <= b(38) and not w38909;
w38918 <= not w38914 and w38917;
w38919 <= w10811 and not w38918;
w38920 <= not w38916 and w38919;
w38921 <= not w38908 and w38920;
w38922 <= w10273 and not w38915;
w38923 <= not w38921 and not w38922;
w38924 <= not w38412 and w38906;
w38925 <= not w38902 and w38924;
w38926 <= not w38903 and not w38906;
w38927 <= not w38925 and not w38926;
w38928 <= not w38923 and not w38927;
w38929 <= not w38402 and not w38922;
w38930 <= not w38921 and w38929;
w38931 <= not w38928 and not w38930;
w38932 <= not w38403 and not w38918;
w38933 <= not w38916 and w38932;
w38934 <= not w38907 and w38933;
w38935 <= not w38916 and not w38918;
w38936 <= not w38908 and not w38935;
w38937 <= not w38934 and not w38936;
w38938 <= not w38923 and not w38937;
w38939 <= not w38915 and not w38922;
w38940 <= not w38921 and w38939;
w38941 <= not w38938 and not w38940;
w38942 <= not b(39) and not w38941;
w38943 <= not b(38) and not w38931;
w38944 <= not w38421 and w38901;
w38945 <= not w38897 and w38944;
w38946 <= not w38898 and not w38901;
w38947 <= not w38945 and not w38946;
w38948 <= not w38923 and not w38947;
w38949 <= not w38411 and not w38922;
w38950 <= not w38921 and w38949;
w38951 <= not w38948 and not w38950;
w38952 <= not b(37) and not w38951;
w38953 <= not w38430 and w38896;
w38954 <= not w38892 and w38953;
w38955 <= not w38893 and not w38896;
w38956 <= not w38954 and not w38955;
w38957 <= not w38923 and not w38956;
w38958 <= not w38420 and not w38922;
w38959 <= not w38921 and w38958;
w38960 <= not w38957 and not w38959;
w38961 <= not b(36) and not w38960;
w38962 <= not w38439 and w38891;
w38963 <= not w38887 and w38962;
w38964 <= not w38888 and not w38891;
w38965 <= not w38963 and not w38964;
w38966 <= not w38923 and not w38965;
w38967 <= not w38429 and not w38922;
w38968 <= not w38921 and w38967;
w38969 <= not w38966 and not w38968;
w38970 <= not b(35) and not w38969;
w38971 <= not w38448 and w38886;
w38972 <= not w38882 and w38971;
w38973 <= not w38883 and not w38886;
w38974 <= not w38972 and not w38973;
w38975 <= not w38923 and not w38974;
w38976 <= not w38438 and not w38922;
w38977 <= not w38921 and w38976;
w38978 <= not w38975 and not w38977;
w38979 <= not b(34) and not w38978;
w38980 <= not w38457 and w38881;
w38981 <= not w38877 and w38980;
w38982 <= not w38878 and not w38881;
w38983 <= not w38981 and not w38982;
w38984 <= not w38923 and not w38983;
w38985 <= not w38447 and not w38922;
w38986 <= not w38921 and w38985;
w38987 <= not w38984 and not w38986;
w38988 <= not b(33) and not w38987;
w38989 <= not w38466 and w38876;
w38990 <= not w38872 and w38989;
w38991 <= not w38873 and not w38876;
w38992 <= not w38990 and not w38991;
w38993 <= not w38923 and not w38992;
w38994 <= not w38456 and not w38922;
w38995 <= not w38921 and w38994;
w38996 <= not w38993 and not w38995;
w38997 <= not b(32) and not w38996;
w38998 <= not w38475 and w38871;
w38999 <= not w38867 and w38998;
w39000 <= not w38868 and not w38871;
w39001 <= not w38999 and not w39000;
w39002 <= not w38923 and not w39001;
w39003 <= not w38465 and not w38922;
w39004 <= not w38921 and w39003;
w39005 <= not w39002 and not w39004;
w39006 <= not b(31) and not w39005;
w39007 <= not w38484 and w38866;
w39008 <= not w38862 and w39007;
w39009 <= not w38863 and not w38866;
w39010 <= not w39008 and not w39009;
w39011 <= not w38923 and not w39010;
w39012 <= not w38474 and not w38922;
w39013 <= not w38921 and w39012;
w39014 <= not w39011 and not w39013;
w39015 <= not b(30) and not w39014;
w39016 <= not w38493 and w38861;
w39017 <= not w38857 and w39016;
w39018 <= not w38858 and not w38861;
w39019 <= not w39017 and not w39018;
w39020 <= not w38923 and not w39019;
w39021 <= not w38483 and not w38922;
w39022 <= not w38921 and w39021;
w39023 <= not w39020 and not w39022;
w39024 <= not b(29) and not w39023;
w39025 <= not w38502 and w38856;
w39026 <= not w38852 and w39025;
w39027 <= not w38853 and not w38856;
w39028 <= not w39026 and not w39027;
w39029 <= not w38923 and not w39028;
w39030 <= not w38492 and not w38922;
w39031 <= not w38921 and w39030;
w39032 <= not w39029 and not w39031;
w39033 <= not b(28) and not w39032;
w39034 <= not w38511 and w38851;
w39035 <= not w38847 and w39034;
w39036 <= not w38848 and not w38851;
w39037 <= not w39035 and not w39036;
w39038 <= not w38923 and not w39037;
w39039 <= not w38501 and not w38922;
w39040 <= not w38921 and w39039;
w39041 <= not w39038 and not w39040;
w39042 <= not b(27) and not w39041;
w39043 <= not w38520 and w38846;
w39044 <= not w38842 and w39043;
w39045 <= not w38843 and not w38846;
w39046 <= not w39044 and not w39045;
w39047 <= not w38923 and not w39046;
w39048 <= not w38510 and not w38922;
w39049 <= not w38921 and w39048;
w39050 <= not w39047 and not w39049;
w39051 <= not b(26) and not w39050;
w39052 <= not w38529 and w38841;
w39053 <= not w38837 and w39052;
w39054 <= not w38838 and not w38841;
w39055 <= not w39053 and not w39054;
w39056 <= not w38923 and not w39055;
w39057 <= not w38519 and not w38922;
w39058 <= not w38921 and w39057;
w39059 <= not w39056 and not w39058;
w39060 <= not b(25) and not w39059;
w39061 <= not w38538 and w38836;
w39062 <= not w38832 and w39061;
w39063 <= not w38833 and not w38836;
w39064 <= not w39062 and not w39063;
w39065 <= not w38923 and not w39064;
w39066 <= not w38528 and not w38922;
w39067 <= not w38921 and w39066;
w39068 <= not w39065 and not w39067;
w39069 <= not b(24) and not w39068;
w39070 <= not w38547 and w38831;
w39071 <= not w38827 and w39070;
w39072 <= not w38828 and not w38831;
w39073 <= not w39071 and not w39072;
w39074 <= not w38923 and not w39073;
w39075 <= not w38537 and not w38922;
w39076 <= not w38921 and w39075;
w39077 <= not w39074 and not w39076;
w39078 <= not b(23) and not w39077;
w39079 <= not w38556 and w38826;
w39080 <= not w38822 and w39079;
w39081 <= not w38823 and not w38826;
w39082 <= not w39080 and not w39081;
w39083 <= not w38923 and not w39082;
w39084 <= not w38546 and not w38922;
w39085 <= not w38921 and w39084;
w39086 <= not w39083 and not w39085;
w39087 <= not b(22) and not w39086;
w39088 <= not w38565 and w38821;
w39089 <= not w38817 and w39088;
w39090 <= not w38818 and not w38821;
w39091 <= not w39089 and not w39090;
w39092 <= not w38923 and not w39091;
w39093 <= not w38555 and not w38922;
w39094 <= not w38921 and w39093;
w39095 <= not w39092 and not w39094;
w39096 <= not b(21) and not w39095;
w39097 <= not w38574 and w38816;
w39098 <= not w38812 and w39097;
w39099 <= not w38813 and not w38816;
w39100 <= not w39098 and not w39099;
w39101 <= not w38923 and not w39100;
w39102 <= not w38564 and not w38922;
w39103 <= not w38921 and w39102;
w39104 <= not w39101 and not w39103;
w39105 <= not b(20) and not w39104;
w39106 <= not w38583 and w38811;
w39107 <= not w38807 and w39106;
w39108 <= not w38808 and not w38811;
w39109 <= not w39107 and not w39108;
w39110 <= not w38923 and not w39109;
w39111 <= not w38573 and not w38922;
w39112 <= not w38921 and w39111;
w39113 <= not w39110 and not w39112;
w39114 <= not b(19) and not w39113;
w39115 <= not w38592 and w38806;
w39116 <= not w38802 and w39115;
w39117 <= not w38803 and not w38806;
w39118 <= not w39116 and not w39117;
w39119 <= not w38923 and not w39118;
w39120 <= not w38582 and not w38922;
w39121 <= not w38921 and w39120;
w39122 <= not w39119 and not w39121;
w39123 <= not b(18) and not w39122;
w39124 <= not w38601 and w38801;
w39125 <= not w38797 and w39124;
w39126 <= not w38798 and not w38801;
w39127 <= not w39125 and not w39126;
w39128 <= not w38923 and not w39127;
w39129 <= not w38591 and not w38922;
w39130 <= not w38921 and w39129;
w39131 <= not w39128 and not w39130;
w39132 <= not b(17) and not w39131;
w39133 <= not w38610 and w38796;
w39134 <= not w38792 and w39133;
w39135 <= not w38793 and not w38796;
w39136 <= not w39134 and not w39135;
w39137 <= not w38923 and not w39136;
w39138 <= not w38600 and not w38922;
w39139 <= not w38921 and w39138;
w39140 <= not w39137 and not w39139;
w39141 <= not b(16) and not w39140;
w39142 <= not w38619 and w38791;
w39143 <= not w38787 and w39142;
w39144 <= not w38788 and not w38791;
w39145 <= not w39143 and not w39144;
w39146 <= not w38923 and not w39145;
w39147 <= not w38609 and not w38922;
w39148 <= not w38921 and w39147;
w39149 <= not w39146 and not w39148;
w39150 <= not b(15) and not w39149;
w39151 <= not w38628 and w38786;
w39152 <= not w38782 and w39151;
w39153 <= not w38783 and not w38786;
w39154 <= not w39152 and not w39153;
w39155 <= not w38923 and not w39154;
w39156 <= not w38618 and not w38922;
w39157 <= not w38921 and w39156;
w39158 <= not w39155 and not w39157;
w39159 <= not b(14) and not w39158;
w39160 <= not w38637 and w38781;
w39161 <= not w38777 and w39160;
w39162 <= not w38778 and not w38781;
w39163 <= not w39161 and not w39162;
w39164 <= not w38923 and not w39163;
w39165 <= not w38627 and not w38922;
w39166 <= not w38921 and w39165;
w39167 <= not w39164 and not w39166;
w39168 <= not b(13) and not w39167;
w39169 <= not w38646 and w38776;
w39170 <= not w38772 and w39169;
w39171 <= not w38773 and not w38776;
w39172 <= not w39170 and not w39171;
w39173 <= not w38923 and not w39172;
w39174 <= not w38636 and not w38922;
w39175 <= not w38921 and w39174;
w39176 <= not w39173 and not w39175;
w39177 <= not b(12) and not w39176;
w39178 <= not w38655 and w38771;
w39179 <= not w38767 and w39178;
w39180 <= not w38768 and not w38771;
w39181 <= not w39179 and not w39180;
w39182 <= not w38923 and not w39181;
w39183 <= not w38645 and not w38922;
w39184 <= not w38921 and w39183;
w39185 <= not w39182 and not w39184;
w39186 <= not b(11) and not w39185;
w39187 <= not w38664 and w38766;
w39188 <= not w38762 and w39187;
w39189 <= not w38763 and not w38766;
w39190 <= not w39188 and not w39189;
w39191 <= not w38923 and not w39190;
w39192 <= not w38654 and not w38922;
w39193 <= not w38921 and w39192;
w39194 <= not w39191 and not w39193;
w39195 <= not b(10) and not w39194;
w39196 <= not w38673 and w38761;
w39197 <= not w38757 and w39196;
w39198 <= not w38758 and not w38761;
w39199 <= not w39197 and not w39198;
w39200 <= not w38923 and not w39199;
w39201 <= not w38663 and not w38922;
w39202 <= not w38921 and w39201;
w39203 <= not w39200 and not w39202;
w39204 <= not b(9) and not w39203;
w39205 <= not w38682 and w38756;
w39206 <= not w38752 and w39205;
w39207 <= not w38753 and not w38756;
w39208 <= not w39206 and not w39207;
w39209 <= not w38923 and not w39208;
w39210 <= not w38672 and not w38922;
w39211 <= not w38921 and w39210;
w39212 <= not w39209 and not w39211;
w39213 <= not b(8) and not w39212;
w39214 <= not w38691 and w38751;
w39215 <= not w38747 and w39214;
w39216 <= not w38748 and not w38751;
w39217 <= not w39215 and not w39216;
w39218 <= not w38923 and not w39217;
w39219 <= not w38681 and not w38922;
w39220 <= not w38921 and w39219;
w39221 <= not w39218 and not w39220;
w39222 <= not b(7) and not w39221;
w39223 <= not w38700 and w38746;
w39224 <= not w38742 and w39223;
w39225 <= not w38743 and not w38746;
w39226 <= not w39224 and not w39225;
w39227 <= not w38923 and not w39226;
w39228 <= not w38690 and not w38922;
w39229 <= not w38921 and w39228;
w39230 <= not w39227 and not w39229;
w39231 <= not b(6) and not w39230;
w39232 <= not w38709 and w38741;
w39233 <= not w38737 and w39232;
w39234 <= not w38738 and not w38741;
w39235 <= not w39233 and not w39234;
w39236 <= not w38923 and not w39235;
w39237 <= not w38699 and not w38922;
w39238 <= not w38921 and w39237;
w39239 <= not w39236 and not w39238;
w39240 <= not b(5) and not w39239;
w39241 <= not w38717 and w38736;
w39242 <= not w38732 and w39241;
w39243 <= not w38733 and not w38736;
w39244 <= not w39242 and not w39243;
w39245 <= not w38923 and not w39244;
w39246 <= not w38708 and not w38922;
w39247 <= not w38921 and w39246;
w39248 <= not w39245 and not w39247;
w39249 <= not b(4) and not w39248;
w39250 <= not w38727 and w38731;
w39251 <= not w38726 and w39250;
w39252 <= not w38728 and not w38731;
w39253 <= not w39251 and not w39252;
w39254 <= not w38923 and not w39253;
w39255 <= not w38716 and not w38922;
w39256 <= not w38921 and w39255;
w39257 <= not w39254 and not w39256;
w39258 <= not b(3) and not w39257;
w39259 <= w10615 and not w38724;
w39260 <= not w38722 and w39259;
w39261 <= not w38726 and not w39260;
w39262 <= not w38923 and w39261;
w39263 <= not w38721 and not w38922;
w39264 <= not w38921 and w39263;
w39265 <= not w39262 and not w39264;
w39266 <= not b(2) and not w39265;
w39267 <= b(0) and not w38923;
w39268 <= a(25) and not w39267;
w39269 <= w10615 and not w38923;
w39270 <= not w39268 and not w39269;
w39271 <= b(1) and not w39270;
w39272 <= not b(1) and not w39269;
w39273 <= not w39268 and w39272;
w39274 <= not w39271 and not w39273;
w39275 <= not w11168 and not w39274;
w39276 <= not b(1) and not w39270;
w39277 <= not w39275 and not w39276;
w39278 <= b(2) and not w39264;
w39279 <= not w39262 and w39278;
w39280 <= not w39266 and not w39279;
w39281 <= not w39277 and w39280;
w39282 <= not w39266 and not w39281;
w39283 <= b(3) and not w39256;
w39284 <= not w39254 and w39283;
w39285 <= not w39258 and not w39284;
w39286 <= not w39282 and w39285;
w39287 <= not w39258 and not w39286;
w39288 <= b(4) and not w39247;
w39289 <= not w39245 and w39288;
w39290 <= not w39249 and not w39289;
w39291 <= not w39287 and w39290;
w39292 <= not w39249 and not w39291;
w39293 <= b(5) and not w39238;
w39294 <= not w39236 and w39293;
w39295 <= not w39240 and not w39294;
w39296 <= not w39292 and w39295;
w39297 <= not w39240 and not w39296;
w39298 <= b(6) and not w39229;
w39299 <= not w39227 and w39298;
w39300 <= not w39231 and not w39299;
w39301 <= not w39297 and w39300;
w39302 <= not w39231 and not w39301;
w39303 <= b(7) and not w39220;
w39304 <= not w39218 and w39303;
w39305 <= not w39222 and not w39304;
w39306 <= not w39302 and w39305;
w39307 <= not w39222 and not w39306;
w39308 <= b(8) and not w39211;
w39309 <= not w39209 and w39308;
w39310 <= not w39213 and not w39309;
w39311 <= not w39307 and w39310;
w39312 <= not w39213 and not w39311;
w39313 <= b(9) and not w39202;
w39314 <= not w39200 and w39313;
w39315 <= not w39204 and not w39314;
w39316 <= not w39312 and w39315;
w39317 <= not w39204 and not w39316;
w39318 <= b(10) and not w39193;
w39319 <= not w39191 and w39318;
w39320 <= not w39195 and not w39319;
w39321 <= not w39317 and w39320;
w39322 <= not w39195 and not w39321;
w39323 <= b(11) and not w39184;
w39324 <= not w39182 and w39323;
w39325 <= not w39186 and not w39324;
w39326 <= not w39322 and w39325;
w39327 <= not w39186 and not w39326;
w39328 <= b(12) and not w39175;
w39329 <= not w39173 and w39328;
w39330 <= not w39177 and not w39329;
w39331 <= not w39327 and w39330;
w39332 <= not w39177 and not w39331;
w39333 <= b(13) and not w39166;
w39334 <= not w39164 and w39333;
w39335 <= not w39168 and not w39334;
w39336 <= not w39332 and w39335;
w39337 <= not w39168 and not w39336;
w39338 <= b(14) and not w39157;
w39339 <= not w39155 and w39338;
w39340 <= not w39159 and not w39339;
w39341 <= not w39337 and w39340;
w39342 <= not w39159 and not w39341;
w39343 <= b(15) and not w39148;
w39344 <= not w39146 and w39343;
w39345 <= not w39150 and not w39344;
w39346 <= not w39342 and w39345;
w39347 <= not w39150 and not w39346;
w39348 <= b(16) and not w39139;
w39349 <= not w39137 and w39348;
w39350 <= not w39141 and not w39349;
w39351 <= not w39347 and w39350;
w39352 <= not w39141 and not w39351;
w39353 <= b(17) and not w39130;
w39354 <= not w39128 and w39353;
w39355 <= not w39132 and not w39354;
w39356 <= not w39352 and w39355;
w39357 <= not w39132 and not w39356;
w39358 <= b(18) and not w39121;
w39359 <= not w39119 and w39358;
w39360 <= not w39123 and not w39359;
w39361 <= not w39357 and w39360;
w39362 <= not w39123 and not w39361;
w39363 <= b(19) and not w39112;
w39364 <= not w39110 and w39363;
w39365 <= not w39114 and not w39364;
w39366 <= not w39362 and w39365;
w39367 <= not w39114 and not w39366;
w39368 <= b(20) and not w39103;
w39369 <= not w39101 and w39368;
w39370 <= not w39105 and not w39369;
w39371 <= not w39367 and w39370;
w39372 <= not w39105 and not w39371;
w39373 <= b(21) and not w39094;
w39374 <= not w39092 and w39373;
w39375 <= not w39096 and not w39374;
w39376 <= not w39372 and w39375;
w39377 <= not w39096 and not w39376;
w39378 <= b(22) and not w39085;
w39379 <= not w39083 and w39378;
w39380 <= not w39087 and not w39379;
w39381 <= not w39377 and w39380;
w39382 <= not w39087 and not w39381;
w39383 <= b(23) and not w39076;
w39384 <= not w39074 and w39383;
w39385 <= not w39078 and not w39384;
w39386 <= not w39382 and w39385;
w39387 <= not w39078 and not w39386;
w39388 <= b(24) and not w39067;
w39389 <= not w39065 and w39388;
w39390 <= not w39069 and not w39389;
w39391 <= not w39387 and w39390;
w39392 <= not w39069 and not w39391;
w39393 <= b(25) and not w39058;
w39394 <= not w39056 and w39393;
w39395 <= not w39060 and not w39394;
w39396 <= not w39392 and w39395;
w39397 <= not w39060 and not w39396;
w39398 <= b(26) and not w39049;
w39399 <= not w39047 and w39398;
w39400 <= not w39051 and not w39399;
w39401 <= not w39397 and w39400;
w39402 <= not w39051 and not w39401;
w39403 <= b(27) and not w39040;
w39404 <= not w39038 and w39403;
w39405 <= not w39042 and not w39404;
w39406 <= not w39402 and w39405;
w39407 <= not w39042 and not w39406;
w39408 <= b(28) and not w39031;
w39409 <= not w39029 and w39408;
w39410 <= not w39033 and not w39409;
w39411 <= not w39407 and w39410;
w39412 <= not w39033 and not w39411;
w39413 <= b(29) and not w39022;
w39414 <= not w39020 and w39413;
w39415 <= not w39024 and not w39414;
w39416 <= not w39412 and w39415;
w39417 <= not w39024 and not w39416;
w39418 <= b(30) and not w39013;
w39419 <= not w39011 and w39418;
w39420 <= not w39015 and not w39419;
w39421 <= not w39417 and w39420;
w39422 <= not w39015 and not w39421;
w39423 <= b(31) and not w39004;
w39424 <= not w39002 and w39423;
w39425 <= not w39006 and not w39424;
w39426 <= not w39422 and w39425;
w39427 <= not w39006 and not w39426;
w39428 <= b(32) and not w38995;
w39429 <= not w38993 and w39428;
w39430 <= not w38997 and not w39429;
w39431 <= not w39427 and w39430;
w39432 <= not w38997 and not w39431;
w39433 <= b(33) and not w38986;
w39434 <= not w38984 and w39433;
w39435 <= not w38988 and not w39434;
w39436 <= not w39432 and w39435;
w39437 <= not w38988 and not w39436;
w39438 <= b(34) and not w38977;
w39439 <= not w38975 and w39438;
w39440 <= not w38979 and not w39439;
w39441 <= not w39437 and w39440;
w39442 <= not w38979 and not w39441;
w39443 <= b(35) and not w38968;
w39444 <= not w38966 and w39443;
w39445 <= not w38970 and not w39444;
w39446 <= not w39442 and w39445;
w39447 <= not w38970 and not w39446;
w39448 <= b(36) and not w38959;
w39449 <= not w38957 and w39448;
w39450 <= not w38961 and not w39449;
w39451 <= not w39447 and w39450;
w39452 <= not w38961 and not w39451;
w39453 <= b(37) and not w38950;
w39454 <= not w38948 and w39453;
w39455 <= not w38952 and not w39454;
w39456 <= not w39452 and w39455;
w39457 <= not w38952 and not w39456;
w39458 <= b(38) and not w38930;
w39459 <= not w38928 and w39458;
w39460 <= not w38943 and not w39459;
w39461 <= not w39457 and w39460;
w39462 <= not w38943 and not w39461;
w39463 <= b(39) and not w38940;
w39464 <= not w38938 and w39463;
w39465 <= not w38942 and not w39464;
w39466 <= not w39462 and w39465;
w39467 <= not w38942 and not w39466;
w39468 <= w11362 and not w39467;
w39469 <= not w38931 and not w39468;
w39470 <= not w38952 and w39460;
w39471 <= not w39456 and w39470;
w39472 <= not w39457 and not w39460;
w39473 <= not w39471 and not w39472;
w39474 <= w11362 and not w39473;
w39475 <= not w39467 and w39474;
w39476 <= not w39469 and not w39475;
w39477 <= not w38941 and not w39468;
w39478 <= not w38943 and w39465;
w39479 <= not w39461 and w39478;
w39480 <= not w39462 and not w39465;
w39481 <= not w39479 and not w39480;
w39482 <= w39468 and not w39481;
w39483 <= not w39477 and not w39482;
w39484 <= not b(40) and not w39483;
w39485 <= not b(39) and not w39476;
w39486 <= not w38951 and not w39468;
w39487 <= not w38961 and w39455;
w39488 <= not w39451 and w39487;
w39489 <= not w39452 and not w39455;
w39490 <= not w39488 and not w39489;
w39491 <= w11362 and not w39490;
w39492 <= not w39467 and w39491;
w39493 <= not w39486 and not w39492;
w39494 <= not b(38) and not w39493;
w39495 <= not w38960 and not w39468;
w39496 <= not w38970 and w39450;
w39497 <= not w39446 and w39496;
w39498 <= not w39447 and not w39450;
w39499 <= not w39497 and not w39498;
w39500 <= w11362 and not w39499;
w39501 <= not w39467 and w39500;
w39502 <= not w39495 and not w39501;
w39503 <= not b(37) and not w39502;
w39504 <= not w38969 and not w39468;
w39505 <= not w38979 and w39445;
w39506 <= not w39441 and w39505;
w39507 <= not w39442 and not w39445;
w39508 <= not w39506 and not w39507;
w39509 <= w11362 and not w39508;
w39510 <= not w39467 and w39509;
w39511 <= not w39504 and not w39510;
w39512 <= not b(36) and not w39511;
w39513 <= not w38978 and not w39468;
w39514 <= not w38988 and w39440;
w39515 <= not w39436 and w39514;
w39516 <= not w39437 and not w39440;
w39517 <= not w39515 and not w39516;
w39518 <= w11362 and not w39517;
w39519 <= not w39467 and w39518;
w39520 <= not w39513 and not w39519;
w39521 <= not b(35) and not w39520;
w39522 <= not w38987 and not w39468;
w39523 <= not w38997 and w39435;
w39524 <= not w39431 and w39523;
w39525 <= not w39432 and not w39435;
w39526 <= not w39524 and not w39525;
w39527 <= w11362 and not w39526;
w39528 <= not w39467 and w39527;
w39529 <= not w39522 and not w39528;
w39530 <= not b(34) and not w39529;
w39531 <= not w38996 and not w39468;
w39532 <= not w39006 and w39430;
w39533 <= not w39426 and w39532;
w39534 <= not w39427 and not w39430;
w39535 <= not w39533 and not w39534;
w39536 <= w11362 and not w39535;
w39537 <= not w39467 and w39536;
w39538 <= not w39531 and not w39537;
w39539 <= not b(33) and not w39538;
w39540 <= not w39005 and not w39468;
w39541 <= not w39015 and w39425;
w39542 <= not w39421 and w39541;
w39543 <= not w39422 and not w39425;
w39544 <= not w39542 and not w39543;
w39545 <= w11362 and not w39544;
w39546 <= not w39467 and w39545;
w39547 <= not w39540 and not w39546;
w39548 <= not b(32) and not w39547;
w39549 <= not w39014 and not w39468;
w39550 <= not w39024 and w39420;
w39551 <= not w39416 and w39550;
w39552 <= not w39417 and not w39420;
w39553 <= not w39551 and not w39552;
w39554 <= w11362 and not w39553;
w39555 <= not w39467 and w39554;
w39556 <= not w39549 and not w39555;
w39557 <= not b(31) and not w39556;
w39558 <= not w39023 and not w39468;
w39559 <= not w39033 and w39415;
w39560 <= not w39411 and w39559;
w39561 <= not w39412 and not w39415;
w39562 <= not w39560 and not w39561;
w39563 <= w11362 and not w39562;
w39564 <= not w39467 and w39563;
w39565 <= not w39558 and not w39564;
w39566 <= not b(30) and not w39565;
w39567 <= not w39032 and not w39468;
w39568 <= not w39042 and w39410;
w39569 <= not w39406 and w39568;
w39570 <= not w39407 and not w39410;
w39571 <= not w39569 and not w39570;
w39572 <= w11362 and not w39571;
w39573 <= not w39467 and w39572;
w39574 <= not w39567 and not w39573;
w39575 <= not b(29) and not w39574;
w39576 <= not w39041 and not w39468;
w39577 <= not w39051 and w39405;
w39578 <= not w39401 and w39577;
w39579 <= not w39402 and not w39405;
w39580 <= not w39578 and not w39579;
w39581 <= w11362 and not w39580;
w39582 <= not w39467 and w39581;
w39583 <= not w39576 and not w39582;
w39584 <= not b(28) and not w39583;
w39585 <= not w39050 and not w39468;
w39586 <= not w39060 and w39400;
w39587 <= not w39396 and w39586;
w39588 <= not w39397 and not w39400;
w39589 <= not w39587 and not w39588;
w39590 <= w11362 and not w39589;
w39591 <= not w39467 and w39590;
w39592 <= not w39585 and not w39591;
w39593 <= not b(27) and not w39592;
w39594 <= not w39059 and not w39468;
w39595 <= not w39069 and w39395;
w39596 <= not w39391 and w39595;
w39597 <= not w39392 and not w39395;
w39598 <= not w39596 and not w39597;
w39599 <= w11362 and not w39598;
w39600 <= not w39467 and w39599;
w39601 <= not w39594 and not w39600;
w39602 <= not b(26) and not w39601;
w39603 <= not w39068 and not w39468;
w39604 <= not w39078 and w39390;
w39605 <= not w39386 and w39604;
w39606 <= not w39387 and not w39390;
w39607 <= not w39605 and not w39606;
w39608 <= w11362 and not w39607;
w39609 <= not w39467 and w39608;
w39610 <= not w39603 and not w39609;
w39611 <= not b(25) and not w39610;
w39612 <= not w39077 and not w39468;
w39613 <= not w39087 and w39385;
w39614 <= not w39381 and w39613;
w39615 <= not w39382 and not w39385;
w39616 <= not w39614 and not w39615;
w39617 <= w11362 and not w39616;
w39618 <= not w39467 and w39617;
w39619 <= not w39612 and not w39618;
w39620 <= not b(24) and not w39619;
w39621 <= not w39086 and not w39468;
w39622 <= not w39096 and w39380;
w39623 <= not w39376 and w39622;
w39624 <= not w39377 and not w39380;
w39625 <= not w39623 and not w39624;
w39626 <= w11362 and not w39625;
w39627 <= not w39467 and w39626;
w39628 <= not w39621 and not w39627;
w39629 <= not b(23) and not w39628;
w39630 <= not w39095 and not w39468;
w39631 <= not w39105 and w39375;
w39632 <= not w39371 and w39631;
w39633 <= not w39372 and not w39375;
w39634 <= not w39632 and not w39633;
w39635 <= w11362 and not w39634;
w39636 <= not w39467 and w39635;
w39637 <= not w39630 and not w39636;
w39638 <= not b(22) and not w39637;
w39639 <= not w39104 and not w39468;
w39640 <= not w39114 and w39370;
w39641 <= not w39366 and w39640;
w39642 <= not w39367 and not w39370;
w39643 <= not w39641 and not w39642;
w39644 <= w11362 and not w39643;
w39645 <= not w39467 and w39644;
w39646 <= not w39639 and not w39645;
w39647 <= not b(21) and not w39646;
w39648 <= not w39113 and not w39468;
w39649 <= not w39123 and w39365;
w39650 <= not w39361 and w39649;
w39651 <= not w39362 and not w39365;
w39652 <= not w39650 and not w39651;
w39653 <= w11362 and not w39652;
w39654 <= not w39467 and w39653;
w39655 <= not w39648 and not w39654;
w39656 <= not b(20) and not w39655;
w39657 <= not w39122 and not w39468;
w39658 <= not w39132 and w39360;
w39659 <= not w39356 and w39658;
w39660 <= not w39357 and not w39360;
w39661 <= not w39659 and not w39660;
w39662 <= w11362 and not w39661;
w39663 <= not w39467 and w39662;
w39664 <= not w39657 and not w39663;
w39665 <= not b(19) and not w39664;
w39666 <= not w39131 and not w39468;
w39667 <= not w39141 and w39355;
w39668 <= not w39351 and w39667;
w39669 <= not w39352 and not w39355;
w39670 <= not w39668 and not w39669;
w39671 <= w11362 and not w39670;
w39672 <= not w39467 and w39671;
w39673 <= not w39666 and not w39672;
w39674 <= not b(18) and not w39673;
w39675 <= not w39140 and not w39468;
w39676 <= not w39150 and w39350;
w39677 <= not w39346 and w39676;
w39678 <= not w39347 and not w39350;
w39679 <= not w39677 and not w39678;
w39680 <= w11362 and not w39679;
w39681 <= not w39467 and w39680;
w39682 <= not w39675 and not w39681;
w39683 <= not b(17) and not w39682;
w39684 <= not w39149 and not w39468;
w39685 <= not w39159 and w39345;
w39686 <= not w39341 and w39685;
w39687 <= not w39342 and not w39345;
w39688 <= not w39686 and not w39687;
w39689 <= w11362 and not w39688;
w39690 <= not w39467 and w39689;
w39691 <= not w39684 and not w39690;
w39692 <= not b(16) and not w39691;
w39693 <= not w39158 and not w39468;
w39694 <= not w39168 and w39340;
w39695 <= not w39336 and w39694;
w39696 <= not w39337 and not w39340;
w39697 <= not w39695 and not w39696;
w39698 <= w11362 and not w39697;
w39699 <= not w39467 and w39698;
w39700 <= not w39693 and not w39699;
w39701 <= not b(15) and not w39700;
w39702 <= not w39167 and not w39468;
w39703 <= not w39177 and w39335;
w39704 <= not w39331 and w39703;
w39705 <= not w39332 and not w39335;
w39706 <= not w39704 and not w39705;
w39707 <= w11362 and not w39706;
w39708 <= not w39467 and w39707;
w39709 <= not w39702 and not w39708;
w39710 <= not b(14) and not w39709;
w39711 <= not w39176 and not w39468;
w39712 <= not w39186 and w39330;
w39713 <= not w39326 and w39712;
w39714 <= not w39327 and not w39330;
w39715 <= not w39713 and not w39714;
w39716 <= w11362 and not w39715;
w39717 <= not w39467 and w39716;
w39718 <= not w39711 and not w39717;
w39719 <= not b(13) and not w39718;
w39720 <= not w39185 and not w39468;
w39721 <= not w39195 and w39325;
w39722 <= not w39321 and w39721;
w39723 <= not w39322 and not w39325;
w39724 <= not w39722 and not w39723;
w39725 <= w11362 and not w39724;
w39726 <= not w39467 and w39725;
w39727 <= not w39720 and not w39726;
w39728 <= not b(12) and not w39727;
w39729 <= not w39194 and not w39468;
w39730 <= not w39204 and w39320;
w39731 <= not w39316 and w39730;
w39732 <= not w39317 and not w39320;
w39733 <= not w39731 and not w39732;
w39734 <= w11362 and not w39733;
w39735 <= not w39467 and w39734;
w39736 <= not w39729 and not w39735;
w39737 <= not b(11) and not w39736;
w39738 <= not w39203 and not w39468;
w39739 <= not w39213 and w39315;
w39740 <= not w39311 and w39739;
w39741 <= not w39312 and not w39315;
w39742 <= not w39740 and not w39741;
w39743 <= w11362 and not w39742;
w39744 <= not w39467 and w39743;
w39745 <= not w39738 and not w39744;
w39746 <= not b(10) and not w39745;
w39747 <= not w39212 and not w39468;
w39748 <= not w39222 and w39310;
w39749 <= not w39306 and w39748;
w39750 <= not w39307 and not w39310;
w39751 <= not w39749 and not w39750;
w39752 <= w11362 and not w39751;
w39753 <= not w39467 and w39752;
w39754 <= not w39747 and not w39753;
w39755 <= not b(9) and not w39754;
w39756 <= not w39221 and not w39468;
w39757 <= not w39231 and w39305;
w39758 <= not w39301 and w39757;
w39759 <= not w39302 and not w39305;
w39760 <= not w39758 and not w39759;
w39761 <= w11362 and not w39760;
w39762 <= not w39467 and w39761;
w39763 <= not w39756 and not w39762;
w39764 <= not b(8) and not w39763;
w39765 <= not w39230 and not w39468;
w39766 <= not w39240 and w39300;
w39767 <= not w39296 and w39766;
w39768 <= not w39297 and not w39300;
w39769 <= not w39767 and not w39768;
w39770 <= w11362 and not w39769;
w39771 <= not w39467 and w39770;
w39772 <= not w39765 and not w39771;
w39773 <= not b(7) and not w39772;
w39774 <= not w39239 and not w39468;
w39775 <= not w39249 and w39295;
w39776 <= not w39291 and w39775;
w39777 <= not w39292 and not w39295;
w39778 <= not w39776 and not w39777;
w39779 <= w11362 and not w39778;
w39780 <= not w39467 and w39779;
w39781 <= not w39774 and not w39780;
w39782 <= not b(6) and not w39781;
w39783 <= not w39248 and not w39468;
w39784 <= not w39258 and w39290;
w39785 <= not w39286 and w39784;
w39786 <= not w39287 and not w39290;
w39787 <= not w39785 and not w39786;
w39788 <= w11362 and not w39787;
w39789 <= not w39467 and w39788;
w39790 <= not w39783 and not w39789;
w39791 <= not b(5) and not w39790;
w39792 <= not w39257 and not w39468;
w39793 <= not w39266 and w39285;
w39794 <= not w39281 and w39793;
w39795 <= not w39282 and not w39285;
w39796 <= not w39794 and not w39795;
w39797 <= w11362 and not w39796;
w39798 <= not w39467 and w39797;
w39799 <= not w39792 and not w39798;
w39800 <= not b(4) and not w39799;
w39801 <= not w39265 and not w39468;
w39802 <= not w39276 and w39280;
w39803 <= not w39275 and w39802;
w39804 <= not w39277 and not w39280;
w39805 <= not w39803 and not w39804;
w39806 <= w11362 and not w39805;
w39807 <= not w39467 and w39806;
w39808 <= not w39801 and not w39807;
w39809 <= not b(3) and not w39808;
w39810 <= not w39270 and not w39468;
w39811 <= w11168 and not w39273;
w39812 <= not w39271 and w39811;
w39813 <= w11362 and not w39812;
w39814 <= not w39275 and w39813;
w39815 <= not w39467 and w39814;
w39816 <= not w39810 and not w39815;
w39817 <= not b(2) and not w39816;
w39818 <= w11716 and not w39467;
w39819 <= a(24) and not w39818;
w39820 <= w11721 and not w39467;
w39821 <= not w39819 and not w39820;
w39822 <= b(1) and not w39821;
w39823 <= not b(1) and not w39820;
w39824 <= not w39819 and w39823;
w39825 <= not w39822 and not w39824;
w39826 <= not w11728 and not w39825;
w39827 <= not b(1) and not w39821;
w39828 <= not w39826 and not w39827;
w39829 <= b(2) and not w39815;
w39830 <= not w39810 and w39829;
w39831 <= not w39817 and not w39830;
w39832 <= not w39828 and w39831;
w39833 <= not w39817 and not w39832;
w39834 <= b(3) and not w39807;
w39835 <= not w39801 and w39834;
w39836 <= not w39809 and not w39835;
w39837 <= not w39833 and w39836;
w39838 <= not w39809 and not w39837;
w39839 <= b(4) and not w39798;
w39840 <= not w39792 and w39839;
w39841 <= not w39800 and not w39840;
w39842 <= not w39838 and w39841;
w39843 <= not w39800 and not w39842;
w39844 <= b(5) and not w39789;
w39845 <= not w39783 and w39844;
w39846 <= not w39791 and not w39845;
w39847 <= not w39843 and w39846;
w39848 <= not w39791 and not w39847;
w39849 <= b(6) and not w39780;
w39850 <= not w39774 and w39849;
w39851 <= not w39782 and not w39850;
w39852 <= not w39848 and w39851;
w39853 <= not w39782 and not w39852;
w39854 <= b(7) and not w39771;
w39855 <= not w39765 and w39854;
w39856 <= not w39773 and not w39855;
w39857 <= not w39853 and w39856;
w39858 <= not w39773 and not w39857;
w39859 <= b(8) and not w39762;
w39860 <= not w39756 and w39859;
w39861 <= not w39764 and not w39860;
w39862 <= not w39858 and w39861;
w39863 <= not w39764 and not w39862;
w39864 <= b(9) and not w39753;
w39865 <= not w39747 and w39864;
w39866 <= not w39755 and not w39865;
w39867 <= not w39863 and w39866;
w39868 <= not w39755 and not w39867;
w39869 <= b(10) and not w39744;
w39870 <= not w39738 and w39869;
w39871 <= not w39746 and not w39870;
w39872 <= not w39868 and w39871;
w39873 <= not w39746 and not w39872;
w39874 <= b(11) and not w39735;
w39875 <= not w39729 and w39874;
w39876 <= not w39737 and not w39875;
w39877 <= not w39873 and w39876;
w39878 <= not w39737 and not w39877;
w39879 <= b(12) and not w39726;
w39880 <= not w39720 and w39879;
w39881 <= not w39728 and not w39880;
w39882 <= not w39878 and w39881;
w39883 <= not w39728 and not w39882;
w39884 <= b(13) and not w39717;
w39885 <= not w39711 and w39884;
w39886 <= not w39719 and not w39885;
w39887 <= not w39883 and w39886;
w39888 <= not w39719 and not w39887;
w39889 <= b(14) and not w39708;
w39890 <= not w39702 and w39889;
w39891 <= not w39710 and not w39890;
w39892 <= not w39888 and w39891;
w39893 <= not w39710 and not w39892;
w39894 <= b(15) and not w39699;
w39895 <= not w39693 and w39894;
w39896 <= not w39701 and not w39895;
w39897 <= not w39893 and w39896;
w39898 <= not w39701 and not w39897;
w39899 <= b(16) and not w39690;
w39900 <= not w39684 and w39899;
w39901 <= not w39692 and not w39900;
w39902 <= not w39898 and w39901;
w39903 <= not w39692 and not w39902;
w39904 <= b(17) and not w39681;
w39905 <= not w39675 and w39904;
w39906 <= not w39683 and not w39905;
w39907 <= not w39903 and w39906;
w39908 <= not w39683 and not w39907;
w39909 <= b(18) and not w39672;
w39910 <= not w39666 and w39909;
w39911 <= not w39674 and not w39910;
w39912 <= not w39908 and w39911;
w39913 <= not w39674 and not w39912;
w39914 <= b(19) and not w39663;
w39915 <= not w39657 and w39914;
w39916 <= not w39665 and not w39915;
w39917 <= not w39913 and w39916;
w39918 <= not w39665 and not w39917;
w39919 <= b(20) and not w39654;
w39920 <= not w39648 and w39919;
w39921 <= not w39656 and not w39920;
w39922 <= not w39918 and w39921;
w39923 <= not w39656 and not w39922;
w39924 <= b(21) and not w39645;
w39925 <= not w39639 and w39924;
w39926 <= not w39647 and not w39925;
w39927 <= not w39923 and w39926;
w39928 <= not w39647 and not w39927;
w39929 <= b(22) and not w39636;
w39930 <= not w39630 and w39929;
w39931 <= not w39638 and not w39930;
w39932 <= not w39928 and w39931;
w39933 <= not w39638 and not w39932;
w39934 <= b(23) and not w39627;
w39935 <= not w39621 and w39934;
w39936 <= not w39629 and not w39935;
w39937 <= not w39933 and w39936;
w39938 <= not w39629 and not w39937;
w39939 <= b(24) and not w39618;
w39940 <= not w39612 and w39939;
w39941 <= not w39620 and not w39940;
w39942 <= not w39938 and w39941;
w39943 <= not w39620 and not w39942;
w39944 <= b(25) and not w39609;
w39945 <= not w39603 and w39944;
w39946 <= not w39611 and not w39945;
w39947 <= not w39943 and w39946;
w39948 <= not w39611 and not w39947;
w39949 <= b(26) and not w39600;
w39950 <= not w39594 and w39949;
w39951 <= not w39602 and not w39950;
w39952 <= not w39948 and w39951;
w39953 <= not w39602 and not w39952;
w39954 <= b(27) and not w39591;
w39955 <= not w39585 and w39954;
w39956 <= not w39593 and not w39955;
w39957 <= not w39953 and w39956;
w39958 <= not w39593 and not w39957;
w39959 <= b(28) and not w39582;
w39960 <= not w39576 and w39959;
w39961 <= not w39584 and not w39960;
w39962 <= not w39958 and w39961;
w39963 <= not w39584 and not w39962;
w39964 <= b(29) and not w39573;
w39965 <= not w39567 and w39964;
w39966 <= not w39575 and not w39965;
w39967 <= not w39963 and w39966;
w39968 <= not w39575 and not w39967;
w39969 <= b(30) and not w39564;
w39970 <= not w39558 and w39969;
w39971 <= not w39566 and not w39970;
w39972 <= not w39968 and w39971;
w39973 <= not w39566 and not w39972;
w39974 <= b(31) and not w39555;
w39975 <= not w39549 and w39974;
w39976 <= not w39557 and not w39975;
w39977 <= not w39973 and w39976;
w39978 <= not w39557 and not w39977;
w39979 <= b(32) and not w39546;
w39980 <= not w39540 and w39979;
w39981 <= not w39548 and not w39980;
w39982 <= not w39978 and w39981;
w39983 <= not w39548 and not w39982;
w39984 <= b(33) and not w39537;
w39985 <= not w39531 and w39984;
w39986 <= not w39539 and not w39985;
w39987 <= not w39983 and w39986;
w39988 <= not w39539 and not w39987;
w39989 <= b(34) and not w39528;
w39990 <= not w39522 and w39989;
w39991 <= not w39530 and not w39990;
w39992 <= not w39988 and w39991;
w39993 <= not w39530 and not w39992;
w39994 <= b(35) and not w39519;
w39995 <= not w39513 and w39994;
w39996 <= not w39521 and not w39995;
w39997 <= not w39993 and w39996;
w39998 <= not w39521 and not w39997;
w39999 <= b(36) and not w39510;
w40000 <= not w39504 and w39999;
w40001 <= not w39512 and not w40000;
w40002 <= not w39998 and w40001;
w40003 <= not w39512 and not w40002;
w40004 <= b(37) and not w39501;
w40005 <= not w39495 and w40004;
w40006 <= not w39503 and not w40005;
w40007 <= not w40003 and w40006;
w40008 <= not w39503 and not w40007;
w40009 <= b(38) and not w39492;
w40010 <= not w39486 and w40009;
w40011 <= not w39494 and not w40010;
w40012 <= not w40008 and w40011;
w40013 <= not w39494 and not w40012;
w40014 <= b(39) and not w39475;
w40015 <= not w39469 and w40014;
w40016 <= not w39485 and not w40015;
w40017 <= not w40013 and w40016;
w40018 <= not w39485 and not w40017;
w40019 <= b(40) and not w39477;
w40020 <= not w39482 and w40019;
w40021 <= not w39484 and not w40020;
w40022 <= not w40018 and w40021;
w40023 <= not w39484 and not w40022;
w40024 <= w11927 and not w40023;
w40025 <= not w39476 and not w40024;
w40026 <= not w39494 and w40016;
w40027 <= not w40012 and w40026;
w40028 <= not w40013 and not w40016;
w40029 <= not w40027 and not w40028;
w40030 <= w11927 and not w40029;
w40031 <= not w40023 and w40030;
w40032 <= not w40025 and not w40031;
w40033 <= not b(40) and not w40032;
w40034 <= not w39493 and not w40024;
w40035 <= not w39503 and w40011;
w40036 <= not w40007 and w40035;
w40037 <= not w40008 and not w40011;
w40038 <= not w40036 and not w40037;
w40039 <= w11927 and not w40038;
w40040 <= not w40023 and w40039;
w40041 <= not w40034 and not w40040;
w40042 <= not b(39) and not w40041;
w40043 <= not w39502 and not w40024;
w40044 <= not w39512 and w40006;
w40045 <= not w40002 and w40044;
w40046 <= not w40003 and not w40006;
w40047 <= not w40045 and not w40046;
w40048 <= w11927 and not w40047;
w40049 <= not w40023 and w40048;
w40050 <= not w40043 and not w40049;
w40051 <= not b(38) and not w40050;
w40052 <= not w39511 and not w40024;
w40053 <= not w39521 and w40001;
w40054 <= not w39997 and w40053;
w40055 <= not w39998 and not w40001;
w40056 <= not w40054 and not w40055;
w40057 <= w11927 and not w40056;
w40058 <= not w40023 and w40057;
w40059 <= not w40052 and not w40058;
w40060 <= not b(37) and not w40059;
w40061 <= not w39520 and not w40024;
w40062 <= not w39530 and w39996;
w40063 <= not w39992 and w40062;
w40064 <= not w39993 and not w39996;
w40065 <= not w40063 and not w40064;
w40066 <= w11927 and not w40065;
w40067 <= not w40023 and w40066;
w40068 <= not w40061 and not w40067;
w40069 <= not b(36) and not w40068;
w40070 <= not w39529 and not w40024;
w40071 <= not w39539 and w39991;
w40072 <= not w39987 and w40071;
w40073 <= not w39988 and not w39991;
w40074 <= not w40072 and not w40073;
w40075 <= w11927 and not w40074;
w40076 <= not w40023 and w40075;
w40077 <= not w40070 and not w40076;
w40078 <= not b(35) and not w40077;
w40079 <= not w39538 and not w40024;
w40080 <= not w39548 and w39986;
w40081 <= not w39982 and w40080;
w40082 <= not w39983 and not w39986;
w40083 <= not w40081 and not w40082;
w40084 <= w11927 and not w40083;
w40085 <= not w40023 and w40084;
w40086 <= not w40079 and not w40085;
w40087 <= not b(34) and not w40086;
w40088 <= not w39547 and not w40024;
w40089 <= not w39557 and w39981;
w40090 <= not w39977 and w40089;
w40091 <= not w39978 and not w39981;
w40092 <= not w40090 and not w40091;
w40093 <= w11927 and not w40092;
w40094 <= not w40023 and w40093;
w40095 <= not w40088 and not w40094;
w40096 <= not b(33) and not w40095;
w40097 <= not w39556 and not w40024;
w40098 <= not w39566 and w39976;
w40099 <= not w39972 and w40098;
w40100 <= not w39973 and not w39976;
w40101 <= not w40099 and not w40100;
w40102 <= w11927 and not w40101;
w40103 <= not w40023 and w40102;
w40104 <= not w40097 and not w40103;
w40105 <= not b(32) and not w40104;
w40106 <= not w39565 and not w40024;
w40107 <= not w39575 and w39971;
w40108 <= not w39967 and w40107;
w40109 <= not w39968 and not w39971;
w40110 <= not w40108 and not w40109;
w40111 <= w11927 and not w40110;
w40112 <= not w40023 and w40111;
w40113 <= not w40106 and not w40112;
w40114 <= not b(31) and not w40113;
w40115 <= not w39574 and not w40024;
w40116 <= not w39584 and w39966;
w40117 <= not w39962 and w40116;
w40118 <= not w39963 and not w39966;
w40119 <= not w40117 and not w40118;
w40120 <= w11927 and not w40119;
w40121 <= not w40023 and w40120;
w40122 <= not w40115 and not w40121;
w40123 <= not b(30) and not w40122;
w40124 <= not w39583 and not w40024;
w40125 <= not w39593 and w39961;
w40126 <= not w39957 and w40125;
w40127 <= not w39958 and not w39961;
w40128 <= not w40126 and not w40127;
w40129 <= w11927 and not w40128;
w40130 <= not w40023 and w40129;
w40131 <= not w40124 and not w40130;
w40132 <= not b(29) and not w40131;
w40133 <= not w39592 and not w40024;
w40134 <= not w39602 and w39956;
w40135 <= not w39952 and w40134;
w40136 <= not w39953 and not w39956;
w40137 <= not w40135 and not w40136;
w40138 <= w11927 and not w40137;
w40139 <= not w40023 and w40138;
w40140 <= not w40133 and not w40139;
w40141 <= not b(28) and not w40140;
w40142 <= not w39601 and not w40024;
w40143 <= not w39611 and w39951;
w40144 <= not w39947 and w40143;
w40145 <= not w39948 and not w39951;
w40146 <= not w40144 and not w40145;
w40147 <= w11927 and not w40146;
w40148 <= not w40023 and w40147;
w40149 <= not w40142 and not w40148;
w40150 <= not b(27) and not w40149;
w40151 <= not w39610 and not w40024;
w40152 <= not w39620 and w39946;
w40153 <= not w39942 and w40152;
w40154 <= not w39943 and not w39946;
w40155 <= not w40153 and not w40154;
w40156 <= w11927 and not w40155;
w40157 <= not w40023 and w40156;
w40158 <= not w40151 and not w40157;
w40159 <= not b(26) and not w40158;
w40160 <= not w39619 and not w40024;
w40161 <= not w39629 and w39941;
w40162 <= not w39937 and w40161;
w40163 <= not w39938 and not w39941;
w40164 <= not w40162 and not w40163;
w40165 <= w11927 and not w40164;
w40166 <= not w40023 and w40165;
w40167 <= not w40160 and not w40166;
w40168 <= not b(25) and not w40167;
w40169 <= not w39628 and not w40024;
w40170 <= not w39638 and w39936;
w40171 <= not w39932 and w40170;
w40172 <= not w39933 and not w39936;
w40173 <= not w40171 and not w40172;
w40174 <= w11927 and not w40173;
w40175 <= not w40023 and w40174;
w40176 <= not w40169 and not w40175;
w40177 <= not b(24) and not w40176;
w40178 <= not w39637 and not w40024;
w40179 <= not w39647 and w39931;
w40180 <= not w39927 and w40179;
w40181 <= not w39928 and not w39931;
w40182 <= not w40180 and not w40181;
w40183 <= w11927 and not w40182;
w40184 <= not w40023 and w40183;
w40185 <= not w40178 and not w40184;
w40186 <= not b(23) and not w40185;
w40187 <= not w39646 and not w40024;
w40188 <= not w39656 and w39926;
w40189 <= not w39922 and w40188;
w40190 <= not w39923 and not w39926;
w40191 <= not w40189 and not w40190;
w40192 <= w11927 and not w40191;
w40193 <= not w40023 and w40192;
w40194 <= not w40187 and not w40193;
w40195 <= not b(22) and not w40194;
w40196 <= not w39655 and not w40024;
w40197 <= not w39665 and w39921;
w40198 <= not w39917 and w40197;
w40199 <= not w39918 and not w39921;
w40200 <= not w40198 and not w40199;
w40201 <= w11927 and not w40200;
w40202 <= not w40023 and w40201;
w40203 <= not w40196 and not w40202;
w40204 <= not b(21) and not w40203;
w40205 <= not w39664 and not w40024;
w40206 <= not w39674 and w39916;
w40207 <= not w39912 and w40206;
w40208 <= not w39913 and not w39916;
w40209 <= not w40207 and not w40208;
w40210 <= w11927 and not w40209;
w40211 <= not w40023 and w40210;
w40212 <= not w40205 and not w40211;
w40213 <= not b(20) and not w40212;
w40214 <= not w39673 and not w40024;
w40215 <= not w39683 and w39911;
w40216 <= not w39907 and w40215;
w40217 <= not w39908 and not w39911;
w40218 <= not w40216 and not w40217;
w40219 <= w11927 and not w40218;
w40220 <= not w40023 and w40219;
w40221 <= not w40214 and not w40220;
w40222 <= not b(19) and not w40221;
w40223 <= not w39682 and not w40024;
w40224 <= not w39692 and w39906;
w40225 <= not w39902 and w40224;
w40226 <= not w39903 and not w39906;
w40227 <= not w40225 and not w40226;
w40228 <= w11927 and not w40227;
w40229 <= not w40023 and w40228;
w40230 <= not w40223 and not w40229;
w40231 <= not b(18) and not w40230;
w40232 <= not w39691 and not w40024;
w40233 <= not w39701 and w39901;
w40234 <= not w39897 and w40233;
w40235 <= not w39898 and not w39901;
w40236 <= not w40234 and not w40235;
w40237 <= w11927 and not w40236;
w40238 <= not w40023 and w40237;
w40239 <= not w40232 and not w40238;
w40240 <= not b(17) and not w40239;
w40241 <= not w39700 and not w40024;
w40242 <= not w39710 and w39896;
w40243 <= not w39892 and w40242;
w40244 <= not w39893 and not w39896;
w40245 <= not w40243 and not w40244;
w40246 <= w11927 and not w40245;
w40247 <= not w40023 and w40246;
w40248 <= not w40241 and not w40247;
w40249 <= not b(16) and not w40248;
w40250 <= not w39709 and not w40024;
w40251 <= not w39719 and w39891;
w40252 <= not w39887 and w40251;
w40253 <= not w39888 and not w39891;
w40254 <= not w40252 and not w40253;
w40255 <= w11927 and not w40254;
w40256 <= not w40023 and w40255;
w40257 <= not w40250 and not w40256;
w40258 <= not b(15) and not w40257;
w40259 <= not w39718 and not w40024;
w40260 <= not w39728 and w39886;
w40261 <= not w39882 and w40260;
w40262 <= not w39883 and not w39886;
w40263 <= not w40261 and not w40262;
w40264 <= w11927 and not w40263;
w40265 <= not w40023 and w40264;
w40266 <= not w40259 and not w40265;
w40267 <= not b(14) and not w40266;
w40268 <= not w39727 and not w40024;
w40269 <= not w39737 and w39881;
w40270 <= not w39877 and w40269;
w40271 <= not w39878 and not w39881;
w40272 <= not w40270 and not w40271;
w40273 <= w11927 and not w40272;
w40274 <= not w40023 and w40273;
w40275 <= not w40268 and not w40274;
w40276 <= not b(13) and not w40275;
w40277 <= not w39736 and not w40024;
w40278 <= not w39746 and w39876;
w40279 <= not w39872 and w40278;
w40280 <= not w39873 and not w39876;
w40281 <= not w40279 and not w40280;
w40282 <= w11927 and not w40281;
w40283 <= not w40023 and w40282;
w40284 <= not w40277 and not w40283;
w40285 <= not b(12) and not w40284;
w40286 <= not w39745 and not w40024;
w40287 <= not w39755 and w39871;
w40288 <= not w39867 and w40287;
w40289 <= not w39868 and not w39871;
w40290 <= not w40288 and not w40289;
w40291 <= w11927 and not w40290;
w40292 <= not w40023 and w40291;
w40293 <= not w40286 and not w40292;
w40294 <= not b(11) and not w40293;
w40295 <= not w39754 and not w40024;
w40296 <= not w39764 and w39866;
w40297 <= not w39862 and w40296;
w40298 <= not w39863 and not w39866;
w40299 <= not w40297 and not w40298;
w40300 <= w11927 and not w40299;
w40301 <= not w40023 and w40300;
w40302 <= not w40295 and not w40301;
w40303 <= not b(10) and not w40302;
w40304 <= not w39763 and not w40024;
w40305 <= not w39773 and w39861;
w40306 <= not w39857 and w40305;
w40307 <= not w39858 and not w39861;
w40308 <= not w40306 and not w40307;
w40309 <= w11927 and not w40308;
w40310 <= not w40023 and w40309;
w40311 <= not w40304 and not w40310;
w40312 <= not b(9) and not w40311;
w40313 <= not w39772 and not w40024;
w40314 <= not w39782 and w39856;
w40315 <= not w39852 and w40314;
w40316 <= not w39853 and not w39856;
w40317 <= not w40315 and not w40316;
w40318 <= w11927 and not w40317;
w40319 <= not w40023 and w40318;
w40320 <= not w40313 and not w40319;
w40321 <= not b(8) and not w40320;
w40322 <= not w39781 and not w40024;
w40323 <= not w39791 and w39851;
w40324 <= not w39847 and w40323;
w40325 <= not w39848 and not w39851;
w40326 <= not w40324 and not w40325;
w40327 <= w11927 and not w40326;
w40328 <= not w40023 and w40327;
w40329 <= not w40322 and not w40328;
w40330 <= not b(7) and not w40329;
w40331 <= not w39790 and not w40024;
w40332 <= not w39800 and w39846;
w40333 <= not w39842 and w40332;
w40334 <= not w39843 and not w39846;
w40335 <= not w40333 and not w40334;
w40336 <= w11927 and not w40335;
w40337 <= not w40023 and w40336;
w40338 <= not w40331 and not w40337;
w40339 <= not b(6) and not w40338;
w40340 <= not w39799 and not w40024;
w40341 <= not w39809 and w39841;
w40342 <= not w39837 and w40341;
w40343 <= not w39838 and not w39841;
w40344 <= not w40342 and not w40343;
w40345 <= w11927 and not w40344;
w40346 <= not w40023 and w40345;
w40347 <= not w40340 and not w40346;
w40348 <= not b(5) and not w40347;
w40349 <= not w39808 and not w40024;
w40350 <= not w39817 and w39836;
w40351 <= not w39832 and w40350;
w40352 <= not w39833 and not w39836;
w40353 <= not w40351 and not w40352;
w40354 <= w11927 and not w40353;
w40355 <= not w40023 and w40354;
w40356 <= not w40349 and not w40355;
w40357 <= not b(4) and not w40356;
w40358 <= not w39816 and not w40024;
w40359 <= not w39827 and w39831;
w40360 <= not w39826 and w40359;
w40361 <= not w39828 and not w39831;
w40362 <= not w40360 and not w40361;
w40363 <= w11927 and not w40362;
w40364 <= not w40023 and w40363;
w40365 <= not w40358 and not w40364;
w40366 <= not b(3) and not w40365;
w40367 <= not w39821 and not w40024;
w40368 <= w11728 and not w39824;
w40369 <= not w39822 and w40368;
w40370 <= w11927 and not w40369;
w40371 <= not w39826 and w40370;
w40372 <= not w40023 and w40371;
w40373 <= not w40367 and not w40372;
w40374 <= not b(2) and not w40373;
w40375 <= w12282 and not w40023;
w40376 <= a(23) and not w40375;
w40377 <= w12287 and not w40023;
w40378 <= not w40376 and not w40377;
w40379 <= b(1) and not w40378;
w40380 <= not b(1) and not w40377;
w40381 <= not w40376 and w40380;
w40382 <= not w40379 and not w40381;
w40383 <= not w12294 and not w40382;
w40384 <= not b(1) and not w40378;
w40385 <= not w40383 and not w40384;
w40386 <= b(2) and not w40372;
w40387 <= not w40367 and w40386;
w40388 <= not w40374 and not w40387;
w40389 <= not w40385 and w40388;
w40390 <= not w40374 and not w40389;
w40391 <= b(3) and not w40364;
w40392 <= not w40358 and w40391;
w40393 <= not w40366 and not w40392;
w40394 <= not w40390 and w40393;
w40395 <= not w40366 and not w40394;
w40396 <= b(4) and not w40355;
w40397 <= not w40349 and w40396;
w40398 <= not w40357 and not w40397;
w40399 <= not w40395 and w40398;
w40400 <= not w40357 and not w40399;
w40401 <= b(5) and not w40346;
w40402 <= not w40340 and w40401;
w40403 <= not w40348 and not w40402;
w40404 <= not w40400 and w40403;
w40405 <= not w40348 and not w40404;
w40406 <= b(6) and not w40337;
w40407 <= not w40331 and w40406;
w40408 <= not w40339 and not w40407;
w40409 <= not w40405 and w40408;
w40410 <= not w40339 and not w40409;
w40411 <= b(7) and not w40328;
w40412 <= not w40322 and w40411;
w40413 <= not w40330 and not w40412;
w40414 <= not w40410 and w40413;
w40415 <= not w40330 and not w40414;
w40416 <= b(8) and not w40319;
w40417 <= not w40313 and w40416;
w40418 <= not w40321 and not w40417;
w40419 <= not w40415 and w40418;
w40420 <= not w40321 and not w40419;
w40421 <= b(9) and not w40310;
w40422 <= not w40304 and w40421;
w40423 <= not w40312 and not w40422;
w40424 <= not w40420 and w40423;
w40425 <= not w40312 and not w40424;
w40426 <= b(10) and not w40301;
w40427 <= not w40295 and w40426;
w40428 <= not w40303 and not w40427;
w40429 <= not w40425 and w40428;
w40430 <= not w40303 and not w40429;
w40431 <= b(11) and not w40292;
w40432 <= not w40286 and w40431;
w40433 <= not w40294 and not w40432;
w40434 <= not w40430 and w40433;
w40435 <= not w40294 and not w40434;
w40436 <= b(12) and not w40283;
w40437 <= not w40277 and w40436;
w40438 <= not w40285 and not w40437;
w40439 <= not w40435 and w40438;
w40440 <= not w40285 and not w40439;
w40441 <= b(13) and not w40274;
w40442 <= not w40268 and w40441;
w40443 <= not w40276 and not w40442;
w40444 <= not w40440 and w40443;
w40445 <= not w40276 and not w40444;
w40446 <= b(14) and not w40265;
w40447 <= not w40259 and w40446;
w40448 <= not w40267 and not w40447;
w40449 <= not w40445 and w40448;
w40450 <= not w40267 and not w40449;
w40451 <= b(15) and not w40256;
w40452 <= not w40250 and w40451;
w40453 <= not w40258 and not w40452;
w40454 <= not w40450 and w40453;
w40455 <= not w40258 and not w40454;
w40456 <= b(16) and not w40247;
w40457 <= not w40241 and w40456;
w40458 <= not w40249 and not w40457;
w40459 <= not w40455 and w40458;
w40460 <= not w40249 and not w40459;
w40461 <= b(17) and not w40238;
w40462 <= not w40232 and w40461;
w40463 <= not w40240 and not w40462;
w40464 <= not w40460 and w40463;
w40465 <= not w40240 and not w40464;
w40466 <= b(18) and not w40229;
w40467 <= not w40223 and w40466;
w40468 <= not w40231 and not w40467;
w40469 <= not w40465 and w40468;
w40470 <= not w40231 and not w40469;
w40471 <= b(19) and not w40220;
w40472 <= not w40214 and w40471;
w40473 <= not w40222 and not w40472;
w40474 <= not w40470 and w40473;
w40475 <= not w40222 and not w40474;
w40476 <= b(20) and not w40211;
w40477 <= not w40205 and w40476;
w40478 <= not w40213 and not w40477;
w40479 <= not w40475 and w40478;
w40480 <= not w40213 and not w40479;
w40481 <= b(21) and not w40202;
w40482 <= not w40196 and w40481;
w40483 <= not w40204 and not w40482;
w40484 <= not w40480 and w40483;
w40485 <= not w40204 and not w40484;
w40486 <= b(22) and not w40193;
w40487 <= not w40187 and w40486;
w40488 <= not w40195 and not w40487;
w40489 <= not w40485 and w40488;
w40490 <= not w40195 and not w40489;
w40491 <= b(23) and not w40184;
w40492 <= not w40178 and w40491;
w40493 <= not w40186 and not w40492;
w40494 <= not w40490 and w40493;
w40495 <= not w40186 and not w40494;
w40496 <= b(24) and not w40175;
w40497 <= not w40169 and w40496;
w40498 <= not w40177 and not w40497;
w40499 <= not w40495 and w40498;
w40500 <= not w40177 and not w40499;
w40501 <= b(25) and not w40166;
w40502 <= not w40160 and w40501;
w40503 <= not w40168 and not w40502;
w40504 <= not w40500 and w40503;
w40505 <= not w40168 and not w40504;
w40506 <= b(26) and not w40157;
w40507 <= not w40151 and w40506;
w40508 <= not w40159 and not w40507;
w40509 <= not w40505 and w40508;
w40510 <= not w40159 and not w40509;
w40511 <= b(27) and not w40148;
w40512 <= not w40142 and w40511;
w40513 <= not w40150 and not w40512;
w40514 <= not w40510 and w40513;
w40515 <= not w40150 and not w40514;
w40516 <= b(28) and not w40139;
w40517 <= not w40133 and w40516;
w40518 <= not w40141 and not w40517;
w40519 <= not w40515 and w40518;
w40520 <= not w40141 and not w40519;
w40521 <= b(29) and not w40130;
w40522 <= not w40124 and w40521;
w40523 <= not w40132 and not w40522;
w40524 <= not w40520 and w40523;
w40525 <= not w40132 and not w40524;
w40526 <= b(30) and not w40121;
w40527 <= not w40115 and w40526;
w40528 <= not w40123 and not w40527;
w40529 <= not w40525 and w40528;
w40530 <= not w40123 and not w40529;
w40531 <= b(31) and not w40112;
w40532 <= not w40106 and w40531;
w40533 <= not w40114 and not w40532;
w40534 <= not w40530 and w40533;
w40535 <= not w40114 and not w40534;
w40536 <= b(32) and not w40103;
w40537 <= not w40097 and w40536;
w40538 <= not w40105 and not w40537;
w40539 <= not w40535 and w40538;
w40540 <= not w40105 and not w40539;
w40541 <= b(33) and not w40094;
w40542 <= not w40088 and w40541;
w40543 <= not w40096 and not w40542;
w40544 <= not w40540 and w40543;
w40545 <= not w40096 and not w40544;
w40546 <= b(34) and not w40085;
w40547 <= not w40079 and w40546;
w40548 <= not w40087 and not w40547;
w40549 <= not w40545 and w40548;
w40550 <= not w40087 and not w40549;
w40551 <= b(35) and not w40076;
w40552 <= not w40070 and w40551;
w40553 <= not w40078 and not w40552;
w40554 <= not w40550 and w40553;
w40555 <= not w40078 and not w40554;
w40556 <= b(36) and not w40067;
w40557 <= not w40061 and w40556;
w40558 <= not w40069 and not w40557;
w40559 <= not w40555 and w40558;
w40560 <= not w40069 and not w40559;
w40561 <= b(37) and not w40058;
w40562 <= not w40052 and w40561;
w40563 <= not w40060 and not w40562;
w40564 <= not w40560 and w40563;
w40565 <= not w40060 and not w40564;
w40566 <= b(38) and not w40049;
w40567 <= not w40043 and w40566;
w40568 <= not w40051 and not w40567;
w40569 <= not w40565 and w40568;
w40570 <= not w40051 and not w40569;
w40571 <= b(39) and not w40040;
w40572 <= not w40034 and w40571;
w40573 <= not w40042 and not w40572;
w40574 <= not w40570 and w40573;
w40575 <= not w40042 and not w40574;
w40576 <= b(40) and not w40031;
w40577 <= not w40025 and w40576;
w40578 <= not w40033 and not w40577;
w40579 <= not w40575 and w40578;
w40580 <= not w40033 and not w40579;
w40581 <= not w39483 and not w40024;
w40582 <= not w39485 and w40021;
w40583 <= not w40017 and w40582;
w40584 <= not w40018 and not w40021;
w40585 <= not w40583 and not w40584;
w40586 <= w40024 and not w40585;
w40587 <= not w40581 and not w40586;
w40588 <= not b(41) and not w40587;
w40589 <= b(41) and not w40581;
w40590 <= not w40586 and w40589;
w40591 <= w12504 and not w40590;
w40592 <= not w40588 and w40591;
w40593 <= not w40580 and w40592;
w40594 <= w11927 and not w40587;
w40595 <= not w40593 and not w40594;
w40596 <= not w40042 and w40578;
w40597 <= not w40574 and w40596;
w40598 <= not w40575 and not w40578;
w40599 <= not w40597 and not w40598;
w40600 <= not w40595 and not w40599;
w40601 <= not w40032 and not w40594;
w40602 <= not w40593 and w40601;
w40603 <= not w40600 and not w40602;
w40604 <= not w40033 and not w40590;
w40605 <= not w40588 and w40604;
w40606 <= not w40579 and w40605;
w40607 <= not w40588 and not w40590;
w40608 <= not w40580 and not w40607;
w40609 <= not w40606 and not w40608;
w40610 <= not w40595 and not w40609;
w40611 <= not w40587 and not w40594;
w40612 <= not w40593 and w40611;
w40613 <= not w40610 and not w40612;
w40614 <= not b(42) and not w40613;
w40615 <= not b(41) and not w40603;
w40616 <= not w40051 and w40573;
w40617 <= not w40569 and w40616;
w40618 <= not w40570 and not w40573;
w40619 <= not w40617 and not w40618;
w40620 <= not w40595 and not w40619;
w40621 <= not w40041 and not w40594;
w40622 <= not w40593 and w40621;
w40623 <= not w40620 and not w40622;
w40624 <= not b(40) and not w40623;
w40625 <= not w40060 and w40568;
w40626 <= not w40564 and w40625;
w40627 <= not w40565 and not w40568;
w40628 <= not w40626 and not w40627;
w40629 <= not w40595 and not w40628;
w40630 <= not w40050 and not w40594;
w40631 <= not w40593 and w40630;
w40632 <= not w40629 and not w40631;
w40633 <= not b(39) and not w40632;
w40634 <= not w40069 and w40563;
w40635 <= not w40559 and w40634;
w40636 <= not w40560 and not w40563;
w40637 <= not w40635 and not w40636;
w40638 <= not w40595 and not w40637;
w40639 <= not w40059 and not w40594;
w40640 <= not w40593 and w40639;
w40641 <= not w40638 and not w40640;
w40642 <= not b(38) and not w40641;
w40643 <= not w40078 and w40558;
w40644 <= not w40554 and w40643;
w40645 <= not w40555 and not w40558;
w40646 <= not w40644 and not w40645;
w40647 <= not w40595 and not w40646;
w40648 <= not w40068 and not w40594;
w40649 <= not w40593 and w40648;
w40650 <= not w40647 and not w40649;
w40651 <= not b(37) and not w40650;
w40652 <= not w40087 and w40553;
w40653 <= not w40549 and w40652;
w40654 <= not w40550 and not w40553;
w40655 <= not w40653 and not w40654;
w40656 <= not w40595 and not w40655;
w40657 <= not w40077 and not w40594;
w40658 <= not w40593 and w40657;
w40659 <= not w40656 and not w40658;
w40660 <= not b(36) and not w40659;
w40661 <= not w40096 and w40548;
w40662 <= not w40544 and w40661;
w40663 <= not w40545 and not w40548;
w40664 <= not w40662 and not w40663;
w40665 <= not w40595 and not w40664;
w40666 <= not w40086 and not w40594;
w40667 <= not w40593 and w40666;
w40668 <= not w40665 and not w40667;
w40669 <= not b(35) and not w40668;
w40670 <= not w40105 and w40543;
w40671 <= not w40539 and w40670;
w40672 <= not w40540 and not w40543;
w40673 <= not w40671 and not w40672;
w40674 <= not w40595 and not w40673;
w40675 <= not w40095 and not w40594;
w40676 <= not w40593 and w40675;
w40677 <= not w40674 and not w40676;
w40678 <= not b(34) and not w40677;
w40679 <= not w40114 and w40538;
w40680 <= not w40534 and w40679;
w40681 <= not w40535 and not w40538;
w40682 <= not w40680 and not w40681;
w40683 <= not w40595 and not w40682;
w40684 <= not w40104 and not w40594;
w40685 <= not w40593 and w40684;
w40686 <= not w40683 and not w40685;
w40687 <= not b(33) and not w40686;
w40688 <= not w40123 and w40533;
w40689 <= not w40529 and w40688;
w40690 <= not w40530 and not w40533;
w40691 <= not w40689 and not w40690;
w40692 <= not w40595 and not w40691;
w40693 <= not w40113 and not w40594;
w40694 <= not w40593 and w40693;
w40695 <= not w40692 and not w40694;
w40696 <= not b(32) and not w40695;
w40697 <= not w40132 and w40528;
w40698 <= not w40524 and w40697;
w40699 <= not w40525 and not w40528;
w40700 <= not w40698 and not w40699;
w40701 <= not w40595 and not w40700;
w40702 <= not w40122 and not w40594;
w40703 <= not w40593 and w40702;
w40704 <= not w40701 and not w40703;
w40705 <= not b(31) and not w40704;
w40706 <= not w40141 and w40523;
w40707 <= not w40519 and w40706;
w40708 <= not w40520 and not w40523;
w40709 <= not w40707 and not w40708;
w40710 <= not w40595 and not w40709;
w40711 <= not w40131 and not w40594;
w40712 <= not w40593 and w40711;
w40713 <= not w40710 and not w40712;
w40714 <= not b(30) and not w40713;
w40715 <= not w40150 and w40518;
w40716 <= not w40514 and w40715;
w40717 <= not w40515 and not w40518;
w40718 <= not w40716 and not w40717;
w40719 <= not w40595 and not w40718;
w40720 <= not w40140 and not w40594;
w40721 <= not w40593 and w40720;
w40722 <= not w40719 and not w40721;
w40723 <= not b(29) and not w40722;
w40724 <= not w40159 and w40513;
w40725 <= not w40509 and w40724;
w40726 <= not w40510 and not w40513;
w40727 <= not w40725 and not w40726;
w40728 <= not w40595 and not w40727;
w40729 <= not w40149 and not w40594;
w40730 <= not w40593 and w40729;
w40731 <= not w40728 and not w40730;
w40732 <= not b(28) and not w40731;
w40733 <= not w40168 and w40508;
w40734 <= not w40504 and w40733;
w40735 <= not w40505 and not w40508;
w40736 <= not w40734 and not w40735;
w40737 <= not w40595 and not w40736;
w40738 <= not w40158 and not w40594;
w40739 <= not w40593 and w40738;
w40740 <= not w40737 and not w40739;
w40741 <= not b(27) and not w40740;
w40742 <= not w40177 and w40503;
w40743 <= not w40499 and w40742;
w40744 <= not w40500 and not w40503;
w40745 <= not w40743 and not w40744;
w40746 <= not w40595 and not w40745;
w40747 <= not w40167 and not w40594;
w40748 <= not w40593 and w40747;
w40749 <= not w40746 and not w40748;
w40750 <= not b(26) and not w40749;
w40751 <= not w40186 and w40498;
w40752 <= not w40494 and w40751;
w40753 <= not w40495 and not w40498;
w40754 <= not w40752 and not w40753;
w40755 <= not w40595 and not w40754;
w40756 <= not w40176 and not w40594;
w40757 <= not w40593 and w40756;
w40758 <= not w40755 and not w40757;
w40759 <= not b(25) and not w40758;
w40760 <= not w40195 and w40493;
w40761 <= not w40489 and w40760;
w40762 <= not w40490 and not w40493;
w40763 <= not w40761 and not w40762;
w40764 <= not w40595 and not w40763;
w40765 <= not w40185 and not w40594;
w40766 <= not w40593 and w40765;
w40767 <= not w40764 and not w40766;
w40768 <= not b(24) and not w40767;
w40769 <= not w40204 and w40488;
w40770 <= not w40484 and w40769;
w40771 <= not w40485 and not w40488;
w40772 <= not w40770 and not w40771;
w40773 <= not w40595 and not w40772;
w40774 <= not w40194 and not w40594;
w40775 <= not w40593 and w40774;
w40776 <= not w40773 and not w40775;
w40777 <= not b(23) and not w40776;
w40778 <= not w40213 and w40483;
w40779 <= not w40479 and w40778;
w40780 <= not w40480 and not w40483;
w40781 <= not w40779 and not w40780;
w40782 <= not w40595 and not w40781;
w40783 <= not w40203 and not w40594;
w40784 <= not w40593 and w40783;
w40785 <= not w40782 and not w40784;
w40786 <= not b(22) and not w40785;
w40787 <= not w40222 and w40478;
w40788 <= not w40474 and w40787;
w40789 <= not w40475 and not w40478;
w40790 <= not w40788 and not w40789;
w40791 <= not w40595 and not w40790;
w40792 <= not w40212 and not w40594;
w40793 <= not w40593 and w40792;
w40794 <= not w40791 and not w40793;
w40795 <= not b(21) and not w40794;
w40796 <= not w40231 and w40473;
w40797 <= not w40469 and w40796;
w40798 <= not w40470 and not w40473;
w40799 <= not w40797 and not w40798;
w40800 <= not w40595 and not w40799;
w40801 <= not w40221 and not w40594;
w40802 <= not w40593 and w40801;
w40803 <= not w40800 and not w40802;
w40804 <= not b(20) and not w40803;
w40805 <= not w40240 and w40468;
w40806 <= not w40464 and w40805;
w40807 <= not w40465 and not w40468;
w40808 <= not w40806 and not w40807;
w40809 <= not w40595 and not w40808;
w40810 <= not w40230 and not w40594;
w40811 <= not w40593 and w40810;
w40812 <= not w40809 and not w40811;
w40813 <= not b(19) and not w40812;
w40814 <= not w40249 and w40463;
w40815 <= not w40459 and w40814;
w40816 <= not w40460 and not w40463;
w40817 <= not w40815 and not w40816;
w40818 <= not w40595 and not w40817;
w40819 <= not w40239 and not w40594;
w40820 <= not w40593 and w40819;
w40821 <= not w40818 and not w40820;
w40822 <= not b(18) and not w40821;
w40823 <= not w40258 and w40458;
w40824 <= not w40454 and w40823;
w40825 <= not w40455 and not w40458;
w40826 <= not w40824 and not w40825;
w40827 <= not w40595 and not w40826;
w40828 <= not w40248 and not w40594;
w40829 <= not w40593 and w40828;
w40830 <= not w40827 and not w40829;
w40831 <= not b(17) and not w40830;
w40832 <= not w40267 and w40453;
w40833 <= not w40449 and w40832;
w40834 <= not w40450 and not w40453;
w40835 <= not w40833 and not w40834;
w40836 <= not w40595 and not w40835;
w40837 <= not w40257 and not w40594;
w40838 <= not w40593 and w40837;
w40839 <= not w40836 and not w40838;
w40840 <= not b(16) and not w40839;
w40841 <= not w40276 and w40448;
w40842 <= not w40444 and w40841;
w40843 <= not w40445 and not w40448;
w40844 <= not w40842 and not w40843;
w40845 <= not w40595 and not w40844;
w40846 <= not w40266 and not w40594;
w40847 <= not w40593 and w40846;
w40848 <= not w40845 and not w40847;
w40849 <= not b(15) and not w40848;
w40850 <= not w40285 and w40443;
w40851 <= not w40439 and w40850;
w40852 <= not w40440 and not w40443;
w40853 <= not w40851 and not w40852;
w40854 <= not w40595 and not w40853;
w40855 <= not w40275 and not w40594;
w40856 <= not w40593 and w40855;
w40857 <= not w40854 and not w40856;
w40858 <= not b(14) and not w40857;
w40859 <= not w40294 and w40438;
w40860 <= not w40434 and w40859;
w40861 <= not w40435 and not w40438;
w40862 <= not w40860 and not w40861;
w40863 <= not w40595 and not w40862;
w40864 <= not w40284 and not w40594;
w40865 <= not w40593 and w40864;
w40866 <= not w40863 and not w40865;
w40867 <= not b(13) and not w40866;
w40868 <= not w40303 and w40433;
w40869 <= not w40429 and w40868;
w40870 <= not w40430 and not w40433;
w40871 <= not w40869 and not w40870;
w40872 <= not w40595 and not w40871;
w40873 <= not w40293 and not w40594;
w40874 <= not w40593 and w40873;
w40875 <= not w40872 and not w40874;
w40876 <= not b(12) and not w40875;
w40877 <= not w40312 and w40428;
w40878 <= not w40424 and w40877;
w40879 <= not w40425 and not w40428;
w40880 <= not w40878 and not w40879;
w40881 <= not w40595 and not w40880;
w40882 <= not w40302 and not w40594;
w40883 <= not w40593 and w40882;
w40884 <= not w40881 and not w40883;
w40885 <= not b(11) and not w40884;
w40886 <= not w40321 and w40423;
w40887 <= not w40419 and w40886;
w40888 <= not w40420 and not w40423;
w40889 <= not w40887 and not w40888;
w40890 <= not w40595 and not w40889;
w40891 <= not w40311 and not w40594;
w40892 <= not w40593 and w40891;
w40893 <= not w40890 and not w40892;
w40894 <= not b(10) and not w40893;
w40895 <= not w40330 and w40418;
w40896 <= not w40414 and w40895;
w40897 <= not w40415 and not w40418;
w40898 <= not w40896 and not w40897;
w40899 <= not w40595 and not w40898;
w40900 <= not w40320 and not w40594;
w40901 <= not w40593 and w40900;
w40902 <= not w40899 and not w40901;
w40903 <= not b(9) and not w40902;
w40904 <= not w40339 and w40413;
w40905 <= not w40409 and w40904;
w40906 <= not w40410 and not w40413;
w40907 <= not w40905 and not w40906;
w40908 <= not w40595 and not w40907;
w40909 <= not w40329 and not w40594;
w40910 <= not w40593 and w40909;
w40911 <= not w40908 and not w40910;
w40912 <= not b(8) and not w40911;
w40913 <= not w40348 and w40408;
w40914 <= not w40404 and w40913;
w40915 <= not w40405 and not w40408;
w40916 <= not w40914 and not w40915;
w40917 <= not w40595 and not w40916;
w40918 <= not w40338 and not w40594;
w40919 <= not w40593 and w40918;
w40920 <= not w40917 and not w40919;
w40921 <= not b(7) and not w40920;
w40922 <= not w40357 and w40403;
w40923 <= not w40399 and w40922;
w40924 <= not w40400 and not w40403;
w40925 <= not w40923 and not w40924;
w40926 <= not w40595 and not w40925;
w40927 <= not w40347 and not w40594;
w40928 <= not w40593 and w40927;
w40929 <= not w40926 and not w40928;
w40930 <= not b(6) and not w40929;
w40931 <= not w40366 and w40398;
w40932 <= not w40394 and w40931;
w40933 <= not w40395 and not w40398;
w40934 <= not w40932 and not w40933;
w40935 <= not w40595 and not w40934;
w40936 <= not w40356 and not w40594;
w40937 <= not w40593 and w40936;
w40938 <= not w40935 and not w40937;
w40939 <= not b(5) and not w40938;
w40940 <= not w40374 and w40393;
w40941 <= not w40389 and w40940;
w40942 <= not w40390 and not w40393;
w40943 <= not w40941 and not w40942;
w40944 <= not w40595 and not w40943;
w40945 <= not w40365 and not w40594;
w40946 <= not w40593 and w40945;
w40947 <= not w40944 and not w40946;
w40948 <= not b(4) and not w40947;
w40949 <= not w40384 and w40388;
w40950 <= not w40383 and w40949;
w40951 <= not w40385 and not w40388;
w40952 <= not w40950 and not w40951;
w40953 <= not w40595 and not w40952;
w40954 <= not w40373 and not w40594;
w40955 <= not w40593 and w40954;
w40956 <= not w40953 and not w40955;
w40957 <= not b(3) and not w40956;
w40958 <= w12294 and not w40381;
w40959 <= not w40379 and w40958;
w40960 <= not w40383 and not w40959;
w40961 <= not w40595 and w40960;
w40962 <= not w40378 and not w40594;
w40963 <= not w40593 and w40962;
w40964 <= not w40961 and not w40963;
w40965 <= not b(2) and not w40964;
w40966 <= b(0) and not w40595;
w40967 <= a(22) and not w40966;
w40968 <= w12294 and not w40595;
w40969 <= not w40967 and not w40968;
w40970 <= b(1) and not w40969;
w40971 <= not b(1) and not w40968;
w40972 <= not w40967 and w40971;
w40973 <= not w40970 and not w40972;
w40974 <= not w12888 and not w40973;
w40975 <= not b(1) and not w40969;
w40976 <= not w40974 and not w40975;
w40977 <= b(2) and not w40963;
w40978 <= not w40961 and w40977;
w40979 <= not w40965 and not w40978;
w40980 <= not w40976 and w40979;
w40981 <= not w40965 and not w40980;
w40982 <= b(3) and not w40955;
w40983 <= not w40953 and w40982;
w40984 <= not w40957 and not w40983;
w40985 <= not w40981 and w40984;
w40986 <= not w40957 and not w40985;
w40987 <= b(4) and not w40946;
w40988 <= not w40944 and w40987;
w40989 <= not w40948 and not w40988;
w40990 <= not w40986 and w40989;
w40991 <= not w40948 and not w40990;
w40992 <= b(5) and not w40937;
w40993 <= not w40935 and w40992;
w40994 <= not w40939 and not w40993;
w40995 <= not w40991 and w40994;
w40996 <= not w40939 and not w40995;
w40997 <= b(6) and not w40928;
w40998 <= not w40926 and w40997;
w40999 <= not w40930 and not w40998;
w41000 <= not w40996 and w40999;
w41001 <= not w40930 and not w41000;
w41002 <= b(7) and not w40919;
w41003 <= not w40917 and w41002;
w41004 <= not w40921 and not w41003;
w41005 <= not w41001 and w41004;
w41006 <= not w40921 and not w41005;
w41007 <= b(8) and not w40910;
w41008 <= not w40908 and w41007;
w41009 <= not w40912 and not w41008;
w41010 <= not w41006 and w41009;
w41011 <= not w40912 and not w41010;
w41012 <= b(9) and not w40901;
w41013 <= not w40899 and w41012;
w41014 <= not w40903 and not w41013;
w41015 <= not w41011 and w41014;
w41016 <= not w40903 and not w41015;
w41017 <= b(10) and not w40892;
w41018 <= not w40890 and w41017;
w41019 <= not w40894 and not w41018;
w41020 <= not w41016 and w41019;
w41021 <= not w40894 and not w41020;
w41022 <= b(11) and not w40883;
w41023 <= not w40881 and w41022;
w41024 <= not w40885 and not w41023;
w41025 <= not w41021 and w41024;
w41026 <= not w40885 and not w41025;
w41027 <= b(12) and not w40874;
w41028 <= not w40872 and w41027;
w41029 <= not w40876 and not w41028;
w41030 <= not w41026 and w41029;
w41031 <= not w40876 and not w41030;
w41032 <= b(13) and not w40865;
w41033 <= not w40863 and w41032;
w41034 <= not w40867 and not w41033;
w41035 <= not w41031 and w41034;
w41036 <= not w40867 and not w41035;
w41037 <= b(14) and not w40856;
w41038 <= not w40854 and w41037;
w41039 <= not w40858 and not w41038;
w41040 <= not w41036 and w41039;
w41041 <= not w40858 and not w41040;
w41042 <= b(15) and not w40847;
w41043 <= not w40845 and w41042;
w41044 <= not w40849 and not w41043;
w41045 <= not w41041 and w41044;
w41046 <= not w40849 and not w41045;
w41047 <= b(16) and not w40838;
w41048 <= not w40836 and w41047;
w41049 <= not w40840 and not w41048;
w41050 <= not w41046 and w41049;
w41051 <= not w40840 and not w41050;
w41052 <= b(17) and not w40829;
w41053 <= not w40827 and w41052;
w41054 <= not w40831 and not w41053;
w41055 <= not w41051 and w41054;
w41056 <= not w40831 and not w41055;
w41057 <= b(18) and not w40820;
w41058 <= not w40818 and w41057;
w41059 <= not w40822 and not w41058;
w41060 <= not w41056 and w41059;
w41061 <= not w40822 and not w41060;
w41062 <= b(19) and not w40811;
w41063 <= not w40809 and w41062;
w41064 <= not w40813 and not w41063;
w41065 <= not w41061 and w41064;
w41066 <= not w40813 and not w41065;
w41067 <= b(20) and not w40802;
w41068 <= not w40800 and w41067;
w41069 <= not w40804 and not w41068;
w41070 <= not w41066 and w41069;
w41071 <= not w40804 and not w41070;
w41072 <= b(21) and not w40793;
w41073 <= not w40791 and w41072;
w41074 <= not w40795 and not w41073;
w41075 <= not w41071 and w41074;
w41076 <= not w40795 and not w41075;
w41077 <= b(22) and not w40784;
w41078 <= not w40782 and w41077;
w41079 <= not w40786 and not w41078;
w41080 <= not w41076 and w41079;
w41081 <= not w40786 and not w41080;
w41082 <= b(23) and not w40775;
w41083 <= not w40773 and w41082;
w41084 <= not w40777 and not w41083;
w41085 <= not w41081 and w41084;
w41086 <= not w40777 and not w41085;
w41087 <= b(24) and not w40766;
w41088 <= not w40764 and w41087;
w41089 <= not w40768 and not w41088;
w41090 <= not w41086 and w41089;
w41091 <= not w40768 and not w41090;
w41092 <= b(25) and not w40757;
w41093 <= not w40755 and w41092;
w41094 <= not w40759 and not w41093;
w41095 <= not w41091 and w41094;
w41096 <= not w40759 and not w41095;
w41097 <= b(26) and not w40748;
w41098 <= not w40746 and w41097;
w41099 <= not w40750 and not w41098;
w41100 <= not w41096 and w41099;
w41101 <= not w40750 and not w41100;
w41102 <= b(27) and not w40739;
w41103 <= not w40737 and w41102;
w41104 <= not w40741 and not w41103;
w41105 <= not w41101 and w41104;
w41106 <= not w40741 and not w41105;
w41107 <= b(28) and not w40730;
w41108 <= not w40728 and w41107;
w41109 <= not w40732 and not w41108;
w41110 <= not w41106 and w41109;
w41111 <= not w40732 and not w41110;
w41112 <= b(29) and not w40721;
w41113 <= not w40719 and w41112;
w41114 <= not w40723 and not w41113;
w41115 <= not w41111 and w41114;
w41116 <= not w40723 and not w41115;
w41117 <= b(30) and not w40712;
w41118 <= not w40710 and w41117;
w41119 <= not w40714 and not w41118;
w41120 <= not w41116 and w41119;
w41121 <= not w40714 and not w41120;
w41122 <= b(31) and not w40703;
w41123 <= not w40701 and w41122;
w41124 <= not w40705 and not w41123;
w41125 <= not w41121 and w41124;
w41126 <= not w40705 and not w41125;
w41127 <= b(32) and not w40694;
w41128 <= not w40692 and w41127;
w41129 <= not w40696 and not w41128;
w41130 <= not w41126 and w41129;
w41131 <= not w40696 and not w41130;
w41132 <= b(33) and not w40685;
w41133 <= not w40683 and w41132;
w41134 <= not w40687 and not w41133;
w41135 <= not w41131 and w41134;
w41136 <= not w40687 and not w41135;
w41137 <= b(34) and not w40676;
w41138 <= not w40674 and w41137;
w41139 <= not w40678 and not w41138;
w41140 <= not w41136 and w41139;
w41141 <= not w40678 and not w41140;
w41142 <= b(35) and not w40667;
w41143 <= not w40665 and w41142;
w41144 <= not w40669 and not w41143;
w41145 <= not w41141 and w41144;
w41146 <= not w40669 and not w41145;
w41147 <= b(36) and not w40658;
w41148 <= not w40656 and w41147;
w41149 <= not w40660 and not w41148;
w41150 <= not w41146 and w41149;
w41151 <= not w40660 and not w41150;
w41152 <= b(37) and not w40649;
w41153 <= not w40647 and w41152;
w41154 <= not w40651 and not w41153;
w41155 <= not w41151 and w41154;
w41156 <= not w40651 and not w41155;
w41157 <= b(38) and not w40640;
w41158 <= not w40638 and w41157;
w41159 <= not w40642 and not w41158;
w41160 <= not w41156 and w41159;
w41161 <= not w40642 and not w41160;
w41162 <= b(39) and not w40631;
w41163 <= not w40629 and w41162;
w41164 <= not w40633 and not w41163;
w41165 <= not w41161 and w41164;
w41166 <= not w40633 and not w41165;
w41167 <= b(40) and not w40622;
w41168 <= not w40620 and w41167;
w41169 <= not w40624 and not w41168;
w41170 <= not w41166 and w41169;
w41171 <= not w40624 and not w41170;
w41172 <= b(41) and not w40602;
w41173 <= not w40600 and w41172;
w41174 <= not w40615 and not w41173;
w41175 <= not w41171 and w41174;
w41176 <= not w40615 and not w41175;
w41177 <= b(42) and not w40612;
w41178 <= not w40610 and w41177;
w41179 <= not w40614 and not w41178;
w41180 <= not w41176 and w41179;
w41181 <= not w40614 and not w41180;
w41182 <= w13098 and not w41181;
w41183 <= not w40603 and not w41182;
w41184 <= not w40624 and w41174;
w41185 <= not w41170 and w41184;
w41186 <= not w41171 and not w41174;
w41187 <= not w41185 and not w41186;
w41188 <= w13098 and not w41187;
w41189 <= not w41181 and w41188;
w41190 <= not w41183 and not w41189;
w41191 <= not b(42) and not w41190;
w41192 <= not w40623 and not w41182;
w41193 <= not w40633 and w41169;
w41194 <= not w41165 and w41193;
w41195 <= not w41166 and not w41169;
w41196 <= not w41194 and not w41195;
w41197 <= w13098 and not w41196;
w41198 <= not w41181 and w41197;
w41199 <= not w41192 and not w41198;
w41200 <= not b(41) and not w41199;
w41201 <= not w40632 and not w41182;
w41202 <= not w40642 and w41164;
w41203 <= not w41160 and w41202;
w41204 <= not w41161 and not w41164;
w41205 <= not w41203 and not w41204;
w41206 <= w13098 and not w41205;
w41207 <= not w41181 and w41206;
w41208 <= not w41201 and not w41207;
w41209 <= not b(40) and not w41208;
w41210 <= not w40641 and not w41182;
w41211 <= not w40651 and w41159;
w41212 <= not w41155 and w41211;
w41213 <= not w41156 and not w41159;
w41214 <= not w41212 and not w41213;
w41215 <= w13098 and not w41214;
w41216 <= not w41181 and w41215;
w41217 <= not w41210 and not w41216;
w41218 <= not b(39) and not w41217;
w41219 <= not w40650 and not w41182;
w41220 <= not w40660 and w41154;
w41221 <= not w41150 and w41220;
w41222 <= not w41151 and not w41154;
w41223 <= not w41221 and not w41222;
w41224 <= w13098 and not w41223;
w41225 <= not w41181 and w41224;
w41226 <= not w41219 and not w41225;
w41227 <= not b(38) and not w41226;
w41228 <= not w40659 and not w41182;
w41229 <= not w40669 and w41149;
w41230 <= not w41145 and w41229;
w41231 <= not w41146 and not w41149;
w41232 <= not w41230 and not w41231;
w41233 <= w13098 and not w41232;
w41234 <= not w41181 and w41233;
w41235 <= not w41228 and not w41234;
w41236 <= not b(37) and not w41235;
w41237 <= not w40668 and not w41182;
w41238 <= not w40678 and w41144;
w41239 <= not w41140 and w41238;
w41240 <= not w41141 and not w41144;
w41241 <= not w41239 and not w41240;
w41242 <= w13098 and not w41241;
w41243 <= not w41181 and w41242;
w41244 <= not w41237 and not w41243;
w41245 <= not b(36) and not w41244;
w41246 <= not w40677 and not w41182;
w41247 <= not w40687 and w41139;
w41248 <= not w41135 and w41247;
w41249 <= not w41136 and not w41139;
w41250 <= not w41248 and not w41249;
w41251 <= w13098 and not w41250;
w41252 <= not w41181 and w41251;
w41253 <= not w41246 and not w41252;
w41254 <= not b(35) and not w41253;
w41255 <= not w40686 and not w41182;
w41256 <= not w40696 and w41134;
w41257 <= not w41130 and w41256;
w41258 <= not w41131 and not w41134;
w41259 <= not w41257 and not w41258;
w41260 <= w13098 and not w41259;
w41261 <= not w41181 and w41260;
w41262 <= not w41255 and not w41261;
w41263 <= not b(34) and not w41262;
w41264 <= not w40695 and not w41182;
w41265 <= not w40705 and w41129;
w41266 <= not w41125 and w41265;
w41267 <= not w41126 and not w41129;
w41268 <= not w41266 and not w41267;
w41269 <= w13098 and not w41268;
w41270 <= not w41181 and w41269;
w41271 <= not w41264 and not w41270;
w41272 <= not b(33) and not w41271;
w41273 <= not w40704 and not w41182;
w41274 <= not w40714 and w41124;
w41275 <= not w41120 and w41274;
w41276 <= not w41121 and not w41124;
w41277 <= not w41275 and not w41276;
w41278 <= w13098 and not w41277;
w41279 <= not w41181 and w41278;
w41280 <= not w41273 and not w41279;
w41281 <= not b(32) and not w41280;
w41282 <= not w40713 and not w41182;
w41283 <= not w40723 and w41119;
w41284 <= not w41115 and w41283;
w41285 <= not w41116 and not w41119;
w41286 <= not w41284 and not w41285;
w41287 <= w13098 and not w41286;
w41288 <= not w41181 and w41287;
w41289 <= not w41282 and not w41288;
w41290 <= not b(31) and not w41289;
w41291 <= not w40722 and not w41182;
w41292 <= not w40732 and w41114;
w41293 <= not w41110 and w41292;
w41294 <= not w41111 and not w41114;
w41295 <= not w41293 and not w41294;
w41296 <= w13098 and not w41295;
w41297 <= not w41181 and w41296;
w41298 <= not w41291 and not w41297;
w41299 <= not b(30) and not w41298;
w41300 <= not w40731 and not w41182;
w41301 <= not w40741 and w41109;
w41302 <= not w41105 and w41301;
w41303 <= not w41106 and not w41109;
w41304 <= not w41302 and not w41303;
w41305 <= w13098 and not w41304;
w41306 <= not w41181 and w41305;
w41307 <= not w41300 and not w41306;
w41308 <= not b(29) and not w41307;
w41309 <= not w40740 and not w41182;
w41310 <= not w40750 and w41104;
w41311 <= not w41100 and w41310;
w41312 <= not w41101 and not w41104;
w41313 <= not w41311 and not w41312;
w41314 <= w13098 and not w41313;
w41315 <= not w41181 and w41314;
w41316 <= not w41309 and not w41315;
w41317 <= not b(28) and not w41316;
w41318 <= not w40749 and not w41182;
w41319 <= not w40759 and w41099;
w41320 <= not w41095 and w41319;
w41321 <= not w41096 and not w41099;
w41322 <= not w41320 and not w41321;
w41323 <= w13098 and not w41322;
w41324 <= not w41181 and w41323;
w41325 <= not w41318 and not w41324;
w41326 <= not b(27) and not w41325;
w41327 <= not w40758 and not w41182;
w41328 <= not w40768 and w41094;
w41329 <= not w41090 and w41328;
w41330 <= not w41091 and not w41094;
w41331 <= not w41329 and not w41330;
w41332 <= w13098 and not w41331;
w41333 <= not w41181 and w41332;
w41334 <= not w41327 and not w41333;
w41335 <= not b(26) and not w41334;
w41336 <= not w40767 and not w41182;
w41337 <= not w40777 and w41089;
w41338 <= not w41085 and w41337;
w41339 <= not w41086 and not w41089;
w41340 <= not w41338 and not w41339;
w41341 <= w13098 and not w41340;
w41342 <= not w41181 and w41341;
w41343 <= not w41336 and not w41342;
w41344 <= not b(25) and not w41343;
w41345 <= not w40776 and not w41182;
w41346 <= not w40786 and w41084;
w41347 <= not w41080 and w41346;
w41348 <= not w41081 and not w41084;
w41349 <= not w41347 and not w41348;
w41350 <= w13098 and not w41349;
w41351 <= not w41181 and w41350;
w41352 <= not w41345 and not w41351;
w41353 <= not b(24) and not w41352;
w41354 <= not w40785 and not w41182;
w41355 <= not w40795 and w41079;
w41356 <= not w41075 and w41355;
w41357 <= not w41076 and not w41079;
w41358 <= not w41356 and not w41357;
w41359 <= w13098 and not w41358;
w41360 <= not w41181 and w41359;
w41361 <= not w41354 and not w41360;
w41362 <= not b(23) and not w41361;
w41363 <= not w40794 and not w41182;
w41364 <= not w40804 and w41074;
w41365 <= not w41070 and w41364;
w41366 <= not w41071 and not w41074;
w41367 <= not w41365 and not w41366;
w41368 <= w13098 and not w41367;
w41369 <= not w41181 and w41368;
w41370 <= not w41363 and not w41369;
w41371 <= not b(22) and not w41370;
w41372 <= not w40803 and not w41182;
w41373 <= not w40813 and w41069;
w41374 <= not w41065 and w41373;
w41375 <= not w41066 and not w41069;
w41376 <= not w41374 and not w41375;
w41377 <= w13098 and not w41376;
w41378 <= not w41181 and w41377;
w41379 <= not w41372 and not w41378;
w41380 <= not b(21) and not w41379;
w41381 <= not w40812 and not w41182;
w41382 <= not w40822 and w41064;
w41383 <= not w41060 and w41382;
w41384 <= not w41061 and not w41064;
w41385 <= not w41383 and not w41384;
w41386 <= w13098 and not w41385;
w41387 <= not w41181 and w41386;
w41388 <= not w41381 and not w41387;
w41389 <= not b(20) and not w41388;
w41390 <= not w40821 and not w41182;
w41391 <= not w40831 and w41059;
w41392 <= not w41055 and w41391;
w41393 <= not w41056 and not w41059;
w41394 <= not w41392 and not w41393;
w41395 <= w13098 and not w41394;
w41396 <= not w41181 and w41395;
w41397 <= not w41390 and not w41396;
w41398 <= not b(19) and not w41397;
w41399 <= not w40830 and not w41182;
w41400 <= not w40840 and w41054;
w41401 <= not w41050 and w41400;
w41402 <= not w41051 and not w41054;
w41403 <= not w41401 and not w41402;
w41404 <= w13098 and not w41403;
w41405 <= not w41181 and w41404;
w41406 <= not w41399 and not w41405;
w41407 <= not b(18) and not w41406;
w41408 <= not w40839 and not w41182;
w41409 <= not w40849 and w41049;
w41410 <= not w41045 and w41409;
w41411 <= not w41046 and not w41049;
w41412 <= not w41410 and not w41411;
w41413 <= w13098 and not w41412;
w41414 <= not w41181 and w41413;
w41415 <= not w41408 and not w41414;
w41416 <= not b(17) and not w41415;
w41417 <= not w40848 and not w41182;
w41418 <= not w40858 and w41044;
w41419 <= not w41040 and w41418;
w41420 <= not w41041 and not w41044;
w41421 <= not w41419 and not w41420;
w41422 <= w13098 and not w41421;
w41423 <= not w41181 and w41422;
w41424 <= not w41417 and not w41423;
w41425 <= not b(16) and not w41424;
w41426 <= not w40857 and not w41182;
w41427 <= not w40867 and w41039;
w41428 <= not w41035 and w41427;
w41429 <= not w41036 and not w41039;
w41430 <= not w41428 and not w41429;
w41431 <= w13098 and not w41430;
w41432 <= not w41181 and w41431;
w41433 <= not w41426 and not w41432;
w41434 <= not b(15) and not w41433;
w41435 <= not w40866 and not w41182;
w41436 <= not w40876 and w41034;
w41437 <= not w41030 and w41436;
w41438 <= not w41031 and not w41034;
w41439 <= not w41437 and not w41438;
w41440 <= w13098 and not w41439;
w41441 <= not w41181 and w41440;
w41442 <= not w41435 and not w41441;
w41443 <= not b(14) and not w41442;
w41444 <= not w40875 and not w41182;
w41445 <= not w40885 and w41029;
w41446 <= not w41025 and w41445;
w41447 <= not w41026 and not w41029;
w41448 <= not w41446 and not w41447;
w41449 <= w13098 and not w41448;
w41450 <= not w41181 and w41449;
w41451 <= not w41444 and not w41450;
w41452 <= not b(13) and not w41451;
w41453 <= not w40884 and not w41182;
w41454 <= not w40894 and w41024;
w41455 <= not w41020 and w41454;
w41456 <= not w41021 and not w41024;
w41457 <= not w41455 and not w41456;
w41458 <= w13098 and not w41457;
w41459 <= not w41181 and w41458;
w41460 <= not w41453 and not w41459;
w41461 <= not b(12) and not w41460;
w41462 <= not w40893 and not w41182;
w41463 <= not w40903 and w41019;
w41464 <= not w41015 and w41463;
w41465 <= not w41016 and not w41019;
w41466 <= not w41464 and not w41465;
w41467 <= w13098 and not w41466;
w41468 <= not w41181 and w41467;
w41469 <= not w41462 and not w41468;
w41470 <= not b(11) and not w41469;
w41471 <= not w40902 and not w41182;
w41472 <= not w40912 and w41014;
w41473 <= not w41010 and w41472;
w41474 <= not w41011 and not w41014;
w41475 <= not w41473 and not w41474;
w41476 <= w13098 and not w41475;
w41477 <= not w41181 and w41476;
w41478 <= not w41471 and not w41477;
w41479 <= not b(10) and not w41478;
w41480 <= not w40911 and not w41182;
w41481 <= not w40921 and w41009;
w41482 <= not w41005 and w41481;
w41483 <= not w41006 and not w41009;
w41484 <= not w41482 and not w41483;
w41485 <= w13098 and not w41484;
w41486 <= not w41181 and w41485;
w41487 <= not w41480 and not w41486;
w41488 <= not b(9) and not w41487;
w41489 <= not w40920 and not w41182;
w41490 <= not w40930 and w41004;
w41491 <= not w41000 and w41490;
w41492 <= not w41001 and not w41004;
w41493 <= not w41491 and not w41492;
w41494 <= w13098 and not w41493;
w41495 <= not w41181 and w41494;
w41496 <= not w41489 and not w41495;
w41497 <= not b(8) and not w41496;
w41498 <= not w40929 and not w41182;
w41499 <= not w40939 and w40999;
w41500 <= not w40995 and w41499;
w41501 <= not w40996 and not w40999;
w41502 <= not w41500 and not w41501;
w41503 <= w13098 and not w41502;
w41504 <= not w41181 and w41503;
w41505 <= not w41498 and not w41504;
w41506 <= not b(7) and not w41505;
w41507 <= not w40938 and not w41182;
w41508 <= not w40948 and w40994;
w41509 <= not w40990 and w41508;
w41510 <= not w40991 and not w40994;
w41511 <= not w41509 and not w41510;
w41512 <= w13098 and not w41511;
w41513 <= not w41181 and w41512;
w41514 <= not w41507 and not w41513;
w41515 <= not b(6) and not w41514;
w41516 <= not w40947 and not w41182;
w41517 <= not w40957 and w40989;
w41518 <= not w40985 and w41517;
w41519 <= not w40986 and not w40989;
w41520 <= not w41518 and not w41519;
w41521 <= w13098 and not w41520;
w41522 <= not w41181 and w41521;
w41523 <= not w41516 and not w41522;
w41524 <= not b(5) and not w41523;
w41525 <= not w40956 and not w41182;
w41526 <= not w40965 and w40984;
w41527 <= not w40980 and w41526;
w41528 <= not w40981 and not w40984;
w41529 <= not w41527 and not w41528;
w41530 <= w13098 and not w41529;
w41531 <= not w41181 and w41530;
w41532 <= not w41525 and not w41531;
w41533 <= not b(4) and not w41532;
w41534 <= not w40964 and not w41182;
w41535 <= not w40975 and w40979;
w41536 <= not w40974 and w41535;
w41537 <= not w40976 and not w40979;
w41538 <= not w41536 and not w41537;
w41539 <= w13098 and not w41538;
w41540 <= not w41181 and w41539;
w41541 <= not w41534 and not w41540;
w41542 <= not b(3) and not w41541;
w41543 <= not w40969 and not w41182;
w41544 <= w12888 and not w40972;
w41545 <= not w40970 and w41544;
w41546 <= w13098 and not w41545;
w41547 <= not w40974 and w41546;
w41548 <= not w41181 and w41547;
w41549 <= not w41543 and not w41548;
w41550 <= not b(2) and not w41549;
w41551 <= w13470 and not w41181;
w41552 <= a(21) and not w41551;
w41553 <= w13475 and not w41181;
w41554 <= not w41552 and not w41553;
w41555 <= b(1) and not w41554;
w41556 <= not b(1) and not w41553;
w41557 <= not w41552 and w41556;
w41558 <= not w41555 and not w41557;
w41559 <= not w13482 and not w41558;
w41560 <= not b(1) and not w41554;
w41561 <= not w41559 and not w41560;
w41562 <= b(2) and not w41548;
w41563 <= not w41543 and w41562;
w41564 <= not w41550 and not w41563;
w41565 <= not w41561 and w41564;
w41566 <= not w41550 and not w41565;
w41567 <= b(3) and not w41540;
w41568 <= not w41534 and w41567;
w41569 <= not w41542 and not w41568;
w41570 <= not w41566 and w41569;
w41571 <= not w41542 and not w41570;
w41572 <= b(4) and not w41531;
w41573 <= not w41525 and w41572;
w41574 <= not w41533 and not w41573;
w41575 <= not w41571 and w41574;
w41576 <= not w41533 and not w41575;
w41577 <= b(5) and not w41522;
w41578 <= not w41516 and w41577;
w41579 <= not w41524 and not w41578;
w41580 <= not w41576 and w41579;
w41581 <= not w41524 and not w41580;
w41582 <= b(6) and not w41513;
w41583 <= not w41507 and w41582;
w41584 <= not w41515 and not w41583;
w41585 <= not w41581 and w41584;
w41586 <= not w41515 and not w41585;
w41587 <= b(7) and not w41504;
w41588 <= not w41498 and w41587;
w41589 <= not w41506 and not w41588;
w41590 <= not w41586 and w41589;
w41591 <= not w41506 and not w41590;
w41592 <= b(8) and not w41495;
w41593 <= not w41489 and w41592;
w41594 <= not w41497 and not w41593;
w41595 <= not w41591 and w41594;
w41596 <= not w41497 and not w41595;
w41597 <= b(9) and not w41486;
w41598 <= not w41480 and w41597;
w41599 <= not w41488 and not w41598;
w41600 <= not w41596 and w41599;
w41601 <= not w41488 and not w41600;
w41602 <= b(10) and not w41477;
w41603 <= not w41471 and w41602;
w41604 <= not w41479 and not w41603;
w41605 <= not w41601 and w41604;
w41606 <= not w41479 and not w41605;
w41607 <= b(11) and not w41468;
w41608 <= not w41462 and w41607;
w41609 <= not w41470 and not w41608;
w41610 <= not w41606 and w41609;
w41611 <= not w41470 and not w41610;
w41612 <= b(12) and not w41459;
w41613 <= not w41453 and w41612;
w41614 <= not w41461 and not w41613;
w41615 <= not w41611 and w41614;
w41616 <= not w41461 and not w41615;
w41617 <= b(13) and not w41450;
w41618 <= not w41444 and w41617;
w41619 <= not w41452 and not w41618;
w41620 <= not w41616 and w41619;
w41621 <= not w41452 and not w41620;
w41622 <= b(14) and not w41441;
w41623 <= not w41435 and w41622;
w41624 <= not w41443 and not w41623;
w41625 <= not w41621 and w41624;
w41626 <= not w41443 and not w41625;
w41627 <= b(15) and not w41432;
w41628 <= not w41426 and w41627;
w41629 <= not w41434 and not w41628;
w41630 <= not w41626 and w41629;
w41631 <= not w41434 and not w41630;
w41632 <= b(16) and not w41423;
w41633 <= not w41417 and w41632;
w41634 <= not w41425 and not w41633;
w41635 <= not w41631 and w41634;
w41636 <= not w41425 and not w41635;
w41637 <= b(17) and not w41414;
w41638 <= not w41408 and w41637;
w41639 <= not w41416 and not w41638;
w41640 <= not w41636 and w41639;
w41641 <= not w41416 and not w41640;
w41642 <= b(18) and not w41405;
w41643 <= not w41399 and w41642;
w41644 <= not w41407 and not w41643;
w41645 <= not w41641 and w41644;
w41646 <= not w41407 and not w41645;
w41647 <= b(19) and not w41396;
w41648 <= not w41390 and w41647;
w41649 <= not w41398 and not w41648;
w41650 <= not w41646 and w41649;
w41651 <= not w41398 and not w41650;
w41652 <= b(20) and not w41387;
w41653 <= not w41381 and w41652;
w41654 <= not w41389 and not w41653;
w41655 <= not w41651 and w41654;
w41656 <= not w41389 and not w41655;
w41657 <= b(21) and not w41378;
w41658 <= not w41372 and w41657;
w41659 <= not w41380 and not w41658;
w41660 <= not w41656 and w41659;
w41661 <= not w41380 and not w41660;
w41662 <= b(22) and not w41369;
w41663 <= not w41363 and w41662;
w41664 <= not w41371 and not w41663;
w41665 <= not w41661 and w41664;
w41666 <= not w41371 and not w41665;
w41667 <= b(23) and not w41360;
w41668 <= not w41354 and w41667;
w41669 <= not w41362 and not w41668;
w41670 <= not w41666 and w41669;
w41671 <= not w41362 and not w41670;
w41672 <= b(24) and not w41351;
w41673 <= not w41345 and w41672;
w41674 <= not w41353 and not w41673;
w41675 <= not w41671 and w41674;
w41676 <= not w41353 and not w41675;
w41677 <= b(25) and not w41342;
w41678 <= not w41336 and w41677;
w41679 <= not w41344 and not w41678;
w41680 <= not w41676 and w41679;
w41681 <= not w41344 and not w41680;
w41682 <= b(26) and not w41333;
w41683 <= not w41327 and w41682;
w41684 <= not w41335 and not w41683;
w41685 <= not w41681 and w41684;
w41686 <= not w41335 and not w41685;
w41687 <= b(27) and not w41324;
w41688 <= not w41318 and w41687;
w41689 <= not w41326 and not w41688;
w41690 <= not w41686 and w41689;
w41691 <= not w41326 and not w41690;
w41692 <= b(28) and not w41315;
w41693 <= not w41309 and w41692;
w41694 <= not w41317 and not w41693;
w41695 <= not w41691 and w41694;
w41696 <= not w41317 and not w41695;
w41697 <= b(29) and not w41306;
w41698 <= not w41300 and w41697;
w41699 <= not w41308 and not w41698;
w41700 <= not w41696 and w41699;
w41701 <= not w41308 and not w41700;
w41702 <= b(30) and not w41297;
w41703 <= not w41291 and w41702;
w41704 <= not w41299 and not w41703;
w41705 <= not w41701 and w41704;
w41706 <= not w41299 and not w41705;
w41707 <= b(31) and not w41288;
w41708 <= not w41282 and w41707;
w41709 <= not w41290 and not w41708;
w41710 <= not w41706 and w41709;
w41711 <= not w41290 and not w41710;
w41712 <= b(32) and not w41279;
w41713 <= not w41273 and w41712;
w41714 <= not w41281 and not w41713;
w41715 <= not w41711 and w41714;
w41716 <= not w41281 and not w41715;
w41717 <= b(33) and not w41270;
w41718 <= not w41264 and w41717;
w41719 <= not w41272 and not w41718;
w41720 <= not w41716 and w41719;
w41721 <= not w41272 and not w41720;
w41722 <= b(34) and not w41261;
w41723 <= not w41255 and w41722;
w41724 <= not w41263 and not w41723;
w41725 <= not w41721 and w41724;
w41726 <= not w41263 and not w41725;
w41727 <= b(35) and not w41252;
w41728 <= not w41246 and w41727;
w41729 <= not w41254 and not w41728;
w41730 <= not w41726 and w41729;
w41731 <= not w41254 and not w41730;
w41732 <= b(36) and not w41243;
w41733 <= not w41237 and w41732;
w41734 <= not w41245 and not w41733;
w41735 <= not w41731 and w41734;
w41736 <= not w41245 and not w41735;
w41737 <= b(37) and not w41234;
w41738 <= not w41228 and w41737;
w41739 <= not w41236 and not w41738;
w41740 <= not w41736 and w41739;
w41741 <= not w41236 and not w41740;
w41742 <= b(38) and not w41225;
w41743 <= not w41219 and w41742;
w41744 <= not w41227 and not w41743;
w41745 <= not w41741 and w41744;
w41746 <= not w41227 and not w41745;
w41747 <= b(39) and not w41216;
w41748 <= not w41210 and w41747;
w41749 <= not w41218 and not w41748;
w41750 <= not w41746 and w41749;
w41751 <= not w41218 and not w41750;
w41752 <= b(40) and not w41207;
w41753 <= not w41201 and w41752;
w41754 <= not w41209 and not w41753;
w41755 <= not w41751 and w41754;
w41756 <= not w41209 and not w41755;
w41757 <= b(41) and not w41198;
w41758 <= not w41192 and w41757;
w41759 <= not w41200 and not w41758;
w41760 <= not w41756 and w41759;
w41761 <= not w41200 and not w41760;
w41762 <= b(42) and not w41189;
w41763 <= not w41183 and w41762;
w41764 <= not w41191 and not w41763;
w41765 <= not w41761 and w41764;
w41766 <= not w41191 and not w41765;
w41767 <= not w40613 and not w41182;
w41768 <= not w40615 and w41179;
w41769 <= not w41175 and w41768;
w41770 <= not w41176 and not w41179;
w41771 <= not w41769 and not w41770;
w41772 <= w41182 and not w41771;
w41773 <= not w41767 and not w41772;
w41774 <= not b(43) and not w41773;
w41775 <= b(43) and not w41767;
w41776 <= not w41772 and w41775;
w41777 <= w13701 and not w41776;
w41778 <= not w41774 and w41777;
w41779 <= not w41766 and w41778;
w41780 <= w13098 and not w41773;
w41781 <= not w41779 and not w41780;
w41782 <= not w41200 and w41764;
w41783 <= not w41760 and w41782;
w41784 <= not w41761 and not w41764;
w41785 <= not w41783 and not w41784;
w41786 <= not w41781 and not w41785;
w41787 <= not w41190 and not w41780;
w41788 <= not w41779 and w41787;
w41789 <= not w41786 and not w41788;
w41790 <= not b(43) and not w41789;
w41791 <= not w41209 and w41759;
w41792 <= not w41755 and w41791;
w41793 <= not w41756 and not w41759;
w41794 <= not w41792 and not w41793;
w41795 <= not w41781 and not w41794;
w41796 <= not w41199 and not w41780;
w41797 <= not w41779 and w41796;
w41798 <= not w41795 and not w41797;
w41799 <= not b(42) and not w41798;
w41800 <= not w41218 and w41754;
w41801 <= not w41750 and w41800;
w41802 <= not w41751 and not w41754;
w41803 <= not w41801 and not w41802;
w41804 <= not w41781 and not w41803;
w41805 <= not w41208 and not w41780;
w41806 <= not w41779 and w41805;
w41807 <= not w41804 and not w41806;
w41808 <= not b(41) and not w41807;
w41809 <= not w41227 and w41749;
w41810 <= not w41745 and w41809;
w41811 <= not w41746 and not w41749;
w41812 <= not w41810 and not w41811;
w41813 <= not w41781 and not w41812;
w41814 <= not w41217 and not w41780;
w41815 <= not w41779 and w41814;
w41816 <= not w41813 and not w41815;
w41817 <= not b(40) and not w41816;
w41818 <= not w41236 and w41744;
w41819 <= not w41740 and w41818;
w41820 <= not w41741 and not w41744;
w41821 <= not w41819 and not w41820;
w41822 <= not w41781 and not w41821;
w41823 <= not w41226 and not w41780;
w41824 <= not w41779 and w41823;
w41825 <= not w41822 and not w41824;
w41826 <= not b(39) and not w41825;
w41827 <= not w41245 and w41739;
w41828 <= not w41735 and w41827;
w41829 <= not w41736 and not w41739;
w41830 <= not w41828 and not w41829;
w41831 <= not w41781 and not w41830;
w41832 <= not w41235 and not w41780;
w41833 <= not w41779 and w41832;
w41834 <= not w41831 and not w41833;
w41835 <= not b(38) and not w41834;
w41836 <= not w41254 and w41734;
w41837 <= not w41730 and w41836;
w41838 <= not w41731 and not w41734;
w41839 <= not w41837 and not w41838;
w41840 <= not w41781 and not w41839;
w41841 <= not w41244 and not w41780;
w41842 <= not w41779 and w41841;
w41843 <= not w41840 and not w41842;
w41844 <= not b(37) and not w41843;
w41845 <= not w41263 and w41729;
w41846 <= not w41725 and w41845;
w41847 <= not w41726 and not w41729;
w41848 <= not w41846 and not w41847;
w41849 <= not w41781 and not w41848;
w41850 <= not w41253 and not w41780;
w41851 <= not w41779 and w41850;
w41852 <= not w41849 and not w41851;
w41853 <= not b(36) and not w41852;
w41854 <= not w41272 and w41724;
w41855 <= not w41720 and w41854;
w41856 <= not w41721 and not w41724;
w41857 <= not w41855 and not w41856;
w41858 <= not w41781 and not w41857;
w41859 <= not w41262 and not w41780;
w41860 <= not w41779 and w41859;
w41861 <= not w41858 and not w41860;
w41862 <= not b(35) and not w41861;
w41863 <= not w41281 and w41719;
w41864 <= not w41715 and w41863;
w41865 <= not w41716 and not w41719;
w41866 <= not w41864 and not w41865;
w41867 <= not w41781 and not w41866;
w41868 <= not w41271 and not w41780;
w41869 <= not w41779 and w41868;
w41870 <= not w41867 and not w41869;
w41871 <= not b(34) and not w41870;
w41872 <= not w41290 and w41714;
w41873 <= not w41710 and w41872;
w41874 <= not w41711 and not w41714;
w41875 <= not w41873 and not w41874;
w41876 <= not w41781 and not w41875;
w41877 <= not w41280 and not w41780;
w41878 <= not w41779 and w41877;
w41879 <= not w41876 and not w41878;
w41880 <= not b(33) and not w41879;
w41881 <= not w41299 and w41709;
w41882 <= not w41705 and w41881;
w41883 <= not w41706 and not w41709;
w41884 <= not w41882 and not w41883;
w41885 <= not w41781 and not w41884;
w41886 <= not w41289 and not w41780;
w41887 <= not w41779 and w41886;
w41888 <= not w41885 and not w41887;
w41889 <= not b(32) and not w41888;
w41890 <= not w41308 and w41704;
w41891 <= not w41700 and w41890;
w41892 <= not w41701 and not w41704;
w41893 <= not w41891 and not w41892;
w41894 <= not w41781 and not w41893;
w41895 <= not w41298 and not w41780;
w41896 <= not w41779 and w41895;
w41897 <= not w41894 and not w41896;
w41898 <= not b(31) and not w41897;
w41899 <= not w41317 and w41699;
w41900 <= not w41695 and w41899;
w41901 <= not w41696 and not w41699;
w41902 <= not w41900 and not w41901;
w41903 <= not w41781 and not w41902;
w41904 <= not w41307 and not w41780;
w41905 <= not w41779 and w41904;
w41906 <= not w41903 and not w41905;
w41907 <= not b(30) and not w41906;
w41908 <= not w41326 and w41694;
w41909 <= not w41690 and w41908;
w41910 <= not w41691 and not w41694;
w41911 <= not w41909 and not w41910;
w41912 <= not w41781 and not w41911;
w41913 <= not w41316 and not w41780;
w41914 <= not w41779 and w41913;
w41915 <= not w41912 and not w41914;
w41916 <= not b(29) and not w41915;
w41917 <= not w41335 and w41689;
w41918 <= not w41685 and w41917;
w41919 <= not w41686 and not w41689;
w41920 <= not w41918 and not w41919;
w41921 <= not w41781 and not w41920;
w41922 <= not w41325 and not w41780;
w41923 <= not w41779 and w41922;
w41924 <= not w41921 and not w41923;
w41925 <= not b(28) and not w41924;
w41926 <= not w41344 and w41684;
w41927 <= not w41680 and w41926;
w41928 <= not w41681 and not w41684;
w41929 <= not w41927 and not w41928;
w41930 <= not w41781 and not w41929;
w41931 <= not w41334 and not w41780;
w41932 <= not w41779 and w41931;
w41933 <= not w41930 and not w41932;
w41934 <= not b(27) and not w41933;
w41935 <= not w41353 and w41679;
w41936 <= not w41675 and w41935;
w41937 <= not w41676 and not w41679;
w41938 <= not w41936 and not w41937;
w41939 <= not w41781 and not w41938;
w41940 <= not w41343 and not w41780;
w41941 <= not w41779 and w41940;
w41942 <= not w41939 and not w41941;
w41943 <= not b(26) and not w41942;
w41944 <= not w41362 and w41674;
w41945 <= not w41670 and w41944;
w41946 <= not w41671 and not w41674;
w41947 <= not w41945 and not w41946;
w41948 <= not w41781 and not w41947;
w41949 <= not w41352 and not w41780;
w41950 <= not w41779 and w41949;
w41951 <= not w41948 and not w41950;
w41952 <= not b(25) and not w41951;
w41953 <= not w41371 and w41669;
w41954 <= not w41665 and w41953;
w41955 <= not w41666 and not w41669;
w41956 <= not w41954 and not w41955;
w41957 <= not w41781 and not w41956;
w41958 <= not w41361 and not w41780;
w41959 <= not w41779 and w41958;
w41960 <= not w41957 and not w41959;
w41961 <= not b(24) and not w41960;
w41962 <= not w41380 and w41664;
w41963 <= not w41660 and w41962;
w41964 <= not w41661 and not w41664;
w41965 <= not w41963 and not w41964;
w41966 <= not w41781 and not w41965;
w41967 <= not w41370 and not w41780;
w41968 <= not w41779 and w41967;
w41969 <= not w41966 and not w41968;
w41970 <= not b(23) and not w41969;
w41971 <= not w41389 and w41659;
w41972 <= not w41655 and w41971;
w41973 <= not w41656 and not w41659;
w41974 <= not w41972 and not w41973;
w41975 <= not w41781 and not w41974;
w41976 <= not w41379 and not w41780;
w41977 <= not w41779 and w41976;
w41978 <= not w41975 and not w41977;
w41979 <= not b(22) and not w41978;
w41980 <= not w41398 and w41654;
w41981 <= not w41650 and w41980;
w41982 <= not w41651 and not w41654;
w41983 <= not w41981 and not w41982;
w41984 <= not w41781 and not w41983;
w41985 <= not w41388 and not w41780;
w41986 <= not w41779 and w41985;
w41987 <= not w41984 and not w41986;
w41988 <= not b(21) and not w41987;
w41989 <= not w41407 and w41649;
w41990 <= not w41645 and w41989;
w41991 <= not w41646 and not w41649;
w41992 <= not w41990 and not w41991;
w41993 <= not w41781 and not w41992;
w41994 <= not w41397 and not w41780;
w41995 <= not w41779 and w41994;
w41996 <= not w41993 and not w41995;
w41997 <= not b(20) and not w41996;
w41998 <= not w41416 and w41644;
w41999 <= not w41640 and w41998;
w42000 <= not w41641 and not w41644;
w42001 <= not w41999 and not w42000;
w42002 <= not w41781 and not w42001;
w42003 <= not w41406 and not w41780;
w42004 <= not w41779 and w42003;
w42005 <= not w42002 and not w42004;
w42006 <= not b(19) and not w42005;
w42007 <= not w41425 and w41639;
w42008 <= not w41635 and w42007;
w42009 <= not w41636 and not w41639;
w42010 <= not w42008 and not w42009;
w42011 <= not w41781 and not w42010;
w42012 <= not w41415 and not w41780;
w42013 <= not w41779 and w42012;
w42014 <= not w42011 and not w42013;
w42015 <= not b(18) and not w42014;
w42016 <= not w41434 and w41634;
w42017 <= not w41630 and w42016;
w42018 <= not w41631 and not w41634;
w42019 <= not w42017 and not w42018;
w42020 <= not w41781 and not w42019;
w42021 <= not w41424 and not w41780;
w42022 <= not w41779 and w42021;
w42023 <= not w42020 and not w42022;
w42024 <= not b(17) and not w42023;
w42025 <= not w41443 and w41629;
w42026 <= not w41625 and w42025;
w42027 <= not w41626 and not w41629;
w42028 <= not w42026 and not w42027;
w42029 <= not w41781 and not w42028;
w42030 <= not w41433 and not w41780;
w42031 <= not w41779 and w42030;
w42032 <= not w42029 and not w42031;
w42033 <= not b(16) and not w42032;
w42034 <= not w41452 and w41624;
w42035 <= not w41620 and w42034;
w42036 <= not w41621 and not w41624;
w42037 <= not w42035 and not w42036;
w42038 <= not w41781 and not w42037;
w42039 <= not w41442 and not w41780;
w42040 <= not w41779 and w42039;
w42041 <= not w42038 and not w42040;
w42042 <= not b(15) and not w42041;
w42043 <= not w41461 and w41619;
w42044 <= not w41615 and w42043;
w42045 <= not w41616 and not w41619;
w42046 <= not w42044 and not w42045;
w42047 <= not w41781 and not w42046;
w42048 <= not w41451 and not w41780;
w42049 <= not w41779 and w42048;
w42050 <= not w42047 and not w42049;
w42051 <= not b(14) and not w42050;
w42052 <= not w41470 and w41614;
w42053 <= not w41610 and w42052;
w42054 <= not w41611 and not w41614;
w42055 <= not w42053 and not w42054;
w42056 <= not w41781 and not w42055;
w42057 <= not w41460 and not w41780;
w42058 <= not w41779 and w42057;
w42059 <= not w42056 and not w42058;
w42060 <= not b(13) and not w42059;
w42061 <= not w41479 and w41609;
w42062 <= not w41605 and w42061;
w42063 <= not w41606 and not w41609;
w42064 <= not w42062 and not w42063;
w42065 <= not w41781 and not w42064;
w42066 <= not w41469 and not w41780;
w42067 <= not w41779 and w42066;
w42068 <= not w42065 and not w42067;
w42069 <= not b(12) and not w42068;
w42070 <= not w41488 and w41604;
w42071 <= not w41600 and w42070;
w42072 <= not w41601 and not w41604;
w42073 <= not w42071 and not w42072;
w42074 <= not w41781 and not w42073;
w42075 <= not w41478 and not w41780;
w42076 <= not w41779 and w42075;
w42077 <= not w42074 and not w42076;
w42078 <= not b(11) and not w42077;
w42079 <= not w41497 and w41599;
w42080 <= not w41595 and w42079;
w42081 <= not w41596 and not w41599;
w42082 <= not w42080 and not w42081;
w42083 <= not w41781 and not w42082;
w42084 <= not w41487 and not w41780;
w42085 <= not w41779 and w42084;
w42086 <= not w42083 and not w42085;
w42087 <= not b(10) and not w42086;
w42088 <= not w41506 and w41594;
w42089 <= not w41590 and w42088;
w42090 <= not w41591 and not w41594;
w42091 <= not w42089 and not w42090;
w42092 <= not w41781 and not w42091;
w42093 <= not w41496 and not w41780;
w42094 <= not w41779 and w42093;
w42095 <= not w42092 and not w42094;
w42096 <= not b(9) and not w42095;
w42097 <= not w41515 and w41589;
w42098 <= not w41585 and w42097;
w42099 <= not w41586 and not w41589;
w42100 <= not w42098 and not w42099;
w42101 <= not w41781 and not w42100;
w42102 <= not w41505 and not w41780;
w42103 <= not w41779 and w42102;
w42104 <= not w42101 and not w42103;
w42105 <= not b(8) and not w42104;
w42106 <= not w41524 and w41584;
w42107 <= not w41580 and w42106;
w42108 <= not w41581 and not w41584;
w42109 <= not w42107 and not w42108;
w42110 <= not w41781 and not w42109;
w42111 <= not w41514 and not w41780;
w42112 <= not w41779 and w42111;
w42113 <= not w42110 and not w42112;
w42114 <= not b(7) and not w42113;
w42115 <= not w41533 and w41579;
w42116 <= not w41575 and w42115;
w42117 <= not w41576 and not w41579;
w42118 <= not w42116 and not w42117;
w42119 <= not w41781 and not w42118;
w42120 <= not w41523 and not w41780;
w42121 <= not w41779 and w42120;
w42122 <= not w42119 and not w42121;
w42123 <= not b(6) and not w42122;
w42124 <= not w41542 and w41574;
w42125 <= not w41570 and w42124;
w42126 <= not w41571 and not w41574;
w42127 <= not w42125 and not w42126;
w42128 <= not w41781 and not w42127;
w42129 <= not w41532 and not w41780;
w42130 <= not w41779 and w42129;
w42131 <= not w42128 and not w42130;
w42132 <= not b(5) and not w42131;
w42133 <= not w41550 and w41569;
w42134 <= not w41565 and w42133;
w42135 <= not w41566 and not w41569;
w42136 <= not w42134 and not w42135;
w42137 <= not w41781 and not w42136;
w42138 <= not w41541 and not w41780;
w42139 <= not w41779 and w42138;
w42140 <= not w42137 and not w42139;
w42141 <= not b(4) and not w42140;
w42142 <= not w41560 and w41564;
w42143 <= not w41559 and w42142;
w42144 <= not w41561 and not w41564;
w42145 <= not w42143 and not w42144;
w42146 <= not w41781 and not w42145;
w42147 <= not w41549 and not w41780;
w42148 <= not w41779 and w42147;
w42149 <= not w42146 and not w42148;
w42150 <= not b(3) and not w42149;
w42151 <= w13482 and not w41557;
w42152 <= not w41555 and w42151;
w42153 <= not w41559 and not w42152;
w42154 <= not w41781 and w42153;
w42155 <= not w41554 and not w41780;
w42156 <= not w41779 and w42155;
w42157 <= not w42154 and not w42156;
w42158 <= not b(2) and not w42157;
w42159 <= b(0) and not w41781;
w42160 <= a(20) and not w42159;
w42161 <= w13482 and not w41781;
w42162 <= not w42160 and not w42161;
w42163 <= b(1) and not w42162;
w42164 <= not b(1) and not w42161;
w42165 <= not w42160 and w42164;
w42166 <= not w42163 and not w42165;
w42167 <= not w14092 and not w42166;
w42168 <= not b(1) and not w42162;
w42169 <= not w42167 and not w42168;
w42170 <= b(2) and not w42156;
w42171 <= not w42154 and w42170;
w42172 <= not w42158 and not w42171;
w42173 <= not w42169 and w42172;
w42174 <= not w42158 and not w42173;
w42175 <= b(3) and not w42148;
w42176 <= not w42146 and w42175;
w42177 <= not w42150 and not w42176;
w42178 <= not w42174 and w42177;
w42179 <= not w42150 and not w42178;
w42180 <= b(4) and not w42139;
w42181 <= not w42137 and w42180;
w42182 <= not w42141 and not w42181;
w42183 <= not w42179 and w42182;
w42184 <= not w42141 and not w42183;
w42185 <= b(5) and not w42130;
w42186 <= not w42128 and w42185;
w42187 <= not w42132 and not w42186;
w42188 <= not w42184 and w42187;
w42189 <= not w42132 and not w42188;
w42190 <= b(6) and not w42121;
w42191 <= not w42119 and w42190;
w42192 <= not w42123 and not w42191;
w42193 <= not w42189 and w42192;
w42194 <= not w42123 and not w42193;
w42195 <= b(7) and not w42112;
w42196 <= not w42110 and w42195;
w42197 <= not w42114 and not w42196;
w42198 <= not w42194 and w42197;
w42199 <= not w42114 and not w42198;
w42200 <= b(8) and not w42103;
w42201 <= not w42101 and w42200;
w42202 <= not w42105 and not w42201;
w42203 <= not w42199 and w42202;
w42204 <= not w42105 and not w42203;
w42205 <= b(9) and not w42094;
w42206 <= not w42092 and w42205;
w42207 <= not w42096 and not w42206;
w42208 <= not w42204 and w42207;
w42209 <= not w42096 and not w42208;
w42210 <= b(10) and not w42085;
w42211 <= not w42083 and w42210;
w42212 <= not w42087 and not w42211;
w42213 <= not w42209 and w42212;
w42214 <= not w42087 and not w42213;
w42215 <= b(11) and not w42076;
w42216 <= not w42074 and w42215;
w42217 <= not w42078 and not w42216;
w42218 <= not w42214 and w42217;
w42219 <= not w42078 and not w42218;
w42220 <= b(12) and not w42067;
w42221 <= not w42065 and w42220;
w42222 <= not w42069 and not w42221;
w42223 <= not w42219 and w42222;
w42224 <= not w42069 and not w42223;
w42225 <= b(13) and not w42058;
w42226 <= not w42056 and w42225;
w42227 <= not w42060 and not w42226;
w42228 <= not w42224 and w42227;
w42229 <= not w42060 and not w42228;
w42230 <= b(14) and not w42049;
w42231 <= not w42047 and w42230;
w42232 <= not w42051 and not w42231;
w42233 <= not w42229 and w42232;
w42234 <= not w42051 and not w42233;
w42235 <= b(15) and not w42040;
w42236 <= not w42038 and w42235;
w42237 <= not w42042 and not w42236;
w42238 <= not w42234 and w42237;
w42239 <= not w42042 and not w42238;
w42240 <= b(16) and not w42031;
w42241 <= not w42029 and w42240;
w42242 <= not w42033 and not w42241;
w42243 <= not w42239 and w42242;
w42244 <= not w42033 and not w42243;
w42245 <= b(17) and not w42022;
w42246 <= not w42020 and w42245;
w42247 <= not w42024 and not w42246;
w42248 <= not w42244 and w42247;
w42249 <= not w42024 and not w42248;
w42250 <= b(18) and not w42013;
w42251 <= not w42011 and w42250;
w42252 <= not w42015 and not w42251;
w42253 <= not w42249 and w42252;
w42254 <= not w42015 and not w42253;
w42255 <= b(19) and not w42004;
w42256 <= not w42002 and w42255;
w42257 <= not w42006 and not w42256;
w42258 <= not w42254 and w42257;
w42259 <= not w42006 and not w42258;
w42260 <= b(20) and not w41995;
w42261 <= not w41993 and w42260;
w42262 <= not w41997 and not w42261;
w42263 <= not w42259 and w42262;
w42264 <= not w41997 and not w42263;
w42265 <= b(21) and not w41986;
w42266 <= not w41984 and w42265;
w42267 <= not w41988 and not w42266;
w42268 <= not w42264 and w42267;
w42269 <= not w41988 and not w42268;
w42270 <= b(22) and not w41977;
w42271 <= not w41975 and w42270;
w42272 <= not w41979 and not w42271;
w42273 <= not w42269 and w42272;
w42274 <= not w41979 and not w42273;
w42275 <= b(23) and not w41968;
w42276 <= not w41966 and w42275;
w42277 <= not w41970 and not w42276;
w42278 <= not w42274 and w42277;
w42279 <= not w41970 and not w42278;
w42280 <= b(24) and not w41959;
w42281 <= not w41957 and w42280;
w42282 <= not w41961 and not w42281;
w42283 <= not w42279 and w42282;
w42284 <= not w41961 and not w42283;
w42285 <= b(25) and not w41950;
w42286 <= not w41948 and w42285;
w42287 <= not w41952 and not w42286;
w42288 <= not w42284 and w42287;
w42289 <= not w41952 and not w42288;
w42290 <= b(26) and not w41941;
w42291 <= not w41939 and w42290;
w42292 <= not w41943 and not w42291;
w42293 <= not w42289 and w42292;
w42294 <= not w41943 and not w42293;
w42295 <= b(27) and not w41932;
w42296 <= not w41930 and w42295;
w42297 <= not w41934 and not w42296;
w42298 <= not w42294 and w42297;
w42299 <= not w41934 and not w42298;
w42300 <= b(28) and not w41923;
w42301 <= not w41921 and w42300;
w42302 <= not w41925 and not w42301;
w42303 <= not w42299 and w42302;
w42304 <= not w41925 and not w42303;
w42305 <= b(29) and not w41914;
w42306 <= not w41912 and w42305;
w42307 <= not w41916 and not w42306;
w42308 <= not w42304 and w42307;
w42309 <= not w41916 and not w42308;
w42310 <= b(30) and not w41905;
w42311 <= not w41903 and w42310;
w42312 <= not w41907 and not w42311;
w42313 <= not w42309 and w42312;
w42314 <= not w41907 and not w42313;
w42315 <= b(31) and not w41896;
w42316 <= not w41894 and w42315;
w42317 <= not w41898 and not w42316;
w42318 <= not w42314 and w42317;
w42319 <= not w41898 and not w42318;
w42320 <= b(32) and not w41887;
w42321 <= not w41885 and w42320;
w42322 <= not w41889 and not w42321;
w42323 <= not w42319 and w42322;
w42324 <= not w41889 and not w42323;
w42325 <= b(33) and not w41878;
w42326 <= not w41876 and w42325;
w42327 <= not w41880 and not w42326;
w42328 <= not w42324 and w42327;
w42329 <= not w41880 and not w42328;
w42330 <= b(34) and not w41869;
w42331 <= not w41867 and w42330;
w42332 <= not w41871 and not w42331;
w42333 <= not w42329 and w42332;
w42334 <= not w41871 and not w42333;
w42335 <= b(35) and not w41860;
w42336 <= not w41858 and w42335;
w42337 <= not w41862 and not w42336;
w42338 <= not w42334 and w42337;
w42339 <= not w41862 and not w42338;
w42340 <= b(36) and not w41851;
w42341 <= not w41849 and w42340;
w42342 <= not w41853 and not w42341;
w42343 <= not w42339 and w42342;
w42344 <= not w41853 and not w42343;
w42345 <= b(37) and not w41842;
w42346 <= not w41840 and w42345;
w42347 <= not w41844 and not w42346;
w42348 <= not w42344 and w42347;
w42349 <= not w41844 and not w42348;
w42350 <= b(38) and not w41833;
w42351 <= not w41831 and w42350;
w42352 <= not w41835 and not w42351;
w42353 <= not w42349 and w42352;
w42354 <= not w41835 and not w42353;
w42355 <= b(39) and not w41824;
w42356 <= not w41822 and w42355;
w42357 <= not w41826 and not w42356;
w42358 <= not w42354 and w42357;
w42359 <= not w41826 and not w42358;
w42360 <= b(40) and not w41815;
w42361 <= not w41813 and w42360;
w42362 <= not w41817 and not w42361;
w42363 <= not w42359 and w42362;
w42364 <= not w41817 and not w42363;
w42365 <= b(41) and not w41806;
w42366 <= not w41804 and w42365;
w42367 <= not w41808 and not w42366;
w42368 <= not w42364 and w42367;
w42369 <= not w41808 and not w42368;
w42370 <= b(42) and not w41797;
w42371 <= not w41795 and w42370;
w42372 <= not w41799 and not w42371;
w42373 <= not w42369 and w42372;
w42374 <= not w41799 and not w42373;
w42375 <= b(43) and not w41788;
w42376 <= not w41786 and w42375;
w42377 <= not w41790 and not w42376;
w42378 <= not w42374 and w42377;
w42379 <= not w41790 and not w42378;
w42380 <= not w41191 and not w41776;
w42381 <= not w41774 and w42380;
w42382 <= not w41765 and w42381;
w42383 <= not w41774 and not w41776;
w42384 <= not w41766 and not w42383;
w42385 <= not w42382 and not w42384;
w42386 <= not w41781 and not w42385;
w42387 <= not w41773 and not w41780;
w42388 <= not w41779 and w42387;
w42389 <= not w42386 and not w42388;
w42390 <= not b(44) and not w42389;
w42391 <= b(44) and not w42388;
w42392 <= not w42386 and w42391;
w42393 <= w14319 and not w42392;
w42394 <= not w42390 and w42393;
w42395 <= not w42379 and w42394;
w42396 <= w13701 and not w42389;
w42397 <= not w42395 and not w42396;
w42398 <= not w41799 and w42377;
w42399 <= not w42373 and w42398;
w42400 <= not w42374 and not w42377;
w42401 <= not w42399 and not w42400;
w42402 <= not w42397 and not w42401;
w42403 <= not w41789 and not w42396;
w42404 <= not w42395 and w42403;
w42405 <= not w42402 and not w42404;
w42406 <= not w41790 and not w42392;
w42407 <= not w42390 and w42406;
w42408 <= not w42378 and w42407;
w42409 <= not w42390 and not w42392;
w42410 <= not w42379 and not w42409;
w42411 <= not w42408 and not w42410;
w42412 <= not w42397 and not w42411;
w42413 <= not w42389 and not w42396;
w42414 <= not w42395 and w42413;
w42415 <= not w42412 and not w42414;
w42416 <= not b(45) and not w42415;
w42417 <= not b(44) and not w42405;
w42418 <= not w41808 and w42372;
w42419 <= not w42368 and w42418;
w42420 <= not w42369 and not w42372;
w42421 <= not w42419 and not w42420;
w42422 <= not w42397 and not w42421;
w42423 <= not w41798 and not w42396;
w42424 <= not w42395 and w42423;
w42425 <= not w42422 and not w42424;
w42426 <= not b(43) and not w42425;
w42427 <= not w41817 and w42367;
w42428 <= not w42363 and w42427;
w42429 <= not w42364 and not w42367;
w42430 <= not w42428 and not w42429;
w42431 <= not w42397 and not w42430;
w42432 <= not w41807 and not w42396;
w42433 <= not w42395 and w42432;
w42434 <= not w42431 and not w42433;
w42435 <= not b(42) and not w42434;
w42436 <= not w41826 and w42362;
w42437 <= not w42358 and w42436;
w42438 <= not w42359 and not w42362;
w42439 <= not w42437 and not w42438;
w42440 <= not w42397 and not w42439;
w42441 <= not w41816 and not w42396;
w42442 <= not w42395 and w42441;
w42443 <= not w42440 and not w42442;
w42444 <= not b(41) and not w42443;
w42445 <= not w41835 and w42357;
w42446 <= not w42353 and w42445;
w42447 <= not w42354 and not w42357;
w42448 <= not w42446 and not w42447;
w42449 <= not w42397 and not w42448;
w42450 <= not w41825 and not w42396;
w42451 <= not w42395 and w42450;
w42452 <= not w42449 and not w42451;
w42453 <= not b(40) and not w42452;
w42454 <= not w41844 and w42352;
w42455 <= not w42348 and w42454;
w42456 <= not w42349 and not w42352;
w42457 <= not w42455 and not w42456;
w42458 <= not w42397 and not w42457;
w42459 <= not w41834 and not w42396;
w42460 <= not w42395 and w42459;
w42461 <= not w42458 and not w42460;
w42462 <= not b(39) and not w42461;
w42463 <= not w41853 and w42347;
w42464 <= not w42343 and w42463;
w42465 <= not w42344 and not w42347;
w42466 <= not w42464 and not w42465;
w42467 <= not w42397 and not w42466;
w42468 <= not w41843 and not w42396;
w42469 <= not w42395 and w42468;
w42470 <= not w42467 and not w42469;
w42471 <= not b(38) and not w42470;
w42472 <= not w41862 and w42342;
w42473 <= not w42338 and w42472;
w42474 <= not w42339 and not w42342;
w42475 <= not w42473 and not w42474;
w42476 <= not w42397 and not w42475;
w42477 <= not w41852 and not w42396;
w42478 <= not w42395 and w42477;
w42479 <= not w42476 and not w42478;
w42480 <= not b(37) and not w42479;
w42481 <= not w41871 and w42337;
w42482 <= not w42333 and w42481;
w42483 <= not w42334 and not w42337;
w42484 <= not w42482 and not w42483;
w42485 <= not w42397 and not w42484;
w42486 <= not w41861 and not w42396;
w42487 <= not w42395 and w42486;
w42488 <= not w42485 and not w42487;
w42489 <= not b(36) and not w42488;
w42490 <= not w41880 and w42332;
w42491 <= not w42328 and w42490;
w42492 <= not w42329 and not w42332;
w42493 <= not w42491 and not w42492;
w42494 <= not w42397 and not w42493;
w42495 <= not w41870 and not w42396;
w42496 <= not w42395 and w42495;
w42497 <= not w42494 and not w42496;
w42498 <= not b(35) and not w42497;
w42499 <= not w41889 and w42327;
w42500 <= not w42323 and w42499;
w42501 <= not w42324 and not w42327;
w42502 <= not w42500 and not w42501;
w42503 <= not w42397 and not w42502;
w42504 <= not w41879 and not w42396;
w42505 <= not w42395 and w42504;
w42506 <= not w42503 and not w42505;
w42507 <= not b(34) and not w42506;
w42508 <= not w41898 and w42322;
w42509 <= not w42318 and w42508;
w42510 <= not w42319 and not w42322;
w42511 <= not w42509 and not w42510;
w42512 <= not w42397 and not w42511;
w42513 <= not w41888 and not w42396;
w42514 <= not w42395 and w42513;
w42515 <= not w42512 and not w42514;
w42516 <= not b(33) and not w42515;
w42517 <= not w41907 and w42317;
w42518 <= not w42313 and w42517;
w42519 <= not w42314 and not w42317;
w42520 <= not w42518 and not w42519;
w42521 <= not w42397 and not w42520;
w42522 <= not w41897 and not w42396;
w42523 <= not w42395 and w42522;
w42524 <= not w42521 and not w42523;
w42525 <= not b(32) and not w42524;
w42526 <= not w41916 and w42312;
w42527 <= not w42308 and w42526;
w42528 <= not w42309 and not w42312;
w42529 <= not w42527 and not w42528;
w42530 <= not w42397 and not w42529;
w42531 <= not w41906 and not w42396;
w42532 <= not w42395 and w42531;
w42533 <= not w42530 and not w42532;
w42534 <= not b(31) and not w42533;
w42535 <= not w41925 and w42307;
w42536 <= not w42303 and w42535;
w42537 <= not w42304 and not w42307;
w42538 <= not w42536 and not w42537;
w42539 <= not w42397 and not w42538;
w42540 <= not w41915 and not w42396;
w42541 <= not w42395 and w42540;
w42542 <= not w42539 and not w42541;
w42543 <= not b(30) and not w42542;
w42544 <= not w41934 and w42302;
w42545 <= not w42298 and w42544;
w42546 <= not w42299 and not w42302;
w42547 <= not w42545 and not w42546;
w42548 <= not w42397 and not w42547;
w42549 <= not w41924 and not w42396;
w42550 <= not w42395 and w42549;
w42551 <= not w42548 and not w42550;
w42552 <= not b(29) and not w42551;
w42553 <= not w41943 and w42297;
w42554 <= not w42293 and w42553;
w42555 <= not w42294 and not w42297;
w42556 <= not w42554 and not w42555;
w42557 <= not w42397 and not w42556;
w42558 <= not w41933 and not w42396;
w42559 <= not w42395 and w42558;
w42560 <= not w42557 and not w42559;
w42561 <= not b(28) and not w42560;
w42562 <= not w41952 and w42292;
w42563 <= not w42288 and w42562;
w42564 <= not w42289 and not w42292;
w42565 <= not w42563 and not w42564;
w42566 <= not w42397 and not w42565;
w42567 <= not w41942 and not w42396;
w42568 <= not w42395 and w42567;
w42569 <= not w42566 and not w42568;
w42570 <= not b(27) and not w42569;
w42571 <= not w41961 and w42287;
w42572 <= not w42283 and w42571;
w42573 <= not w42284 and not w42287;
w42574 <= not w42572 and not w42573;
w42575 <= not w42397 and not w42574;
w42576 <= not w41951 and not w42396;
w42577 <= not w42395 and w42576;
w42578 <= not w42575 and not w42577;
w42579 <= not b(26) and not w42578;
w42580 <= not w41970 and w42282;
w42581 <= not w42278 and w42580;
w42582 <= not w42279 and not w42282;
w42583 <= not w42581 and not w42582;
w42584 <= not w42397 and not w42583;
w42585 <= not w41960 and not w42396;
w42586 <= not w42395 and w42585;
w42587 <= not w42584 and not w42586;
w42588 <= not b(25) and not w42587;
w42589 <= not w41979 and w42277;
w42590 <= not w42273 and w42589;
w42591 <= not w42274 and not w42277;
w42592 <= not w42590 and not w42591;
w42593 <= not w42397 and not w42592;
w42594 <= not w41969 and not w42396;
w42595 <= not w42395 and w42594;
w42596 <= not w42593 and not w42595;
w42597 <= not b(24) and not w42596;
w42598 <= not w41988 and w42272;
w42599 <= not w42268 and w42598;
w42600 <= not w42269 and not w42272;
w42601 <= not w42599 and not w42600;
w42602 <= not w42397 and not w42601;
w42603 <= not w41978 and not w42396;
w42604 <= not w42395 and w42603;
w42605 <= not w42602 and not w42604;
w42606 <= not b(23) and not w42605;
w42607 <= not w41997 and w42267;
w42608 <= not w42263 and w42607;
w42609 <= not w42264 and not w42267;
w42610 <= not w42608 and not w42609;
w42611 <= not w42397 and not w42610;
w42612 <= not w41987 and not w42396;
w42613 <= not w42395 and w42612;
w42614 <= not w42611 and not w42613;
w42615 <= not b(22) and not w42614;
w42616 <= not w42006 and w42262;
w42617 <= not w42258 and w42616;
w42618 <= not w42259 and not w42262;
w42619 <= not w42617 and not w42618;
w42620 <= not w42397 and not w42619;
w42621 <= not w41996 and not w42396;
w42622 <= not w42395 and w42621;
w42623 <= not w42620 and not w42622;
w42624 <= not b(21) and not w42623;
w42625 <= not w42015 and w42257;
w42626 <= not w42253 and w42625;
w42627 <= not w42254 and not w42257;
w42628 <= not w42626 and not w42627;
w42629 <= not w42397 and not w42628;
w42630 <= not w42005 and not w42396;
w42631 <= not w42395 and w42630;
w42632 <= not w42629 and not w42631;
w42633 <= not b(20) and not w42632;
w42634 <= not w42024 and w42252;
w42635 <= not w42248 and w42634;
w42636 <= not w42249 and not w42252;
w42637 <= not w42635 and not w42636;
w42638 <= not w42397 and not w42637;
w42639 <= not w42014 and not w42396;
w42640 <= not w42395 and w42639;
w42641 <= not w42638 and not w42640;
w42642 <= not b(19) and not w42641;
w42643 <= not w42033 and w42247;
w42644 <= not w42243 and w42643;
w42645 <= not w42244 and not w42247;
w42646 <= not w42644 and not w42645;
w42647 <= not w42397 and not w42646;
w42648 <= not w42023 and not w42396;
w42649 <= not w42395 and w42648;
w42650 <= not w42647 and not w42649;
w42651 <= not b(18) and not w42650;
w42652 <= not w42042 and w42242;
w42653 <= not w42238 and w42652;
w42654 <= not w42239 and not w42242;
w42655 <= not w42653 and not w42654;
w42656 <= not w42397 and not w42655;
w42657 <= not w42032 and not w42396;
w42658 <= not w42395 and w42657;
w42659 <= not w42656 and not w42658;
w42660 <= not b(17) and not w42659;
w42661 <= not w42051 and w42237;
w42662 <= not w42233 and w42661;
w42663 <= not w42234 and not w42237;
w42664 <= not w42662 and not w42663;
w42665 <= not w42397 and not w42664;
w42666 <= not w42041 and not w42396;
w42667 <= not w42395 and w42666;
w42668 <= not w42665 and not w42667;
w42669 <= not b(16) and not w42668;
w42670 <= not w42060 and w42232;
w42671 <= not w42228 and w42670;
w42672 <= not w42229 and not w42232;
w42673 <= not w42671 and not w42672;
w42674 <= not w42397 and not w42673;
w42675 <= not w42050 and not w42396;
w42676 <= not w42395 and w42675;
w42677 <= not w42674 and not w42676;
w42678 <= not b(15) and not w42677;
w42679 <= not w42069 and w42227;
w42680 <= not w42223 and w42679;
w42681 <= not w42224 and not w42227;
w42682 <= not w42680 and not w42681;
w42683 <= not w42397 and not w42682;
w42684 <= not w42059 and not w42396;
w42685 <= not w42395 and w42684;
w42686 <= not w42683 and not w42685;
w42687 <= not b(14) and not w42686;
w42688 <= not w42078 and w42222;
w42689 <= not w42218 and w42688;
w42690 <= not w42219 and not w42222;
w42691 <= not w42689 and not w42690;
w42692 <= not w42397 and not w42691;
w42693 <= not w42068 and not w42396;
w42694 <= not w42395 and w42693;
w42695 <= not w42692 and not w42694;
w42696 <= not b(13) and not w42695;
w42697 <= not w42087 and w42217;
w42698 <= not w42213 and w42697;
w42699 <= not w42214 and not w42217;
w42700 <= not w42698 and not w42699;
w42701 <= not w42397 and not w42700;
w42702 <= not w42077 and not w42396;
w42703 <= not w42395 and w42702;
w42704 <= not w42701 and not w42703;
w42705 <= not b(12) and not w42704;
w42706 <= not w42096 and w42212;
w42707 <= not w42208 and w42706;
w42708 <= not w42209 and not w42212;
w42709 <= not w42707 and not w42708;
w42710 <= not w42397 and not w42709;
w42711 <= not w42086 and not w42396;
w42712 <= not w42395 and w42711;
w42713 <= not w42710 and not w42712;
w42714 <= not b(11) and not w42713;
w42715 <= not w42105 and w42207;
w42716 <= not w42203 and w42715;
w42717 <= not w42204 and not w42207;
w42718 <= not w42716 and not w42717;
w42719 <= not w42397 and not w42718;
w42720 <= not w42095 and not w42396;
w42721 <= not w42395 and w42720;
w42722 <= not w42719 and not w42721;
w42723 <= not b(10) and not w42722;
w42724 <= not w42114 and w42202;
w42725 <= not w42198 and w42724;
w42726 <= not w42199 and not w42202;
w42727 <= not w42725 and not w42726;
w42728 <= not w42397 and not w42727;
w42729 <= not w42104 and not w42396;
w42730 <= not w42395 and w42729;
w42731 <= not w42728 and not w42730;
w42732 <= not b(9) and not w42731;
w42733 <= not w42123 and w42197;
w42734 <= not w42193 and w42733;
w42735 <= not w42194 and not w42197;
w42736 <= not w42734 and not w42735;
w42737 <= not w42397 and not w42736;
w42738 <= not w42113 and not w42396;
w42739 <= not w42395 and w42738;
w42740 <= not w42737 and not w42739;
w42741 <= not b(8) and not w42740;
w42742 <= not w42132 and w42192;
w42743 <= not w42188 and w42742;
w42744 <= not w42189 and not w42192;
w42745 <= not w42743 and not w42744;
w42746 <= not w42397 and not w42745;
w42747 <= not w42122 and not w42396;
w42748 <= not w42395 and w42747;
w42749 <= not w42746 and not w42748;
w42750 <= not b(7) and not w42749;
w42751 <= not w42141 and w42187;
w42752 <= not w42183 and w42751;
w42753 <= not w42184 and not w42187;
w42754 <= not w42752 and not w42753;
w42755 <= not w42397 and not w42754;
w42756 <= not w42131 and not w42396;
w42757 <= not w42395 and w42756;
w42758 <= not w42755 and not w42757;
w42759 <= not b(6) and not w42758;
w42760 <= not w42150 and w42182;
w42761 <= not w42178 and w42760;
w42762 <= not w42179 and not w42182;
w42763 <= not w42761 and not w42762;
w42764 <= not w42397 and not w42763;
w42765 <= not w42140 and not w42396;
w42766 <= not w42395 and w42765;
w42767 <= not w42764 and not w42766;
w42768 <= not b(5) and not w42767;
w42769 <= not w42158 and w42177;
w42770 <= not w42173 and w42769;
w42771 <= not w42174 and not w42177;
w42772 <= not w42770 and not w42771;
w42773 <= not w42397 and not w42772;
w42774 <= not w42149 and not w42396;
w42775 <= not w42395 and w42774;
w42776 <= not w42773 and not w42775;
w42777 <= not b(4) and not w42776;
w42778 <= not w42168 and w42172;
w42779 <= not w42167 and w42778;
w42780 <= not w42169 and not w42172;
w42781 <= not w42779 and not w42780;
w42782 <= not w42397 and not w42781;
w42783 <= not w42157 and not w42396;
w42784 <= not w42395 and w42783;
w42785 <= not w42782 and not w42784;
w42786 <= not b(3) and not w42785;
w42787 <= w14092 and not w42165;
w42788 <= not w42163 and w42787;
w42789 <= not w42167 and not w42788;
w42790 <= not w42397 and w42789;
w42791 <= not w42162 and not w42396;
w42792 <= not w42395 and w42791;
w42793 <= not w42790 and not w42792;
w42794 <= not b(2) and not w42793;
w42795 <= b(0) and not w42397;
w42796 <= a(19) and not w42795;
w42797 <= w14092 and not w42397;
w42798 <= not w42796 and not w42797;
w42799 <= b(1) and not w42798;
w42800 <= not b(1) and not w42797;
w42801 <= not w42796 and w42800;
w42802 <= not w42799 and not w42801;
w42803 <= not w14730 and not w42802;
w42804 <= not b(1) and not w42798;
w42805 <= not w42803 and not w42804;
w42806 <= b(2) and not w42792;
w42807 <= not w42790 and w42806;
w42808 <= not w42794 and not w42807;
w42809 <= not w42805 and w42808;
w42810 <= not w42794 and not w42809;
w42811 <= b(3) and not w42784;
w42812 <= not w42782 and w42811;
w42813 <= not w42786 and not w42812;
w42814 <= not w42810 and w42813;
w42815 <= not w42786 and not w42814;
w42816 <= b(4) and not w42775;
w42817 <= not w42773 and w42816;
w42818 <= not w42777 and not w42817;
w42819 <= not w42815 and w42818;
w42820 <= not w42777 and not w42819;
w42821 <= b(5) and not w42766;
w42822 <= not w42764 and w42821;
w42823 <= not w42768 and not w42822;
w42824 <= not w42820 and w42823;
w42825 <= not w42768 and not w42824;
w42826 <= b(6) and not w42757;
w42827 <= not w42755 and w42826;
w42828 <= not w42759 and not w42827;
w42829 <= not w42825 and w42828;
w42830 <= not w42759 and not w42829;
w42831 <= b(7) and not w42748;
w42832 <= not w42746 and w42831;
w42833 <= not w42750 and not w42832;
w42834 <= not w42830 and w42833;
w42835 <= not w42750 and not w42834;
w42836 <= b(8) and not w42739;
w42837 <= not w42737 and w42836;
w42838 <= not w42741 and not w42837;
w42839 <= not w42835 and w42838;
w42840 <= not w42741 and not w42839;
w42841 <= b(9) and not w42730;
w42842 <= not w42728 and w42841;
w42843 <= not w42732 and not w42842;
w42844 <= not w42840 and w42843;
w42845 <= not w42732 and not w42844;
w42846 <= b(10) and not w42721;
w42847 <= not w42719 and w42846;
w42848 <= not w42723 and not w42847;
w42849 <= not w42845 and w42848;
w42850 <= not w42723 and not w42849;
w42851 <= b(11) and not w42712;
w42852 <= not w42710 and w42851;
w42853 <= not w42714 and not w42852;
w42854 <= not w42850 and w42853;
w42855 <= not w42714 and not w42854;
w42856 <= b(12) and not w42703;
w42857 <= not w42701 and w42856;
w42858 <= not w42705 and not w42857;
w42859 <= not w42855 and w42858;
w42860 <= not w42705 and not w42859;
w42861 <= b(13) and not w42694;
w42862 <= not w42692 and w42861;
w42863 <= not w42696 and not w42862;
w42864 <= not w42860 and w42863;
w42865 <= not w42696 and not w42864;
w42866 <= b(14) and not w42685;
w42867 <= not w42683 and w42866;
w42868 <= not w42687 and not w42867;
w42869 <= not w42865 and w42868;
w42870 <= not w42687 and not w42869;
w42871 <= b(15) and not w42676;
w42872 <= not w42674 and w42871;
w42873 <= not w42678 and not w42872;
w42874 <= not w42870 and w42873;
w42875 <= not w42678 and not w42874;
w42876 <= b(16) and not w42667;
w42877 <= not w42665 and w42876;
w42878 <= not w42669 and not w42877;
w42879 <= not w42875 and w42878;
w42880 <= not w42669 and not w42879;
w42881 <= b(17) and not w42658;
w42882 <= not w42656 and w42881;
w42883 <= not w42660 and not w42882;
w42884 <= not w42880 and w42883;
w42885 <= not w42660 and not w42884;
w42886 <= b(18) and not w42649;
w42887 <= not w42647 and w42886;
w42888 <= not w42651 and not w42887;
w42889 <= not w42885 and w42888;
w42890 <= not w42651 and not w42889;
w42891 <= b(19) and not w42640;
w42892 <= not w42638 and w42891;
w42893 <= not w42642 and not w42892;
w42894 <= not w42890 and w42893;
w42895 <= not w42642 and not w42894;
w42896 <= b(20) and not w42631;
w42897 <= not w42629 and w42896;
w42898 <= not w42633 and not w42897;
w42899 <= not w42895 and w42898;
w42900 <= not w42633 and not w42899;
w42901 <= b(21) and not w42622;
w42902 <= not w42620 and w42901;
w42903 <= not w42624 and not w42902;
w42904 <= not w42900 and w42903;
w42905 <= not w42624 and not w42904;
w42906 <= b(22) and not w42613;
w42907 <= not w42611 and w42906;
w42908 <= not w42615 and not w42907;
w42909 <= not w42905 and w42908;
w42910 <= not w42615 and not w42909;
w42911 <= b(23) and not w42604;
w42912 <= not w42602 and w42911;
w42913 <= not w42606 and not w42912;
w42914 <= not w42910 and w42913;
w42915 <= not w42606 and not w42914;
w42916 <= b(24) and not w42595;
w42917 <= not w42593 and w42916;
w42918 <= not w42597 and not w42917;
w42919 <= not w42915 and w42918;
w42920 <= not w42597 and not w42919;
w42921 <= b(25) and not w42586;
w42922 <= not w42584 and w42921;
w42923 <= not w42588 and not w42922;
w42924 <= not w42920 and w42923;
w42925 <= not w42588 and not w42924;
w42926 <= b(26) and not w42577;
w42927 <= not w42575 and w42926;
w42928 <= not w42579 and not w42927;
w42929 <= not w42925 and w42928;
w42930 <= not w42579 and not w42929;
w42931 <= b(27) and not w42568;
w42932 <= not w42566 and w42931;
w42933 <= not w42570 and not w42932;
w42934 <= not w42930 and w42933;
w42935 <= not w42570 and not w42934;
w42936 <= b(28) and not w42559;
w42937 <= not w42557 and w42936;
w42938 <= not w42561 and not w42937;
w42939 <= not w42935 and w42938;
w42940 <= not w42561 and not w42939;
w42941 <= b(29) and not w42550;
w42942 <= not w42548 and w42941;
w42943 <= not w42552 and not w42942;
w42944 <= not w42940 and w42943;
w42945 <= not w42552 and not w42944;
w42946 <= b(30) and not w42541;
w42947 <= not w42539 and w42946;
w42948 <= not w42543 and not w42947;
w42949 <= not w42945 and w42948;
w42950 <= not w42543 and not w42949;
w42951 <= b(31) and not w42532;
w42952 <= not w42530 and w42951;
w42953 <= not w42534 and not w42952;
w42954 <= not w42950 and w42953;
w42955 <= not w42534 and not w42954;
w42956 <= b(32) and not w42523;
w42957 <= not w42521 and w42956;
w42958 <= not w42525 and not w42957;
w42959 <= not w42955 and w42958;
w42960 <= not w42525 and not w42959;
w42961 <= b(33) and not w42514;
w42962 <= not w42512 and w42961;
w42963 <= not w42516 and not w42962;
w42964 <= not w42960 and w42963;
w42965 <= not w42516 and not w42964;
w42966 <= b(34) and not w42505;
w42967 <= not w42503 and w42966;
w42968 <= not w42507 and not w42967;
w42969 <= not w42965 and w42968;
w42970 <= not w42507 and not w42969;
w42971 <= b(35) and not w42496;
w42972 <= not w42494 and w42971;
w42973 <= not w42498 and not w42972;
w42974 <= not w42970 and w42973;
w42975 <= not w42498 and not w42974;
w42976 <= b(36) and not w42487;
w42977 <= not w42485 and w42976;
w42978 <= not w42489 and not w42977;
w42979 <= not w42975 and w42978;
w42980 <= not w42489 and not w42979;
w42981 <= b(37) and not w42478;
w42982 <= not w42476 and w42981;
w42983 <= not w42480 and not w42982;
w42984 <= not w42980 and w42983;
w42985 <= not w42480 and not w42984;
w42986 <= b(38) and not w42469;
w42987 <= not w42467 and w42986;
w42988 <= not w42471 and not w42987;
w42989 <= not w42985 and w42988;
w42990 <= not w42471 and not w42989;
w42991 <= b(39) and not w42460;
w42992 <= not w42458 and w42991;
w42993 <= not w42462 and not w42992;
w42994 <= not w42990 and w42993;
w42995 <= not w42462 and not w42994;
w42996 <= b(40) and not w42451;
w42997 <= not w42449 and w42996;
w42998 <= not w42453 and not w42997;
w42999 <= not w42995 and w42998;
w43000 <= not w42453 and not w42999;
w43001 <= b(41) and not w42442;
w43002 <= not w42440 and w43001;
w43003 <= not w42444 and not w43002;
w43004 <= not w43000 and w43003;
w43005 <= not w42444 and not w43004;
w43006 <= b(42) and not w42433;
w43007 <= not w42431 and w43006;
w43008 <= not w42435 and not w43007;
w43009 <= not w43005 and w43008;
w43010 <= not w42435 and not w43009;
w43011 <= b(43) and not w42424;
w43012 <= not w42422 and w43011;
w43013 <= not w42426 and not w43012;
w43014 <= not w43010 and w43013;
w43015 <= not w42426 and not w43014;
w43016 <= b(44) and not w42404;
w43017 <= not w42402 and w43016;
w43018 <= not w42417 and not w43017;
w43019 <= not w43015 and w43018;
w43020 <= not w42417 and not w43019;
w43021 <= b(45) and not w42414;
w43022 <= not w42412 and w43021;
w43023 <= not w42416 and not w43022;
w43024 <= not w43020 and w43023;
w43025 <= not w42416 and not w43024;
w43026 <= w14955 and not w43025;
w43027 <= not w42405 and not w43026;
w43028 <= not w42426 and w43018;
w43029 <= not w43014 and w43028;
w43030 <= not w43015 and not w43018;
w43031 <= not w43029 and not w43030;
w43032 <= w14955 and not w43031;
w43033 <= not w43025 and w43032;
w43034 <= not w43027 and not w43033;
w43035 <= not b(45) and not w43034;
w43036 <= not w42425 and not w43026;
w43037 <= not w42435 and w43013;
w43038 <= not w43009 and w43037;
w43039 <= not w43010 and not w43013;
w43040 <= not w43038 and not w43039;
w43041 <= w14955 and not w43040;
w43042 <= not w43025 and w43041;
w43043 <= not w43036 and not w43042;
w43044 <= not b(44) and not w43043;
w43045 <= not w42434 and not w43026;
w43046 <= not w42444 and w43008;
w43047 <= not w43004 and w43046;
w43048 <= not w43005 and not w43008;
w43049 <= not w43047 and not w43048;
w43050 <= w14955 and not w43049;
w43051 <= not w43025 and w43050;
w43052 <= not w43045 and not w43051;
w43053 <= not b(43) and not w43052;
w43054 <= not w42443 and not w43026;
w43055 <= not w42453 and w43003;
w43056 <= not w42999 and w43055;
w43057 <= not w43000 and not w43003;
w43058 <= not w43056 and not w43057;
w43059 <= w14955 and not w43058;
w43060 <= not w43025 and w43059;
w43061 <= not w43054 and not w43060;
w43062 <= not b(42) and not w43061;
w43063 <= not w42452 and not w43026;
w43064 <= not w42462 and w42998;
w43065 <= not w42994 and w43064;
w43066 <= not w42995 and not w42998;
w43067 <= not w43065 and not w43066;
w43068 <= w14955 and not w43067;
w43069 <= not w43025 and w43068;
w43070 <= not w43063 and not w43069;
w43071 <= not b(41) and not w43070;
w43072 <= not w42461 and not w43026;
w43073 <= not w42471 and w42993;
w43074 <= not w42989 and w43073;
w43075 <= not w42990 and not w42993;
w43076 <= not w43074 and not w43075;
w43077 <= w14955 and not w43076;
w43078 <= not w43025 and w43077;
w43079 <= not w43072 and not w43078;
w43080 <= not b(40) and not w43079;
w43081 <= not w42470 and not w43026;
w43082 <= not w42480 and w42988;
w43083 <= not w42984 and w43082;
w43084 <= not w42985 and not w42988;
w43085 <= not w43083 and not w43084;
w43086 <= w14955 and not w43085;
w43087 <= not w43025 and w43086;
w43088 <= not w43081 and not w43087;
w43089 <= not b(39) and not w43088;
w43090 <= not w42479 and not w43026;
w43091 <= not w42489 and w42983;
w43092 <= not w42979 and w43091;
w43093 <= not w42980 and not w42983;
w43094 <= not w43092 and not w43093;
w43095 <= w14955 and not w43094;
w43096 <= not w43025 and w43095;
w43097 <= not w43090 and not w43096;
w43098 <= not b(38) and not w43097;
w43099 <= not w42488 and not w43026;
w43100 <= not w42498 and w42978;
w43101 <= not w42974 and w43100;
w43102 <= not w42975 and not w42978;
w43103 <= not w43101 and not w43102;
w43104 <= w14955 and not w43103;
w43105 <= not w43025 and w43104;
w43106 <= not w43099 and not w43105;
w43107 <= not b(37) and not w43106;
w43108 <= not w42497 and not w43026;
w43109 <= not w42507 and w42973;
w43110 <= not w42969 and w43109;
w43111 <= not w42970 and not w42973;
w43112 <= not w43110 and not w43111;
w43113 <= w14955 and not w43112;
w43114 <= not w43025 and w43113;
w43115 <= not w43108 and not w43114;
w43116 <= not b(36) and not w43115;
w43117 <= not w42506 and not w43026;
w43118 <= not w42516 and w42968;
w43119 <= not w42964 and w43118;
w43120 <= not w42965 and not w42968;
w43121 <= not w43119 and not w43120;
w43122 <= w14955 and not w43121;
w43123 <= not w43025 and w43122;
w43124 <= not w43117 and not w43123;
w43125 <= not b(35) and not w43124;
w43126 <= not w42515 and not w43026;
w43127 <= not w42525 and w42963;
w43128 <= not w42959 and w43127;
w43129 <= not w42960 and not w42963;
w43130 <= not w43128 and not w43129;
w43131 <= w14955 and not w43130;
w43132 <= not w43025 and w43131;
w43133 <= not w43126 and not w43132;
w43134 <= not b(34) and not w43133;
w43135 <= not w42524 and not w43026;
w43136 <= not w42534 and w42958;
w43137 <= not w42954 and w43136;
w43138 <= not w42955 and not w42958;
w43139 <= not w43137 and not w43138;
w43140 <= w14955 and not w43139;
w43141 <= not w43025 and w43140;
w43142 <= not w43135 and not w43141;
w43143 <= not b(33) and not w43142;
w43144 <= not w42533 and not w43026;
w43145 <= not w42543 and w42953;
w43146 <= not w42949 and w43145;
w43147 <= not w42950 and not w42953;
w43148 <= not w43146 and not w43147;
w43149 <= w14955 and not w43148;
w43150 <= not w43025 and w43149;
w43151 <= not w43144 and not w43150;
w43152 <= not b(32) and not w43151;
w43153 <= not w42542 and not w43026;
w43154 <= not w42552 and w42948;
w43155 <= not w42944 and w43154;
w43156 <= not w42945 and not w42948;
w43157 <= not w43155 and not w43156;
w43158 <= w14955 and not w43157;
w43159 <= not w43025 and w43158;
w43160 <= not w43153 and not w43159;
w43161 <= not b(31) and not w43160;
w43162 <= not w42551 and not w43026;
w43163 <= not w42561 and w42943;
w43164 <= not w42939 and w43163;
w43165 <= not w42940 and not w42943;
w43166 <= not w43164 and not w43165;
w43167 <= w14955 and not w43166;
w43168 <= not w43025 and w43167;
w43169 <= not w43162 and not w43168;
w43170 <= not b(30) and not w43169;
w43171 <= not w42560 and not w43026;
w43172 <= not w42570 and w42938;
w43173 <= not w42934 and w43172;
w43174 <= not w42935 and not w42938;
w43175 <= not w43173 and not w43174;
w43176 <= w14955 and not w43175;
w43177 <= not w43025 and w43176;
w43178 <= not w43171 and not w43177;
w43179 <= not b(29) and not w43178;
w43180 <= not w42569 and not w43026;
w43181 <= not w42579 and w42933;
w43182 <= not w42929 and w43181;
w43183 <= not w42930 and not w42933;
w43184 <= not w43182 and not w43183;
w43185 <= w14955 and not w43184;
w43186 <= not w43025 and w43185;
w43187 <= not w43180 and not w43186;
w43188 <= not b(28) and not w43187;
w43189 <= not w42578 and not w43026;
w43190 <= not w42588 and w42928;
w43191 <= not w42924 and w43190;
w43192 <= not w42925 and not w42928;
w43193 <= not w43191 and not w43192;
w43194 <= w14955 and not w43193;
w43195 <= not w43025 and w43194;
w43196 <= not w43189 and not w43195;
w43197 <= not b(27) and not w43196;
w43198 <= not w42587 and not w43026;
w43199 <= not w42597 and w42923;
w43200 <= not w42919 and w43199;
w43201 <= not w42920 and not w42923;
w43202 <= not w43200 and not w43201;
w43203 <= w14955 and not w43202;
w43204 <= not w43025 and w43203;
w43205 <= not w43198 and not w43204;
w43206 <= not b(26) and not w43205;
w43207 <= not w42596 and not w43026;
w43208 <= not w42606 and w42918;
w43209 <= not w42914 and w43208;
w43210 <= not w42915 and not w42918;
w43211 <= not w43209 and not w43210;
w43212 <= w14955 and not w43211;
w43213 <= not w43025 and w43212;
w43214 <= not w43207 and not w43213;
w43215 <= not b(25) and not w43214;
w43216 <= not w42605 and not w43026;
w43217 <= not w42615 and w42913;
w43218 <= not w42909 and w43217;
w43219 <= not w42910 and not w42913;
w43220 <= not w43218 and not w43219;
w43221 <= w14955 and not w43220;
w43222 <= not w43025 and w43221;
w43223 <= not w43216 and not w43222;
w43224 <= not b(24) and not w43223;
w43225 <= not w42614 and not w43026;
w43226 <= not w42624 and w42908;
w43227 <= not w42904 and w43226;
w43228 <= not w42905 and not w42908;
w43229 <= not w43227 and not w43228;
w43230 <= w14955 and not w43229;
w43231 <= not w43025 and w43230;
w43232 <= not w43225 and not w43231;
w43233 <= not b(23) and not w43232;
w43234 <= not w42623 and not w43026;
w43235 <= not w42633 and w42903;
w43236 <= not w42899 and w43235;
w43237 <= not w42900 and not w42903;
w43238 <= not w43236 and not w43237;
w43239 <= w14955 and not w43238;
w43240 <= not w43025 and w43239;
w43241 <= not w43234 and not w43240;
w43242 <= not b(22) and not w43241;
w43243 <= not w42632 and not w43026;
w43244 <= not w42642 and w42898;
w43245 <= not w42894 and w43244;
w43246 <= not w42895 and not w42898;
w43247 <= not w43245 and not w43246;
w43248 <= w14955 and not w43247;
w43249 <= not w43025 and w43248;
w43250 <= not w43243 and not w43249;
w43251 <= not b(21) and not w43250;
w43252 <= not w42641 and not w43026;
w43253 <= not w42651 and w42893;
w43254 <= not w42889 and w43253;
w43255 <= not w42890 and not w42893;
w43256 <= not w43254 and not w43255;
w43257 <= w14955 and not w43256;
w43258 <= not w43025 and w43257;
w43259 <= not w43252 and not w43258;
w43260 <= not b(20) and not w43259;
w43261 <= not w42650 and not w43026;
w43262 <= not w42660 and w42888;
w43263 <= not w42884 and w43262;
w43264 <= not w42885 and not w42888;
w43265 <= not w43263 and not w43264;
w43266 <= w14955 and not w43265;
w43267 <= not w43025 and w43266;
w43268 <= not w43261 and not w43267;
w43269 <= not b(19) and not w43268;
w43270 <= not w42659 and not w43026;
w43271 <= not w42669 and w42883;
w43272 <= not w42879 and w43271;
w43273 <= not w42880 and not w42883;
w43274 <= not w43272 and not w43273;
w43275 <= w14955 and not w43274;
w43276 <= not w43025 and w43275;
w43277 <= not w43270 and not w43276;
w43278 <= not b(18) and not w43277;
w43279 <= not w42668 and not w43026;
w43280 <= not w42678 and w42878;
w43281 <= not w42874 and w43280;
w43282 <= not w42875 and not w42878;
w43283 <= not w43281 and not w43282;
w43284 <= w14955 and not w43283;
w43285 <= not w43025 and w43284;
w43286 <= not w43279 and not w43285;
w43287 <= not b(17) and not w43286;
w43288 <= not w42677 and not w43026;
w43289 <= not w42687 and w42873;
w43290 <= not w42869 and w43289;
w43291 <= not w42870 and not w42873;
w43292 <= not w43290 and not w43291;
w43293 <= w14955 and not w43292;
w43294 <= not w43025 and w43293;
w43295 <= not w43288 and not w43294;
w43296 <= not b(16) and not w43295;
w43297 <= not w42686 and not w43026;
w43298 <= not w42696 and w42868;
w43299 <= not w42864 and w43298;
w43300 <= not w42865 and not w42868;
w43301 <= not w43299 and not w43300;
w43302 <= w14955 and not w43301;
w43303 <= not w43025 and w43302;
w43304 <= not w43297 and not w43303;
w43305 <= not b(15) and not w43304;
w43306 <= not w42695 and not w43026;
w43307 <= not w42705 and w42863;
w43308 <= not w42859 and w43307;
w43309 <= not w42860 and not w42863;
w43310 <= not w43308 and not w43309;
w43311 <= w14955 and not w43310;
w43312 <= not w43025 and w43311;
w43313 <= not w43306 and not w43312;
w43314 <= not b(14) and not w43313;
w43315 <= not w42704 and not w43026;
w43316 <= not w42714 and w42858;
w43317 <= not w42854 and w43316;
w43318 <= not w42855 and not w42858;
w43319 <= not w43317 and not w43318;
w43320 <= w14955 and not w43319;
w43321 <= not w43025 and w43320;
w43322 <= not w43315 and not w43321;
w43323 <= not b(13) and not w43322;
w43324 <= not w42713 and not w43026;
w43325 <= not w42723 and w42853;
w43326 <= not w42849 and w43325;
w43327 <= not w42850 and not w42853;
w43328 <= not w43326 and not w43327;
w43329 <= w14955 and not w43328;
w43330 <= not w43025 and w43329;
w43331 <= not w43324 and not w43330;
w43332 <= not b(12) and not w43331;
w43333 <= not w42722 and not w43026;
w43334 <= not w42732 and w42848;
w43335 <= not w42844 and w43334;
w43336 <= not w42845 and not w42848;
w43337 <= not w43335 and not w43336;
w43338 <= w14955 and not w43337;
w43339 <= not w43025 and w43338;
w43340 <= not w43333 and not w43339;
w43341 <= not b(11) and not w43340;
w43342 <= not w42731 and not w43026;
w43343 <= not w42741 and w42843;
w43344 <= not w42839 and w43343;
w43345 <= not w42840 and not w42843;
w43346 <= not w43344 and not w43345;
w43347 <= w14955 and not w43346;
w43348 <= not w43025 and w43347;
w43349 <= not w43342 and not w43348;
w43350 <= not b(10) and not w43349;
w43351 <= not w42740 and not w43026;
w43352 <= not w42750 and w42838;
w43353 <= not w42834 and w43352;
w43354 <= not w42835 and not w42838;
w43355 <= not w43353 and not w43354;
w43356 <= w14955 and not w43355;
w43357 <= not w43025 and w43356;
w43358 <= not w43351 and not w43357;
w43359 <= not b(9) and not w43358;
w43360 <= not w42749 and not w43026;
w43361 <= not w42759 and w42833;
w43362 <= not w42829 and w43361;
w43363 <= not w42830 and not w42833;
w43364 <= not w43362 and not w43363;
w43365 <= w14955 and not w43364;
w43366 <= not w43025 and w43365;
w43367 <= not w43360 and not w43366;
w43368 <= not b(8) and not w43367;
w43369 <= not w42758 and not w43026;
w43370 <= not w42768 and w42828;
w43371 <= not w42824 and w43370;
w43372 <= not w42825 and not w42828;
w43373 <= not w43371 and not w43372;
w43374 <= w14955 and not w43373;
w43375 <= not w43025 and w43374;
w43376 <= not w43369 and not w43375;
w43377 <= not b(7) and not w43376;
w43378 <= not w42767 and not w43026;
w43379 <= not w42777 and w42823;
w43380 <= not w42819 and w43379;
w43381 <= not w42820 and not w42823;
w43382 <= not w43380 and not w43381;
w43383 <= w14955 and not w43382;
w43384 <= not w43025 and w43383;
w43385 <= not w43378 and not w43384;
w43386 <= not b(6) and not w43385;
w43387 <= not w42776 and not w43026;
w43388 <= not w42786 and w42818;
w43389 <= not w42814 and w43388;
w43390 <= not w42815 and not w42818;
w43391 <= not w43389 and not w43390;
w43392 <= w14955 and not w43391;
w43393 <= not w43025 and w43392;
w43394 <= not w43387 and not w43393;
w43395 <= not b(5) and not w43394;
w43396 <= not w42785 and not w43026;
w43397 <= not w42794 and w42813;
w43398 <= not w42809 and w43397;
w43399 <= not w42810 and not w42813;
w43400 <= not w43398 and not w43399;
w43401 <= w14955 and not w43400;
w43402 <= not w43025 and w43401;
w43403 <= not w43396 and not w43402;
w43404 <= not b(4) and not w43403;
w43405 <= not w42793 and not w43026;
w43406 <= not w42804 and w42808;
w43407 <= not w42803 and w43406;
w43408 <= not w42805 and not w42808;
w43409 <= not w43407 and not w43408;
w43410 <= w14955 and not w43409;
w43411 <= not w43025 and w43410;
w43412 <= not w43405 and not w43411;
w43413 <= not b(3) and not w43412;
w43414 <= not w42798 and not w43026;
w43415 <= w14730 and not w42801;
w43416 <= not w42799 and w43415;
w43417 <= w14955 and not w43416;
w43418 <= not w42803 and w43417;
w43419 <= not w43025 and w43418;
w43420 <= not w43414 and not w43419;
w43421 <= not b(2) and not w43420;
w43422 <= w15355 and not w43025;
w43423 <= a(18) and not w43422;
w43424 <= w15360 and not w43025;
w43425 <= not w43423 and not w43424;
w43426 <= b(1) and not w43425;
w43427 <= not b(1) and not w43424;
w43428 <= not w43423 and w43427;
w43429 <= not w43426 and not w43428;
w43430 <= not w15367 and not w43429;
w43431 <= not b(1) and not w43425;
w43432 <= not w43430 and not w43431;
w43433 <= b(2) and not w43419;
w43434 <= not w43414 and w43433;
w43435 <= not w43421 and not w43434;
w43436 <= not w43432 and w43435;
w43437 <= not w43421 and not w43436;
w43438 <= b(3) and not w43411;
w43439 <= not w43405 and w43438;
w43440 <= not w43413 and not w43439;
w43441 <= not w43437 and w43440;
w43442 <= not w43413 and not w43441;
w43443 <= b(4) and not w43402;
w43444 <= not w43396 and w43443;
w43445 <= not w43404 and not w43444;
w43446 <= not w43442 and w43445;
w43447 <= not w43404 and not w43446;
w43448 <= b(5) and not w43393;
w43449 <= not w43387 and w43448;
w43450 <= not w43395 and not w43449;
w43451 <= not w43447 and w43450;
w43452 <= not w43395 and not w43451;
w43453 <= b(6) and not w43384;
w43454 <= not w43378 and w43453;
w43455 <= not w43386 and not w43454;
w43456 <= not w43452 and w43455;
w43457 <= not w43386 and not w43456;
w43458 <= b(7) and not w43375;
w43459 <= not w43369 and w43458;
w43460 <= not w43377 and not w43459;
w43461 <= not w43457 and w43460;
w43462 <= not w43377 and not w43461;
w43463 <= b(8) and not w43366;
w43464 <= not w43360 and w43463;
w43465 <= not w43368 and not w43464;
w43466 <= not w43462 and w43465;
w43467 <= not w43368 and not w43466;
w43468 <= b(9) and not w43357;
w43469 <= not w43351 and w43468;
w43470 <= not w43359 and not w43469;
w43471 <= not w43467 and w43470;
w43472 <= not w43359 and not w43471;
w43473 <= b(10) and not w43348;
w43474 <= not w43342 and w43473;
w43475 <= not w43350 and not w43474;
w43476 <= not w43472 and w43475;
w43477 <= not w43350 and not w43476;
w43478 <= b(11) and not w43339;
w43479 <= not w43333 and w43478;
w43480 <= not w43341 and not w43479;
w43481 <= not w43477 and w43480;
w43482 <= not w43341 and not w43481;
w43483 <= b(12) and not w43330;
w43484 <= not w43324 and w43483;
w43485 <= not w43332 and not w43484;
w43486 <= not w43482 and w43485;
w43487 <= not w43332 and not w43486;
w43488 <= b(13) and not w43321;
w43489 <= not w43315 and w43488;
w43490 <= not w43323 and not w43489;
w43491 <= not w43487 and w43490;
w43492 <= not w43323 and not w43491;
w43493 <= b(14) and not w43312;
w43494 <= not w43306 and w43493;
w43495 <= not w43314 and not w43494;
w43496 <= not w43492 and w43495;
w43497 <= not w43314 and not w43496;
w43498 <= b(15) and not w43303;
w43499 <= not w43297 and w43498;
w43500 <= not w43305 and not w43499;
w43501 <= not w43497 and w43500;
w43502 <= not w43305 and not w43501;
w43503 <= b(16) and not w43294;
w43504 <= not w43288 and w43503;
w43505 <= not w43296 and not w43504;
w43506 <= not w43502 and w43505;
w43507 <= not w43296 and not w43506;
w43508 <= b(17) and not w43285;
w43509 <= not w43279 and w43508;
w43510 <= not w43287 and not w43509;
w43511 <= not w43507 and w43510;
w43512 <= not w43287 and not w43511;
w43513 <= b(18) and not w43276;
w43514 <= not w43270 and w43513;
w43515 <= not w43278 and not w43514;
w43516 <= not w43512 and w43515;
w43517 <= not w43278 and not w43516;
w43518 <= b(19) and not w43267;
w43519 <= not w43261 and w43518;
w43520 <= not w43269 and not w43519;
w43521 <= not w43517 and w43520;
w43522 <= not w43269 and not w43521;
w43523 <= b(20) and not w43258;
w43524 <= not w43252 and w43523;
w43525 <= not w43260 and not w43524;
w43526 <= not w43522 and w43525;
w43527 <= not w43260 and not w43526;
w43528 <= b(21) and not w43249;
w43529 <= not w43243 and w43528;
w43530 <= not w43251 and not w43529;
w43531 <= not w43527 and w43530;
w43532 <= not w43251 and not w43531;
w43533 <= b(22) and not w43240;
w43534 <= not w43234 and w43533;
w43535 <= not w43242 and not w43534;
w43536 <= not w43532 and w43535;
w43537 <= not w43242 and not w43536;
w43538 <= b(23) and not w43231;
w43539 <= not w43225 and w43538;
w43540 <= not w43233 and not w43539;
w43541 <= not w43537 and w43540;
w43542 <= not w43233 and not w43541;
w43543 <= b(24) and not w43222;
w43544 <= not w43216 and w43543;
w43545 <= not w43224 and not w43544;
w43546 <= not w43542 and w43545;
w43547 <= not w43224 and not w43546;
w43548 <= b(25) and not w43213;
w43549 <= not w43207 and w43548;
w43550 <= not w43215 and not w43549;
w43551 <= not w43547 and w43550;
w43552 <= not w43215 and not w43551;
w43553 <= b(26) and not w43204;
w43554 <= not w43198 and w43553;
w43555 <= not w43206 and not w43554;
w43556 <= not w43552 and w43555;
w43557 <= not w43206 and not w43556;
w43558 <= b(27) and not w43195;
w43559 <= not w43189 and w43558;
w43560 <= not w43197 and not w43559;
w43561 <= not w43557 and w43560;
w43562 <= not w43197 and not w43561;
w43563 <= b(28) and not w43186;
w43564 <= not w43180 and w43563;
w43565 <= not w43188 and not w43564;
w43566 <= not w43562 and w43565;
w43567 <= not w43188 and not w43566;
w43568 <= b(29) and not w43177;
w43569 <= not w43171 and w43568;
w43570 <= not w43179 and not w43569;
w43571 <= not w43567 and w43570;
w43572 <= not w43179 and not w43571;
w43573 <= b(30) and not w43168;
w43574 <= not w43162 and w43573;
w43575 <= not w43170 and not w43574;
w43576 <= not w43572 and w43575;
w43577 <= not w43170 and not w43576;
w43578 <= b(31) and not w43159;
w43579 <= not w43153 and w43578;
w43580 <= not w43161 and not w43579;
w43581 <= not w43577 and w43580;
w43582 <= not w43161 and not w43581;
w43583 <= b(32) and not w43150;
w43584 <= not w43144 and w43583;
w43585 <= not w43152 and not w43584;
w43586 <= not w43582 and w43585;
w43587 <= not w43152 and not w43586;
w43588 <= b(33) and not w43141;
w43589 <= not w43135 and w43588;
w43590 <= not w43143 and not w43589;
w43591 <= not w43587 and w43590;
w43592 <= not w43143 and not w43591;
w43593 <= b(34) and not w43132;
w43594 <= not w43126 and w43593;
w43595 <= not w43134 and not w43594;
w43596 <= not w43592 and w43595;
w43597 <= not w43134 and not w43596;
w43598 <= b(35) and not w43123;
w43599 <= not w43117 and w43598;
w43600 <= not w43125 and not w43599;
w43601 <= not w43597 and w43600;
w43602 <= not w43125 and not w43601;
w43603 <= b(36) and not w43114;
w43604 <= not w43108 and w43603;
w43605 <= not w43116 and not w43604;
w43606 <= not w43602 and w43605;
w43607 <= not w43116 and not w43606;
w43608 <= b(37) and not w43105;
w43609 <= not w43099 and w43608;
w43610 <= not w43107 and not w43609;
w43611 <= not w43607 and w43610;
w43612 <= not w43107 and not w43611;
w43613 <= b(38) and not w43096;
w43614 <= not w43090 and w43613;
w43615 <= not w43098 and not w43614;
w43616 <= not w43612 and w43615;
w43617 <= not w43098 and not w43616;
w43618 <= b(39) and not w43087;
w43619 <= not w43081 and w43618;
w43620 <= not w43089 and not w43619;
w43621 <= not w43617 and w43620;
w43622 <= not w43089 and not w43621;
w43623 <= b(40) and not w43078;
w43624 <= not w43072 and w43623;
w43625 <= not w43080 and not w43624;
w43626 <= not w43622 and w43625;
w43627 <= not w43080 and not w43626;
w43628 <= b(41) and not w43069;
w43629 <= not w43063 and w43628;
w43630 <= not w43071 and not w43629;
w43631 <= not w43627 and w43630;
w43632 <= not w43071 and not w43631;
w43633 <= b(42) and not w43060;
w43634 <= not w43054 and w43633;
w43635 <= not w43062 and not w43634;
w43636 <= not w43632 and w43635;
w43637 <= not w43062 and not w43636;
w43638 <= b(43) and not w43051;
w43639 <= not w43045 and w43638;
w43640 <= not w43053 and not w43639;
w43641 <= not w43637 and w43640;
w43642 <= not w43053 and not w43641;
w43643 <= b(44) and not w43042;
w43644 <= not w43036 and w43643;
w43645 <= not w43044 and not w43644;
w43646 <= not w43642 and w43645;
w43647 <= not w43044 and not w43646;
w43648 <= b(45) and not w43033;
w43649 <= not w43027 and w43648;
w43650 <= not w43035 and not w43649;
w43651 <= not w43647 and w43650;
w43652 <= not w43035 and not w43651;
w43653 <= not w42415 and not w43026;
w43654 <= not w42417 and w43023;
w43655 <= not w43019 and w43654;
w43656 <= not w43020 and not w43023;
w43657 <= not w43655 and not w43656;
w43658 <= w43026 and not w43657;
w43659 <= not w43653 and not w43658;
w43660 <= not b(46) and not w43659;
w43661 <= b(46) and not w43653;
w43662 <= not w43658 and w43661;
w43663 <= w15602 and not w43662;
w43664 <= not w43660 and w43663;
w43665 <= not w43652 and w43664;
w43666 <= w14955 and not w43659;
w43667 <= not w43665 and not w43666;
w43668 <= not w43044 and w43650;
w43669 <= not w43646 and w43668;
w43670 <= not w43647 and not w43650;
w43671 <= not w43669 and not w43670;
w43672 <= not w43667 and not w43671;
w43673 <= not w43034 and not w43666;
w43674 <= not w43665 and w43673;
w43675 <= not w43672 and not w43674;
w43676 <= not b(46) and not w43675;
w43677 <= not w43053 and w43645;
w43678 <= not w43641 and w43677;
w43679 <= not w43642 and not w43645;
w43680 <= not w43678 and not w43679;
w43681 <= not w43667 and not w43680;
w43682 <= not w43043 and not w43666;
w43683 <= not w43665 and w43682;
w43684 <= not w43681 and not w43683;
w43685 <= not b(45) and not w43684;
w43686 <= not w43062 and w43640;
w43687 <= not w43636 and w43686;
w43688 <= not w43637 and not w43640;
w43689 <= not w43687 and not w43688;
w43690 <= not w43667 and not w43689;
w43691 <= not w43052 and not w43666;
w43692 <= not w43665 and w43691;
w43693 <= not w43690 and not w43692;
w43694 <= not b(44) and not w43693;
w43695 <= not w43071 and w43635;
w43696 <= not w43631 and w43695;
w43697 <= not w43632 and not w43635;
w43698 <= not w43696 and not w43697;
w43699 <= not w43667 and not w43698;
w43700 <= not w43061 and not w43666;
w43701 <= not w43665 and w43700;
w43702 <= not w43699 and not w43701;
w43703 <= not b(43) and not w43702;
w43704 <= not w43080 and w43630;
w43705 <= not w43626 and w43704;
w43706 <= not w43627 and not w43630;
w43707 <= not w43705 and not w43706;
w43708 <= not w43667 and not w43707;
w43709 <= not w43070 and not w43666;
w43710 <= not w43665 and w43709;
w43711 <= not w43708 and not w43710;
w43712 <= not b(42) and not w43711;
w43713 <= not w43089 and w43625;
w43714 <= not w43621 and w43713;
w43715 <= not w43622 and not w43625;
w43716 <= not w43714 and not w43715;
w43717 <= not w43667 and not w43716;
w43718 <= not w43079 and not w43666;
w43719 <= not w43665 and w43718;
w43720 <= not w43717 and not w43719;
w43721 <= not b(41) and not w43720;
w43722 <= not w43098 and w43620;
w43723 <= not w43616 and w43722;
w43724 <= not w43617 and not w43620;
w43725 <= not w43723 and not w43724;
w43726 <= not w43667 and not w43725;
w43727 <= not w43088 and not w43666;
w43728 <= not w43665 and w43727;
w43729 <= not w43726 and not w43728;
w43730 <= not b(40) and not w43729;
w43731 <= not w43107 and w43615;
w43732 <= not w43611 and w43731;
w43733 <= not w43612 and not w43615;
w43734 <= not w43732 and not w43733;
w43735 <= not w43667 and not w43734;
w43736 <= not w43097 and not w43666;
w43737 <= not w43665 and w43736;
w43738 <= not w43735 and not w43737;
w43739 <= not b(39) and not w43738;
w43740 <= not w43116 and w43610;
w43741 <= not w43606 and w43740;
w43742 <= not w43607 and not w43610;
w43743 <= not w43741 and not w43742;
w43744 <= not w43667 and not w43743;
w43745 <= not w43106 and not w43666;
w43746 <= not w43665 and w43745;
w43747 <= not w43744 and not w43746;
w43748 <= not b(38) and not w43747;
w43749 <= not w43125 and w43605;
w43750 <= not w43601 and w43749;
w43751 <= not w43602 and not w43605;
w43752 <= not w43750 and not w43751;
w43753 <= not w43667 and not w43752;
w43754 <= not w43115 and not w43666;
w43755 <= not w43665 and w43754;
w43756 <= not w43753 and not w43755;
w43757 <= not b(37) and not w43756;
w43758 <= not w43134 and w43600;
w43759 <= not w43596 and w43758;
w43760 <= not w43597 and not w43600;
w43761 <= not w43759 and not w43760;
w43762 <= not w43667 and not w43761;
w43763 <= not w43124 and not w43666;
w43764 <= not w43665 and w43763;
w43765 <= not w43762 and not w43764;
w43766 <= not b(36) and not w43765;
w43767 <= not w43143 and w43595;
w43768 <= not w43591 and w43767;
w43769 <= not w43592 and not w43595;
w43770 <= not w43768 and not w43769;
w43771 <= not w43667 and not w43770;
w43772 <= not w43133 and not w43666;
w43773 <= not w43665 and w43772;
w43774 <= not w43771 and not w43773;
w43775 <= not b(35) and not w43774;
w43776 <= not w43152 and w43590;
w43777 <= not w43586 and w43776;
w43778 <= not w43587 and not w43590;
w43779 <= not w43777 and not w43778;
w43780 <= not w43667 and not w43779;
w43781 <= not w43142 and not w43666;
w43782 <= not w43665 and w43781;
w43783 <= not w43780 and not w43782;
w43784 <= not b(34) and not w43783;
w43785 <= not w43161 and w43585;
w43786 <= not w43581 and w43785;
w43787 <= not w43582 and not w43585;
w43788 <= not w43786 and not w43787;
w43789 <= not w43667 and not w43788;
w43790 <= not w43151 and not w43666;
w43791 <= not w43665 and w43790;
w43792 <= not w43789 and not w43791;
w43793 <= not b(33) and not w43792;
w43794 <= not w43170 and w43580;
w43795 <= not w43576 and w43794;
w43796 <= not w43577 and not w43580;
w43797 <= not w43795 and not w43796;
w43798 <= not w43667 and not w43797;
w43799 <= not w43160 and not w43666;
w43800 <= not w43665 and w43799;
w43801 <= not w43798 and not w43800;
w43802 <= not b(32) and not w43801;
w43803 <= not w43179 and w43575;
w43804 <= not w43571 and w43803;
w43805 <= not w43572 and not w43575;
w43806 <= not w43804 and not w43805;
w43807 <= not w43667 and not w43806;
w43808 <= not w43169 and not w43666;
w43809 <= not w43665 and w43808;
w43810 <= not w43807 and not w43809;
w43811 <= not b(31) and not w43810;
w43812 <= not w43188 and w43570;
w43813 <= not w43566 and w43812;
w43814 <= not w43567 and not w43570;
w43815 <= not w43813 and not w43814;
w43816 <= not w43667 and not w43815;
w43817 <= not w43178 and not w43666;
w43818 <= not w43665 and w43817;
w43819 <= not w43816 and not w43818;
w43820 <= not b(30) and not w43819;
w43821 <= not w43197 and w43565;
w43822 <= not w43561 and w43821;
w43823 <= not w43562 and not w43565;
w43824 <= not w43822 and not w43823;
w43825 <= not w43667 and not w43824;
w43826 <= not w43187 and not w43666;
w43827 <= not w43665 and w43826;
w43828 <= not w43825 and not w43827;
w43829 <= not b(29) and not w43828;
w43830 <= not w43206 and w43560;
w43831 <= not w43556 and w43830;
w43832 <= not w43557 and not w43560;
w43833 <= not w43831 and not w43832;
w43834 <= not w43667 and not w43833;
w43835 <= not w43196 and not w43666;
w43836 <= not w43665 and w43835;
w43837 <= not w43834 and not w43836;
w43838 <= not b(28) and not w43837;
w43839 <= not w43215 and w43555;
w43840 <= not w43551 and w43839;
w43841 <= not w43552 and not w43555;
w43842 <= not w43840 and not w43841;
w43843 <= not w43667 and not w43842;
w43844 <= not w43205 and not w43666;
w43845 <= not w43665 and w43844;
w43846 <= not w43843 and not w43845;
w43847 <= not b(27) and not w43846;
w43848 <= not w43224 and w43550;
w43849 <= not w43546 and w43848;
w43850 <= not w43547 and not w43550;
w43851 <= not w43849 and not w43850;
w43852 <= not w43667 and not w43851;
w43853 <= not w43214 and not w43666;
w43854 <= not w43665 and w43853;
w43855 <= not w43852 and not w43854;
w43856 <= not b(26) and not w43855;
w43857 <= not w43233 and w43545;
w43858 <= not w43541 and w43857;
w43859 <= not w43542 and not w43545;
w43860 <= not w43858 and not w43859;
w43861 <= not w43667 and not w43860;
w43862 <= not w43223 and not w43666;
w43863 <= not w43665 and w43862;
w43864 <= not w43861 and not w43863;
w43865 <= not b(25) and not w43864;
w43866 <= not w43242 and w43540;
w43867 <= not w43536 and w43866;
w43868 <= not w43537 and not w43540;
w43869 <= not w43867 and not w43868;
w43870 <= not w43667 and not w43869;
w43871 <= not w43232 and not w43666;
w43872 <= not w43665 and w43871;
w43873 <= not w43870 and not w43872;
w43874 <= not b(24) and not w43873;
w43875 <= not w43251 and w43535;
w43876 <= not w43531 and w43875;
w43877 <= not w43532 and not w43535;
w43878 <= not w43876 and not w43877;
w43879 <= not w43667 and not w43878;
w43880 <= not w43241 and not w43666;
w43881 <= not w43665 and w43880;
w43882 <= not w43879 and not w43881;
w43883 <= not b(23) and not w43882;
w43884 <= not w43260 and w43530;
w43885 <= not w43526 and w43884;
w43886 <= not w43527 and not w43530;
w43887 <= not w43885 and not w43886;
w43888 <= not w43667 and not w43887;
w43889 <= not w43250 and not w43666;
w43890 <= not w43665 and w43889;
w43891 <= not w43888 and not w43890;
w43892 <= not b(22) and not w43891;
w43893 <= not w43269 and w43525;
w43894 <= not w43521 and w43893;
w43895 <= not w43522 and not w43525;
w43896 <= not w43894 and not w43895;
w43897 <= not w43667 and not w43896;
w43898 <= not w43259 and not w43666;
w43899 <= not w43665 and w43898;
w43900 <= not w43897 and not w43899;
w43901 <= not b(21) and not w43900;
w43902 <= not w43278 and w43520;
w43903 <= not w43516 and w43902;
w43904 <= not w43517 and not w43520;
w43905 <= not w43903 and not w43904;
w43906 <= not w43667 and not w43905;
w43907 <= not w43268 and not w43666;
w43908 <= not w43665 and w43907;
w43909 <= not w43906 and not w43908;
w43910 <= not b(20) and not w43909;
w43911 <= not w43287 and w43515;
w43912 <= not w43511 and w43911;
w43913 <= not w43512 and not w43515;
w43914 <= not w43912 and not w43913;
w43915 <= not w43667 and not w43914;
w43916 <= not w43277 and not w43666;
w43917 <= not w43665 and w43916;
w43918 <= not w43915 and not w43917;
w43919 <= not b(19) and not w43918;
w43920 <= not w43296 and w43510;
w43921 <= not w43506 and w43920;
w43922 <= not w43507 and not w43510;
w43923 <= not w43921 and not w43922;
w43924 <= not w43667 and not w43923;
w43925 <= not w43286 and not w43666;
w43926 <= not w43665 and w43925;
w43927 <= not w43924 and not w43926;
w43928 <= not b(18) and not w43927;
w43929 <= not w43305 and w43505;
w43930 <= not w43501 and w43929;
w43931 <= not w43502 and not w43505;
w43932 <= not w43930 and not w43931;
w43933 <= not w43667 and not w43932;
w43934 <= not w43295 and not w43666;
w43935 <= not w43665 and w43934;
w43936 <= not w43933 and not w43935;
w43937 <= not b(17) and not w43936;
w43938 <= not w43314 and w43500;
w43939 <= not w43496 and w43938;
w43940 <= not w43497 and not w43500;
w43941 <= not w43939 and not w43940;
w43942 <= not w43667 and not w43941;
w43943 <= not w43304 and not w43666;
w43944 <= not w43665 and w43943;
w43945 <= not w43942 and not w43944;
w43946 <= not b(16) and not w43945;
w43947 <= not w43323 and w43495;
w43948 <= not w43491 and w43947;
w43949 <= not w43492 and not w43495;
w43950 <= not w43948 and not w43949;
w43951 <= not w43667 and not w43950;
w43952 <= not w43313 and not w43666;
w43953 <= not w43665 and w43952;
w43954 <= not w43951 and not w43953;
w43955 <= not b(15) and not w43954;
w43956 <= not w43332 and w43490;
w43957 <= not w43486 and w43956;
w43958 <= not w43487 and not w43490;
w43959 <= not w43957 and not w43958;
w43960 <= not w43667 and not w43959;
w43961 <= not w43322 and not w43666;
w43962 <= not w43665 and w43961;
w43963 <= not w43960 and not w43962;
w43964 <= not b(14) and not w43963;
w43965 <= not w43341 and w43485;
w43966 <= not w43481 and w43965;
w43967 <= not w43482 and not w43485;
w43968 <= not w43966 and not w43967;
w43969 <= not w43667 and not w43968;
w43970 <= not w43331 and not w43666;
w43971 <= not w43665 and w43970;
w43972 <= not w43969 and not w43971;
w43973 <= not b(13) and not w43972;
w43974 <= not w43350 and w43480;
w43975 <= not w43476 and w43974;
w43976 <= not w43477 and not w43480;
w43977 <= not w43975 and not w43976;
w43978 <= not w43667 and not w43977;
w43979 <= not w43340 and not w43666;
w43980 <= not w43665 and w43979;
w43981 <= not w43978 and not w43980;
w43982 <= not b(12) and not w43981;
w43983 <= not w43359 and w43475;
w43984 <= not w43471 and w43983;
w43985 <= not w43472 and not w43475;
w43986 <= not w43984 and not w43985;
w43987 <= not w43667 and not w43986;
w43988 <= not w43349 and not w43666;
w43989 <= not w43665 and w43988;
w43990 <= not w43987 and not w43989;
w43991 <= not b(11) and not w43990;
w43992 <= not w43368 and w43470;
w43993 <= not w43466 and w43992;
w43994 <= not w43467 and not w43470;
w43995 <= not w43993 and not w43994;
w43996 <= not w43667 and not w43995;
w43997 <= not w43358 and not w43666;
w43998 <= not w43665 and w43997;
w43999 <= not w43996 and not w43998;
w44000 <= not b(10) and not w43999;
w44001 <= not w43377 and w43465;
w44002 <= not w43461 and w44001;
w44003 <= not w43462 and not w43465;
w44004 <= not w44002 and not w44003;
w44005 <= not w43667 and not w44004;
w44006 <= not w43367 and not w43666;
w44007 <= not w43665 and w44006;
w44008 <= not w44005 and not w44007;
w44009 <= not b(9) and not w44008;
w44010 <= not w43386 and w43460;
w44011 <= not w43456 and w44010;
w44012 <= not w43457 and not w43460;
w44013 <= not w44011 and not w44012;
w44014 <= not w43667 and not w44013;
w44015 <= not w43376 and not w43666;
w44016 <= not w43665 and w44015;
w44017 <= not w44014 and not w44016;
w44018 <= not b(8) and not w44017;
w44019 <= not w43395 and w43455;
w44020 <= not w43451 and w44019;
w44021 <= not w43452 and not w43455;
w44022 <= not w44020 and not w44021;
w44023 <= not w43667 and not w44022;
w44024 <= not w43385 and not w43666;
w44025 <= not w43665 and w44024;
w44026 <= not w44023 and not w44025;
w44027 <= not b(7) and not w44026;
w44028 <= not w43404 and w43450;
w44029 <= not w43446 and w44028;
w44030 <= not w43447 and not w43450;
w44031 <= not w44029 and not w44030;
w44032 <= not w43667 and not w44031;
w44033 <= not w43394 and not w43666;
w44034 <= not w43665 and w44033;
w44035 <= not w44032 and not w44034;
w44036 <= not b(6) and not w44035;
w44037 <= not w43413 and w43445;
w44038 <= not w43441 and w44037;
w44039 <= not w43442 and not w43445;
w44040 <= not w44038 and not w44039;
w44041 <= not w43667 and not w44040;
w44042 <= not w43403 and not w43666;
w44043 <= not w43665 and w44042;
w44044 <= not w44041 and not w44043;
w44045 <= not b(5) and not w44044;
w44046 <= not w43421 and w43440;
w44047 <= not w43436 and w44046;
w44048 <= not w43437 and not w43440;
w44049 <= not w44047 and not w44048;
w44050 <= not w43667 and not w44049;
w44051 <= not w43412 and not w43666;
w44052 <= not w43665 and w44051;
w44053 <= not w44050 and not w44052;
w44054 <= not b(4) and not w44053;
w44055 <= not w43431 and w43435;
w44056 <= not w43430 and w44055;
w44057 <= not w43432 and not w43435;
w44058 <= not w44056 and not w44057;
w44059 <= not w43667 and not w44058;
w44060 <= not w43420 and not w43666;
w44061 <= not w43665 and w44060;
w44062 <= not w44059 and not w44061;
w44063 <= not b(3) and not w44062;
w44064 <= w15367 and not w43428;
w44065 <= not w43426 and w44064;
w44066 <= not w43430 and not w44065;
w44067 <= not w43667 and w44066;
w44068 <= not w43425 and not w43666;
w44069 <= not w43665 and w44068;
w44070 <= not w44067 and not w44069;
w44071 <= not b(2) and not w44070;
w44072 <= b(0) and not w43667;
w44073 <= a(17) and not w44072;
w44074 <= w15367 and not w43667;
w44075 <= not w44073 and not w44074;
w44076 <= b(1) and not w44075;
w44077 <= not b(1) and not w44074;
w44078 <= not w44073 and w44077;
w44079 <= not w44076 and not w44078;
w44080 <= not w16020 and not w44079;
w44081 <= not b(1) and not w44075;
w44082 <= not w44080 and not w44081;
w44083 <= b(2) and not w44069;
w44084 <= not w44067 and w44083;
w44085 <= not w44071 and not w44084;
w44086 <= not w44082 and w44085;
w44087 <= not w44071 and not w44086;
w44088 <= b(3) and not w44061;
w44089 <= not w44059 and w44088;
w44090 <= not w44063 and not w44089;
w44091 <= not w44087 and w44090;
w44092 <= not w44063 and not w44091;
w44093 <= b(4) and not w44052;
w44094 <= not w44050 and w44093;
w44095 <= not w44054 and not w44094;
w44096 <= not w44092 and w44095;
w44097 <= not w44054 and not w44096;
w44098 <= b(5) and not w44043;
w44099 <= not w44041 and w44098;
w44100 <= not w44045 and not w44099;
w44101 <= not w44097 and w44100;
w44102 <= not w44045 and not w44101;
w44103 <= b(6) and not w44034;
w44104 <= not w44032 and w44103;
w44105 <= not w44036 and not w44104;
w44106 <= not w44102 and w44105;
w44107 <= not w44036 and not w44106;
w44108 <= b(7) and not w44025;
w44109 <= not w44023 and w44108;
w44110 <= not w44027 and not w44109;
w44111 <= not w44107 and w44110;
w44112 <= not w44027 and not w44111;
w44113 <= b(8) and not w44016;
w44114 <= not w44014 and w44113;
w44115 <= not w44018 and not w44114;
w44116 <= not w44112 and w44115;
w44117 <= not w44018 and not w44116;
w44118 <= b(9) and not w44007;
w44119 <= not w44005 and w44118;
w44120 <= not w44009 and not w44119;
w44121 <= not w44117 and w44120;
w44122 <= not w44009 and not w44121;
w44123 <= b(10) and not w43998;
w44124 <= not w43996 and w44123;
w44125 <= not w44000 and not w44124;
w44126 <= not w44122 and w44125;
w44127 <= not w44000 and not w44126;
w44128 <= b(11) and not w43989;
w44129 <= not w43987 and w44128;
w44130 <= not w43991 and not w44129;
w44131 <= not w44127 and w44130;
w44132 <= not w43991 and not w44131;
w44133 <= b(12) and not w43980;
w44134 <= not w43978 and w44133;
w44135 <= not w43982 and not w44134;
w44136 <= not w44132 and w44135;
w44137 <= not w43982 and not w44136;
w44138 <= b(13) and not w43971;
w44139 <= not w43969 and w44138;
w44140 <= not w43973 and not w44139;
w44141 <= not w44137 and w44140;
w44142 <= not w43973 and not w44141;
w44143 <= b(14) and not w43962;
w44144 <= not w43960 and w44143;
w44145 <= not w43964 and not w44144;
w44146 <= not w44142 and w44145;
w44147 <= not w43964 and not w44146;
w44148 <= b(15) and not w43953;
w44149 <= not w43951 and w44148;
w44150 <= not w43955 and not w44149;
w44151 <= not w44147 and w44150;
w44152 <= not w43955 and not w44151;
w44153 <= b(16) and not w43944;
w44154 <= not w43942 and w44153;
w44155 <= not w43946 and not w44154;
w44156 <= not w44152 and w44155;
w44157 <= not w43946 and not w44156;
w44158 <= b(17) and not w43935;
w44159 <= not w43933 and w44158;
w44160 <= not w43937 and not w44159;
w44161 <= not w44157 and w44160;
w44162 <= not w43937 and not w44161;
w44163 <= b(18) and not w43926;
w44164 <= not w43924 and w44163;
w44165 <= not w43928 and not w44164;
w44166 <= not w44162 and w44165;
w44167 <= not w43928 and not w44166;
w44168 <= b(19) and not w43917;
w44169 <= not w43915 and w44168;
w44170 <= not w43919 and not w44169;
w44171 <= not w44167 and w44170;
w44172 <= not w43919 and not w44171;
w44173 <= b(20) and not w43908;
w44174 <= not w43906 and w44173;
w44175 <= not w43910 and not w44174;
w44176 <= not w44172 and w44175;
w44177 <= not w43910 and not w44176;
w44178 <= b(21) and not w43899;
w44179 <= not w43897 and w44178;
w44180 <= not w43901 and not w44179;
w44181 <= not w44177 and w44180;
w44182 <= not w43901 and not w44181;
w44183 <= b(22) and not w43890;
w44184 <= not w43888 and w44183;
w44185 <= not w43892 and not w44184;
w44186 <= not w44182 and w44185;
w44187 <= not w43892 and not w44186;
w44188 <= b(23) and not w43881;
w44189 <= not w43879 and w44188;
w44190 <= not w43883 and not w44189;
w44191 <= not w44187 and w44190;
w44192 <= not w43883 and not w44191;
w44193 <= b(24) and not w43872;
w44194 <= not w43870 and w44193;
w44195 <= not w43874 and not w44194;
w44196 <= not w44192 and w44195;
w44197 <= not w43874 and not w44196;
w44198 <= b(25) and not w43863;
w44199 <= not w43861 and w44198;
w44200 <= not w43865 and not w44199;
w44201 <= not w44197 and w44200;
w44202 <= not w43865 and not w44201;
w44203 <= b(26) and not w43854;
w44204 <= not w43852 and w44203;
w44205 <= not w43856 and not w44204;
w44206 <= not w44202 and w44205;
w44207 <= not w43856 and not w44206;
w44208 <= b(27) and not w43845;
w44209 <= not w43843 and w44208;
w44210 <= not w43847 and not w44209;
w44211 <= not w44207 and w44210;
w44212 <= not w43847 and not w44211;
w44213 <= b(28) and not w43836;
w44214 <= not w43834 and w44213;
w44215 <= not w43838 and not w44214;
w44216 <= not w44212 and w44215;
w44217 <= not w43838 and not w44216;
w44218 <= b(29) and not w43827;
w44219 <= not w43825 and w44218;
w44220 <= not w43829 and not w44219;
w44221 <= not w44217 and w44220;
w44222 <= not w43829 and not w44221;
w44223 <= b(30) and not w43818;
w44224 <= not w43816 and w44223;
w44225 <= not w43820 and not w44224;
w44226 <= not w44222 and w44225;
w44227 <= not w43820 and not w44226;
w44228 <= b(31) and not w43809;
w44229 <= not w43807 and w44228;
w44230 <= not w43811 and not w44229;
w44231 <= not w44227 and w44230;
w44232 <= not w43811 and not w44231;
w44233 <= b(32) and not w43800;
w44234 <= not w43798 and w44233;
w44235 <= not w43802 and not w44234;
w44236 <= not w44232 and w44235;
w44237 <= not w43802 and not w44236;
w44238 <= b(33) and not w43791;
w44239 <= not w43789 and w44238;
w44240 <= not w43793 and not w44239;
w44241 <= not w44237 and w44240;
w44242 <= not w43793 and not w44241;
w44243 <= b(34) and not w43782;
w44244 <= not w43780 and w44243;
w44245 <= not w43784 and not w44244;
w44246 <= not w44242 and w44245;
w44247 <= not w43784 and not w44246;
w44248 <= b(35) and not w43773;
w44249 <= not w43771 and w44248;
w44250 <= not w43775 and not w44249;
w44251 <= not w44247 and w44250;
w44252 <= not w43775 and not w44251;
w44253 <= b(36) and not w43764;
w44254 <= not w43762 and w44253;
w44255 <= not w43766 and not w44254;
w44256 <= not w44252 and w44255;
w44257 <= not w43766 and not w44256;
w44258 <= b(37) and not w43755;
w44259 <= not w43753 and w44258;
w44260 <= not w43757 and not w44259;
w44261 <= not w44257 and w44260;
w44262 <= not w43757 and not w44261;
w44263 <= b(38) and not w43746;
w44264 <= not w43744 and w44263;
w44265 <= not w43748 and not w44264;
w44266 <= not w44262 and w44265;
w44267 <= not w43748 and not w44266;
w44268 <= b(39) and not w43737;
w44269 <= not w43735 and w44268;
w44270 <= not w43739 and not w44269;
w44271 <= not w44267 and w44270;
w44272 <= not w43739 and not w44271;
w44273 <= b(40) and not w43728;
w44274 <= not w43726 and w44273;
w44275 <= not w43730 and not w44274;
w44276 <= not w44272 and w44275;
w44277 <= not w43730 and not w44276;
w44278 <= b(41) and not w43719;
w44279 <= not w43717 and w44278;
w44280 <= not w43721 and not w44279;
w44281 <= not w44277 and w44280;
w44282 <= not w43721 and not w44281;
w44283 <= b(42) and not w43710;
w44284 <= not w43708 and w44283;
w44285 <= not w43712 and not w44284;
w44286 <= not w44282 and w44285;
w44287 <= not w43712 and not w44286;
w44288 <= b(43) and not w43701;
w44289 <= not w43699 and w44288;
w44290 <= not w43703 and not w44289;
w44291 <= not w44287 and w44290;
w44292 <= not w43703 and not w44291;
w44293 <= b(44) and not w43692;
w44294 <= not w43690 and w44293;
w44295 <= not w43694 and not w44294;
w44296 <= not w44292 and w44295;
w44297 <= not w43694 and not w44296;
w44298 <= b(45) and not w43683;
w44299 <= not w43681 and w44298;
w44300 <= not w43685 and not w44299;
w44301 <= not w44297 and w44300;
w44302 <= not w43685 and not w44301;
w44303 <= b(46) and not w43674;
w44304 <= not w43672 and w44303;
w44305 <= not w43676 and not w44304;
w44306 <= not w44302 and w44305;
w44307 <= not w43676 and not w44306;
w44308 <= not w43035 and not w43662;
w44309 <= not w43660 and w44308;
w44310 <= not w43651 and w44309;
w44311 <= not w43660 and not w43662;
w44312 <= not w43652 and not w44311;
w44313 <= not w44310 and not w44312;
w44314 <= not w43667 and not w44313;
w44315 <= not w43659 and not w43666;
w44316 <= not w43665 and w44315;
w44317 <= not w44314 and not w44316;
w44318 <= not b(47) and not w44317;
w44319 <= b(47) and not w44316;
w44320 <= not w44314 and w44319;
w44321 <= w81 and not w44320;
w44322 <= not w44318 and w44321;
w44323 <= not w44307 and w44322;
w44324 <= w15602 and not w44317;
w44325 <= not w44323 and not w44324;
w44326 <= not w43685 and w44305;
w44327 <= not w44301 and w44326;
w44328 <= not w44302 and not w44305;
w44329 <= not w44327 and not w44328;
w44330 <= not w44325 and not w44329;
w44331 <= not w43675 and not w44324;
w44332 <= not w44323 and w44331;
w44333 <= not w44330 and not w44332;
w44334 <= not w43676 and not w44320;
w44335 <= not w44318 and w44334;
w44336 <= not w44306 and w44335;
w44337 <= not w44318 and not w44320;
w44338 <= not w44307 and not w44337;
w44339 <= not w44336 and not w44338;
w44340 <= not w44325 and not w44339;
w44341 <= not w44317 and not w44324;
w44342 <= not w44323 and w44341;
w44343 <= not w44340 and not w44342;
w44344 <= not b(48) and not w44343;
w44345 <= not b(47) and not w44333;
w44346 <= not w43694 and w44300;
w44347 <= not w44296 and w44346;
w44348 <= not w44297 and not w44300;
w44349 <= not w44347 and not w44348;
w44350 <= not w44325 and not w44349;
w44351 <= not w43684 and not w44324;
w44352 <= not w44323 and w44351;
w44353 <= not w44350 and not w44352;
w44354 <= not b(46) and not w44353;
w44355 <= not w43703 and w44295;
w44356 <= not w44291 and w44355;
w44357 <= not w44292 and not w44295;
w44358 <= not w44356 and not w44357;
w44359 <= not w44325 and not w44358;
w44360 <= not w43693 and not w44324;
w44361 <= not w44323 and w44360;
w44362 <= not w44359 and not w44361;
w44363 <= not b(45) and not w44362;
w44364 <= not w43712 and w44290;
w44365 <= not w44286 and w44364;
w44366 <= not w44287 and not w44290;
w44367 <= not w44365 and not w44366;
w44368 <= not w44325 and not w44367;
w44369 <= not w43702 and not w44324;
w44370 <= not w44323 and w44369;
w44371 <= not w44368 and not w44370;
w44372 <= not b(44) and not w44371;
w44373 <= not w43721 and w44285;
w44374 <= not w44281 and w44373;
w44375 <= not w44282 and not w44285;
w44376 <= not w44374 and not w44375;
w44377 <= not w44325 and not w44376;
w44378 <= not w43711 and not w44324;
w44379 <= not w44323 and w44378;
w44380 <= not w44377 and not w44379;
w44381 <= not b(43) and not w44380;
w44382 <= not w43730 and w44280;
w44383 <= not w44276 and w44382;
w44384 <= not w44277 and not w44280;
w44385 <= not w44383 and not w44384;
w44386 <= not w44325 and not w44385;
w44387 <= not w43720 and not w44324;
w44388 <= not w44323 and w44387;
w44389 <= not w44386 and not w44388;
w44390 <= not b(42) and not w44389;
w44391 <= not w43739 and w44275;
w44392 <= not w44271 and w44391;
w44393 <= not w44272 and not w44275;
w44394 <= not w44392 and not w44393;
w44395 <= not w44325 and not w44394;
w44396 <= not w43729 and not w44324;
w44397 <= not w44323 and w44396;
w44398 <= not w44395 and not w44397;
w44399 <= not b(41) and not w44398;
w44400 <= not w43748 and w44270;
w44401 <= not w44266 and w44400;
w44402 <= not w44267 and not w44270;
w44403 <= not w44401 and not w44402;
w44404 <= not w44325 and not w44403;
w44405 <= not w43738 and not w44324;
w44406 <= not w44323 and w44405;
w44407 <= not w44404 and not w44406;
w44408 <= not b(40) and not w44407;
w44409 <= not w43757 and w44265;
w44410 <= not w44261 and w44409;
w44411 <= not w44262 and not w44265;
w44412 <= not w44410 and not w44411;
w44413 <= not w44325 and not w44412;
w44414 <= not w43747 and not w44324;
w44415 <= not w44323 and w44414;
w44416 <= not w44413 and not w44415;
w44417 <= not b(39) and not w44416;
w44418 <= not w43766 and w44260;
w44419 <= not w44256 and w44418;
w44420 <= not w44257 and not w44260;
w44421 <= not w44419 and not w44420;
w44422 <= not w44325 and not w44421;
w44423 <= not w43756 and not w44324;
w44424 <= not w44323 and w44423;
w44425 <= not w44422 and not w44424;
w44426 <= not b(38) and not w44425;
w44427 <= not w43775 and w44255;
w44428 <= not w44251 and w44427;
w44429 <= not w44252 and not w44255;
w44430 <= not w44428 and not w44429;
w44431 <= not w44325 and not w44430;
w44432 <= not w43765 and not w44324;
w44433 <= not w44323 and w44432;
w44434 <= not w44431 and not w44433;
w44435 <= not b(37) and not w44434;
w44436 <= not w43784 and w44250;
w44437 <= not w44246 and w44436;
w44438 <= not w44247 and not w44250;
w44439 <= not w44437 and not w44438;
w44440 <= not w44325 and not w44439;
w44441 <= not w43774 and not w44324;
w44442 <= not w44323 and w44441;
w44443 <= not w44440 and not w44442;
w44444 <= not b(36) and not w44443;
w44445 <= not w43793 and w44245;
w44446 <= not w44241 and w44445;
w44447 <= not w44242 and not w44245;
w44448 <= not w44446 and not w44447;
w44449 <= not w44325 and not w44448;
w44450 <= not w43783 and not w44324;
w44451 <= not w44323 and w44450;
w44452 <= not w44449 and not w44451;
w44453 <= not b(35) and not w44452;
w44454 <= not w43802 and w44240;
w44455 <= not w44236 and w44454;
w44456 <= not w44237 and not w44240;
w44457 <= not w44455 and not w44456;
w44458 <= not w44325 and not w44457;
w44459 <= not w43792 and not w44324;
w44460 <= not w44323 and w44459;
w44461 <= not w44458 and not w44460;
w44462 <= not b(34) and not w44461;
w44463 <= not w43811 and w44235;
w44464 <= not w44231 and w44463;
w44465 <= not w44232 and not w44235;
w44466 <= not w44464 and not w44465;
w44467 <= not w44325 and not w44466;
w44468 <= not w43801 and not w44324;
w44469 <= not w44323 and w44468;
w44470 <= not w44467 and not w44469;
w44471 <= not b(33) and not w44470;
w44472 <= not w43820 and w44230;
w44473 <= not w44226 and w44472;
w44474 <= not w44227 and not w44230;
w44475 <= not w44473 and not w44474;
w44476 <= not w44325 and not w44475;
w44477 <= not w43810 and not w44324;
w44478 <= not w44323 and w44477;
w44479 <= not w44476 and not w44478;
w44480 <= not b(32) and not w44479;
w44481 <= not w43829 and w44225;
w44482 <= not w44221 and w44481;
w44483 <= not w44222 and not w44225;
w44484 <= not w44482 and not w44483;
w44485 <= not w44325 and not w44484;
w44486 <= not w43819 and not w44324;
w44487 <= not w44323 and w44486;
w44488 <= not w44485 and not w44487;
w44489 <= not b(31) and not w44488;
w44490 <= not w43838 and w44220;
w44491 <= not w44216 and w44490;
w44492 <= not w44217 and not w44220;
w44493 <= not w44491 and not w44492;
w44494 <= not w44325 and not w44493;
w44495 <= not w43828 and not w44324;
w44496 <= not w44323 and w44495;
w44497 <= not w44494 and not w44496;
w44498 <= not b(30) and not w44497;
w44499 <= not w43847 and w44215;
w44500 <= not w44211 and w44499;
w44501 <= not w44212 and not w44215;
w44502 <= not w44500 and not w44501;
w44503 <= not w44325 and not w44502;
w44504 <= not w43837 and not w44324;
w44505 <= not w44323 and w44504;
w44506 <= not w44503 and not w44505;
w44507 <= not b(29) and not w44506;
w44508 <= not w43856 and w44210;
w44509 <= not w44206 and w44508;
w44510 <= not w44207 and not w44210;
w44511 <= not w44509 and not w44510;
w44512 <= not w44325 and not w44511;
w44513 <= not w43846 and not w44324;
w44514 <= not w44323 and w44513;
w44515 <= not w44512 and not w44514;
w44516 <= not b(28) and not w44515;
w44517 <= not w43865 and w44205;
w44518 <= not w44201 and w44517;
w44519 <= not w44202 and not w44205;
w44520 <= not w44518 and not w44519;
w44521 <= not w44325 and not w44520;
w44522 <= not w43855 and not w44324;
w44523 <= not w44323 and w44522;
w44524 <= not w44521 and not w44523;
w44525 <= not b(27) and not w44524;
w44526 <= not w43874 and w44200;
w44527 <= not w44196 and w44526;
w44528 <= not w44197 and not w44200;
w44529 <= not w44527 and not w44528;
w44530 <= not w44325 and not w44529;
w44531 <= not w43864 and not w44324;
w44532 <= not w44323 and w44531;
w44533 <= not w44530 and not w44532;
w44534 <= not b(26) and not w44533;
w44535 <= not w43883 and w44195;
w44536 <= not w44191 and w44535;
w44537 <= not w44192 and not w44195;
w44538 <= not w44536 and not w44537;
w44539 <= not w44325 and not w44538;
w44540 <= not w43873 and not w44324;
w44541 <= not w44323 and w44540;
w44542 <= not w44539 and not w44541;
w44543 <= not b(25) and not w44542;
w44544 <= not w43892 and w44190;
w44545 <= not w44186 and w44544;
w44546 <= not w44187 and not w44190;
w44547 <= not w44545 and not w44546;
w44548 <= not w44325 and not w44547;
w44549 <= not w43882 and not w44324;
w44550 <= not w44323 and w44549;
w44551 <= not w44548 and not w44550;
w44552 <= not b(24) and not w44551;
w44553 <= not w43901 and w44185;
w44554 <= not w44181 and w44553;
w44555 <= not w44182 and not w44185;
w44556 <= not w44554 and not w44555;
w44557 <= not w44325 and not w44556;
w44558 <= not w43891 and not w44324;
w44559 <= not w44323 and w44558;
w44560 <= not w44557 and not w44559;
w44561 <= not b(23) and not w44560;
w44562 <= not w43910 and w44180;
w44563 <= not w44176 and w44562;
w44564 <= not w44177 and not w44180;
w44565 <= not w44563 and not w44564;
w44566 <= not w44325 and not w44565;
w44567 <= not w43900 and not w44324;
w44568 <= not w44323 and w44567;
w44569 <= not w44566 and not w44568;
w44570 <= not b(22) and not w44569;
w44571 <= not w43919 and w44175;
w44572 <= not w44171 and w44571;
w44573 <= not w44172 and not w44175;
w44574 <= not w44572 and not w44573;
w44575 <= not w44325 and not w44574;
w44576 <= not w43909 and not w44324;
w44577 <= not w44323 and w44576;
w44578 <= not w44575 and not w44577;
w44579 <= not b(21) and not w44578;
w44580 <= not w43928 and w44170;
w44581 <= not w44166 and w44580;
w44582 <= not w44167 and not w44170;
w44583 <= not w44581 and not w44582;
w44584 <= not w44325 and not w44583;
w44585 <= not w43918 and not w44324;
w44586 <= not w44323 and w44585;
w44587 <= not w44584 and not w44586;
w44588 <= not b(20) and not w44587;
w44589 <= not w43937 and w44165;
w44590 <= not w44161 and w44589;
w44591 <= not w44162 and not w44165;
w44592 <= not w44590 and not w44591;
w44593 <= not w44325 and not w44592;
w44594 <= not w43927 and not w44324;
w44595 <= not w44323 and w44594;
w44596 <= not w44593 and not w44595;
w44597 <= not b(19) and not w44596;
w44598 <= not w43946 and w44160;
w44599 <= not w44156 and w44598;
w44600 <= not w44157 and not w44160;
w44601 <= not w44599 and not w44600;
w44602 <= not w44325 and not w44601;
w44603 <= not w43936 and not w44324;
w44604 <= not w44323 and w44603;
w44605 <= not w44602 and not w44604;
w44606 <= not b(18) and not w44605;
w44607 <= not w43955 and w44155;
w44608 <= not w44151 and w44607;
w44609 <= not w44152 and not w44155;
w44610 <= not w44608 and not w44609;
w44611 <= not w44325 and not w44610;
w44612 <= not w43945 and not w44324;
w44613 <= not w44323 and w44612;
w44614 <= not w44611 and not w44613;
w44615 <= not b(17) and not w44614;
w44616 <= not w43964 and w44150;
w44617 <= not w44146 and w44616;
w44618 <= not w44147 and not w44150;
w44619 <= not w44617 and not w44618;
w44620 <= not w44325 and not w44619;
w44621 <= not w43954 and not w44324;
w44622 <= not w44323 and w44621;
w44623 <= not w44620 and not w44622;
w44624 <= not b(16) and not w44623;
w44625 <= not w43973 and w44145;
w44626 <= not w44141 and w44625;
w44627 <= not w44142 and not w44145;
w44628 <= not w44626 and not w44627;
w44629 <= not w44325 and not w44628;
w44630 <= not w43963 and not w44324;
w44631 <= not w44323 and w44630;
w44632 <= not w44629 and not w44631;
w44633 <= not b(15) and not w44632;
w44634 <= not w43982 and w44140;
w44635 <= not w44136 and w44634;
w44636 <= not w44137 and not w44140;
w44637 <= not w44635 and not w44636;
w44638 <= not w44325 and not w44637;
w44639 <= not w43972 and not w44324;
w44640 <= not w44323 and w44639;
w44641 <= not w44638 and not w44640;
w44642 <= not b(14) and not w44641;
w44643 <= not w43991 and w44135;
w44644 <= not w44131 and w44643;
w44645 <= not w44132 and not w44135;
w44646 <= not w44644 and not w44645;
w44647 <= not w44325 and not w44646;
w44648 <= not w43981 and not w44324;
w44649 <= not w44323 and w44648;
w44650 <= not w44647 and not w44649;
w44651 <= not b(13) and not w44650;
w44652 <= not w44000 and w44130;
w44653 <= not w44126 and w44652;
w44654 <= not w44127 and not w44130;
w44655 <= not w44653 and not w44654;
w44656 <= not w44325 and not w44655;
w44657 <= not w43990 and not w44324;
w44658 <= not w44323 and w44657;
w44659 <= not w44656 and not w44658;
w44660 <= not b(12) and not w44659;
w44661 <= not w44009 and w44125;
w44662 <= not w44121 and w44661;
w44663 <= not w44122 and not w44125;
w44664 <= not w44662 and not w44663;
w44665 <= not w44325 and not w44664;
w44666 <= not w43999 and not w44324;
w44667 <= not w44323 and w44666;
w44668 <= not w44665 and not w44667;
w44669 <= not b(11) and not w44668;
w44670 <= not w44018 and w44120;
w44671 <= not w44116 and w44670;
w44672 <= not w44117 and not w44120;
w44673 <= not w44671 and not w44672;
w44674 <= not w44325 and not w44673;
w44675 <= not w44008 and not w44324;
w44676 <= not w44323 and w44675;
w44677 <= not w44674 and not w44676;
w44678 <= not b(10) and not w44677;
w44679 <= not w44027 and w44115;
w44680 <= not w44111 and w44679;
w44681 <= not w44112 and not w44115;
w44682 <= not w44680 and not w44681;
w44683 <= not w44325 and not w44682;
w44684 <= not w44017 and not w44324;
w44685 <= not w44323 and w44684;
w44686 <= not w44683 and not w44685;
w44687 <= not b(9) and not w44686;
w44688 <= not w44036 and w44110;
w44689 <= not w44106 and w44688;
w44690 <= not w44107 and not w44110;
w44691 <= not w44689 and not w44690;
w44692 <= not w44325 and not w44691;
w44693 <= not w44026 and not w44324;
w44694 <= not w44323 and w44693;
w44695 <= not w44692 and not w44694;
w44696 <= not b(8) and not w44695;
w44697 <= not w44045 and w44105;
w44698 <= not w44101 and w44697;
w44699 <= not w44102 and not w44105;
w44700 <= not w44698 and not w44699;
w44701 <= not w44325 and not w44700;
w44702 <= not w44035 and not w44324;
w44703 <= not w44323 and w44702;
w44704 <= not w44701 and not w44703;
w44705 <= not b(7) and not w44704;
w44706 <= not w44054 and w44100;
w44707 <= not w44096 and w44706;
w44708 <= not w44097 and not w44100;
w44709 <= not w44707 and not w44708;
w44710 <= not w44325 and not w44709;
w44711 <= not w44044 and not w44324;
w44712 <= not w44323 and w44711;
w44713 <= not w44710 and not w44712;
w44714 <= not b(6) and not w44713;
w44715 <= not w44063 and w44095;
w44716 <= not w44091 and w44715;
w44717 <= not w44092 and not w44095;
w44718 <= not w44716 and not w44717;
w44719 <= not w44325 and not w44718;
w44720 <= not w44053 and not w44324;
w44721 <= not w44323 and w44720;
w44722 <= not w44719 and not w44721;
w44723 <= not b(5) and not w44722;
w44724 <= not w44071 and w44090;
w44725 <= not w44086 and w44724;
w44726 <= not w44087 and not w44090;
w44727 <= not w44725 and not w44726;
w44728 <= not w44325 and not w44727;
w44729 <= not w44062 and not w44324;
w44730 <= not w44323 and w44729;
w44731 <= not w44728 and not w44730;
w44732 <= not b(4) and not w44731;
w44733 <= not w44081 and w44085;
w44734 <= not w44080 and w44733;
w44735 <= not w44082 and not w44085;
w44736 <= not w44734 and not w44735;
w44737 <= not w44325 and not w44736;
w44738 <= not w44070 and not w44324;
w44739 <= not w44323 and w44738;
w44740 <= not w44737 and not w44739;
w44741 <= not b(3) and not w44740;
w44742 <= w16020 and not w44078;
w44743 <= not w44076 and w44742;
w44744 <= not w44080 and not w44743;
w44745 <= not w44325 and w44744;
w44746 <= not w44075 and not w44324;
w44747 <= not w44323 and w44746;
w44748 <= not w44745 and not w44747;
w44749 <= not b(2) and not w44748;
w44750 <= b(0) and not w44325;
w44751 <= a(16) and not w44750;
w44752 <= w16020 and not w44325;
w44753 <= not w44751 and not w44752;
w44754 <= b(1) and not w44753;
w44755 <= not b(1) and not w44752;
w44756 <= not w44751 and w44755;
w44757 <= not w44754 and not w44756;
w44758 <= not w16699 and not w44757;
w44759 <= not b(1) and not w44753;
w44760 <= not w44758 and not w44759;
w44761 <= b(2) and not w44747;
w44762 <= not w44745 and w44761;
w44763 <= not w44749 and not w44762;
w44764 <= not w44760 and w44763;
w44765 <= not w44749 and not w44764;
w44766 <= b(3) and not w44739;
w44767 <= not w44737 and w44766;
w44768 <= not w44741 and not w44767;
w44769 <= not w44765 and w44768;
w44770 <= not w44741 and not w44769;
w44771 <= b(4) and not w44730;
w44772 <= not w44728 and w44771;
w44773 <= not w44732 and not w44772;
w44774 <= not w44770 and w44773;
w44775 <= not w44732 and not w44774;
w44776 <= b(5) and not w44721;
w44777 <= not w44719 and w44776;
w44778 <= not w44723 and not w44777;
w44779 <= not w44775 and w44778;
w44780 <= not w44723 and not w44779;
w44781 <= b(6) and not w44712;
w44782 <= not w44710 and w44781;
w44783 <= not w44714 and not w44782;
w44784 <= not w44780 and w44783;
w44785 <= not w44714 and not w44784;
w44786 <= b(7) and not w44703;
w44787 <= not w44701 and w44786;
w44788 <= not w44705 and not w44787;
w44789 <= not w44785 and w44788;
w44790 <= not w44705 and not w44789;
w44791 <= b(8) and not w44694;
w44792 <= not w44692 and w44791;
w44793 <= not w44696 and not w44792;
w44794 <= not w44790 and w44793;
w44795 <= not w44696 and not w44794;
w44796 <= b(9) and not w44685;
w44797 <= not w44683 and w44796;
w44798 <= not w44687 and not w44797;
w44799 <= not w44795 and w44798;
w44800 <= not w44687 and not w44799;
w44801 <= b(10) and not w44676;
w44802 <= not w44674 and w44801;
w44803 <= not w44678 and not w44802;
w44804 <= not w44800 and w44803;
w44805 <= not w44678 and not w44804;
w44806 <= b(11) and not w44667;
w44807 <= not w44665 and w44806;
w44808 <= not w44669 and not w44807;
w44809 <= not w44805 and w44808;
w44810 <= not w44669 and not w44809;
w44811 <= b(12) and not w44658;
w44812 <= not w44656 and w44811;
w44813 <= not w44660 and not w44812;
w44814 <= not w44810 and w44813;
w44815 <= not w44660 and not w44814;
w44816 <= b(13) and not w44649;
w44817 <= not w44647 and w44816;
w44818 <= not w44651 and not w44817;
w44819 <= not w44815 and w44818;
w44820 <= not w44651 and not w44819;
w44821 <= b(14) and not w44640;
w44822 <= not w44638 and w44821;
w44823 <= not w44642 and not w44822;
w44824 <= not w44820 and w44823;
w44825 <= not w44642 and not w44824;
w44826 <= b(15) and not w44631;
w44827 <= not w44629 and w44826;
w44828 <= not w44633 and not w44827;
w44829 <= not w44825 and w44828;
w44830 <= not w44633 and not w44829;
w44831 <= b(16) and not w44622;
w44832 <= not w44620 and w44831;
w44833 <= not w44624 and not w44832;
w44834 <= not w44830 and w44833;
w44835 <= not w44624 and not w44834;
w44836 <= b(17) and not w44613;
w44837 <= not w44611 and w44836;
w44838 <= not w44615 and not w44837;
w44839 <= not w44835 and w44838;
w44840 <= not w44615 and not w44839;
w44841 <= b(18) and not w44604;
w44842 <= not w44602 and w44841;
w44843 <= not w44606 and not w44842;
w44844 <= not w44840 and w44843;
w44845 <= not w44606 and not w44844;
w44846 <= b(19) and not w44595;
w44847 <= not w44593 and w44846;
w44848 <= not w44597 and not w44847;
w44849 <= not w44845 and w44848;
w44850 <= not w44597 and not w44849;
w44851 <= b(20) and not w44586;
w44852 <= not w44584 and w44851;
w44853 <= not w44588 and not w44852;
w44854 <= not w44850 and w44853;
w44855 <= not w44588 and not w44854;
w44856 <= b(21) and not w44577;
w44857 <= not w44575 and w44856;
w44858 <= not w44579 and not w44857;
w44859 <= not w44855 and w44858;
w44860 <= not w44579 and not w44859;
w44861 <= b(22) and not w44568;
w44862 <= not w44566 and w44861;
w44863 <= not w44570 and not w44862;
w44864 <= not w44860 and w44863;
w44865 <= not w44570 and not w44864;
w44866 <= b(23) and not w44559;
w44867 <= not w44557 and w44866;
w44868 <= not w44561 and not w44867;
w44869 <= not w44865 and w44868;
w44870 <= not w44561 and not w44869;
w44871 <= b(24) and not w44550;
w44872 <= not w44548 and w44871;
w44873 <= not w44552 and not w44872;
w44874 <= not w44870 and w44873;
w44875 <= not w44552 and not w44874;
w44876 <= b(25) and not w44541;
w44877 <= not w44539 and w44876;
w44878 <= not w44543 and not w44877;
w44879 <= not w44875 and w44878;
w44880 <= not w44543 and not w44879;
w44881 <= b(26) and not w44532;
w44882 <= not w44530 and w44881;
w44883 <= not w44534 and not w44882;
w44884 <= not w44880 and w44883;
w44885 <= not w44534 and not w44884;
w44886 <= b(27) and not w44523;
w44887 <= not w44521 and w44886;
w44888 <= not w44525 and not w44887;
w44889 <= not w44885 and w44888;
w44890 <= not w44525 and not w44889;
w44891 <= b(28) and not w44514;
w44892 <= not w44512 and w44891;
w44893 <= not w44516 and not w44892;
w44894 <= not w44890 and w44893;
w44895 <= not w44516 and not w44894;
w44896 <= b(29) and not w44505;
w44897 <= not w44503 and w44896;
w44898 <= not w44507 and not w44897;
w44899 <= not w44895 and w44898;
w44900 <= not w44507 and not w44899;
w44901 <= b(30) and not w44496;
w44902 <= not w44494 and w44901;
w44903 <= not w44498 and not w44902;
w44904 <= not w44900 and w44903;
w44905 <= not w44498 and not w44904;
w44906 <= b(31) and not w44487;
w44907 <= not w44485 and w44906;
w44908 <= not w44489 and not w44907;
w44909 <= not w44905 and w44908;
w44910 <= not w44489 and not w44909;
w44911 <= b(32) and not w44478;
w44912 <= not w44476 and w44911;
w44913 <= not w44480 and not w44912;
w44914 <= not w44910 and w44913;
w44915 <= not w44480 and not w44914;
w44916 <= b(33) and not w44469;
w44917 <= not w44467 and w44916;
w44918 <= not w44471 and not w44917;
w44919 <= not w44915 and w44918;
w44920 <= not w44471 and not w44919;
w44921 <= b(34) and not w44460;
w44922 <= not w44458 and w44921;
w44923 <= not w44462 and not w44922;
w44924 <= not w44920 and w44923;
w44925 <= not w44462 and not w44924;
w44926 <= b(35) and not w44451;
w44927 <= not w44449 and w44926;
w44928 <= not w44453 and not w44927;
w44929 <= not w44925 and w44928;
w44930 <= not w44453 and not w44929;
w44931 <= b(36) and not w44442;
w44932 <= not w44440 and w44931;
w44933 <= not w44444 and not w44932;
w44934 <= not w44930 and w44933;
w44935 <= not w44444 and not w44934;
w44936 <= b(37) and not w44433;
w44937 <= not w44431 and w44936;
w44938 <= not w44435 and not w44937;
w44939 <= not w44935 and w44938;
w44940 <= not w44435 and not w44939;
w44941 <= b(38) and not w44424;
w44942 <= not w44422 and w44941;
w44943 <= not w44426 and not w44942;
w44944 <= not w44940 and w44943;
w44945 <= not w44426 and not w44944;
w44946 <= b(39) and not w44415;
w44947 <= not w44413 and w44946;
w44948 <= not w44417 and not w44947;
w44949 <= not w44945 and w44948;
w44950 <= not w44417 and not w44949;
w44951 <= b(40) and not w44406;
w44952 <= not w44404 and w44951;
w44953 <= not w44408 and not w44952;
w44954 <= not w44950 and w44953;
w44955 <= not w44408 and not w44954;
w44956 <= b(41) and not w44397;
w44957 <= not w44395 and w44956;
w44958 <= not w44399 and not w44957;
w44959 <= not w44955 and w44958;
w44960 <= not w44399 and not w44959;
w44961 <= b(42) and not w44388;
w44962 <= not w44386 and w44961;
w44963 <= not w44390 and not w44962;
w44964 <= not w44960 and w44963;
w44965 <= not w44390 and not w44964;
w44966 <= b(43) and not w44379;
w44967 <= not w44377 and w44966;
w44968 <= not w44381 and not w44967;
w44969 <= not w44965 and w44968;
w44970 <= not w44381 and not w44969;
w44971 <= b(44) and not w44370;
w44972 <= not w44368 and w44971;
w44973 <= not w44372 and not w44972;
w44974 <= not w44970 and w44973;
w44975 <= not w44372 and not w44974;
w44976 <= b(45) and not w44361;
w44977 <= not w44359 and w44976;
w44978 <= not w44363 and not w44977;
w44979 <= not w44975 and w44978;
w44980 <= not w44363 and not w44979;
w44981 <= b(46) and not w44352;
w44982 <= not w44350 and w44981;
w44983 <= not w44354 and not w44982;
w44984 <= not w44980 and w44983;
w44985 <= not w44354 and not w44984;
w44986 <= b(47) and not w44332;
w44987 <= not w44330 and w44986;
w44988 <= not w44345 and not w44987;
w44989 <= not w44985 and w44988;
w44990 <= not w44345 and not w44989;
w44991 <= b(48) and not w44342;
w44992 <= not w44340 and w44991;
w44993 <= not w44344 and not w44992;
w44994 <= not w44990 and w44993;
w44995 <= not w44344 and not w44994;
w44996 <= w151 and not w44995;
w44997 <= not w44333 and not w44996;
w44998 <= not w44354 and w44988;
w44999 <= not w44984 and w44998;
w45000 <= not w44985 and not w44988;
w45001 <= not w44999 and not w45000;
w45002 <= w151 and not w45001;
w45003 <= not w44995 and w45002;
w45004 <= not w44997 and not w45003;
w45005 <= not b(48) and not w45004;
w45006 <= not w44353 and not w44996;
w45007 <= not w44363 and w44983;
w45008 <= not w44979 and w45007;
w45009 <= not w44980 and not w44983;
w45010 <= not w45008 and not w45009;
w45011 <= w151 and not w45010;
w45012 <= not w44995 and w45011;
w45013 <= not w45006 and not w45012;
w45014 <= not b(47) and not w45013;
w45015 <= not w44362 and not w44996;
w45016 <= not w44372 and w44978;
w45017 <= not w44974 and w45016;
w45018 <= not w44975 and not w44978;
w45019 <= not w45017 and not w45018;
w45020 <= w151 and not w45019;
w45021 <= not w44995 and w45020;
w45022 <= not w45015 and not w45021;
w45023 <= not b(46) and not w45022;
w45024 <= not w44371 and not w44996;
w45025 <= not w44381 and w44973;
w45026 <= not w44969 and w45025;
w45027 <= not w44970 and not w44973;
w45028 <= not w45026 and not w45027;
w45029 <= w151 and not w45028;
w45030 <= not w44995 and w45029;
w45031 <= not w45024 and not w45030;
w45032 <= not b(45) and not w45031;
w45033 <= not w44380 and not w44996;
w45034 <= not w44390 and w44968;
w45035 <= not w44964 and w45034;
w45036 <= not w44965 and not w44968;
w45037 <= not w45035 and not w45036;
w45038 <= w151 and not w45037;
w45039 <= not w44995 and w45038;
w45040 <= not w45033 and not w45039;
w45041 <= not b(44) and not w45040;
w45042 <= not w44389 and not w44996;
w45043 <= not w44399 and w44963;
w45044 <= not w44959 and w45043;
w45045 <= not w44960 and not w44963;
w45046 <= not w45044 and not w45045;
w45047 <= w151 and not w45046;
w45048 <= not w44995 and w45047;
w45049 <= not w45042 and not w45048;
w45050 <= not b(43) and not w45049;
w45051 <= not w44398 and not w44996;
w45052 <= not w44408 and w44958;
w45053 <= not w44954 and w45052;
w45054 <= not w44955 and not w44958;
w45055 <= not w45053 and not w45054;
w45056 <= w151 and not w45055;
w45057 <= not w44995 and w45056;
w45058 <= not w45051 and not w45057;
w45059 <= not b(42) and not w45058;
w45060 <= not w44407 and not w44996;
w45061 <= not w44417 and w44953;
w45062 <= not w44949 and w45061;
w45063 <= not w44950 and not w44953;
w45064 <= not w45062 and not w45063;
w45065 <= w151 and not w45064;
w45066 <= not w44995 and w45065;
w45067 <= not w45060 and not w45066;
w45068 <= not b(41) and not w45067;
w45069 <= not w44416 and not w44996;
w45070 <= not w44426 and w44948;
w45071 <= not w44944 and w45070;
w45072 <= not w44945 and not w44948;
w45073 <= not w45071 and not w45072;
w45074 <= w151 and not w45073;
w45075 <= not w44995 and w45074;
w45076 <= not w45069 and not w45075;
w45077 <= not b(40) and not w45076;
w45078 <= not w44425 and not w44996;
w45079 <= not w44435 and w44943;
w45080 <= not w44939 and w45079;
w45081 <= not w44940 and not w44943;
w45082 <= not w45080 and not w45081;
w45083 <= w151 and not w45082;
w45084 <= not w44995 and w45083;
w45085 <= not w45078 and not w45084;
w45086 <= not b(39) and not w45085;
w45087 <= not w44434 and not w44996;
w45088 <= not w44444 and w44938;
w45089 <= not w44934 and w45088;
w45090 <= not w44935 and not w44938;
w45091 <= not w45089 and not w45090;
w45092 <= w151 and not w45091;
w45093 <= not w44995 and w45092;
w45094 <= not w45087 and not w45093;
w45095 <= not b(38) and not w45094;
w45096 <= not w44443 and not w44996;
w45097 <= not w44453 and w44933;
w45098 <= not w44929 and w45097;
w45099 <= not w44930 and not w44933;
w45100 <= not w45098 and not w45099;
w45101 <= w151 and not w45100;
w45102 <= not w44995 and w45101;
w45103 <= not w45096 and not w45102;
w45104 <= not b(37) and not w45103;
w45105 <= not w44452 and not w44996;
w45106 <= not w44462 and w44928;
w45107 <= not w44924 and w45106;
w45108 <= not w44925 and not w44928;
w45109 <= not w45107 and not w45108;
w45110 <= w151 and not w45109;
w45111 <= not w44995 and w45110;
w45112 <= not w45105 and not w45111;
w45113 <= not b(36) and not w45112;
w45114 <= not w44461 and not w44996;
w45115 <= not w44471 and w44923;
w45116 <= not w44919 and w45115;
w45117 <= not w44920 and not w44923;
w45118 <= not w45116 and not w45117;
w45119 <= w151 and not w45118;
w45120 <= not w44995 and w45119;
w45121 <= not w45114 and not w45120;
w45122 <= not b(35) and not w45121;
w45123 <= not w44470 and not w44996;
w45124 <= not w44480 and w44918;
w45125 <= not w44914 and w45124;
w45126 <= not w44915 and not w44918;
w45127 <= not w45125 and not w45126;
w45128 <= w151 and not w45127;
w45129 <= not w44995 and w45128;
w45130 <= not w45123 and not w45129;
w45131 <= not b(34) and not w45130;
w45132 <= not w44479 and not w44996;
w45133 <= not w44489 and w44913;
w45134 <= not w44909 and w45133;
w45135 <= not w44910 and not w44913;
w45136 <= not w45134 and not w45135;
w45137 <= w151 and not w45136;
w45138 <= not w44995 and w45137;
w45139 <= not w45132 and not w45138;
w45140 <= not b(33) and not w45139;
w45141 <= not w44488 and not w44996;
w45142 <= not w44498 and w44908;
w45143 <= not w44904 and w45142;
w45144 <= not w44905 and not w44908;
w45145 <= not w45143 and not w45144;
w45146 <= w151 and not w45145;
w45147 <= not w44995 and w45146;
w45148 <= not w45141 and not w45147;
w45149 <= not b(32) and not w45148;
w45150 <= not w44497 and not w44996;
w45151 <= not w44507 and w44903;
w45152 <= not w44899 and w45151;
w45153 <= not w44900 and not w44903;
w45154 <= not w45152 and not w45153;
w45155 <= w151 and not w45154;
w45156 <= not w44995 and w45155;
w45157 <= not w45150 and not w45156;
w45158 <= not b(31) and not w45157;
w45159 <= not w44506 and not w44996;
w45160 <= not w44516 and w44898;
w45161 <= not w44894 and w45160;
w45162 <= not w44895 and not w44898;
w45163 <= not w45161 and not w45162;
w45164 <= w151 and not w45163;
w45165 <= not w44995 and w45164;
w45166 <= not w45159 and not w45165;
w45167 <= not b(30) and not w45166;
w45168 <= not w44515 and not w44996;
w45169 <= not w44525 and w44893;
w45170 <= not w44889 and w45169;
w45171 <= not w44890 and not w44893;
w45172 <= not w45170 and not w45171;
w45173 <= w151 and not w45172;
w45174 <= not w44995 and w45173;
w45175 <= not w45168 and not w45174;
w45176 <= not b(29) and not w45175;
w45177 <= not w44524 and not w44996;
w45178 <= not w44534 and w44888;
w45179 <= not w44884 and w45178;
w45180 <= not w44885 and not w44888;
w45181 <= not w45179 and not w45180;
w45182 <= w151 and not w45181;
w45183 <= not w44995 and w45182;
w45184 <= not w45177 and not w45183;
w45185 <= not b(28) and not w45184;
w45186 <= not w44533 and not w44996;
w45187 <= not w44543 and w44883;
w45188 <= not w44879 and w45187;
w45189 <= not w44880 and not w44883;
w45190 <= not w45188 and not w45189;
w45191 <= w151 and not w45190;
w45192 <= not w44995 and w45191;
w45193 <= not w45186 and not w45192;
w45194 <= not b(27) and not w45193;
w45195 <= not w44542 and not w44996;
w45196 <= not w44552 and w44878;
w45197 <= not w44874 and w45196;
w45198 <= not w44875 and not w44878;
w45199 <= not w45197 and not w45198;
w45200 <= w151 and not w45199;
w45201 <= not w44995 and w45200;
w45202 <= not w45195 and not w45201;
w45203 <= not b(26) and not w45202;
w45204 <= not w44551 and not w44996;
w45205 <= not w44561 and w44873;
w45206 <= not w44869 and w45205;
w45207 <= not w44870 and not w44873;
w45208 <= not w45206 and not w45207;
w45209 <= w151 and not w45208;
w45210 <= not w44995 and w45209;
w45211 <= not w45204 and not w45210;
w45212 <= not b(25) and not w45211;
w45213 <= not w44560 and not w44996;
w45214 <= not w44570 and w44868;
w45215 <= not w44864 and w45214;
w45216 <= not w44865 and not w44868;
w45217 <= not w45215 and not w45216;
w45218 <= w151 and not w45217;
w45219 <= not w44995 and w45218;
w45220 <= not w45213 and not w45219;
w45221 <= not b(24) and not w45220;
w45222 <= not w44569 and not w44996;
w45223 <= not w44579 and w44863;
w45224 <= not w44859 and w45223;
w45225 <= not w44860 and not w44863;
w45226 <= not w45224 and not w45225;
w45227 <= w151 and not w45226;
w45228 <= not w44995 and w45227;
w45229 <= not w45222 and not w45228;
w45230 <= not b(23) and not w45229;
w45231 <= not w44578 and not w44996;
w45232 <= not w44588 and w44858;
w45233 <= not w44854 and w45232;
w45234 <= not w44855 and not w44858;
w45235 <= not w45233 and not w45234;
w45236 <= w151 and not w45235;
w45237 <= not w44995 and w45236;
w45238 <= not w45231 and not w45237;
w45239 <= not b(22) and not w45238;
w45240 <= not w44587 and not w44996;
w45241 <= not w44597 and w44853;
w45242 <= not w44849 and w45241;
w45243 <= not w44850 and not w44853;
w45244 <= not w45242 and not w45243;
w45245 <= w151 and not w45244;
w45246 <= not w44995 and w45245;
w45247 <= not w45240 and not w45246;
w45248 <= not b(21) and not w45247;
w45249 <= not w44596 and not w44996;
w45250 <= not w44606 and w44848;
w45251 <= not w44844 and w45250;
w45252 <= not w44845 and not w44848;
w45253 <= not w45251 and not w45252;
w45254 <= w151 and not w45253;
w45255 <= not w44995 and w45254;
w45256 <= not w45249 and not w45255;
w45257 <= not b(20) and not w45256;
w45258 <= not w44605 and not w44996;
w45259 <= not w44615 and w44843;
w45260 <= not w44839 and w45259;
w45261 <= not w44840 and not w44843;
w45262 <= not w45260 and not w45261;
w45263 <= w151 and not w45262;
w45264 <= not w44995 and w45263;
w45265 <= not w45258 and not w45264;
w45266 <= not b(19) and not w45265;
w45267 <= not w44614 and not w44996;
w45268 <= not w44624 and w44838;
w45269 <= not w44834 and w45268;
w45270 <= not w44835 and not w44838;
w45271 <= not w45269 and not w45270;
w45272 <= w151 and not w45271;
w45273 <= not w44995 and w45272;
w45274 <= not w45267 and not w45273;
w45275 <= not b(18) and not w45274;
w45276 <= not w44623 and not w44996;
w45277 <= not w44633 and w44833;
w45278 <= not w44829 and w45277;
w45279 <= not w44830 and not w44833;
w45280 <= not w45278 and not w45279;
w45281 <= w151 and not w45280;
w45282 <= not w44995 and w45281;
w45283 <= not w45276 and not w45282;
w45284 <= not b(17) and not w45283;
w45285 <= not w44632 and not w44996;
w45286 <= not w44642 and w44828;
w45287 <= not w44824 and w45286;
w45288 <= not w44825 and not w44828;
w45289 <= not w45287 and not w45288;
w45290 <= w151 and not w45289;
w45291 <= not w44995 and w45290;
w45292 <= not w45285 and not w45291;
w45293 <= not b(16) and not w45292;
w45294 <= not w44641 and not w44996;
w45295 <= not w44651 and w44823;
w45296 <= not w44819 and w45295;
w45297 <= not w44820 and not w44823;
w45298 <= not w45296 and not w45297;
w45299 <= w151 and not w45298;
w45300 <= not w44995 and w45299;
w45301 <= not w45294 and not w45300;
w45302 <= not b(15) and not w45301;
w45303 <= not w44650 and not w44996;
w45304 <= not w44660 and w44818;
w45305 <= not w44814 and w45304;
w45306 <= not w44815 and not w44818;
w45307 <= not w45305 and not w45306;
w45308 <= w151 and not w45307;
w45309 <= not w44995 and w45308;
w45310 <= not w45303 and not w45309;
w45311 <= not b(14) and not w45310;
w45312 <= not w44659 and not w44996;
w45313 <= not w44669 and w44813;
w45314 <= not w44809 and w45313;
w45315 <= not w44810 and not w44813;
w45316 <= not w45314 and not w45315;
w45317 <= w151 and not w45316;
w45318 <= not w44995 and w45317;
w45319 <= not w45312 and not w45318;
w45320 <= not b(13) and not w45319;
w45321 <= not w44668 and not w44996;
w45322 <= not w44678 and w44808;
w45323 <= not w44804 and w45322;
w45324 <= not w44805 and not w44808;
w45325 <= not w45323 and not w45324;
w45326 <= w151 and not w45325;
w45327 <= not w44995 and w45326;
w45328 <= not w45321 and not w45327;
w45329 <= not b(12) and not w45328;
w45330 <= not w44677 and not w44996;
w45331 <= not w44687 and w44803;
w45332 <= not w44799 and w45331;
w45333 <= not w44800 and not w44803;
w45334 <= not w45332 and not w45333;
w45335 <= w151 and not w45334;
w45336 <= not w44995 and w45335;
w45337 <= not w45330 and not w45336;
w45338 <= not b(11) and not w45337;
w45339 <= not w44686 and not w44996;
w45340 <= not w44696 and w44798;
w45341 <= not w44794 and w45340;
w45342 <= not w44795 and not w44798;
w45343 <= not w45341 and not w45342;
w45344 <= w151 and not w45343;
w45345 <= not w44995 and w45344;
w45346 <= not w45339 and not w45345;
w45347 <= not b(10) and not w45346;
w45348 <= not w44695 and not w44996;
w45349 <= not w44705 and w44793;
w45350 <= not w44789 and w45349;
w45351 <= not w44790 and not w44793;
w45352 <= not w45350 and not w45351;
w45353 <= w151 and not w45352;
w45354 <= not w44995 and w45353;
w45355 <= not w45348 and not w45354;
w45356 <= not b(9) and not w45355;
w45357 <= not w44704 and not w44996;
w45358 <= not w44714 and w44788;
w45359 <= not w44784 and w45358;
w45360 <= not w44785 and not w44788;
w45361 <= not w45359 and not w45360;
w45362 <= w151 and not w45361;
w45363 <= not w44995 and w45362;
w45364 <= not w45357 and not w45363;
w45365 <= not b(8) and not w45364;
w45366 <= not w44713 and not w44996;
w45367 <= not w44723 and w44783;
w45368 <= not w44779 and w45367;
w45369 <= not w44780 and not w44783;
w45370 <= not w45368 and not w45369;
w45371 <= w151 and not w45370;
w45372 <= not w44995 and w45371;
w45373 <= not w45366 and not w45372;
w45374 <= not b(7) and not w45373;
w45375 <= not w44722 and not w44996;
w45376 <= not w44732 and w44778;
w45377 <= not w44774 and w45376;
w45378 <= not w44775 and not w44778;
w45379 <= not w45377 and not w45378;
w45380 <= w151 and not w45379;
w45381 <= not w44995 and w45380;
w45382 <= not w45375 and not w45381;
w45383 <= not b(6) and not w45382;
w45384 <= not w44731 and not w44996;
w45385 <= not w44741 and w44773;
w45386 <= not w44769 and w45385;
w45387 <= not w44770 and not w44773;
w45388 <= not w45386 and not w45387;
w45389 <= w151 and not w45388;
w45390 <= not w44995 and w45389;
w45391 <= not w45384 and not w45390;
w45392 <= not b(5) and not w45391;
w45393 <= not w44740 and not w44996;
w45394 <= not w44749 and w44768;
w45395 <= not w44764 and w45394;
w45396 <= not w44765 and not w44768;
w45397 <= not w45395 and not w45396;
w45398 <= w151 and not w45397;
w45399 <= not w44995 and w45398;
w45400 <= not w45393 and not w45399;
w45401 <= not b(4) and not w45400;
w45402 <= not w44748 and not w44996;
w45403 <= not w44759 and w44763;
w45404 <= not w44758 and w45403;
w45405 <= not w44760 and not w44763;
w45406 <= not w45404 and not w45405;
w45407 <= w151 and not w45406;
w45408 <= not w44995 and w45407;
w45409 <= not w45402 and not w45408;
w45410 <= not b(3) and not w45409;
w45411 <= not w44753 and not w44996;
w45412 <= w16699 and not w44756;
w45413 <= not w44754 and w45412;
w45414 <= w151 and not w45413;
w45415 <= not w44758 and w45414;
w45416 <= not w44995 and w45415;
w45417 <= not w45411 and not w45416;
w45418 <= not b(2) and not w45417;
w45419 <= w17364 and not w44995;
w45420 <= a(15) and not w45419;
w45421 <= w17368 and not w44995;
w45422 <= not w45420 and not w45421;
w45423 <= b(1) and not w45422;
w45424 <= not b(1) and not w45421;
w45425 <= not w45420 and w45424;
w45426 <= not w45423 and not w45425;
w45427 <= not w17375 and not w45426;
w45428 <= not b(1) and not w45422;
w45429 <= not w45427 and not w45428;
w45430 <= b(2) and not w45416;
w45431 <= not w45411 and w45430;
w45432 <= not w45418 and not w45431;
w45433 <= not w45429 and w45432;
w45434 <= not w45418 and not w45433;
w45435 <= b(3) and not w45408;
w45436 <= not w45402 and w45435;
w45437 <= not w45410 and not w45436;
w45438 <= not w45434 and w45437;
w45439 <= not w45410 and not w45438;
w45440 <= b(4) and not w45399;
w45441 <= not w45393 and w45440;
w45442 <= not w45401 and not w45441;
w45443 <= not w45439 and w45442;
w45444 <= not w45401 and not w45443;
w45445 <= b(5) and not w45390;
w45446 <= not w45384 and w45445;
w45447 <= not w45392 and not w45446;
w45448 <= not w45444 and w45447;
w45449 <= not w45392 and not w45448;
w45450 <= b(6) and not w45381;
w45451 <= not w45375 and w45450;
w45452 <= not w45383 and not w45451;
w45453 <= not w45449 and w45452;
w45454 <= not w45383 and not w45453;
w45455 <= b(7) and not w45372;
w45456 <= not w45366 and w45455;
w45457 <= not w45374 and not w45456;
w45458 <= not w45454 and w45457;
w45459 <= not w45374 and not w45458;
w45460 <= b(8) and not w45363;
w45461 <= not w45357 and w45460;
w45462 <= not w45365 and not w45461;
w45463 <= not w45459 and w45462;
w45464 <= not w45365 and not w45463;
w45465 <= b(9) and not w45354;
w45466 <= not w45348 and w45465;
w45467 <= not w45356 and not w45466;
w45468 <= not w45464 and w45467;
w45469 <= not w45356 and not w45468;
w45470 <= b(10) and not w45345;
w45471 <= not w45339 and w45470;
w45472 <= not w45347 and not w45471;
w45473 <= not w45469 and w45472;
w45474 <= not w45347 and not w45473;
w45475 <= b(11) and not w45336;
w45476 <= not w45330 and w45475;
w45477 <= not w45338 and not w45476;
w45478 <= not w45474 and w45477;
w45479 <= not w45338 and not w45478;
w45480 <= b(12) and not w45327;
w45481 <= not w45321 and w45480;
w45482 <= not w45329 and not w45481;
w45483 <= not w45479 and w45482;
w45484 <= not w45329 and not w45483;
w45485 <= b(13) and not w45318;
w45486 <= not w45312 and w45485;
w45487 <= not w45320 and not w45486;
w45488 <= not w45484 and w45487;
w45489 <= not w45320 and not w45488;
w45490 <= b(14) and not w45309;
w45491 <= not w45303 and w45490;
w45492 <= not w45311 and not w45491;
w45493 <= not w45489 and w45492;
w45494 <= not w45311 and not w45493;
w45495 <= b(15) and not w45300;
w45496 <= not w45294 and w45495;
w45497 <= not w45302 and not w45496;
w45498 <= not w45494 and w45497;
w45499 <= not w45302 and not w45498;
w45500 <= b(16) and not w45291;
w45501 <= not w45285 and w45500;
w45502 <= not w45293 and not w45501;
w45503 <= not w45499 and w45502;
w45504 <= not w45293 and not w45503;
w45505 <= b(17) and not w45282;
w45506 <= not w45276 and w45505;
w45507 <= not w45284 and not w45506;
w45508 <= not w45504 and w45507;
w45509 <= not w45284 and not w45508;
w45510 <= b(18) and not w45273;
w45511 <= not w45267 and w45510;
w45512 <= not w45275 and not w45511;
w45513 <= not w45509 and w45512;
w45514 <= not w45275 and not w45513;
w45515 <= b(19) and not w45264;
w45516 <= not w45258 and w45515;
w45517 <= not w45266 and not w45516;
w45518 <= not w45514 and w45517;
w45519 <= not w45266 and not w45518;
w45520 <= b(20) and not w45255;
w45521 <= not w45249 and w45520;
w45522 <= not w45257 and not w45521;
w45523 <= not w45519 and w45522;
w45524 <= not w45257 and not w45523;
w45525 <= b(21) and not w45246;
w45526 <= not w45240 and w45525;
w45527 <= not w45248 and not w45526;
w45528 <= not w45524 and w45527;
w45529 <= not w45248 and not w45528;
w45530 <= b(22) and not w45237;
w45531 <= not w45231 and w45530;
w45532 <= not w45239 and not w45531;
w45533 <= not w45529 and w45532;
w45534 <= not w45239 and not w45533;
w45535 <= b(23) and not w45228;
w45536 <= not w45222 and w45535;
w45537 <= not w45230 and not w45536;
w45538 <= not w45534 and w45537;
w45539 <= not w45230 and not w45538;
w45540 <= b(24) and not w45219;
w45541 <= not w45213 and w45540;
w45542 <= not w45221 and not w45541;
w45543 <= not w45539 and w45542;
w45544 <= not w45221 and not w45543;
w45545 <= b(25) and not w45210;
w45546 <= not w45204 and w45545;
w45547 <= not w45212 and not w45546;
w45548 <= not w45544 and w45547;
w45549 <= not w45212 and not w45548;
w45550 <= b(26) and not w45201;
w45551 <= not w45195 and w45550;
w45552 <= not w45203 and not w45551;
w45553 <= not w45549 and w45552;
w45554 <= not w45203 and not w45553;
w45555 <= b(27) and not w45192;
w45556 <= not w45186 and w45555;
w45557 <= not w45194 and not w45556;
w45558 <= not w45554 and w45557;
w45559 <= not w45194 and not w45558;
w45560 <= b(28) and not w45183;
w45561 <= not w45177 and w45560;
w45562 <= not w45185 and not w45561;
w45563 <= not w45559 and w45562;
w45564 <= not w45185 and not w45563;
w45565 <= b(29) and not w45174;
w45566 <= not w45168 and w45565;
w45567 <= not w45176 and not w45566;
w45568 <= not w45564 and w45567;
w45569 <= not w45176 and not w45568;
w45570 <= b(30) and not w45165;
w45571 <= not w45159 and w45570;
w45572 <= not w45167 and not w45571;
w45573 <= not w45569 and w45572;
w45574 <= not w45167 and not w45573;
w45575 <= b(31) and not w45156;
w45576 <= not w45150 and w45575;
w45577 <= not w45158 and not w45576;
w45578 <= not w45574 and w45577;
w45579 <= not w45158 and not w45578;
w45580 <= b(32) and not w45147;
w45581 <= not w45141 and w45580;
w45582 <= not w45149 and not w45581;
w45583 <= not w45579 and w45582;
w45584 <= not w45149 and not w45583;
w45585 <= b(33) and not w45138;
w45586 <= not w45132 and w45585;
w45587 <= not w45140 and not w45586;
w45588 <= not w45584 and w45587;
w45589 <= not w45140 and not w45588;
w45590 <= b(34) and not w45129;
w45591 <= not w45123 and w45590;
w45592 <= not w45131 and not w45591;
w45593 <= not w45589 and w45592;
w45594 <= not w45131 and not w45593;
w45595 <= b(35) and not w45120;
w45596 <= not w45114 and w45595;
w45597 <= not w45122 and not w45596;
w45598 <= not w45594 and w45597;
w45599 <= not w45122 and not w45598;
w45600 <= b(36) and not w45111;
w45601 <= not w45105 and w45600;
w45602 <= not w45113 and not w45601;
w45603 <= not w45599 and w45602;
w45604 <= not w45113 and not w45603;
w45605 <= b(37) and not w45102;
w45606 <= not w45096 and w45605;
w45607 <= not w45104 and not w45606;
w45608 <= not w45604 and w45607;
w45609 <= not w45104 and not w45608;
w45610 <= b(38) and not w45093;
w45611 <= not w45087 and w45610;
w45612 <= not w45095 and not w45611;
w45613 <= not w45609 and w45612;
w45614 <= not w45095 and not w45613;
w45615 <= b(39) and not w45084;
w45616 <= not w45078 and w45615;
w45617 <= not w45086 and not w45616;
w45618 <= not w45614 and w45617;
w45619 <= not w45086 and not w45618;
w45620 <= b(40) and not w45075;
w45621 <= not w45069 and w45620;
w45622 <= not w45077 and not w45621;
w45623 <= not w45619 and w45622;
w45624 <= not w45077 and not w45623;
w45625 <= b(41) and not w45066;
w45626 <= not w45060 and w45625;
w45627 <= not w45068 and not w45626;
w45628 <= not w45624 and w45627;
w45629 <= not w45068 and not w45628;
w45630 <= b(42) and not w45057;
w45631 <= not w45051 and w45630;
w45632 <= not w45059 and not w45631;
w45633 <= not w45629 and w45632;
w45634 <= not w45059 and not w45633;
w45635 <= b(43) and not w45048;
w45636 <= not w45042 and w45635;
w45637 <= not w45050 and not w45636;
w45638 <= not w45634 and w45637;
w45639 <= not w45050 and not w45638;
w45640 <= b(44) and not w45039;
w45641 <= not w45033 and w45640;
w45642 <= not w45041 and not w45641;
w45643 <= not w45639 and w45642;
w45644 <= not w45041 and not w45643;
w45645 <= b(45) and not w45030;
w45646 <= not w45024 and w45645;
w45647 <= not w45032 and not w45646;
w45648 <= not w45644 and w45647;
w45649 <= not w45032 and not w45648;
w45650 <= b(46) and not w45021;
w45651 <= not w45015 and w45650;
w45652 <= not w45023 and not w45651;
w45653 <= not w45649 and w45652;
w45654 <= not w45023 and not w45653;
w45655 <= b(47) and not w45012;
w45656 <= not w45006 and w45655;
w45657 <= not w45014 and not w45656;
w45658 <= not w45654 and w45657;
w45659 <= not w45014 and not w45658;
w45660 <= b(48) and not w45003;
w45661 <= not w44997 and w45660;
w45662 <= not w45005 and not w45661;
w45663 <= not w45659 and w45662;
w45664 <= not w45005 and not w45663;
w45665 <= not w44343 and not w44996;
w45666 <= not w44345 and w44993;
w45667 <= not w44989 and w45666;
w45668 <= not w44990 and not w44993;
w45669 <= not w45667 and not w45668;
w45670 <= w44996 and not w45669;
w45671 <= not w45665 and not w45670;
w45672 <= not b(49) and not w45671;
w45673 <= b(49) and not w45665;
w45674 <= not w45670 and w45673;
w45675 <= w17625 and not w45674;
w45676 <= not w45672 and w45675;
w45677 <= not w45664 and w45676;
w45678 <= w151 and not w45671;
w45679 <= not w45677 and not w45678;
w45680 <= not w45014 and w45662;
w45681 <= not w45658 and w45680;
w45682 <= not w45659 and not w45662;
w45683 <= not w45681 and not w45682;
w45684 <= not w45679 and not w45683;
w45685 <= not w45004 and not w45678;
w45686 <= not w45677 and w45685;
w45687 <= not w45684 and not w45686;
w45688 <= not b(49) and not w45687;
w45689 <= not w45023 and w45657;
w45690 <= not w45653 and w45689;
w45691 <= not w45654 and not w45657;
w45692 <= not w45690 and not w45691;
w45693 <= not w45679 and not w45692;
w45694 <= not w45013 and not w45678;
w45695 <= not w45677 and w45694;
w45696 <= not w45693 and not w45695;
w45697 <= not b(48) and not w45696;
w45698 <= not w45032 and w45652;
w45699 <= not w45648 and w45698;
w45700 <= not w45649 and not w45652;
w45701 <= not w45699 and not w45700;
w45702 <= not w45679 and not w45701;
w45703 <= not w45022 and not w45678;
w45704 <= not w45677 and w45703;
w45705 <= not w45702 and not w45704;
w45706 <= not b(47) and not w45705;
w45707 <= not w45041 and w45647;
w45708 <= not w45643 and w45707;
w45709 <= not w45644 and not w45647;
w45710 <= not w45708 and not w45709;
w45711 <= not w45679 and not w45710;
w45712 <= not w45031 and not w45678;
w45713 <= not w45677 and w45712;
w45714 <= not w45711 and not w45713;
w45715 <= not b(46) and not w45714;
w45716 <= not w45050 and w45642;
w45717 <= not w45638 and w45716;
w45718 <= not w45639 and not w45642;
w45719 <= not w45717 and not w45718;
w45720 <= not w45679 and not w45719;
w45721 <= not w45040 and not w45678;
w45722 <= not w45677 and w45721;
w45723 <= not w45720 and not w45722;
w45724 <= not b(45) and not w45723;
w45725 <= not w45059 and w45637;
w45726 <= not w45633 and w45725;
w45727 <= not w45634 and not w45637;
w45728 <= not w45726 and not w45727;
w45729 <= not w45679 and not w45728;
w45730 <= not w45049 and not w45678;
w45731 <= not w45677 and w45730;
w45732 <= not w45729 and not w45731;
w45733 <= not b(44) and not w45732;
w45734 <= not w45068 and w45632;
w45735 <= not w45628 and w45734;
w45736 <= not w45629 and not w45632;
w45737 <= not w45735 and not w45736;
w45738 <= not w45679 and not w45737;
w45739 <= not w45058 and not w45678;
w45740 <= not w45677 and w45739;
w45741 <= not w45738 and not w45740;
w45742 <= not b(43) and not w45741;
w45743 <= not w45077 and w45627;
w45744 <= not w45623 and w45743;
w45745 <= not w45624 and not w45627;
w45746 <= not w45744 and not w45745;
w45747 <= not w45679 and not w45746;
w45748 <= not w45067 and not w45678;
w45749 <= not w45677 and w45748;
w45750 <= not w45747 and not w45749;
w45751 <= not b(42) and not w45750;
w45752 <= not w45086 and w45622;
w45753 <= not w45618 and w45752;
w45754 <= not w45619 and not w45622;
w45755 <= not w45753 and not w45754;
w45756 <= not w45679 and not w45755;
w45757 <= not w45076 and not w45678;
w45758 <= not w45677 and w45757;
w45759 <= not w45756 and not w45758;
w45760 <= not b(41) and not w45759;
w45761 <= not w45095 and w45617;
w45762 <= not w45613 and w45761;
w45763 <= not w45614 and not w45617;
w45764 <= not w45762 and not w45763;
w45765 <= not w45679 and not w45764;
w45766 <= not w45085 and not w45678;
w45767 <= not w45677 and w45766;
w45768 <= not w45765 and not w45767;
w45769 <= not b(40) and not w45768;
w45770 <= not w45104 and w45612;
w45771 <= not w45608 and w45770;
w45772 <= not w45609 and not w45612;
w45773 <= not w45771 and not w45772;
w45774 <= not w45679 and not w45773;
w45775 <= not w45094 and not w45678;
w45776 <= not w45677 and w45775;
w45777 <= not w45774 and not w45776;
w45778 <= not b(39) and not w45777;
w45779 <= not w45113 and w45607;
w45780 <= not w45603 and w45779;
w45781 <= not w45604 and not w45607;
w45782 <= not w45780 and not w45781;
w45783 <= not w45679 and not w45782;
w45784 <= not w45103 and not w45678;
w45785 <= not w45677 and w45784;
w45786 <= not w45783 and not w45785;
w45787 <= not b(38) and not w45786;
w45788 <= not w45122 and w45602;
w45789 <= not w45598 and w45788;
w45790 <= not w45599 and not w45602;
w45791 <= not w45789 and not w45790;
w45792 <= not w45679 and not w45791;
w45793 <= not w45112 and not w45678;
w45794 <= not w45677 and w45793;
w45795 <= not w45792 and not w45794;
w45796 <= not b(37) and not w45795;
w45797 <= not w45131 and w45597;
w45798 <= not w45593 and w45797;
w45799 <= not w45594 and not w45597;
w45800 <= not w45798 and not w45799;
w45801 <= not w45679 and not w45800;
w45802 <= not w45121 and not w45678;
w45803 <= not w45677 and w45802;
w45804 <= not w45801 and not w45803;
w45805 <= not b(36) and not w45804;
w45806 <= not w45140 and w45592;
w45807 <= not w45588 and w45806;
w45808 <= not w45589 and not w45592;
w45809 <= not w45807 and not w45808;
w45810 <= not w45679 and not w45809;
w45811 <= not w45130 and not w45678;
w45812 <= not w45677 and w45811;
w45813 <= not w45810 and not w45812;
w45814 <= not b(35) and not w45813;
w45815 <= not w45149 and w45587;
w45816 <= not w45583 and w45815;
w45817 <= not w45584 and not w45587;
w45818 <= not w45816 and not w45817;
w45819 <= not w45679 and not w45818;
w45820 <= not w45139 and not w45678;
w45821 <= not w45677 and w45820;
w45822 <= not w45819 and not w45821;
w45823 <= not b(34) and not w45822;
w45824 <= not w45158 and w45582;
w45825 <= not w45578 and w45824;
w45826 <= not w45579 and not w45582;
w45827 <= not w45825 and not w45826;
w45828 <= not w45679 and not w45827;
w45829 <= not w45148 and not w45678;
w45830 <= not w45677 and w45829;
w45831 <= not w45828 and not w45830;
w45832 <= not b(33) and not w45831;
w45833 <= not w45167 and w45577;
w45834 <= not w45573 and w45833;
w45835 <= not w45574 and not w45577;
w45836 <= not w45834 and not w45835;
w45837 <= not w45679 and not w45836;
w45838 <= not w45157 and not w45678;
w45839 <= not w45677 and w45838;
w45840 <= not w45837 and not w45839;
w45841 <= not b(32) and not w45840;
w45842 <= not w45176 and w45572;
w45843 <= not w45568 and w45842;
w45844 <= not w45569 and not w45572;
w45845 <= not w45843 and not w45844;
w45846 <= not w45679 and not w45845;
w45847 <= not w45166 and not w45678;
w45848 <= not w45677 and w45847;
w45849 <= not w45846 and not w45848;
w45850 <= not b(31) and not w45849;
w45851 <= not w45185 and w45567;
w45852 <= not w45563 and w45851;
w45853 <= not w45564 and not w45567;
w45854 <= not w45852 and not w45853;
w45855 <= not w45679 and not w45854;
w45856 <= not w45175 and not w45678;
w45857 <= not w45677 and w45856;
w45858 <= not w45855 and not w45857;
w45859 <= not b(30) and not w45858;
w45860 <= not w45194 and w45562;
w45861 <= not w45558 and w45860;
w45862 <= not w45559 and not w45562;
w45863 <= not w45861 and not w45862;
w45864 <= not w45679 and not w45863;
w45865 <= not w45184 and not w45678;
w45866 <= not w45677 and w45865;
w45867 <= not w45864 and not w45866;
w45868 <= not b(29) and not w45867;
w45869 <= not w45203 and w45557;
w45870 <= not w45553 and w45869;
w45871 <= not w45554 and not w45557;
w45872 <= not w45870 and not w45871;
w45873 <= not w45679 and not w45872;
w45874 <= not w45193 and not w45678;
w45875 <= not w45677 and w45874;
w45876 <= not w45873 and not w45875;
w45877 <= not b(28) and not w45876;
w45878 <= not w45212 and w45552;
w45879 <= not w45548 and w45878;
w45880 <= not w45549 and not w45552;
w45881 <= not w45879 and not w45880;
w45882 <= not w45679 and not w45881;
w45883 <= not w45202 and not w45678;
w45884 <= not w45677 and w45883;
w45885 <= not w45882 and not w45884;
w45886 <= not b(27) and not w45885;
w45887 <= not w45221 and w45547;
w45888 <= not w45543 and w45887;
w45889 <= not w45544 and not w45547;
w45890 <= not w45888 and not w45889;
w45891 <= not w45679 and not w45890;
w45892 <= not w45211 and not w45678;
w45893 <= not w45677 and w45892;
w45894 <= not w45891 and not w45893;
w45895 <= not b(26) and not w45894;
w45896 <= not w45230 and w45542;
w45897 <= not w45538 and w45896;
w45898 <= not w45539 and not w45542;
w45899 <= not w45897 and not w45898;
w45900 <= not w45679 and not w45899;
w45901 <= not w45220 and not w45678;
w45902 <= not w45677 and w45901;
w45903 <= not w45900 and not w45902;
w45904 <= not b(25) and not w45903;
w45905 <= not w45239 and w45537;
w45906 <= not w45533 and w45905;
w45907 <= not w45534 and not w45537;
w45908 <= not w45906 and not w45907;
w45909 <= not w45679 and not w45908;
w45910 <= not w45229 and not w45678;
w45911 <= not w45677 and w45910;
w45912 <= not w45909 and not w45911;
w45913 <= not b(24) and not w45912;
w45914 <= not w45248 and w45532;
w45915 <= not w45528 and w45914;
w45916 <= not w45529 and not w45532;
w45917 <= not w45915 and not w45916;
w45918 <= not w45679 and not w45917;
w45919 <= not w45238 and not w45678;
w45920 <= not w45677 and w45919;
w45921 <= not w45918 and not w45920;
w45922 <= not b(23) and not w45921;
w45923 <= not w45257 and w45527;
w45924 <= not w45523 and w45923;
w45925 <= not w45524 and not w45527;
w45926 <= not w45924 and not w45925;
w45927 <= not w45679 and not w45926;
w45928 <= not w45247 and not w45678;
w45929 <= not w45677 and w45928;
w45930 <= not w45927 and not w45929;
w45931 <= not b(22) and not w45930;
w45932 <= not w45266 and w45522;
w45933 <= not w45518 and w45932;
w45934 <= not w45519 and not w45522;
w45935 <= not w45933 and not w45934;
w45936 <= not w45679 and not w45935;
w45937 <= not w45256 and not w45678;
w45938 <= not w45677 and w45937;
w45939 <= not w45936 and not w45938;
w45940 <= not b(21) and not w45939;
w45941 <= not w45275 and w45517;
w45942 <= not w45513 and w45941;
w45943 <= not w45514 and not w45517;
w45944 <= not w45942 and not w45943;
w45945 <= not w45679 and not w45944;
w45946 <= not w45265 and not w45678;
w45947 <= not w45677 and w45946;
w45948 <= not w45945 and not w45947;
w45949 <= not b(20) and not w45948;
w45950 <= not w45284 and w45512;
w45951 <= not w45508 and w45950;
w45952 <= not w45509 and not w45512;
w45953 <= not w45951 and not w45952;
w45954 <= not w45679 and not w45953;
w45955 <= not w45274 and not w45678;
w45956 <= not w45677 and w45955;
w45957 <= not w45954 and not w45956;
w45958 <= not b(19) and not w45957;
w45959 <= not w45293 and w45507;
w45960 <= not w45503 and w45959;
w45961 <= not w45504 and not w45507;
w45962 <= not w45960 and not w45961;
w45963 <= not w45679 and not w45962;
w45964 <= not w45283 and not w45678;
w45965 <= not w45677 and w45964;
w45966 <= not w45963 and not w45965;
w45967 <= not b(18) and not w45966;
w45968 <= not w45302 and w45502;
w45969 <= not w45498 and w45968;
w45970 <= not w45499 and not w45502;
w45971 <= not w45969 and not w45970;
w45972 <= not w45679 and not w45971;
w45973 <= not w45292 and not w45678;
w45974 <= not w45677 and w45973;
w45975 <= not w45972 and not w45974;
w45976 <= not b(17) and not w45975;
w45977 <= not w45311 and w45497;
w45978 <= not w45493 and w45977;
w45979 <= not w45494 and not w45497;
w45980 <= not w45978 and not w45979;
w45981 <= not w45679 and not w45980;
w45982 <= not w45301 and not w45678;
w45983 <= not w45677 and w45982;
w45984 <= not w45981 and not w45983;
w45985 <= not b(16) and not w45984;
w45986 <= not w45320 and w45492;
w45987 <= not w45488 and w45986;
w45988 <= not w45489 and not w45492;
w45989 <= not w45987 and not w45988;
w45990 <= not w45679 and not w45989;
w45991 <= not w45310 and not w45678;
w45992 <= not w45677 and w45991;
w45993 <= not w45990 and not w45992;
w45994 <= not b(15) and not w45993;
w45995 <= not w45329 and w45487;
w45996 <= not w45483 and w45995;
w45997 <= not w45484 and not w45487;
w45998 <= not w45996 and not w45997;
w45999 <= not w45679 and not w45998;
w46000 <= not w45319 and not w45678;
w46001 <= not w45677 and w46000;
w46002 <= not w45999 and not w46001;
w46003 <= not b(14) and not w46002;
w46004 <= not w45338 and w45482;
w46005 <= not w45478 and w46004;
w46006 <= not w45479 and not w45482;
w46007 <= not w46005 and not w46006;
w46008 <= not w45679 and not w46007;
w46009 <= not w45328 and not w45678;
w46010 <= not w45677 and w46009;
w46011 <= not w46008 and not w46010;
w46012 <= not b(13) and not w46011;
w46013 <= not w45347 and w45477;
w46014 <= not w45473 and w46013;
w46015 <= not w45474 and not w45477;
w46016 <= not w46014 and not w46015;
w46017 <= not w45679 and not w46016;
w46018 <= not w45337 and not w45678;
w46019 <= not w45677 and w46018;
w46020 <= not w46017 and not w46019;
w46021 <= not b(12) and not w46020;
w46022 <= not w45356 and w45472;
w46023 <= not w45468 and w46022;
w46024 <= not w45469 and not w45472;
w46025 <= not w46023 and not w46024;
w46026 <= not w45679 and not w46025;
w46027 <= not w45346 and not w45678;
w46028 <= not w45677 and w46027;
w46029 <= not w46026 and not w46028;
w46030 <= not b(11) and not w46029;
w46031 <= not w45365 and w45467;
w46032 <= not w45463 and w46031;
w46033 <= not w45464 and not w45467;
w46034 <= not w46032 and not w46033;
w46035 <= not w45679 and not w46034;
w46036 <= not w45355 and not w45678;
w46037 <= not w45677 and w46036;
w46038 <= not w46035 and not w46037;
w46039 <= not b(10) and not w46038;
w46040 <= not w45374 and w45462;
w46041 <= not w45458 and w46040;
w46042 <= not w45459 and not w45462;
w46043 <= not w46041 and not w46042;
w46044 <= not w45679 and not w46043;
w46045 <= not w45364 and not w45678;
w46046 <= not w45677 and w46045;
w46047 <= not w46044 and not w46046;
w46048 <= not b(9) and not w46047;
w46049 <= not w45383 and w45457;
w46050 <= not w45453 and w46049;
w46051 <= not w45454 and not w45457;
w46052 <= not w46050 and not w46051;
w46053 <= not w45679 and not w46052;
w46054 <= not w45373 and not w45678;
w46055 <= not w45677 and w46054;
w46056 <= not w46053 and not w46055;
w46057 <= not b(8) and not w46056;
w46058 <= not w45392 and w45452;
w46059 <= not w45448 and w46058;
w46060 <= not w45449 and not w45452;
w46061 <= not w46059 and not w46060;
w46062 <= not w45679 and not w46061;
w46063 <= not w45382 and not w45678;
w46064 <= not w45677 and w46063;
w46065 <= not w46062 and not w46064;
w46066 <= not b(7) and not w46065;
w46067 <= not w45401 and w45447;
w46068 <= not w45443 and w46067;
w46069 <= not w45444 and not w45447;
w46070 <= not w46068 and not w46069;
w46071 <= not w45679 and not w46070;
w46072 <= not w45391 and not w45678;
w46073 <= not w45677 and w46072;
w46074 <= not w46071 and not w46073;
w46075 <= not b(6) and not w46074;
w46076 <= not w45410 and w45442;
w46077 <= not w45438 and w46076;
w46078 <= not w45439 and not w45442;
w46079 <= not w46077 and not w46078;
w46080 <= not w45679 and not w46079;
w46081 <= not w45400 and not w45678;
w46082 <= not w45677 and w46081;
w46083 <= not w46080 and not w46082;
w46084 <= not b(5) and not w46083;
w46085 <= not w45418 and w45437;
w46086 <= not w45433 and w46085;
w46087 <= not w45434 and not w45437;
w46088 <= not w46086 and not w46087;
w46089 <= not w45679 and not w46088;
w46090 <= not w45409 and not w45678;
w46091 <= not w45677 and w46090;
w46092 <= not w46089 and not w46091;
w46093 <= not b(4) and not w46092;
w46094 <= not w45428 and w45432;
w46095 <= not w45427 and w46094;
w46096 <= not w45429 and not w45432;
w46097 <= not w46095 and not w46096;
w46098 <= not w45679 and not w46097;
w46099 <= not w45417 and not w45678;
w46100 <= not w45677 and w46099;
w46101 <= not w46098 and not w46100;
w46102 <= not b(3) and not w46101;
w46103 <= w17375 and not w45425;
w46104 <= not w45423 and w46103;
w46105 <= not w45427 and not w46104;
w46106 <= not w45679 and w46105;
w46107 <= not w45422 and not w45678;
w46108 <= not w45677 and w46107;
w46109 <= not w46106 and not w46108;
w46110 <= not b(2) and not w46109;
w46111 <= b(0) and not w45679;
w46112 <= a(14) and not w46111;
w46113 <= w17375 and not w45679;
w46114 <= not w46112 and not w46113;
w46115 <= b(1) and not w46114;
w46116 <= not b(1) and not w46113;
w46117 <= not w46112 and w46116;
w46118 <= not w46115 and not w46117;
w46119 <= not w18070 and not w46118;
w46120 <= not b(1) and not w46114;
w46121 <= not w46119 and not w46120;
w46122 <= b(2) and not w46108;
w46123 <= not w46106 and w46122;
w46124 <= not w46110 and not w46123;
w46125 <= not w46121 and w46124;
w46126 <= not w46110 and not w46125;
w46127 <= b(3) and not w46100;
w46128 <= not w46098 and w46127;
w46129 <= not w46102 and not w46128;
w46130 <= not w46126 and w46129;
w46131 <= not w46102 and not w46130;
w46132 <= b(4) and not w46091;
w46133 <= not w46089 and w46132;
w46134 <= not w46093 and not w46133;
w46135 <= not w46131 and w46134;
w46136 <= not w46093 and not w46135;
w46137 <= b(5) and not w46082;
w46138 <= not w46080 and w46137;
w46139 <= not w46084 and not w46138;
w46140 <= not w46136 and w46139;
w46141 <= not w46084 and not w46140;
w46142 <= b(6) and not w46073;
w46143 <= not w46071 and w46142;
w46144 <= not w46075 and not w46143;
w46145 <= not w46141 and w46144;
w46146 <= not w46075 and not w46145;
w46147 <= b(7) and not w46064;
w46148 <= not w46062 and w46147;
w46149 <= not w46066 and not w46148;
w46150 <= not w46146 and w46149;
w46151 <= not w46066 and not w46150;
w46152 <= b(8) and not w46055;
w46153 <= not w46053 and w46152;
w46154 <= not w46057 and not w46153;
w46155 <= not w46151 and w46154;
w46156 <= not w46057 and not w46155;
w46157 <= b(9) and not w46046;
w46158 <= not w46044 and w46157;
w46159 <= not w46048 and not w46158;
w46160 <= not w46156 and w46159;
w46161 <= not w46048 and not w46160;
w46162 <= b(10) and not w46037;
w46163 <= not w46035 and w46162;
w46164 <= not w46039 and not w46163;
w46165 <= not w46161 and w46164;
w46166 <= not w46039 and not w46165;
w46167 <= b(11) and not w46028;
w46168 <= not w46026 and w46167;
w46169 <= not w46030 and not w46168;
w46170 <= not w46166 and w46169;
w46171 <= not w46030 and not w46170;
w46172 <= b(12) and not w46019;
w46173 <= not w46017 and w46172;
w46174 <= not w46021 and not w46173;
w46175 <= not w46171 and w46174;
w46176 <= not w46021 and not w46175;
w46177 <= b(13) and not w46010;
w46178 <= not w46008 and w46177;
w46179 <= not w46012 and not w46178;
w46180 <= not w46176 and w46179;
w46181 <= not w46012 and not w46180;
w46182 <= b(14) and not w46001;
w46183 <= not w45999 and w46182;
w46184 <= not w46003 and not w46183;
w46185 <= not w46181 and w46184;
w46186 <= not w46003 and not w46185;
w46187 <= b(15) and not w45992;
w46188 <= not w45990 and w46187;
w46189 <= not w45994 and not w46188;
w46190 <= not w46186 and w46189;
w46191 <= not w45994 and not w46190;
w46192 <= b(16) and not w45983;
w46193 <= not w45981 and w46192;
w46194 <= not w45985 and not w46193;
w46195 <= not w46191 and w46194;
w46196 <= not w45985 and not w46195;
w46197 <= b(17) and not w45974;
w46198 <= not w45972 and w46197;
w46199 <= not w45976 and not w46198;
w46200 <= not w46196 and w46199;
w46201 <= not w45976 and not w46200;
w46202 <= b(18) and not w45965;
w46203 <= not w45963 and w46202;
w46204 <= not w45967 and not w46203;
w46205 <= not w46201 and w46204;
w46206 <= not w45967 and not w46205;
w46207 <= b(19) and not w45956;
w46208 <= not w45954 and w46207;
w46209 <= not w45958 and not w46208;
w46210 <= not w46206 and w46209;
w46211 <= not w45958 and not w46210;
w46212 <= b(20) and not w45947;
w46213 <= not w45945 and w46212;
w46214 <= not w45949 and not w46213;
w46215 <= not w46211 and w46214;
w46216 <= not w45949 and not w46215;
w46217 <= b(21) and not w45938;
w46218 <= not w45936 and w46217;
w46219 <= not w45940 and not w46218;
w46220 <= not w46216 and w46219;
w46221 <= not w45940 and not w46220;
w46222 <= b(22) and not w45929;
w46223 <= not w45927 and w46222;
w46224 <= not w45931 and not w46223;
w46225 <= not w46221 and w46224;
w46226 <= not w45931 and not w46225;
w46227 <= b(23) and not w45920;
w46228 <= not w45918 and w46227;
w46229 <= not w45922 and not w46228;
w46230 <= not w46226 and w46229;
w46231 <= not w45922 and not w46230;
w46232 <= b(24) and not w45911;
w46233 <= not w45909 and w46232;
w46234 <= not w45913 and not w46233;
w46235 <= not w46231 and w46234;
w46236 <= not w45913 and not w46235;
w46237 <= b(25) and not w45902;
w46238 <= not w45900 and w46237;
w46239 <= not w45904 and not w46238;
w46240 <= not w46236 and w46239;
w46241 <= not w45904 and not w46240;
w46242 <= b(26) and not w45893;
w46243 <= not w45891 and w46242;
w46244 <= not w45895 and not w46243;
w46245 <= not w46241 and w46244;
w46246 <= not w45895 and not w46245;
w46247 <= b(27) and not w45884;
w46248 <= not w45882 and w46247;
w46249 <= not w45886 and not w46248;
w46250 <= not w46246 and w46249;
w46251 <= not w45886 and not w46250;
w46252 <= b(28) and not w45875;
w46253 <= not w45873 and w46252;
w46254 <= not w45877 and not w46253;
w46255 <= not w46251 and w46254;
w46256 <= not w45877 and not w46255;
w46257 <= b(29) and not w45866;
w46258 <= not w45864 and w46257;
w46259 <= not w45868 and not w46258;
w46260 <= not w46256 and w46259;
w46261 <= not w45868 and not w46260;
w46262 <= b(30) and not w45857;
w46263 <= not w45855 and w46262;
w46264 <= not w45859 and not w46263;
w46265 <= not w46261 and w46264;
w46266 <= not w45859 and not w46265;
w46267 <= b(31) and not w45848;
w46268 <= not w45846 and w46267;
w46269 <= not w45850 and not w46268;
w46270 <= not w46266 and w46269;
w46271 <= not w45850 and not w46270;
w46272 <= b(32) and not w45839;
w46273 <= not w45837 and w46272;
w46274 <= not w45841 and not w46273;
w46275 <= not w46271 and w46274;
w46276 <= not w45841 and not w46275;
w46277 <= b(33) and not w45830;
w46278 <= not w45828 and w46277;
w46279 <= not w45832 and not w46278;
w46280 <= not w46276 and w46279;
w46281 <= not w45832 and not w46280;
w46282 <= b(34) and not w45821;
w46283 <= not w45819 and w46282;
w46284 <= not w45823 and not w46283;
w46285 <= not w46281 and w46284;
w46286 <= not w45823 and not w46285;
w46287 <= b(35) and not w45812;
w46288 <= not w45810 and w46287;
w46289 <= not w45814 and not w46288;
w46290 <= not w46286 and w46289;
w46291 <= not w45814 and not w46290;
w46292 <= b(36) and not w45803;
w46293 <= not w45801 and w46292;
w46294 <= not w45805 and not w46293;
w46295 <= not w46291 and w46294;
w46296 <= not w45805 and not w46295;
w46297 <= b(37) and not w45794;
w46298 <= not w45792 and w46297;
w46299 <= not w45796 and not w46298;
w46300 <= not w46296 and w46299;
w46301 <= not w45796 and not w46300;
w46302 <= b(38) and not w45785;
w46303 <= not w45783 and w46302;
w46304 <= not w45787 and not w46303;
w46305 <= not w46301 and w46304;
w46306 <= not w45787 and not w46305;
w46307 <= b(39) and not w45776;
w46308 <= not w45774 and w46307;
w46309 <= not w45778 and not w46308;
w46310 <= not w46306 and w46309;
w46311 <= not w45778 and not w46310;
w46312 <= b(40) and not w45767;
w46313 <= not w45765 and w46312;
w46314 <= not w45769 and not w46313;
w46315 <= not w46311 and w46314;
w46316 <= not w45769 and not w46315;
w46317 <= b(41) and not w45758;
w46318 <= not w45756 and w46317;
w46319 <= not w45760 and not w46318;
w46320 <= not w46316 and w46319;
w46321 <= not w45760 and not w46320;
w46322 <= b(42) and not w45749;
w46323 <= not w45747 and w46322;
w46324 <= not w45751 and not w46323;
w46325 <= not w46321 and w46324;
w46326 <= not w45751 and not w46325;
w46327 <= b(43) and not w45740;
w46328 <= not w45738 and w46327;
w46329 <= not w45742 and not w46328;
w46330 <= not w46326 and w46329;
w46331 <= not w45742 and not w46330;
w46332 <= b(44) and not w45731;
w46333 <= not w45729 and w46332;
w46334 <= not w45733 and not w46333;
w46335 <= not w46331 and w46334;
w46336 <= not w45733 and not w46335;
w46337 <= b(45) and not w45722;
w46338 <= not w45720 and w46337;
w46339 <= not w45724 and not w46338;
w46340 <= not w46336 and w46339;
w46341 <= not w45724 and not w46340;
w46342 <= b(46) and not w45713;
w46343 <= not w45711 and w46342;
w46344 <= not w45715 and not w46343;
w46345 <= not w46341 and w46344;
w46346 <= not w45715 and not w46345;
w46347 <= b(47) and not w45704;
w46348 <= not w45702 and w46347;
w46349 <= not w45706 and not w46348;
w46350 <= not w46346 and w46349;
w46351 <= not w45706 and not w46350;
w46352 <= b(48) and not w45695;
w46353 <= not w45693 and w46352;
w46354 <= not w45697 and not w46353;
w46355 <= not w46351 and w46354;
w46356 <= not w45697 and not w46355;
w46357 <= b(49) and not w45686;
w46358 <= not w45684 and w46357;
w46359 <= not w45688 and not w46358;
w46360 <= not w46356 and w46359;
w46361 <= not w45688 and not w46360;
w46362 <= not w45005 and not w45674;
w46363 <= not w45672 and w46362;
w46364 <= not w45663 and w46363;
w46365 <= not w45672 and not w45674;
w46366 <= not w45664 and not w46365;
w46367 <= not w46364 and not w46366;
w46368 <= not w45679 and not w46367;
w46369 <= not w45671 and not w45678;
w46370 <= not w45677 and w46369;
w46371 <= not w46368 and not w46370;
w46372 <= not b(50) and not w46371;
w46373 <= b(50) and not w46370;
w46374 <= not w46368 and w46373;
w46375 <= w18328 and not w46374;
w46376 <= not w46372 and w46375;
w46377 <= not w46361 and w46376;
w46378 <= w17625 and not w46371;
w46379 <= not w46377 and not w46378;
w46380 <= not w45697 and w46359;
w46381 <= not w46355 and w46380;
w46382 <= not w46356 and not w46359;
w46383 <= not w46381 and not w46382;
w46384 <= not w46379 and not w46383;
w46385 <= not w45687 and not w46378;
w46386 <= not w46377 and w46385;
w46387 <= not w46384 and not w46386;
w46388 <= not w45688 and not w46374;
w46389 <= not w46372 and w46388;
w46390 <= not w46360 and w46389;
w46391 <= not w46372 and not w46374;
w46392 <= not w46361 and not w46391;
w46393 <= not w46390 and not w46392;
w46394 <= not w46379 and not w46393;
w46395 <= not w46371 and not w46378;
w46396 <= not w46377 and w46395;
w46397 <= not w46394 and not w46396;
w46398 <= not b(51) and not w46397;
w46399 <= not b(50) and not w46387;
w46400 <= not w45706 and w46354;
w46401 <= not w46350 and w46400;
w46402 <= not w46351 and not w46354;
w46403 <= not w46401 and not w46402;
w46404 <= not w46379 and not w46403;
w46405 <= not w45696 and not w46378;
w46406 <= not w46377 and w46405;
w46407 <= not w46404 and not w46406;
w46408 <= not b(49) and not w46407;
w46409 <= not w45715 and w46349;
w46410 <= not w46345 and w46409;
w46411 <= not w46346 and not w46349;
w46412 <= not w46410 and not w46411;
w46413 <= not w46379 and not w46412;
w46414 <= not w45705 and not w46378;
w46415 <= not w46377 and w46414;
w46416 <= not w46413 and not w46415;
w46417 <= not b(48) and not w46416;
w46418 <= not w45724 and w46344;
w46419 <= not w46340 and w46418;
w46420 <= not w46341 and not w46344;
w46421 <= not w46419 and not w46420;
w46422 <= not w46379 and not w46421;
w46423 <= not w45714 and not w46378;
w46424 <= not w46377 and w46423;
w46425 <= not w46422 and not w46424;
w46426 <= not b(47) and not w46425;
w46427 <= not w45733 and w46339;
w46428 <= not w46335 and w46427;
w46429 <= not w46336 and not w46339;
w46430 <= not w46428 and not w46429;
w46431 <= not w46379 and not w46430;
w46432 <= not w45723 and not w46378;
w46433 <= not w46377 and w46432;
w46434 <= not w46431 and not w46433;
w46435 <= not b(46) and not w46434;
w46436 <= not w45742 and w46334;
w46437 <= not w46330 and w46436;
w46438 <= not w46331 and not w46334;
w46439 <= not w46437 and not w46438;
w46440 <= not w46379 and not w46439;
w46441 <= not w45732 and not w46378;
w46442 <= not w46377 and w46441;
w46443 <= not w46440 and not w46442;
w46444 <= not b(45) and not w46443;
w46445 <= not w45751 and w46329;
w46446 <= not w46325 and w46445;
w46447 <= not w46326 and not w46329;
w46448 <= not w46446 and not w46447;
w46449 <= not w46379 and not w46448;
w46450 <= not w45741 and not w46378;
w46451 <= not w46377 and w46450;
w46452 <= not w46449 and not w46451;
w46453 <= not b(44) and not w46452;
w46454 <= not w45760 and w46324;
w46455 <= not w46320 and w46454;
w46456 <= not w46321 and not w46324;
w46457 <= not w46455 and not w46456;
w46458 <= not w46379 and not w46457;
w46459 <= not w45750 and not w46378;
w46460 <= not w46377 and w46459;
w46461 <= not w46458 and not w46460;
w46462 <= not b(43) and not w46461;
w46463 <= not w45769 and w46319;
w46464 <= not w46315 and w46463;
w46465 <= not w46316 and not w46319;
w46466 <= not w46464 and not w46465;
w46467 <= not w46379 and not w46466;
w46468 <= not w45759 and not w46378;
w46469 <= not w46377 and w46468;
w46470 <= not w46467 and not w46469;
w46471 <= not b(42) and not w46470;
w46472 <= not w45778 and w46314;
w46473 <= not w46310 and w46472;
w46474 <= not w46311 and not w46314;
w46475 <= not w46473 and not w46474;
w46476 <= not w46379 and not w46475;
w46477 <= not w45768 and not w46378;
w46478 <= not w46377 and w46477;
w46479 <= not w46476 and not w46478;
w46480 <= not b(41) and not w46479;
w46481 <= not w45787 and w46309;
w46482 <= not w46305 and w46481;
w46483 <= not w46306 and not w46309;
w46484 <= not w46482 and not w46483;
w46485 <= not w46379 and not w46484;
w46486 <= not w45777 and not w46378;
w46487 <= not w46377 and w46486;
w46488 <= not w46485 and not w46487;
w46489 <= not b(40) and not w46488;
w46490 <= not w45796 and w46304;
w46491 <= not w46300 and w46490;
w46492 <= not w46301 and not w46304;
w46493 <= not w46491 and not w46492;
w46494 <= not w46379 and not w46493;
w46495 <= not w45786 and not w46378;
w46496 <= not w46377 and w46495;
w46497 <= not w46494 and not w46496;
w46498 <= not b(39) and not w46497;
w46499 <= not w45805 and w46299;
w46500 <= not w46295 and w46499;
w46501 <= not w46296 and not w46299;
w46502 <= not w46500 and not w46501;
w46503 <= not w46379 and not w46502;
w46504 <= not w45795 and not w46378;
w46505 <= not w46377 and w46504;
w46506 <= not w46503 and not w46505;
w46507 <= not b(38) and not w46506;
w46508 <= not w45814 and w46294;
w46509 <= not w46290 and w46508;
w46510 <= not w46291 and not w46294;
w46511 <= not w46509 and not w46510;
w46512 <= not w46379 and not w46511;
w46513 <= not w45804 and not w46378;
w46514 <= not w46377 and w46513;
w46515 <= not w46512 and not w46514;
w46516 <= not b(37) and not w46515;
w46517 <= not w45823 and w46289;
w46518 <= not w46285 and w46517;
w46519 <= not w46286 and not w46289;
w46520 <= not w46518 and not w46519;
w46521 <= not w46379 and not w46520;
w46522 <= not w45813 and not w46378;
w46523 <= not w46377 and w46522;
w46524 <= not w46521 and not w46523;
w46525 <= not b(36) and not w46524;
w46526 <= not w45832 and w46284;
w46527 <= not w46280 and w46526;
w46528 <= not w46281 and not w46284;
w46529 <= not w46527 and not w46528;
w46530 <= not w46379 and not w46529;
w46531 <= not w45822 and not w46378;
w46532 <= not w46377 and w46531;
w46533 <= not w46530 and not w46532;
w46534 <= not b(35) and not w46533;
w46535 <= not w45841 and w46279;
w46536 <= not w46275 and w46535;
w46537 <= not w46276 and not w46279;
w46538 <= not w46536 and not w46537;
w46539 <= not w46379 and not w46538;
w46540 <= not w45831 and not w46378;
w46541 <= not w46377 and w46540;
w46542 <= not w46539 and not w46541;
w46543 <= not b(34) and not w46542;
w46544 <= not w45850 and w46274;
w46545 <= not w46270 and w46544;
w46546 <= not w46271 and not w46274;
w46547 <= not w46545 and not w46546;
w46548 <= not w46379 and not w46547;
w46549 <= not w45840 and not w46378;
w46550 <= not w46377 and w46549;
w46551 <= not w46548 and not w46550;
w46552 <= not b(33) and not w46551;
w46553 <= not w45859 and w46269;
w46554 <= not w46265 and w46553;
w46555 <= not w46266 and not w46269;
w46556 <= not w46554 and not w46555;
w46557 <= not w46379 and not w46556;
w46558 <= not w45849 and not w46378;
w46559 <= not w46377 and w46558;
w46560 <= not w46557 and not w46559;
w46561 <= not b(32) and not w46560;
w46562 <= not w45868 and w46264;
w46563 <= not w46260 and w46562;
w46564 <= not w46261 and not w46264;
w46565 <= not w46563 and not w46564;
w46566 <= not w46379 and not w46565;
w46567 <= not w45858 and not w46378;
w46568 <= not w46377 and w46567;
w46569 <= not w46566 and not w46568;
w46570 <= not b(31) and not w46569;
w46571 <= not w45877 and w46259;
w46572 <= not w46255 and w46571;
w46573 <= not w46256 and not w46259;
w46574 <= not w46572 and not w46573;
w46575 <= not w46379 and not w46574;
w46576 <= not w45867 and not w46378;
w46577 <= not w46377 and w46576;
w46578 <= not w46575 and not w46577;
w46579 <= not b(30) and not w46578;
w46580 <= not w45886 and w46254;
w46581 <= not w46250 and w46580;
w46582 <= not w46251 and not w46254;
w46583 <= not w46581 and not w46582;
w46584 <= not w46379 and not w46583;
w46585 <= not w45876 and not w46378;
w46586 <= not w46377 and w46585;
w46587 <= not w46584 and not w46586;
w46588 <= not b(29) and not w46587;
w46589 <= not w45895 and w46249;
w46590 <= not w46245 and w46589;
w46591 <= not w46246 and not w46249;
w46592 <= not w46590 and not w46591;
w46593 <= not w46379 and not w46592;
w46594 <= not w45885 and not w46378;
w46595 <= not w46377 and w46594;
w46596 <= not w46593 and not w46595;
w46597 <= not b(28) and not w46596;
w46598 <= not w45904 and w46244;
w46599 <= not w46240 and w46598;
w46600 <= not w46241 and not w46244;
w46601 <= not w46599 and not w46600;
w46602 <= not w46379 and not w46601;
w46603 <= not w45894 and not w46378;
w46604 <= not w46377 and w46603;
w46605 <= not w46602 and not w46604;
w46606 <= not b(27) and not w46605;
w46607 <= not w45913 and w46239;
w46608 <= not w46235 and w46607;
w46609 <= not w46236 and not w46239;
w46610 <= not w46608 and not w46609;
w46611 <= not w46379 and not w46610;
w46612 <= not w45903 and not w46378;
w46613 <= not w46377 and w46612;
w46614 <= not w46611 and not w46613;
w46615 <= not b(26) and not w46614;
w46616 <= not w45922 and w46234;
w46617 <= not w46230 and w46616;
w46618 <= not w46231 and not w46234;
w46619 <= not w46617 and not w46618;
w46620 <= not w46379 and not w46619;
w46621 <= not w45912 and not w46378;
w46622 <= not w46377 and w46621;
w46623 <= not w46620 and not w46622;
w46624 <= not b(25) and not w46623;
w46625 <= not w45931 and w46229;
w46626 <= not w46225 and w46625;
w46627 <= not w46226 and not w46229;
w46628 <= not w46626 and not w46627;
w46629 <= not w46379 and not w46628;
w46630 <= not w45921 and not w46378;
w46631 <= not w46377 and w46630;
w46632 <= not w46629 and not w46631;
w46633 <= not b(24) and not w46632;
w46634 <= not w45940 and w46224;
w46635 <= not w46220 and w46634;
w46636 <= not w46221 and not w46224;
w46637 <= not w46635 and not w46636;
w46638 <= not w46379 and not w46637;
w46639 <= not w45930 and not w46378;
w46640 <= not w46377 and w46639;
w46641 <= not w46638 and not w46640;
w46642 <= not b(23) and not w46641;
w46643 <= not w45949 and w46219;
w46644 <= not w46215 and w46643;
w46645 <= not w46216 and not w46219;
w46646 <= not w46644 and not w46645;
w46647 <= not w46379 and not w46646;
w46648 <= not w45939 and not w46378;
w46649 <= not w46377 and w46648;
w46650 <= not w46647 and not w46649;
w46651 <= not b(22) and not w46650;
w46652 <= not w45958 and w46214;
w46653 <= not w46210 and w46652;
w46654 <= not w46211 and not w46214;
w46655 <= not w46653 and not w46654;
w46656 <= not w46379 and not w46655;
w46657 <= not w45948 and not w46378;
w46658 <= not w46377 and w46657;
w46659 <= not w46656 and not w46658;
w46660 <= not b(21) and not w46659;
w46661 <= not w45967 and w46209;
w46662 <= not w46205 and w46661;
w46663 <= not w46206 and not w46209;
w46664 <= not w46662 and not w46663;
w46665 <= not w46379 and not w46664;
w46666 <= not w45957 and not w46378;
w46667 <= not w46377 and w46666;
w46668 <= not w46665 and not w46667;
w46669 <= not b(20) and not w46668;
w46670 <= not w45976 and w46204;
w46671 <= not w46200 and w46670;
w46672 <= not w46201 and not w46204;
w46673 <= not w46671 and not w46672;
w46674 <= not w46379 and not w46673;
w46675 <= not w45966 and not w46378;
w46676 <= not w46377 and w46675;
w46677 <= not w46674 and not w46676;
w46678 <= not b(19) and not w46677;
w46679 <= not w45985 and w46199;
w46680 <= not w46195 and w46679;
w46681 <= not w46196 and not w46199;
w46682 <= not w46680 and not w46681;
w46683 <= not w46379 and not w46682;
w46684 <= not w45975 and not w46378;
w46685 <= not w46377 and w46684;
w46686 <= not w46683 and not w46685;
w46687 <= not b(18) and not w46686;
w46688 <= not w45994 and w46194;
w46689 <= not w46190 and w46688;
w46690 <= not w46191 and not w46194;
w46691 <= not w46689 and not w46690;
w46692 <= not w46379 and not w46691;
w46693 <= not w45984 and not w46378;
w46694 <= not w46377 and w46693;
w46695 <= not w46692 and not w46694;
w46696 <= not b(17) and not w46695;
w46697 <= not w46003 and w46189;
w46698 <= not w46185 and w46697;
w46699 <= not w46186 and not w46189;
w46700 <= not w46698 and not w46699;
w46701 <= not w46379 and not w46700;
w46702 <= not w45993 and not w46378;
w46703 <= not w46377 and w46702;
w46704 <= not w46701 and not w46703;
w46705 <= not b(16) and not w46704;
w46706 <= not w46012 and w46184;
w46707 <= not w46180 and w46706;
w46708 <= not w46181 and not w46184;
w46709 <= not w46707 and not w46708;
w46710 <= not w46379 and not w46709;
w46711 <= not w46002 and not w46378;
w46712 <= not w46377 and w46711;
w46713 <= not w46710 and not w46712;
w46714 <= not b(15) and not w46713;
w46715 <= not w46021 and w46179;
w46716 <= not w46175 and w46715;
w46717 <= not w46176 and not w46179;
w46718 <= not w46716 and not w46717;
w46719 <= not w46379 and not w46718;
w46720 <= not w46011 and not w46378;
w46721 <= not w46377 and w46720;
w46722 <= not w46719 and not w46721;
w46723 <= not b(14) and not w46722;
w46724 <= not w46030 and w46174;
w46725 <= not w46170 and w46724;
w46726 <= not w46171 and not w46174;
w46727 <= not w46725 and not w46726;
w46728 <= not w46379 and not w46727;
w46729 <= not w46020 and not w46378;
w46730 <= not w46377 and w46729;
w46731 <= not w46728 and not w46730;
w46732 <= not b(13) and not w46731;
w46733 <= not w46039 and w46169;
w46734 <= not w46165 and w46733;
w46735 <= not w46166 and not w46169;
w46736 <= not w46734 and not w46735;
w46737 <= not w46379 and not w46736;
w46738 <= not w46029 and not w46378;
w46739 <= not w46377 and w46738;
w46740 <= not w46737 and not w46739;
w46741 <= not b(12) and not w46740;
w46742 <= not w46048 and w46164;
w46743 <= not w46160 and w46742;
w46744 <= not w46161 and not w46164;
w46745 <= not w46743 and not w46744;
w46746 <= not w46379 and not w46745;
w46747 <= not w46038 and not w46378;
w46748 <= not w46377 and w46747;
w46749 <= not w46746 and not w46748;
w46750 <= not b(11) and not w46749;
w46751 <= not w46057 and w46159;
w46752 <= not w46155 and w46751;
w46753 <= not w46156 and not w46159;
w46754 <= not w46752 and not w46753;
w46755 <= not w46379 and not w46754;
w46756 <= not w46047 and not w46378;
w46757 <= not w46377 and w46756;
w46758 <= not w46755 and not w46757;
w46759 <= not b(10) and not w46758;
w46760 <= not w46066 and w46154;
w46761 <= not w46150 and w46760;
w46762 <= not w46151 and not w46154;
w46763 <= not w46761 and not w46762;
w46764 <= not w46379 and not w46763;
w46765 <= not w46056 and not w46378;
w46766 <= not w46377 and w46765;
w46767 <= not w46764 and not w46766;
w46768 <= not b(9) and not w46767;
w46769 <= not w46075 and w46149;
w46770 <= not w46145 and w46769;
w46771 <= not w46146 and not w46149;
w46772 <= not w46770 and not w46771;
w46773 <= not w46379 and not w46772;
w46774 <= not w46065 and not w46378;
w46775 <= not w46377 and w46774;
w46776 <= not w46773 and not w46775;
w46777 <= not b(8) and not w46776;
w46778 <= not w46084 and w46144;
w46779 <= not w46140 and w46778;
w46780 <= not w46141 and not w46144;
w46781 <= not w46779 and not w46780;
w46782 <= not w46379 and not w46781;
w46783 <= not w46074 and not w46378;
w46784 <= not w46377 and w46783;
w46785 <= not w46782 and not w46784;
w46786 <= not b(7) and not w46785;
w46787 <= not w46093 and w46139;
w46788 <= not w46135 and w46787;
w46789 <= not w46136 and not w46139;
w46790 <= not w46788 and not w46789;
w46791 <= not w46379 and not w46790;
w46792 <= not w46083 and not w46378;
w46793 <= not w46377 and w46792;
w46794 <= not w46791 and not w46793;
w46795 <= not b(6) and not w46794;
w46796 <= not w46102 and w46134;
w46797 <= not w46130 and w46796;
w46798 <= not w46131 and not w46134;
w46799 <= not w46797 and not w46798;
w46800 <= not w46379 and not w46799;
w46801 <= not w46092 and not w46378;
w46802 <= not w46377 and w46801;
w46803 <= not w46800 and not w46802;
w46804 <= not b(5) and not w46803;
w46805 <= not w46110 and w46129;
w46806 <= not w46125 and w46805;
w46807 <= not w46126 and not w46129;
w46808 <= not w46806 and not w46807;
w46809 <= not w46379 and not w46808;
w46810 <= not w46101 and not w46378;
w46811 <= not w46377 and w46810;
w46812 <= not w46809 and not w46811;
w46813 <= not b(4) and not w46812;
w46814 <= not w46120 and w46124;
w46815 <= not w46119 and w46814;
w46816 <= not w46121 and not w46124;
w46817 <= not w46815 and not w46816;
w46818 <= not w46379 and not w46817;
w46819 <= not w46109 and not w46378;
w46820 <= not w46377 and w46819;
w46821 <= not w46818 and not w46820;
w46822 <= not b(3) and not w46821;
w46823 <= w18070 and not w46117;
w46824 <= not w46115 and w46823;
w46825 <= not w46119 and not w46824;
w46826 <= not w46379 and w46825;
w46827 <= not w46114 and not w46378;
w46828 <= not w46377 and w46827;
w46829 <= not w46826 and not w46828;
w46830 <= not b(2) and not w46829;
w46831 <= b(0) and not w46379;
w46832 <= a(13) and not w46831;
w46833 <= w18070 and not w46379;
w46834 <= not w46832 and not w46833;
w46835 <= b(1) and not w46834;
w46836 <= not b(1) and not w46833;
w46837 <= not w46832 and w46836;
w46838 <= not w46835 and not w46837;
w46839 <= not w18793 and not w46838;
w46840 <= not b(1) and not w46834;
w46841 <= not w46839 and not w46840;
w46842 <= b(2) and not w46828;
w46843 <= not w46826 and w46842;
w46844 <= not w46830 and not w46843;
w46845 <= not w46841 and w46844;
w46846 <= not w46830 and not w46845;
w46847 <= b(3) and not w46820;
w46848 <= not w46818 and w46847;
w46849 <= not w46822 and not w46848;
w46850 <= not w46846 and w46849;
w46851 <= not w46822 and not w46850;
w46852 <= b(4) and not w46811;
w46853 <= not w46809 and w46852;
w46854 <= not w46813 and not w46853;
w46855 <= not w46851 and w46854;
w46856 <= not w46813 and not w46855;
w46857 <= b(5) and not w46802;
w46858 <= not w46800 and w46857;
w46859 <= not w46804 and not w46858;
w46860 <= not w46856 and w46859;
w46861 <= not w46804 and not w46860;
w46862 <= b(6) and not w46793;
w46863 <= not w46791 and w46862;
w46864 <= not w46795 and not w46863;
w46865 <= not w46861 and w46864;
w46866 <= not w46795 and not w46865;
w46867 <= b(7) and not w46784;
w46868 <= not w46782 and w46867;
w46869 <= not w46786 and not w46868;
w46870 <= not w46866 and w46869;
w46871 <= not w46786 and not w46870;
w46872 <= b(8) and not w46775;
w46873 <= not w46773 and w46872;
w46874 <= not w46777 and not w46873;
w46875 <= not w46871 and w46874;
w46876 <= not w46777 and not w46875;
w46877 <= b(9) and not w46766;
w46878 <= not w46764 and w46877;
w46879 <= not w46768 and not w46878;
w46880 <= not w46876 and w46879;
w46881 <= not w46768 and not w46880;
w46882 <= b(10) and not w46757;
w46883 <= not w46755 and w46882;
w46884 <= not w46759 and not w46883;
w46885 <= not w46881 and w46884;
w46886 <= not w46759 and not w46885;
w46887 <= b(11) and not w46748;
w46888 <= not w46746 and w46887;
w46889 <= not w46750 and not w46888;
w46890 <= not w46886 and w46889;
w46891 <= not w46750 and not w46890;
w46892 <= b(12) and not w46739;
w46893 <= not w46737 and w46892;
w46894 <= not w46741 and not w46893;
w46895 <= not w46891 and w46894;
w46896 <= not w46741 and not w46895;
w46897 <= b(13) and not w46730;
w46898 <= not w46728 and w46897;
w46899 <= not w46732 and not w46898;
w46900 <= not w46896 and w46899;
w46901 <= not w46732 and not w46900;
w46902 <= b(14) and not w46721;
w46903 <= not w46719 and w46902;
w46904 <= not w46723 and not w46903;
w46905 <= not w46901 and w46904;
w46906 <= not w46723 and not w46905;
w46907 <= b(15) and not w46712;
w46908 <= not w46710 and w46907;
w46909 <= not w46714 and not w46908;
w46910 <= not w46906 and w46909;
w46911 <= not w46714 and not w46910;
w46912 <= b(16) and not w46703;
w46913 <= not w46701 and w46912;
w46914 <= not w46705 and not w46913;
w46915 <= not w46911 and w46914;
w46916 <= not w46705 and not w46915;
w46917 <= b(17) and not w46694;
w46918 <= not w46692 and w46917;
w46919 <= not w46696 and not w46918;
w46920 <= not w46916 and w46919;
w46921 <= not w46696 and not w46920;
w46922 <= b(18) and not w46685;
w46923 <= not w46683 and w46922;
w46924 <= not w46687 and not w46923;
w46925 <= not w46921 and w46924;
w46926 <= not w46687 and not w46925;
w46927 <= b(19) and not w46676;
w46928 <= not w46674 and w46927;
w46929 <= not w46678 and not w46928;
w46930 <= not w46926 and w46929;
w46931 <= not w46678 and not w46930;
w46932 <= b(20) and not w46667;
w46933 <= not w46665 and w46932;
w46934 <= not w46669 and not w46933;
w46935 <= not w46931 and w46934;
w46936 <= not w46669 and not w46935;
w46937 <= b(21) and not w46658;
w46938 <= not w46656 and w46937;
w46939 <= not w46660 and not w46938;
w46940 <= not w46936 and w46939;
w46941 <= not w46660 and not w46940;
w46942 <= b(22) and not w46649;
w46943 <= not w46647 and w46942;
w46944 <= not w46651 and not w46943;
w46945 <= not w46941 and w46944;
w46946 <= not w46651 and not w46945;
w46947 <= b(23) and not w46640;
w46948 <= not w46638 and w46947;
w46949 <= not w46642 and not w46948;
w46950 <= not w46946 and w46949;
w46951 <= not w46642 and not w46950;
w46952 <= b(24) and not w46631;
w46953 <= not w46629 and w46952;
w46954 <= not w46633 and not w46953;
w46955 <= not w46951 and w46954;
w46956 <= not w46633 and not w46955;
w46957 <= b(25) and not w46622;
w46958 <= not w46620 and w46957;
w46959 <= not w46624 and not w46958;
w46960 <= not w46956 and w46959;
w46961 <= not w46624 and not w46960;
w46962 <= b(26) and not w46613;
w46963 <= not w46611 and w46962;
w46964 <= not w46615 and not w46963;
w46965 <= not w46961 and w46964;
w46966 <= not w46615 and not w46965;
w46967 <= b(27) and not w46604;
w46968 <= not w46602 and w46967;
w46969 <= not w46606 and not w46968;
w46970 <= not w46966 and w46969;
w46971 <= not w46606 and not w46970;
w46972 <= b(28) and not w46595;
w46973 <= not w46593 and w46972;
w46974 <= not w46597 and not w46973;
w46975 <= not w46971 and w46974;
w46976 <= not w46597 and not w46975;
w46977 <= b(29) and not w46586;
w46978 <= not w46584 and w46977;
w46979 <= not w46588 and not w46978;
w46980 <= not w46976 and w46979;
w46981 <= not w46588 and not w46980;
w46982 <= b(30) and not w46577;
w46983 <= not w46575 and w46982;
w46984 <= not w46579 and not w46983;
w46985 <= not w46981 and w46984;
w46986 <= not w46579 and not w46985;
w46987 <= b(31) and not w46568;
w46988 <= not w46566 and w46987;
w46989 <= not w46570 and not w46988;
w46990 <= not w46986 and w46989;
w46991 <= not w46570 and not w46990;
w46992 <= b(32) and not w46559;
w46993 <= not w46557 and w46992;
w46994 <= not w46561 and not w46993;
w46995 <= not w46991 and w46994;
w46996 <= not w46561 and not w46995;
w46997 <= b(33) and not w46550;
w46998 <= not w46548 and w46997;
w46999 <= not w46552 and not w46998;
w47000 <= not w46996 and w46999;
w47001 <= not w46552 and not w47000;
w47002 <= b(34) and not w46541;
w47003 <= not w46539 and w47002;
w47004 <= not w46543 and not w47003;
w47005 <= not w47001 and w47004;
w47006 <= not w46543 and not w47005;
w47007 <= b(35) and not w46532;
w47008 <= not w46530 and w47007;
w47009 <= not w46534 and not w47008;
w47010 <= not w47006 and w47009;
w47011 <= not w46534 and not w47010;
w47012 <= b(36) and not w46523;
w47013 <= not w46521 and w47012;
w47014 <= not w46525 and not w47013;
w47015 <= not w47011 and w47014;
w47016 <= not w46525 and not w47015;
w47017 <= b(37) and not w46514;
w47018 <= not w46512 and w47017;
w47019 <= not w46516 and not w47018;
w47020 <= not w47016 and w47019;
w47021 <= not w46516 and not w47020;
w47022 <= b(38) and not w46505;
w47023 <= not w46503 and w47022;
w47024 <= not w46507 and not w47023;
w47025 <= not w47021 and w47024;
w47026 <= not w46507 and not w47025;
w47027 <= b(39) and not w46496;
w47028 <= not w46494 and w47027;
w47029 <= not w46498 and not w47028;
w47030 <= not w47026 and w47029;
w47031 <= not w46498 and not w47030;
w47032 <= b(40) and not w46487;
w47033 <= not w46485 and w47032;
w47034 <= not w46489 and not w47033;
w47035 <= not w47031 and w47034;
w47036 <= not w46489 and not w47035;
w47037 <= b(41) and not w46478;
w47038 <= not w46476 and w47037;
w47039 <= not w46480 and not w47038;
w47040 <= not w47036 and w47039;
w47041 <= not w46480 and not w47040;
w47042 <= b(42) and not w46469;
w47043 <= not w46467 and w47042;
w47044 <= not w46471 and not w47043;
w47045 <= not w47041 and w47044;
w47046 <= not w46471 and not w47045;
w47047 <= b(43) and not w46460;
w47048 <= not w46458 and w47047;
w47049 <= not w46462 and not w47048;
w47050 <= not w47046 and w47049;
w47051 <= not w46462 and not w47050;
w47052 <= b(44) and not w46451;
w47053 <= not w46449 and w47052;
w47054 <= not w46453 and not w47053;
w47055 <= not w47051 and w47054;
w47056 <= not w46453 and not w47055;
w47057 <= b(45) and not w46442;
w47058 <= not w46440 and w47057;
w47059 <= not w46444 and not w47058;
w47060 <= not w47056 and w47059;
w47061 <= not w46444 and not w47060;
w47062 <= b(46) and not w46433;
w47063 <= not w46431 and w47062;
w47064 <= not w46435 and not w47063;
w47065 <= not w47061 and w47064;
w47066 <= not w46435 and not w47065;
w47067 <= b(47) and not w46424;
w47068 <= not w46422 and w47067;
w47069 <= not w46426 and not w47068;
w47070 <= not w47066 and w47069;
w47071 <= not w46426 and not w47070;
w47072 <= b(48) and not w46415;
w47073 <= not w46413 and w47072;
w47074 <= not w46417 and not w47073;
w47075 <= not w47071 and w47074;
w47076 <= not w46417 and not w47075;
w47077 <= b(49) and not w46406;
w47078 <= not w46404 and w47077;
w47079 <= not w46408 and not w47078;
w47080 <= not w47076 and w47079;
w47081 <= not w46408 and not w47080;
w47082 <= b(50) and not w46386;
w47083 <= not w46384 and w47082;
w47084 <= not w46399 and not w47083;
w47085 <= not w47081 and w47084;
w47086 <= not w46399 and not w47085;
w47087 <= b(51) and not w46396;
w47088 <= not w46394 and w47087;
w47089 <= not w46398 and not w47088;
w47090 <= not w47086 and w47089;
w47091 <= not w46398 and not w47090;
w47092 <= w31 and not w47091;
w47093 <= not w46387 and not w47092;
w47094 <= not w46408 and w47084;
w47095 <= not w47080 and w47094;
w47096 <= not w47081 and not w47084;
w47097 <= not w47095 and not w47096;
w47098 <= w31 and not w47097;
w47099 <= not w47091 and w47098;
w47100 <= not w47093 and not w47099;
w47101 <= not b(51) and not w47100;
w47102 <= not w46407 and not w47092;
w47103 <= not w46417 and w47079;
w47104 <= not w47075 and w47103;
w47105 <= not w47076 and not w47079;
w47106 <= not w47104 and not w47105;
w47107 <= w31 and not w47106;
w47108 <= not w47091 and w47107;
w47109 <= not w47102 and not w47108;
w47110 <= not b(50) and not w47109;
w47111 <= not w46416 and not w47092;
w47112 <= not w46426 and w47074;
w47113 <= not w47070 and w47112;
w47114 <= not w47071 and not w47074;
w47115 <= not w47113 and not w47114;
w47116 <= w31 and not w47115;
w47117 <= not w47091 and w47116;
w47118 <= not w47111 and not w47117;
w47119 <= not b(49) and not w47118;
w47120 <= not w46425 and not w47092;
w47121 <= not w46435 and w47069;
w47122 <= not w47065 and w47121;
w47123 <= not w47066 and not w47069;
w47124 <= not w47122 and not w47123;
w47125 <= w31 and not w47124;
w47126 <= not w47091 and w47125;
w47127 <= not w47120 and not w47126;
w47128 <= not b(48) and not w47127;
w47129 <= not w46434 and not w47092;
w47130 <= not w46444 and w47064;
w47131 <= not w47060 and w47130;
w47132 <= not w47061 and not w47064;
w47133 <= not w47131 and not w47132;
w47134 <= w31 and not w47133;
w47135 <= not w47091 and w47134;
w47136 <= not w47129 and not w47135;
w47137 <= not b(47) and not w47136;
w47138 <= not w46443 and not w47092;
w47139 <= not w46453 and w47059;
w47140 <= not w47055 and w47139;
w47141 <= not w47056 and not w47059;
w47142 <= not w47140 and not w47141;
w47143 <= w31 and not w47142;
w47144 <= not w47091 and w47143;
w47145 <= not w47138 and not w47144;
w47146 <= not b(46) and not w47145;
w47147 <= not w46452 and not w47092;
w47148 <= not w46462 and w47054;
w47149 <= not w47050 and w47148;
w47150 <= not w47051 and not w47054;
w47151 <= not w47149 and not w47150;
w47152 <= w31 and not w47151;
w47153 <= not w47091 and w47152;
w47154 <= not w47147 and not w47153;
w47155 <= not b(45) and not w47154;
w47156 <= not w46461 and not w47092;
w47157 <= not w46471 and w47049;
w47158 <= not w47045 and w47157;
w47159 <= not w47046 and not w47049;
w47160 <= not w47158 and not w47159;
w47161 <= w31 and not w47160;
w47162 <= not w47091 and w47161;
w47163 <= not w47156 and not w47162;
w47164 <= not b(44) and not w47163;
w47165 <= not w46470 and not w47092;
w47166 <= not w46480 and w47044;
w47167 <= not w47040 and w47166;
w47168 <= not w47041 and not w47044;
w47169 <= not w47167 and not w47168;
w47170 <= w31 and not w47169;
w47171 <= not w47091 and w47170;
w47172 <= not w47165 and not w47171;
w47173 <= not b(43) and not w47172;
w47174 <= not w46479 and not w47092;
w47175 <= not w46489 and w47039;
w47176 <= not w47035 and w47175;
w47177 <= not w47036 and not w47039;
w47178 <= not w47176 and not w47177;
w47179 <= w31 and not w47178;
w47180 <= not w47091 and w47179;
w47181 <= not w47174 and not w47180;
w47182 <= not b(42) and not w47181;
w47183 <= not w46488 and not w47092;
w47184 <= not w46498 and w47034;
w47185 <= not w47030 and w47184;
w47186 <= not w47031 and not w47034;
w47187 <= not w47185 and not w47186;
w47188 <= w31 and not w47187;
w47189 <= not w47091 and w47188;
w47190 <= not w47183 and not w47189;
w47191 <= not b(41) and not w47190;
w47192 <= not w46497 and not w47092;
w47193 <= not w46507 and w47029;
w47194 <= not w47025 and w47193;
w47195 <= not w47026 and not w47029;
w47196 <= not w47194 and not w47195;
w47197 <= w31 and not w47196;
w47198 <= not w47091 and w47197;
w47199 <= not w47192 and not w47198;
w47200 <= not b(40) and not w47199;
w47201 <= not w46506 and not w47092;
w47202 <= not w46516 and w47024;
w47203 <= not w47020 and w47202;
w47204 <= not w47021 and not w47024;
w47205 <= not w47203 and not w47204;
w47206 <= w31 and not w47205;
w47207 <= not w47091 and w47206;
w47208 <= not w47201 and not w47207;
w47209 <= not b(39) and not w47208;
w47210 <= not w46515 and not w47092;
w47211 <= not w46525 and w47019;
w47212 <= not w47015 and w47211;
w47213 <= not w47016 and not w47019;
w47214 <= not w47212 and not w47213;
w47215 <= w31 and not w47214;
w47216 <= not w47091 and w47215;
w47217 <= not w47210 and not w47216;
w47218 <= not b(38) and not w47217;
w47219 <= not w46524 and not w47092;
w47220 <= not w46534 and w47014;
w47221 <= not w47010 and w47220;
w47222 <= not w47011 and not w47014;
w47223 <= not w47221 and not w47222;
w47224 <= w31 and not w47223;
w47225 <= not w47091 and w47224;
w47226 <= not w47219 and not w47225;
w47227 <= not b(37) and not w47226;
w47228 <= not w46533 and not w47092;
w47229 <= not w46543 and w47009;
w47230 <= not w47005 and w47229;
w47231 <= not w47006 and not w47009;
w47232 <= not w47230 and not w47231;
w47233 <= w31 and not w47232;
w47234 <= not w47091 and w47233;
w47235 <= not w47228 and not w47234;
w47236 <= not b(36) and not w47235;
w47237 <= not w46542 and not w47092;
w47238 <= not w46552 and w47004;
w47239 <= not w47000 and w47238;
w47240 <= not w47001 and not w47004;
w47241 <= not w47239 and not w47240;
w47242 <= w31 and not w47241;
w47243 <= not w47091 and w47242;
w47244 <= not w47237 and not w47243;
w47245 <= not b(35) and not w47244;
w47246 <= not w46551 and not w47092;
w47247 <= not w46561 and w46999;
w47248 <= not w46995 and w47247;
w47249 <= not w46996 and not w46999;
w47250 <= not w47248 and not w47249;
w47251 <= w31 and not w47250;
w47252 <= not w47091 and w47251;
w47253 <= not w47246 and not w47252;
w47254 <= not b(34) and not w47253;
w47255 <= not w46560 and not w47092;
w47256 <= not w46570 and w46994;
w47257 <= not w46990 and w47256;
w47258 <= not w46991 and not w46994;
w47259 <= not w47257 and not w47258;
w47260 <= w31 and not w47259;
w47261 <= not w47091 and w47260;
w47262 <= not w47255 and not w47261;
w47263 <= not b(33) and not w47262;
w47264 <= not w46569 and not w47092;
w47265 <= not w46579 and w46989;
w47266 <= not w46985 and w47265;
w47267 <= not w46986 and not w46989;
w47268 <= not w47266 and not w47267;
w47269 <= w31 and not w47268;
w47270 <= not w47091 and w47269;
w47271 <= not w47264 and not w47270;
w47272 <= not b(32) and not w47271;
w47273 <= not w46578 and not w47092;
w47274 <= not w46588 and w46984;
w47275 <= not w46980 and w47274;
w47276 <= not w46981 and not w46984;
w47277 <= not w47275 and not w47276;
w47278 <= w31 and not w47277;
w47279 <= not w47091 and w47278;
w47280 <= not w47273 and not w47279;
w47281 <= not b(31) and not w47280;
w47282 <= not w46587 and not w47092;
w47283 <= not w46597 and w46979;
w47284 <= not w46975 and w47283;
w47285 <= not w46976 and not w46979;
w47286 <= not w47284 and not w47285;
w47287 <= w31 and not w47286;
w47288 <= not w47091 and w47287;
w47289 <= not w47282 and not w47288;
w47290 <= not b(30) and not w47289;
w47291 <= not w46596 and not w47092;
w47292 <= not w46606 and w46974;
w47293 <= not w46970 and w47292;
w47294 <= not w46971 and not w46974;
w47295 <= not w47293 and not w47294;
w47296 <= w31 and not w47295;
w47297 <= not w47091 and w47296;
w47298 <= not w47291 and not w47297;
w47299 <= not b(29) and not w47298;
w47300 <= not w46605 and not w47092;
w47301 <= not w46615 and w46969;
w47302 <= not w46965 and w47301;
w47303 <= not w46966 and not w46969;
w47304 <= not w47302 and not w47303;
w47305 <= w31 and not w47304;
w47306 <= not w47091 and w47305;
w47307 <= not w47300 and not w47306;
w47308 <= not b(28) and not w47307;
w47309 <= not w46614 and not w47092;
w47310 <= not w46624 and w46964;
w47311 <= not w46960 and w47310;
w47312 <= not w46961 and not w46964;
w47313 <= not w47311 and not w47312;
w47314 <= w31 and not w47313;
w47315 <= not w47091 and w47314;
w47316 <= not w47309 and not w47315;
w47317 <= not b(27) and not w47316;
w47318 <= not w46623 and not w47092;
w47319 <= not w46633 and w46959;
w47320 <= not w46955 and w47319;
w47321 <= not w46956 and not w46959;
w47322 <= not w47320 and not w47321;
w47323 <= w31 and not w47322;
w47324 <= not w47091 and w47323;
w47325 <= not w47318 and not w47324;
w47326 <= not b(26) and not w47325;
w47327 <= not w46632 and not w47092;
w47328 <= not w46642 and w46954;
w47329 <= not w46950 and w47328;
w47330 <= not w46951 and not w46954;
w47331 <= not w47329 and not w47330;
w47332 <= w31 and not w47331;
w47333 <= not w47091 and w47332;
w47334 <= not w47327 and not w47333;
w47335 <= not b(25) and not w47334;
w47336 <= not w46641 and not w47092;
w47337 <= not w46651 and w46949;
w47338 <= not w46945 and w47337;
w47339 <= not w46946 and not w46949;
w47340 <= not w47338 and not w47339;
w47341 <= w31 and not w47340;
w47342 <= not w47091 and w47341;
w47343 <= not w47336 and not w47342;
w47344 <= not b(24) and not w47343;
w47345 <= not w46650 and not w47092;
w47346 <= not w46660 and w46944;
w47347 <= not w46940 and w47346;
w47348 <= not w46941 and not w46944;
w47349 <= not w47347 and not w47348;
w47350 <= w31 and not w47349;
w47351 <= not w47091 and w47350;
w47352 <= not w47345 and not w47351;
w47353 <= not b(23) and not w47352;
w47354 <= not w46659 and not w47092;
w47355 <= not w46669 and w46939;
w47356 <= not w46935 and w47355;
w47357 <= not w46936 and not w46939;
w47358 <= not w47356 and not w47357;
w47359 <= w31 and not w47358;
w47360 <= not w47091 and w47359;
w47361 <= not w47354 and not w47360;
w47362 <= not b(22) and not w47361;
w47363 <= not w46668 and not w47092;
w47364 <= not w46678 and w46934;
w47365 <= not w46930 and w47364;
w47366 <= not w46931 and not w46934;
w47367 <= not w47365 and not w47366;
w47368 <= w31 and not w47367;
w47369 <= not w47091 and w47368;
w47370 <= not w47363 and not w47369;
w47371 <= not b(21) and not w47370;
w47372 <= not w46677 and not w47092;
w47373 <= not w46687 and w46929;
w47374 <= not w46925 and w47373;
w47375 <= not w46926 and not w46929;
w47376 <= not w47374 and not w47375;
w47377 <= w31 and not w47376;
w47378 <= not w47091 and w47377;
w47379 <= not w47372 and not w47378;
w47380 <= not b(20) and not w47379;
w47381 <= not w46686 and not w47092;
w47382 <= not w46696 and w46924;
w47383 <= not w46920 and w47382;
w47384 <= not w46921 and not w46924;
w47385 <= not w47383 and not w47384;
w47386 <= w31 and not w47385;
w47387 <= not w47091 and w47386;
w47388 <= not w47381 and not w47387;
w47389 <= not b(19) and not w47388;
w47390 <= not w46695 and not w47092;
w47391 <= not w46705 and w46919;
w47392 <= not w46915 and w47391;
w47393 <= not w46916 and not w46919;
w47394 <= not w47392 and not w47393;
w47395 <= w31 and not w47394;
w47396 <= not w47091 and w47395;
w47397 <= not w47390 and not w47396;
w47398 <= not b(18) and not w47397;
w47399 <= not w46704 and not w47092;
w47400 <= not w46714 and w46914;
w47401 <= not w46910 and w47400;
w47402 <= not w46911 and not w46914;
w47403 <= not w47401 and not w47402;
w47404 <= w31 and not w47403;
w47405 <= not w47091 and w47404;
w47406 <= not w47399 and not w47405;
w47407 <= not b(17) and not w47406;
w47408 <= not w46713 and not w47092;
w47409 <= not w46723 and w46909;
w47410 <= not w46905 and w47409;
w47411 <= not w46906 and not w46909;
w47412 <= not w47410 and not w47411;
w47413 <= w31 and not w47412;
w47414 <= not w47091 and w47413;
w47415 <= not w47408 and not w47414;
w47416 <= not b(16) and not w47415;
w47417 <= not w46722 and not w47092;
w47418 <= not w46732 and w46904;
w47419 <= not w46900 and w47418;
w47420 <= not w46901 and not w46904;
w47421 <= not w47419 and not w47420;
w47422 <= w31 and not w47421;
w47423 <= not w47091 and w47422;
w47424 <= not w47417 and not w47423;
w47425 <= not b(15) and not w47424;
w47426 <= not w46731 and not w47092;
w47427 <= not w46741 and w46899;
w47428 <= not w46895 and w47427;
w47429 <= not w46896 and not w46899;
w47430 <= not w47428 and not w47429;
w47431 <= w31 and not w47430;
w47432 <= not w47091 and w47431;
w47433 <= not w47426 and not w47432;
w47434 <= not b(14) and not w47433;
w47435 <= not w46740 and not w47092;
w47436 <= not w46750 and w46894;
w47437 <= not w46890 and w47436;
w47438 <= not w46891 and not w46894;
w47439 <= not w47437 and not w47438;
w47440 <= w31 and not w47439;
w47441 <= not w47091 and w47440;
w47442 <= not w47435 and not w47441;
w47443 <= not b(13) and not w47442;
w47444 <= not w46749 and not w47092;
w47445 <= not w46759 and w46889;
w47446 <= not w46885 and w47445;
w47447 <= not w46886 and not w46889;
w47448 <= not w47446 and not w47447;
w47449 <= w31 and not w47448;
w47450 <= not w47091 and w47449;
w47451 <= not w47444 and not w47450;
w47452 <= not b(12) and not w47451;
w47453 <= not w46758 and not w47092;
w47454 <= not w46768 and w46884;
w47455 <= not w46880 and w47454;
w47456 <= not w46881 and not w46884;
w47457 <= not w47455 and not w47456;
w47458 <= w31 and not w47457;
w47459 <= not w47091 and w47458;
w47460 <= not w47453 and not w47459;
w47461 <= not b(11) and not w47460;
w47462 <= not w46767 and not w47092;
w47463 <= not w46777 and w46879;
w47464 <= not w46875 and w47463;
w47465 <= not w46876 and not w46879;
w47466 <= not w47464 and not w47465;
w47467 <= w31 and not w47466;
w47468 <= not w47091 and w47467;
w47469 <= not w47462 and not w47468;
w47470 <= not b(10) and not w47469;
w47471 <= not w46776 and not w47092;
w47472 <= not w46786 and w46874;
w47473 <= not w46870 and w47472;
w47474 <= not w46871 and not w46874;
w47475 <= not w47473 and not w47474;
w47476 <= w31 and not w47475;
w47477 <= not w47091 and w47476;
w47478 <= not w47471 and not w47477;
w47479 <= not b(9) and not w47478;
w47480 <= not w46785 and not w47092;
w47481 <= not w46795 and w46869;
w47482 <= not w46865 and w47481;
w47483 <= not w46866 and not w46869;
w47484 <= not w47482 and not w47483;
w47485 <= w31 and not w47484;
w47486 <= not w47091 and w47485;
w47487 <= not w47480 and not w47486;
w47488 <= not b(8) and not w47487;
w47489 <= not w46794 and not w47092;
w47490 <= not w46804 and w46864;
w47491 <= not w46860 and w47490;
w47492 <= not w46861 and not w46864;
w47493 <= not w47491 and not w47492;
w47494 <= w31 and not w47493;
w47495 <= not w47091 and w47494;
w47496 <= not w47489 and not w47495;
w47497 <= not b(7) and not w47496;
w47498 <= not w46803 and not w47092;
w47499 <= not w46813 and w46859;
w47500 <= not w46855 and w47499;
w47501 <= not w46856 and not w46859;
w47502 <= not w47500 and not w47501;
w47503 <= w31 and not w47502;
w47504 <= not w47091 and w47503;
w47505 <= not w47498 and not w47504;
w47506 <= not b(6) and not w47505;
w47507 <= not w46812 and not w47092;
w47508 <= not w46822 and w46854;
w47509 <= not w46850 and w47508;
w47510 <= not w46851 and not w46854;
w47511 <= not w47509 and not w47510;
w47512 <= w31 and not w47511;
w47513 <= not w47091 and w47512;
w47514 <= not w47507 and not w47513;
w47515 <= not b(5) and not w47514;
w47516 <= not w46821 and not w47092;
w47517 <= not w46830 and w46849;
w47518 <= not w46845 and w47517;
w47519 <= not w46846 and not w46849;
w47520 <= not w47518 and not w47519;
w47521 <= w31 and not w47520;
w47522 <= not w47091 and w47521;
w47523 <= not w47516 and not w47522;
w47524 <= not b(4) and not w47523;
w47525 <= not w46829 and not w47092;
w47526 <= not w46840 and w46844;
w47527 <= not w46839 and w47526;
w47528 <= not w46841 and not w46844;
w47529 <= not w47527 and not w47528;
w47530 <= w31 and not w47529;
w47531 <= not w47091 and w47530;
w47532 <= not w47525 and not w47531;
w47533 <= not b(3) and not w47532;
w47534 <= not w46834 and not w47092;
w47535 <= w18793 and not w46837;
w47536 <= not w46835 and w47535;
w47537 <= w31 and not w47536;
w47538 <= not w46839 and w47537;
w47539 <= not w47091 and w47538;
w47540 <= not w47534 and not w47539;
w47541 <= not b(2) and not w47540;
w47542 <= w19499 and not w47091;
w47543 <= a(12) and not w47542;
w47544 <= w19503 and not w47091;
w47545 <= not w47543 and not w47544;
w47546 <= b(1) and not w47545;
w47547 <= not b(1) and not w47544;
w47548 <= not w47543 and w47547;
w47549 <= not w47546 and not w47548;
w47550 <= not w19510 and not w47549;
w47551 <= not b(1) and not w47545;
w47552 <= not w47550 and not w47551;
w47553 <= b(2) and not w47539;
w47554 <= not w47534 and w47553;
w47555 <= not w47541 and not w47554;
w47556 <= not w47552 and w47555;
w47557 <= not w47541 and not w47556;
w47558 <= b(3) and not w47531;
w47559 <= not w47525 and w47558;
w47560 <= not w47533 and not w47559;
w47561 <= not w47557 and w47560;
w47562 <= not w47533 and not w47561;
w47563 <= b(4) and not w47522;
w47564 <= not w47516 and w47563;
w47565 <= not w47524 and not w47564;
w47566 <= not w47562 and w47565;
w47567 <= not w47524 and not w47566;
w47568 <= b(5) and not w47513;
w47569 <= not w47507 and w47568;
w47570 <= not w47515 and not w47569;
w47571 <= not w47567 and w47570;
w47572 <= not w47515 and not w47571;
w47573 <= b(6) and not w47504;
w47574 <= not w47498 and w47573;
w47575 <= not w47506 and not w47574;
w47576 <= not w47572 and w47575;
w47577 <= not w47506 and not w47576;
w47578 <= b(7) and not w47495;
w47579 <= not w47489 and w47578;
w47580 <= not w47497 and not w47579;
w47581 <= not w47577 and w47580;
w47582 <= not w47497 and not w47581;
w47583 <= b(8) and not w47486;
w47584 <= not w47480 and w47583;
w47585 <= not w47488 and not w47584;
w47586 <= not w47582 and w47585;
w47587 <= not w47488 and not w47586;
w47588 <= b(9) and not w47477;
w47589 <= not w47471 and w47588;
w47590 <= not w47479 and not w47589;
w47591 <= not w47587 and w47590;
w47592 <= not w47479 and not w47591;
w47593 <= b(10) and not w47468;
w47594 <= not w47462 and w47593;
w47595 <= not w47470 and not w47594;
w47596 <= not w47592 and w47595;
w47597 <= not w47470 and not w47596;
w47598 <= b(11) and not w47459;
w47599 <= not w47453 and w47598;
w47600 <= not w47461 and not w47599;
w47601 <= not w47597 and w47600;
w47602 <= not w47461 and not w47601;
w47603 <= b(12) and not w47450;
w47604 <= not w47444 and w47603;
w47605 <= not w47452 and not w47604;
w47606 <= not w47602 and w47605;
w47607 <= not w47452 and not w47606;
w47608 <= b(13) and not w47441;
w47609 <= not w47435 and w47608;
w47610 <= not w47443 and not w47609;
w47611 <= not w47607 and w47610;
w47612 <= not w47443 and not w47611;
w47613 <= b(14) and not w47432;
w47614 <= not w47426 and w47613;
w47615 <= not w47434 and not w47614;
w47616 <= not w47612 and w47615;
w47617 <= not w47434 and not w47616;
w47618 <= b(15) and not w47423;
w47619 <= not w47417 and w47618;
w47620 <= not w47425 and not w47619;
w47621 <= not w47617 and w47620;
w47622 <= not w47425 and not w47621;
w47623 <= b(16) and not w47414;
w47624 <= not w47408 and w47623;
w47625 <= not w47416 and not w47624;
w47626 <= not w47622 and w47625;
w47627 <= not w47416 and not w47626;
w47628 <= b(17) and not w47405;
w47629 <= not w47399 and w47628;
w47630 <= not w47407 and not w47629;
w47631 <= not w47627 and w47630;
w47632 <= not w47407 and not w47631;
w47633 <= b(18) and not w47396;
w47634 <= not w47390 and w47633;
w47635 <= not w47398 and not w47634;
w47636 <= not w47632 and w47635;
w47637 <= not w47398 and not w47636;
w47638 <= b(19) and not w47387;
w47639 <= not w47381 and w47638;
w47640 <= not w47389 and not w47639;
w47641 <= not w47637 and w47640;
w47642 <= not w47389 and not w47641;
w47643 <= b(20) and not w47378;
w47644 <= not w47372 and w47643;
w47645 <= not w47380 and not w47644;
w47646 <= not w47642 and w47645;
w47647 <= not w47380 and not w47646;
w47648 <= b(21) and not w47369;
w47649 <= not w47363 and w47648;
w47650 <= not w47371 and not w47649;
w47651 <= not w47647 and w47650;
w47652 <= not w47371 and not w47651;
w47653 <= b(22) and not w47360;
w47654 <= not w47354 and w47653;
w47655 <= not w47362 and not w47654;
w47656 <= not w47652 and w47655;
w47657 <= not w47362 and not w47656;
w47658 <= b(23) and not w47351;
w47659 <= not w47345 and w47658;
w47660 <= not w47353 and not w47659;
w47661 <= not w47657 and w47660;
w47662 <= not w47353 and not w47661;
w47663 <= b(24) and not w47342;
w47664 <= not w47336 and w47663;
w47665 <= not w47344 and not w47664;
w47666 <= not w47662 and w47665;
w47667 <= not w47344 and not w47666;
w47668 <= b(25) and not w47333;
w47669 <= not w47327 and w47668;
w47670 <= not w47335 and not w47669;
w47671 <= not w47667 and w47670;
w47672 <= not w47335 and not w47671;
w47673 <= b(26) and not w47324;
w47674 <= not w47318 and w47673;
w47675 <= not w47326 and not w47674;
w47676 <= not w47672 and w47675;
w47677 <= not w47326 and not w47676;
w47678 <= b(27) and not w47315;
w47679 <= not w47309 and w47678;
w47680 <= not w47317 and not w47679;
w47681 <= not w47677 and w47680;
w47682 <= not w47317 and not w47681;
w47683 <= b(28) and not w47306;
w47684 <= not w47300 and w47683;
w47685 <= not w47308 and not w47684;
w47686 <= not w47682 and w47685;
w47687 <= not w47308 and not w47686;
w47688 <= b(29) and not w47297;
w47689 <= not w47291 and w47688;
w47690 <= not w47299 and not w47689;
w47691 <= not w47687 and w47690;
w47692 <= not w47299 and not w47691;
w47693 <= b(30) and not w47288;
w47694 <= not w47282 and w47693;
w47695 <= not w47290 and not w47694;
w47696 <= not w47692 and w47695;
w47697 <= not w47290 and not w47696;
w47698 <= b(31) and not w47279;
w47699 <= not w47273 and w47698;
w47700 <= not w47281 and not w47699;
w47701 <= not w47697 and w47700;
w47702 <= not w47281 and not w47701;
w47703 <= b(32) and not w47270;
w47704 <= not w47264 and w47703;
w47705 <= not w47272 and not w47704;
w47706 <= not w47702 and w47705;
w47707 <= not w47272 and not w47706;
w47708 <= b(33) and not w47261;
w47709 <= not w47255 and w47708;
w47710 <= not w47263 and not w47709;
w47711 <= not w47707 and w47710;
w47712 <= not w47263 and not w47711;
w47713 <= b(34) and not w47252;
w47714 <= not w47246 and w47713;
w47715 <= not w47254 and not w47714;
w47716 <= not w47712 and w47715;
w47717 <= not w47254 and not w47716;
w47718 <= b(35) and not w47243;
w47719 <= not w47237 and w47718;
w47720 <= not w47245 and not w47719;
w47721 <= not w47717 and w47720;
w47722 <= not w47245 and not w47721;
w47723 <= b(36) and not w47234;
w47724 <= not w47228 and w47723;
w47725 <= not w47236 and not w47724;
w47726 <= not w47722 and w47725;
w47727 <= not w47236 and not w47726;
w47728 <= b(37) and not w47225;
w47729 <= not w47219 and w47728;
w47730 <= not w47227 and not w47729;
w47731 <= not w47727 and w47730;
w47732 <= not w47227 and not w47731;
w47733 <= b(38) and not w47216;
w47734 <= not w47210 and w47733;
w47735 <= not w47218 and not w47734;
w47736 <= not w47732 and w47735;
w47737 <= not w47218 and not w47736;
w47738 <= b(39) and not w47207;
w47739 <= not w47201 and w47738;
w47740 <= not w47209 and not w47739;
w47741 <= not w47737 and w47740;
w47742 <= not w47209 and not w47741;
w47743 <= b(40) and not w47198;
w47744 <= not w47192 and w47743;
w47745 <= not w47200 and not w47744;
w47746 <= not w47742 and w47745;
w47747 <= not w47200 and not w47746;
w47748 <= b(41) and not w47189;
w47749 <= not w47183 and w47748;
w47750 <= not w47191 and not w47749;
w47751 <= not w47747 and w47750;
w47752 <= not w47191 and not w47751;
w47753 <= b(42) and not w47180;
w47754 <= not w47174 and w47753;
w47755 <= not w47182 and not w47754;
w47756 <= not w47752 and w47755;
w47757 <= not w47182 and not w47756;
w47758 <= b(43) and not w47171;
w47759 <= not w47165 and w47758;
w47760 <= not w47173 and not w47759;
w47761 <= not w47757 and w47760;
w47762 <= not w47173 and not w47761;
w47763 <= b(44) and not w47162;
w47764 <= not w47156 and w47763;
w47765 <= not w47164 and not w47764;
w47766 <= not w47762 and w47765;
w47767 <= not w47164 and not w47766;
w47768 <= b(45) and not w47153;
w47769 <= not w47147 and w47768;
w47770 <= not w47155 and not w47769;
w47771 <= not w47767 and w47770;
w47772 <= not w47155 and not w47771;
w47773 <= b(46) and not w47144;
w47774 <= not w47138 and w47773;
w47775 <= not w47146 and not w47774;
w47776 <= not w47772 and w47775;
w47777 <= not w47146 and not w47776;
w47778 <= b(47) and not w47135;
w47779 <= not w47129 and w47778;
w47780 <= not w47137 and not w47779;
w47781 <= not w47777 and w47780;
w47782 <= not w47137 and not w47781;
w47783 <= b(48) and not w47126;
w47784 <= not w47120 and w47783;
w47785 <= not w47128 and not w47784;
w47786 <= not w47782 and w47785;
w47787 <= not w47128 and not w47786;
w47788 <= b(49) and not w47117;
w47789 <= not w47111 and w47788;
w47790 <= not w47119 and not w47789;
w47791 <= not w47787 and w47790;
w47792 <= not w47119 and not w47791;
w47793 <= b(50) and not w47108;
w47794 <= not w47102 and w47793;
w47795 <= not w47110 and not w47794;
w47796 <= not w47792 and w47795;
w47797 <= not w47110 and not w47796;
w47798 <= b(51) and not w47099;
w47799 <= not w47093 and w47798;
w47800 <= not w47101 and not w47799;
w47801 <= not w47797 and w47800;
w47802 <= not w47101 and not w47801;
w47803 <= not w46397 and not w47092;
w47804 <= not w46399 and w47089;
w47805 <= not w47085 and w47804;
w47806 <= not w47086 and not w47089;
w47807 <= not w47805 and not w47806;
w47808 <= w47092 and not w47807;
w47809 <= not w47803 and not w47808;
w47810 <= not b(52) and not w47809;
w47811 <= b(52) and not w47803;
w47812 <= not w47808 and w47811;
w47813 <= w338 and not w47812;
w47814 <= not w47810 and w47813;
w47815 <= not w47802 and w47814;
w47816 <= w31 and not w47809;
w47817 <= not w47815 and not w47816;
w47818 <= not w47110 and w47800;
w47819 <= not w47796 and w47818;
w47820 <= not w47797 and not w47800;
w47821 <= not w47819 and not w47820;
w47822 <= not w47817 and not w47821;
w47823 <= not w47100 and not w47816;
w47824 <= not w47815 and w47823;
w47825 <= not w47822 and not w47824;
w47826 <= not b(52) and not w47825;
w47827 <= not w47119 and w47795;
w47828 <= not w47791 and w47827;
w47829 <= not w47792 and not w47795;
w47830 <= not w47828 and not w47829;
w47831 <= not w47817 and not w47830;
w47832 <= not w47109 and not w47816;
w47833 <= not w47815 and w47832;
w47834 <= not w47831 and not w47833;
w47835 <= not b(51) and not w47834;
w47836 <= not w47128 and w47790;
w47837 <= not w47786 and w47836;
w47838 <= not w47787 and not w47790;
w47839 <= not w47837 and not w47838;
w47840 <= not w47817 and not w47839;
w47841 <= not w47118 and not w47816;
w47842 <= not w47815 and w47841;
w47843 <= not w47840 and not w47842;
w47844 <= not b(50) and not w47843;
w47845 <= not w47137 and w47785;
w47846 <= not w47781 and w47845;
w47847 <= not w47782 and not w47785;
w47848 <= not w47846 and not w47847;
w47849 <= not w47817 and not w47848;
w47850 <= not w47127 and not w47816;
w47851 <= not w47815 and w47850;
w47852 <= not w47849 and not w47851;
w47853 <= not b(49) and not w47852;
w47854 <= not w47146 and w47780;
w47855 <= not w47776 and w47854;
w47856 <= not w47777 and not w47780;
w47857 <= not w47855 and not w47856;
w47858 <= not w47817 and not w47857;
w47859 <= not w47136 and not w47816;
w47860 <= not w47815 and w47859;
w47861 <= not w47858 and not w47860;
w47862 <= not b(48) and not w47861;
w47863 <= not w47155 and w47775;
w47864 <= not w47771 and w47863;
w47865 <= not w47772 and not w47775;
w47866 <= not w47864 and not w47865;
w47867 <= not w47817 and not w47866;
w47868 <= not w47145 and not w47816;
w47869 <= not w47815 and w47868;
w47870 <= not w47867 and not w47869;
w47871 <= not b(47) and not w47870;
w47872 <= not w47164 and w47770;
w47873 <= not w47766 and w47872;
w47874 <= not w47767 and not w47770;
w47875 <= not w47873 and not w47874;
w47876 <= not w47817 and not w47875;
w47877 <= not w47154 and not w47816;
w47878 <= not w47815 and w47877;
w47879 <= not w47876 and not w47878;
w47880 <= not b(46) and not w47879;
w47881 <= not w47173 and w47765;
w47882 <= not w47761 and w47881;
w47883 <= not w47762 and not w47765;
w47884 <= not w47882 and not w47883;
w47885 <= not w47817 and not w47884;
w47886 <= not w47163 and not w47816;
w47887 <= not w47815 and w47886;
w47888 <= not w47885 and not w47887;
w47889 <= not b(45) and not w47888;
w47890 <= not w47182 and w47760;
w47891 <= not w47756 and w47890;
w47892 <= not w47757 and not w47760;
w47893 <= not w47891 and not w47892;
w47894 <= not w47817 and not w47893;
w47895 <= not w47172 and not w47816;
w47896 <= not w47815 and w47895;
w47897 <= not w47894 and not w47896;
w47898 <= not b(44) and not w47897;
w47899 <= not w47191 and w47755;
w47900 <= not w47751 and w47899;
w47901 <= not w47752 and not w47755;
w47902 <= not w47900 and not w47901;
w47903 <= not w47817 and not w47902;
w47904 <= not w47181 and not w47816;
w47905 <= not w47815 and w47904;
w47906 <= not w47903 and not w47905;
w47907 <= not b(43) and not w47906;
w47908 <= not w47200 and w47750;
w47909 <= not w47746 and w47908;
w47910 <= not w47747 and not w47750;
w47911 <= not w47909 and not w47910;
w47912 <= not w47817 and not w47911;
w47913 <= not w47190 and not w47816;
w47914 <= not w47815 and w47913;
w47915 <= not w47912 and not w47914;
w47916 <= not b(42) and not w47915;
w47917 <= not w47209 and w47745;
w47918 <= not w47741 and w47917;
w47919 <= not w47742 and not w47745;
w47920 <= not w47918 and not w47919;
w47921 <= not w47817 and not w47920;
w47922 <= not w47199 and not w47816;
w47923 <= not w47815 and w47922;
w47924 <= not w47921 and not w47923;
w47925 <= not b(41) and not w47924;
w47926 <= not w47218 and w47740;
w47927 <= not w47736 and w47926;
w47928 <= not w47737 and not w47740;
w47929 <= not w47927 and not w47928;
w47930 <= not w47817 and not w47929;
w47931 <= not w47208 and not w47816;
w47932 <= not w47815 and w47931;
w47933 <= not w47930 and not w47932;
w47934 <= not b(40) and not w47933;
w47935 <= not w47227 and w47735;
w47936 <= not w47731 and w47935;
w47937 <= not w47732 and not w47735;
w47938 <= not w47936 and not w47937;
w47939 <= not w47817 and not w47938;
w47940 <= not w47217 and not w47816;
w47941 <= not w47815 and w47940;
w47942 <= not w47939 and not w47941;
w47943 <= not b(39) and not w47942;
w47944 <= not w47236 and w47730;
w47945 <= not w47726 and w47944;
w47946 <= not w47727 and not w47730;
w47947 <= not w47945 and not w47946;
w47948 <= not w47817 and not w47947;
w47949 <= not w47226 and not w47816;
w47950 <= not w47815 and w47949;
w47951 <= not w47948 and not w47950;
w47952 <= not b(38) and not w47951;
w47953 <= not w47245 and w47725;
w47954 <= not w47721 and w47953;
w47955 <= not w47722 and not w47725;
w47956 <= not w47954 and not w47955;
w47957 <= not w47817 and not w47956;
w47958 <= not w47235 and not w47816;
w47959 <= not w47815 and w47958;
w47960 <= not w47957 and not w47959;
w47961 <= not b(37) and not w47960;
w47962 <= not w47254 and w47720;
w47963 <= not w47716 and w47962;
w47964 <= not w47717 and not w47720;
w47965 <= not w47963 and not w47964;
w47966 <= not w47817 and not w47965;
w47967 <= not w47244 and not w47816;
w47968 <= not w47815 and w47967;
w47969 <= not w47966 and not w47968;
w47970 <= not b(36) and not w47969;
w47971 <= not w47263 and w47715;
w47972 <= not w47711 and w47971;
w47973 <= not w47712 and not w47715;
w47974 <= not w47972 and not w47973;
w47975 <= not w47817 and not w47974;
w47976 <= not w47253 and not w47816;
w47977 <= not w47815 and w47976;
w47978 <= not w47975 and not w47977;
w47979 <= not b(35) and not w47978;
w47980 <= not w47272 and w47710;
w47981 <= not w47706 and w47980;
w47982 <= not w47707 and not w47710;
w47983 <= not w47981 and not w47982;
w47984 <= not w47817 and not w47983;
w47985 <= not w47262 and not w47816;
w47986 <= not w47815 and w47985;
w47987 <= not w47984 and not w47986;
w47988 <= not b(34) and not w47987;
w47989 <= not w47281 and w47705;
w47990 <= not w47701 and w47989;
w47991 <= not w47702 and not w47705;
w47992 <= not w47990 and not w47991;
w47993 <= not w47817 and not w47992;
w47994 <= not w47271 and not w47816;
w47995 <= not w47815 and w47994;
w47996 <= not w47993 and not w47995;
w47997 <= not b(33) and not w47996;
w47998 <= not w47290 and w47700;
w47999 <= not w47696 and w47998;
w48000 <= not w47697 and not w47700;
w48001 <= not w47999 and not w48000;
w48002 <= not w47817 and not w48001;
w48003 <= not w47280 and not w47816;
w48004 <= not w47815 and w48003;
w48005 <= not w48002 and not w48004;
w48006 <= not b(32) and not w48005;
w48007 <= not w47299 and w47695;
w48008 <= not w47691 and w48007;
w48009 <= not w47692 and not w47695;
w48010 <= not w48008 and not w48009;
w48011 <= not w47817 and not w48010;
w48012 <= not w47289 and not w47816;
w48013 <= not w47815 and w48012;
w48014 <= not w48011 and not w48013;
w48015 <= not b(31) and not w48014;
w48016 <= not w47308 and w47690;
w48017 <= not w47686 and w48016;
w48018 <= not w47687 and not w47690;
w48019 <= not w48017 and not w48018;
w48020 <= not w47817 and not w48019;
w48021 <= not w47298 and not w47816;
w48022 <= not w47815 and w48021;
w48023 <= not w48020 and not w48022;
w48024 <= not b(30) and not w48023;
w48025 <= not w47317 and w47685;
w48026 <= not w47681 and w48025;
w48027 <= not w47682 and not w47685;
w48028 <= not w48026 and not w48027;
w48029 <= not w47817 and not w48028;
w48030 <= not w47307 and not w47816;
w48031 <= not w47815 and w48030;
w48032 <= not w48029 and not w48031;
w48033 <= not b(29) and not w48032;
w48034 <= not w47326 and w47680;
w48035 <= not w47676 and w48034;
w48036 <= not w47677 and not w47680;
w48037 <= not w48035 and not w48036;
w48038 <= not w47817 and not w48037;
w48039 <= not w47316 and not w47816;
w48040 <= not w47815 and w48039;
w48041 <= not w48038 and not w48040;
w48042 <= not b(28) and not w48041;
w48043 <= not w47335 and w47675;
w48044 <= not w47671 and w48043;
w48045 <= not w47672 and not w47675;
w48046 <= not w48044 and not w48045;
w48047 <= not w47817 and not w48046;
w48048 <= not w47325 and not w47816;
w48049 <= not w47815 and w48048;
w48050 <= not w48047 and not w48049;
w48051 <= not b(27) and not w48050;
w48052 <= not w47344 and w47670;
w48053 <= not w47666 and w48052;
w48054 <= not w47667 and not w47670;
w48055 <= not w48053 and not w48054;
w48056 <= not w47817 and not w48055;
w48057 <= not w47334 and not w47816;
w48058 <= not w47815 and w48057;
w48059 <= not w48056 and not w48058;
w48060 <= not b(26) and not w48059;
w48061 <= not w47353 and w47665;
w48062 <= not w47661 and w48061;
w48063 <= not w47662 and not w47665;
w48064 <= not w48062 and not w48063;
w48065 <= not w47817 and not w48064;
w48066 <= not w47343 and not w47816;
w48067 <= not w47815 and w48066;
w48068 <= not w48065 and not w48067;
w48069 <= not b(25) and not w48068;
w48070 <= not w47362 and w47660;
w48071 <= not w47656 and w48070;
w48072 <= not w47657 and not w47660;
w48073 <= not w48071 and not w48072;
w48074 <= not w47817 and not w48073;
w48075 <= not w47352 and not w47816;
w48076 <= not w47815 and w48075;
w48077 <= not w48074 and not w48076;
w48078 <= not b(24) and not w48077;
w48079 <= not w47371 and w47655;
w48080 <= not w47651 and w48079;
w48081 <= not w47652 and not w47655;
w48082 <= not w48080 and not w48081;
w48083 <= not w47817 and not w48082;
w48084 <= not w47361 and not w47816;
w48085 <= not w47815 and w48084;
w48086 <= not w48083 and not w48085;
w48087 <= not b(23) and not w48086;
w48088 <= not w47380 and w47650;
w48089 <= not w47646 and w48088;
w48090 <= not w47647 and not w47650;
w48091 <= not w48089 and not w48090;
w48092 <= not w47817 and not w48091;
w48093 <= not w47370 and not w47816;
w48094 <= not w47815 and w48093;
w48095 <= not w48092 and not w48094;
w48096 <= not b(22) and not w48095;
w48097 <= not w47389 and w47645;
w48098 <= not w47641 and w48097;
w48099 <= not w47642 and not w47645;
w48100 <= not w48098 and not w48099;
w48101 <= not w47817 and not w48100;
w48102 <= not w47379 and not w47816;
w48103 <= not w47815 and w48102;
w48104 <= not w48101 and not w48103;
w48105 <= not b(21) and not w48104;
w48106 <= not w47398 and w47640;
w48107 <= not w47636 and w48106;
w48108 <= not w47637 and not w47640;
w48109 <= not w48107 and not w48108;
w48110 <= not w47817 and not w48109;
w48111 <= not w47388 and not w47816;
w48112 <= not w47815 and w48111;
w48113 <= not w48110 and not w48112;
w48114 <= not b(20) and not w48113;
w48115 <= not w47407 and w47635;
w48116 <= not w47631 and w48115;
w48117 <= not w47632 and not w47635;
w48118 <= not w48116 and not w48117;
w48119 <= not w47817 and not w48118;
w48120 <= not w47397 and not w47816;
w48121 <= not w47815 and w48120;
w48122 <= not w48119 and not w48121;
w48123 <= not b(19) and not w48122;
w48124 <= not w47416 and w47630;
w48125 <= not w47626 and w48124;
w48126 <= not w47627 and not w47630;
w48127 <= not w48125 and not w48126;
w48128 <= not w47817 and not w48127;
w48129 <= not w47406 and not w47816;
w48130 <= not w47815 and w48129;
w48131 <= not w48128 and not w48130;
w48132 <= not b(18) and not w48131;
w48133 <= not w47425 and w47625;
w48134 <= not w47621 and w48133;
w48135 <= not w47622 and not w47625;
w48136 <= not w48134 and not w48135;
w48137 <= not w47817 and not w48136;
w48138 <= not w47415 and not w47816;
w48139 <= not w47815 and w48138;
w48140 <= not w48137 and not w48139;
w48141 <= not b(17) and not w48140;
w48142 <= not w47434 and w47620;
w48143 <= not w47616 and w48142;
w48144 <= not w47617 and not w47620;
w48145 <= not w48143 and not w48144;
w48146 <= not w47817 and not w48145;
w48147 <= not w47424 and not w47816;
w48148 <= not w47815 and w48147;
w48149 <= not w48146 and not w48148;
w48150 <= not b(16) and not w48149;
w48151 <= not w47443 and w47615;
w48152 <= not w47611 and w48151;
w48153 <= not w47612 and not w47615;
w48154 <= not w48152 and not w48153;
w48155 <= not w47817 and not w48154;
w48156 <= not w47433 and not w47816;
w48157 <= not w47815 and w48156;
w48158 <= not w48155 and not w48157;
w48159 <= not b(15) and not w48158;
w48160 <= not w47452 and w47610;
w48161 <= not w47606 and w48160;
w48162 <= not w47607 and not w47610;
w48163 <= not w48161 and not w48162;
w48164 <= not w47817 and not w48163;
w48165 <= not w47442 and not w47816;
w48166 <= not w47815 and w48165;
w48167 <= not w48164 and not w48166;
w48168 <= not b(14) and not w48167;
w48169 <= not w47461 and w47605;
w48170 <= not w47601 and w48169;
w48171 <= not w47602 and not w47605;
w48172 <= not w48170 and not w48171;
w48173 <= not w47817 and not w48172;
w48174 <= not w47451 and not w47816;
w48175 <= not w47815 and w48174;
w48176 <= not w48173 and not w48175;
w48177 <= not b(13) and not w48176;
w48178 <= not w47470 and w47600;
w48179 <= not w47596 and w48178;
w48180 <= not w47597 and not w47600;
w48181 <= not w48179 and not w48180;
w48182 <= not w47817 and not w48181;
w48183 <= not w47460 and not w47816;
w48184 <= not w47815 and w48183;
w48185 <= not w48182 and not w48184;
w48186 <= not b(12) and not w48185;
w48187 <= not w47479 and w47595;
w48188 <= not w47591 and w48187;
w48189 <= not w47592 and not w47595;
w48190 <= not w48188 and not w48189;
w48191 <= not w47817 and not w48190;
w48192 <= not w47469 and not w47816;
w48193 <= not w47815 and w48192;
w48194 <= not w48191 and not w48193;
w48195 <= not b(11) and not w48194;
w48196 <= not w47488 and w47590;
w48197 <= not w47586 and w48196;
w48198 <= not w47587 and not w47590;
w48199 <= not w48197 and not w48198;
w48200 <= not w47817 and not w48199;
w48201 <= not w47478 and not w47816;
w48202 <= not w47815 and w48201;
w48203 <= not w48200 and not w48202;
w48204 <= not b(10) and not w48203;
w48205 <= not w47497 and w47585;
w48206 <= not w47581 and w48205;
w48207 <= not w47582 and not w47585;
w48208 <= not w48206 and not w48207;
w48209 <= not w47817 and not w48208;
w48210 <= not w47487 and not w47816;
w48211 <= not w47815 and w48210;
w48212 <= not w48209 and not w48211;
w48213 <= not b(9) and not w48212;
w48214 <= not w47506 and w47580;
w48215 <= not w47576 and w48214;
w48216 <= not w47577 and not w47580;
w48217 <= not w48215 and not w48216;
w48218 <= not w47817 and not w48217;
w48219 <= not w47496 and not w47816;
w48220 <= not w47815 and w48219;
w48221 <= not w48218 and not w48220;
w48222 <= not b(8) and not w48221;
w48223 <= not w47515 and w47575;
w48224 <= not w47571 and w48223;
w48225 <= not w47572 and not w47575;
w48226 <= not w48224 and not w48225;
w48227 <= not w47817 and not w48226;
w48228 <= not w47505 and not w47816;
w48229 <= not w47815 and w48228;
w48230 <= not w48227 and not w48229;
w48231 <= not b(7) and not w48230;
w48232 <= not w47524 and w47570;
w48233 <= not w47566 and w48232;
w48234 <= not w47567 and not w47570;
w48235 <= not w48233 and not w48234;
w48236 <= not w47817 and not w48235;
w48237 <= not w47514 and not w47816;
w48238 <= not w47815 and w48237;
w48239 <= not w48236 and not w48238;
w48240 <= not b(6) and not w48239;
w48241 <= not w47533 and w47565;
w48242 <= not w47561 and w48241;
w48243 <= not w47562 and not w47565;
w48244 <= not w48242 and not w48243;
w48245 <= not w47817 and not w48244;
w48246 <= not w47523 and not w47816;
w48247 <= not w47815 and w48246;
w48248 <= not w48245 and not w48247;
w48249 <= not b(5) and not w48248;
w48250 <= not w47541 and w47560;
w48251 <= not w47556 and w48250;
w48252 <= not w47557 and not w47560;
w48253 <= not w48251 and not w48252;
w48254 <= not w47817 and not w48253;
w48255 <= not w47532 and not w47816;
w48256 <= not w47815 and w48255;
w48257 <= not w48254 and not w48256;
w48258 <= not b(4) and not w48257;
w48259 <= not w47551 and w47555;
w48260 <= not w47550 and w48259;
w48261 <= not w47552 and not w47555;
w48262 <= not w48260 and not w48261;
w48263 <= not w47817 and not w48262;
w48264 <= not w47540 and not w47816;
w48265 <= not w47815 and w48264;
w48266 <= not w48263 and not w48265;
w48267 <= not b(3) and not w48266;
w48268 <= w19510 and not w47548;
w48269 <= not w47546 and w48268;
w48270 <= not w47550 and not w48269;
w48271 <= not w47817 and w48270;
w48272 <= not w47545 and not w47816;
w48273 <= not w47815 and w48272;
w48274 <= not w48271 and not w48273;
w48275 <= not b(2) and not w48274;
w48276 <= b(0) and not w47817;
w48277 <= a(11) and not w48276;
w48278 <= w19510 and not w47817;
w48279 <= not w48277 and not w48278;
w48280 <= b(1) and not w48279;
w48281 <= not b(1) and not w48278;
w48282 <= not w48277 and w48281;
w48283 <= not w48280 and not w48282;
w48284 <= not w20245 and not w48283;
w48285 <= not b(1) and not w48279;
w48286 <= not w48284 and not w48285;
w48287 <= b(2) and not w48273;
w48288 <= not w48271 and w48287;
w48289 <= not w48275 and not w48288;
w48290 <= not w48286 and w48289;
w48291 <= not w48275 and not w48290;
w48292 <= b(3) and not w48265;
w48293 <= not w48263 and w48292;
w48294 <= not w48267 and not w48293;
w48295 <= not w48291 and w48294;
w48296 <= not w48267 and not w48295;
w48297 <= b(4) and not w48256;
w48298 <= not w48254 and w48297;
w48299 <= not w48258 and not w48298;
w48300 <= not w48296 and w48299;
w48301 <= not w48258 and not w48300;
w48302 <= b(5) and not w48247;
w48303 <= not w48245 and w48302;
w48304 <= not w48249 and not w48303;
w48305 <= not w48301 and w48304;
w48306 <= not w48249 and not w48305;
w48307 <= b(6) and not w48238;
w48308 <= not w48236 and w48307;
w48309 <= not w48240 and not w48308;
w48310 <= not w48306 and w48309;
w48311 <= not w48240 and not w48310;
w48312 <= b(7) and not w48229;
w48313 <= not w48227 and w48312;
w48314 <= not w48231 and not w48313;
w48315 <= not w48311 and w48314;
w48316 <= not w48231 and not w48315;
w48317 <= b(8) and not w48220;
w48318 <= not w48218 and w48317;
w48319 <= not w48222 and not w48318;
w48320 <= not w48316 and w48319;
w48321 <= not w48222 and not w48320;
w48322 <= b(9) and not w48211;
w48323 <= not w48209 and w48322;
w48324 <= not w48213 and not w48323;
w48325 <= not w48321 and w48324;
w48326 <= not w48213 and not w48325;
w48327 <= b(10) and not w48202;
w48328 <= not w48200 and w48327;
w48329 <= not w48204 and not w48328;
w48330 <= not w48326 and w48329;
w48331 <= not w48204 and not w48330;
w48332 <= b(11) and not w48193;
w48333 <= not w48191 and w48332;
w48334 <= not w48195 and not w48333;
w48335 <= not w48331 and w48334;
w48336 <= not w48195 and not w48335;
w48337 <= b(12) and not w48184;
w48338 <= not w48182 and w48337;
w48339 <= not w48186 and not w48338;
w48340 <= not w48336 and w48339;
w48341 <= not w48186 and not w48340;
w48342 <= b(13) and not w48175;
w48343 <= not w48173 and w48342;
w48344 <= not w48177 and not w48343;
w48345 <= not w48341 and w48344;
w48346 <= not w48177 and not w48345;
w48347 <= b(14) and not w48166;
w48348 <= not w48164 and w48347;
w48349 <= not w48168 and not w48348;
w48350 <= not w48346 and w48349;
w48351 <= not w48168 and not w48350;
w48352 <= b(15) and not w48157;
w48353 <= not w48155 and w48352;
w48354 <= not w48159 and not w48353;
w48355 <= not w48351 and w48354;
w48356 <= not w48159 and not w48355;
w48357 <= b(16) and not w48148;
w48358 <= not w48146 and w48357;
w48359 <= not w48150 and not w48358;
w48360 <= not w48356 and w48359;
w48361 <= not w48150 and not w48360;
w48362 <= b(17) and not w48139;
w48363 <= not w48137 and w48362;
w48364 <= not w48141 and not w48363;
w48365 <= not w48361 and w48364;
w48366 <= not w48141 and not w48365;
w48367 <= b(18) and not w48130;
w48368 <= not w48128 and w48367;
w48369 <= not w48132 and not w48368;
w48370 <= not w48366 and w48369;
w48371 <= not w48132 and not w48370;
w48372 <= b(19) and not w48121;
w48373 <= not w48119 and w48372;
w48374 <= not w48123 and not w48373;
w48375 <= not w48371 and w48374;
w48376 <= not w48123 and not w48375;
w48377 <= b(20) and not w48112;
w48378 <= not w48110 and w48377;
w48379 <= not w48114 and not w48378;
w48380 <= not w48376 and w48379;
w48381 <= not w48114 and not w48380;
w48382 <= b(21) and not w48103;
w48383 <= not w48101 and w48382;
w48384 <= not w48105 and not w48383;
w48385 <= not w48381 and w48384;
w48386 <= not w48105 and not w48385;
w48387 <= b(22) and not w48094;
w48388 <= not w48092 and w48387;
w48389 <= not w48096 and not w48388;
w48390 <= not w48386 and w48389;
w48391 <= not w48096 and not w48390;
w48392 <= b(23) and not w48085;
w48393 <= not w48083 and w48392;
w48394 <= not w48087 and not w48393;
w48395 <= not w48391 and w48394;
w48396 <= not w48087 and not w48395;
w48397 <= b(24) and not w48076;
w48398 <= not w48074 and w48397;
w48399 <= not w48078 and not w48398;
w48400 <= not w48396 and w48399;
w48401 <= not w48078 and not w48400;
w48402 <= b(25) and not w48067;
w48403 <= not w48065 and w48402;
w48404 <= not w48069 and not w48403;
w48405 <= not w48401 and w48404;
w48406 <= not w48069 and not w48405;
w48407 <= b(26) and not w48058;
w48408 <= not w48056 and w48407;
w48409 <= not w48060 and not w48408;
w48410 <= not w48406 and w48409;
w48411 <= not w48060 and not w48410;
w48412 <= b(27) and not w48049;
w48413 <= not w48047 and w48412;
w48414 <= not w48051 and not w48413;
w48415 <= not w48411 and w48414;
w48416 <= not w48051 and not w48415;
w48417 <= b(28) and not w48040;
w48418 <= not w48038 and w48417;
w48419 <= not w48042 and not w48418;
w48420 <= not w48416 and w48419;
w48421 <= not w48042 and not w48420;
w48422 <= b(29) and not w48031;
w48423 <= not w48029 and w48422;
w48424 <= not w48033 and not w48423;
w48425 <= not w48421 and w48424;
w48426 <= not w48033 and not w48425;
w48427 <= b(30) and not w48022;
w48428 <= not w48020 and w48427;
w48429 <= not w48024 and not w48428;
w48430 <= not w48426 and w48429;
w48431 <= not w48024 and not w48430;
w48432 <= b(31) and not w48013;
w48433 <= not w48011 and w48432;
w48434 <= not w48015 and not w48433;
w48435 <= not w48431 and w48434;
w48436 <= not w48015 and not w48435;
w48437 <= b(32) and not w48004;
w48438 <= not w48002 and w48437;
w48439 <= not w48006 and not w48438;
w48440 <= not w48436 and w48439;
w48441 <= not w48006 and not w48440;
w48442 <= b(33) and not w47995;
w48443 <= not w47993 and w48442;
w48444 <= not w47997 and not w48443;
w48445 <= not w48441 and w48444;
w48446 <= not w47997 and not w48445;
w48447 <= b(34) and not w47986;
w48448 <= not w47984 and w48447;
w48449 <= not w47988 and not w48448;
w48450 <= not w48446 and w48449;
w48451 <= not w47988 and not w48450;
w48452 <= b(35) and not w47977;
w48453 <= not w47975 and w48452;
w48454 <= not w47979 and not w48453;
w48455 <= not w48451 and w48454;
w48456 <= not w47979 and not w48455;
w48457 <= b(36) and not w47968;
w48458 <= not w47966 and w48457;
w48459 <= not w47970 and not w48458;
w48460 <= not w48456 and w48459;
w48461 <= not w47970 and not w48460;
w48462 <= b(37) and not w47959;
w48463 <= not w47957 and w48462;
w48464 <= not w47961 and not w48463;
w48465 <= not w48461 and w48464;
w48466 <= not w47961 and not w48465;
w48467 <= b(38) and not w47950;
w48468 <= not w47948 and w48467;
w48469 <= not w47952 and not w48468;
w48470 <= not w48466 and w48469;
w48471 <= not w47952 and not w48470;
w48472 <= b(39) and not w47941;
w48473 <= not w47939 and w48472;
w48474 <= not w47943 and not w48473;
w48475 <= not w48471 and w48474;
w48476 <= not w47943 and not w48475;
w48477 <= b(40) and not w47932;
w48478 <= not w47930 and w48477;
w48479 <= not w47934 and not w48478;
w48480 <= not w48476 and w48479;
w48481 <= not w47934 and not w48480;
w48482 <= b(41) and not w47923;
w48483 <= not w47921 and w48482;
w48484 <= not w47925 and not w48483;
w48485 <= not w48481 and w48484;
w48486 <= not w47925 and not w48485;
w48487 <= b(42) and not w47914;
w48488 <= not w47912 and w48487;
w48489 <= not w47916 and not w48488;
w48490 <= not w48486 and w48489;
w48491 <= not w47916 and not w48490;
w48492 <= b(43) and not w47905;
w48493 <= not w47903 and w48492;
w48494 <= not w47907 and not w48493;
w48495 <= not w48491 and w48494;
w48496 <= not w47907 and not w48495;
w48497 <= b(44) and not w47896;
w48498 <= not w47894 and w48497;
w48499 <= not w47898 and not w48498;
w48500 <= not w48496 and w48499;
w48501 <= not w47898 and not w48500;
w48502 <= b(45) and not w47887;
w48503 <= not w47885 and w48502;
w48504 <= not w47889 and not w48503;
w48505 <= not w48501 and w48504;
w48506 <= not w47889 and not w48505;
w48507 <= b(46) and not w47878;
w48508 <= not w47876 and w48507;
w48509 <= not w47880 and not w48508;
w48510 <= not w48506 and w48509;
w48511 <= not w47880 and not w48510;
w48512 <= b(47) and not w47869;
w48513 <= not w47867 and w48512;
w48514 <= not w47871 and not w48513;
w48515 <= not w48511 and w48514;
w48516 <= not w47871 and not w48515;
w48517 <= b(48) and not w47860;
w48518 <= not w47858 and w48517;
w48519 <= not w47862 and not w48518;
w48520 <= not w48516 and w48519;
w48521 <= not w47862 and not w48520;
w48522 <= b(49) and not w47851;
w48523 <= not w47849 and w48522;
w48524 <= not w47853 and not w48523;
w48525 <= not w48521 and w48524;
w48526 <= not w47853 and not w48525;
w48527 <= b(50) and not w47842;
w48528 <= not w47840 and w48527;
w48529 <= not w47844 and not w48528;
w48530 <= not w48526 and w48529;
w48531 <= not w47844 and not w48530;
w48532 <= b(51) and not w47833;
w48533 <= not w47831 and w48532;
w48534 <= not w47835 and not w48533;
w48535 <= not w48531 and w48534;
w48536 <= not w47835 and not w48535;
w48537 <= b(52) and not w47824;
w48538 <= not w47822 and w48537;
w48539 <= not w47826 and not w48538;
w48540 <= not w48536 and w48539;
w48541 <= not w47826 and not w48540;
w48542 <= not w47101 and not w47812;
w48543 <= not w47810 and w48542;
w48544 <= not w47801 and w48543;
w48545 <= not w47810 and not w47812;
w48546 <= not w47802 and not w48545;
w48547 <= not w48544 and not w48546;
w48548 <= not w47817 and not w48547;
w48549 <= not w47809 and not w47816;
w48550 <= not w47815 and w48549;
w48551 <= not w48548 and not w48550;
w48552 <= not b(53) and not w48551;
w48553 <= b(53) and not w48550;
w48554 <= not w48548 and w48553;
w48555 <= w20518 and not w48554;
w48556 <= not w48552 and w48555;
w48557 <= not w48541 and w48556;
w48558 <= w338 and not w48551;
w48559 <= not w48557 and not w48558;
w48560 <= not w47835 and w48539;
w48561 <= not w48535 and w48560;
w48562 <= not w48536 and not w48539;
w48563 <= not w48561 and not w48562;
w48564 <= not w48559 and not w48563;
w48565 <= not w47825 and not w48558;
w48566 <= not w48557 and w48565;
w48567 <= not w48564 and not w48566;
w48568 <= not w47826 and not w48554;
w48569 <= not w48552 and w48568;
w48570 <= not w48540 and w48569;
w48571 <= not w48552 and not w48554;
w48572 <= not w48541 and not w48571;
w48573 <= not w48570 and not w48572;
w48574 <= not w48559 and not w48573;
w48575 <= not w48551 and not w48558;
w48576 <= not w48557 and w48575;
w48577 <= not w48574 and not w48576;
w48578 <= not b(54) and not w48577;
w48579 <= not b(53) and not w48567;
w48580 <= not w47844 and w48534;
w48581 <= not w48530 and w48580;
w48582 <= not w48531 and not w48534;
w48583 <= not w48581 and not w48582;
w48584 <= not w48559 and not w48583;
w48585 <= not w47834 and not w48558;
w48586 <= not w48557 and w48585;
w48587 <= not w48584 and not w48586;
w48588 <= not b(52) and not w48587;
w48589 <= not w47853 and w48529;
w48590 <= not w48525 and w48589;
w48591 <= not w48526 and not w48529;
w48592 <= not w48590 and not w48591;
w48593 <= not w48559 and not w48592;
w48594 <= not w47843 and not w48558;
w48595 <= not w48557 and w48594;
w48596 <= not w48593 and not w48595;
w48597 <= not b(51) and not w48596;
w48598 <= not w47862 and w48524;
w48599 <= not w48520 and w48598;
w48600 <= not w48521 and not w48524;
w48601 <= not w48599 and not w48600;
w48602 <= not w48559 and not w48601;
w48603 <= not w47852 and not w48558;
w48604 <= not w48557 and w48603;
w48605 <= not w48602 and not w48604;
w48606 <= not b(50) and not w48605;
w48607 <= not w47871 and w48519;
w48608 <= not w48515 and w48607;
w48609 <= not w48516 and not w48519;
w48610 <= not w48608 and not w48609;
w48611 <= not w48559 and not w48610;
w48612 <= not w47861 and not w48558;
w48613 <= not w48557 and w48612;
w48614 <= not w48611 and not w48613;
w48615 <= not b(49) and not w48614;
w48616 <= not w47880 and w48514;
w48617 <= not w48510 and w48616;
w48618 <= not w48511 and not w48514;
w48619 <= not w48617 and not w48618;
w48620 <= not w48559 and not w48619;
w48621 <= not w47870 and not w48558;
w48622 <= not w48557 and w48621;
w48623 <= not w48620 and not w48622;
w48624 <= not b(48) and not w48623;
w48625 <= not w47889 and w48509;
w48626 <= not w48505 and w48625;
w48627 <= not w48506 and not w48509;
w48628 <= not w48626 and not w48627;
w48629 <= not w48559 and not w48628;
w48630 <= not w47879 and not w48558;
w48631 <= not w48557 and w48630;
w48632 <= not w48629 and not w48631;
w48633 <= not b(47) and not w48632;
w48634 <= not w47898 and w48504;
w48635 <= not w48500 and w48634;
w48636 <= not w48501 and not w48504;
w48637 <= not w48635 and not w48636;
w48638 <= not w48559 and not w48637;
w48639 <= not w47888 and not w48558;
w48640 <= not w48557 and w48639;
w48641 <= not w48638 and not w48640;
w48642 <= not b(46) and not w48641;
w48643 <= not w47907 and w48499;
w48644 <= not w48495 and w48643;
w48645 <= not w48496 and not w48499;
w48646 <= not w48644 and not w48645;
w48647 <= not w48559 and not w48646;
w48648 <= not w47897 and not w48558;
w48649 <= not w48557 and w48648;
w48650 <= not w48647 and not w48649;
w48651 <= not b(45) and not w48650;
w48652 <= not w47916 and w48494;
w48653 <= not w48490 and w48652;
w48654 <= not w48491 and not w48494;
w48655 <= not w48653 and not w48654;
w48656 <= not w48559 and not w48655;
w48657 <= not w47906 and not w48558;
w48658 <= not w48557 and w48657;
w48659 <= not w48656 and not w48658;
w48660 <= not b(44) and not w48659;
w48661 <= not w47925 and w48489;
w48662 <= not w48485 and w48661;
w48663 <= not w48486 and not w48489;
w48664 <= not w48662 and not w48663;
w48665 <= not w48559 and not w48664;
w48666 <= not w47915 and not w48558;
w48667 <= not w48557 and w48666;
w48668 <= not w48665 and not w48667;
w48669 <= not b(43) and not w48668;
w48670 <= not w47934 and w48484;
w48671 <= not w48480 and w48670;
w48672 <= not w48481 and not w48484;
w48673 <= not w48671 and not w48672;
w48674 <= not w48559 and not w48673;
w48675 <= not w47924 and not w48558;
w48676 <= not w48557 and w48675;
w48677 <= not w48674 and not w48676;
w48678 <= not b(42) and not w48677;
w48679 <= not w47943 and w48479;
w48680 <= not w48475 and w48679;
w48681 <= not w48476 and not w48479;
w48682 <= not w48680 and not w48681;
w48683 <= not w48559 and not w48682;
w48684 <= not w47933 and not w48558;
w48685 <= not w48557 and w48684;
w48686 <= not w48683 and not w48685;
w48687 <= not b(41) and not w48686;
w48688 <= not w47952 and w48474;
w48689 <= not w48470 and w48688;
w48690 <= not w48471 and not w48474;
w48691 <= not w48689 and not w48690;
w48692 <= not w48559 and not w48691;
w48693 <= not w47942 and not w48558;
w48694 <= not w48557 and w48693;
w48695 <= not w48692 and not w48694;
w48696 <= not b(40) and not w48695;
w48697 <= not w47961 and w48469;
w48698 <= not w48465 and w48697;
w48699 <= not w48466 and not w48469;
w48700 <= not w48698 and not w48699;
w48701 <= not w48559 and not w48700;
w48702 <= not w47951 and not w48558;
w48703 <= not w48557 and w48702;
w48704 <= not w48701 and not w48703;
w48705 <= not b(39) and not w48704;
w48706 <= not w47970 and w48464;
w48707 <= not w48460 and w48706;
w48708 <= not w48461 and not w48464;
w48709 <= not w48707 and not w48708;
w48710 <= not w48559 and not w48709;
w48711 <= not w47960 and not w48558;
w48712 <= not w48557 and w48711;
w48713 <= not w48710 and not w48712;
w48714 <= not b(38) and not w48713;
w48715 <= not w47979 and w48459;
w48716 <= not w48455 and w48715;
w48717 <= not w48456 and not w48459;
w48718 <= not w48716 and not w48717;
w48719 <= not w48559 and not w48718;
w48720 <= not w47969 and not w48558;
w48721 <= not w48557 and w48720;
w48722 <= not w48719 and not w48721;
w48723 <= not b(37) and not w48722;
w48724 <= not w47988 and w48454;
w48725 <= not w48450 and w48724;
w48726 <= not w48451 and not w48454;
w48727 <= not w48725 and not w48726;
w48728 <= not w48559 and not w48727;
w48729 <= not w47978 and not w48558;
w48730 <= not w48557 and w48729;
w48731 <= not w48728 and not w48730;
w48732 <= not b(36) and not w48731;
w48733 <= not w47997 and w48449;
w48734 <= not w48445 and w48733;
w48735 <= not w48446 and not w48449;
w48736 <= not w48734 and not w48735;
w48737 <= not w48559 and not w48736;
w48738 <= not w47987 and not w48558;
w48739 <= not w48557 and w48738;
w48740 <= not w48737 and not w48739;
w48741 <= not b(35) and not w48740;
w48742 <= not w48006 and w48444;
w48743 <= not w48440 and w48742;
w48744 <= not w48441 and not w48444;
w48745 <= not w48743 and not w48744;
w48746 <= not w48559 and not w48745;
w48747 <= not w47996 and not w48558;
w48748 <= not w48557 and w48747;
w48749 <= not w48746 and not w48748;
w48750 <= not b(34) and not w48749;
w48751 <= not w48015 and w48439;
w48752 <= not w48435 and w48751;
w48753 <= not w48436 and not w48439;
w48754 <= not w48752 and not w48753;
w48755 <= not w48559 and not w48754;
w48756 <= not w48005 and not w48558;
w48757 <= not w48557 and w48756;
w48758 <= not w48755 and not w48757;
w48759 <= not b(33) and not w48758;
w48760 <= not w48024 and w48434;
w48761 <= not w48430 and w48760;
w48762 <= not w48431 and not w48434;
w48763 <= not w48761 and not w48762;
w48764 <= not w48559 and not w48763;
w48765 <= not w48014 and not w48558;
w48766 <= not w48557 and w48765;
w48767 <= not w48764 and not w48766;
w48768 <= not b(32) and not w48767;
w48769 <= not w48033 and w48429;
w48770 <= not w48425 and w48769;
w48771 <= not w48426 and not w48429;
w48772 <= not w48770 and not w48771;
w48773 <= not w48559 and not w48772;
w48774 <= not w48023 and not w48558;
w48775 <= not w48557 and w48774;
w48776 <= not w48773 and not w48775;
w48777 <= not b(31) and not w48776;
w48778 <= not w48042 and w48424;
w48779 <= not w48420 and w48778;
w48780 <= not w48421 and not w48424;
w48781 <= not w48779 and not w48780;
w48782 <= not w48559 and not w48781;
w48783 <= not w48032 and not w48558;
w48784 <= not w48557 and w48783;
w48785 <= not w48782 and not w48784;
w48786 <= not b(30) and not w48785;
w48787 <= not w48051 and w48419;
w48788 <= not w48415 and w48787;
w48789 <= not w48416 and not w48419;
w48790 <= not w48788 and not w48789;
w48791 <= not w48559 and not w48790;
w48792 <= not w48041 and not w48558;
w48793 <= not w48557 and w48792;
w48794 <= not w48791 and not w48793;
w48795 <= not b(29) and not w48794;
w48796 <= not w48060 and w48414;
w48797 <= not w48410 and w48796;
w48798 <= not w48411 and not w48414;
w48799 <= not w48797 and not w48798;
w48800 <= not w48559 and not w48799;
w48801 <= not w48050 and not w48558;
w48802 <= not w48557 and w48801;
w48803 <= not w48800 and not w48802;
w48804 <= not b(28) and not w48803;
w48805 <= not w48069 and w48409;
w48806 <= not w48405 and w48805;
w48807 <= not w48406 and not w48409;
w48808 <= not w48806 and not w48807;
w48809 <= not w48559 and not w48808;
w48810 <= not w48059 and not w48558;
w48811 <= not w48557 and w48810;
w48812 <= not w48809 and not w48811;
w48813 <= not b(27) and not w48812;
w48814 <= not w48078 and w48404;
w48815 <= not w48400 and w48814;
w48816 <= not w48401 and not w48404;
w48817 <= not w48815 and not w48816;
w48818 <= not w48559 and not w48817;
w48819 <= not w48068 and not w48558;
w48820 <= not w48557 and w48819;
w48821 <= not w48818 and not w48820;
w48822 <= not b(26) and not w48821;
w48823 <= not w48087 and w48399;
w48824 <= not w48395 and w48823;
w48825 <= not w48396 and not w48399;
w48826 <= not w48824 and not w48825;
w48827 <= not w48559 and not w48826;
w48828 <= not w48077 and not w48558;
w48829 <= not w48557 and w48828;
w48830 <= not w48827 and not w48829;
w48831 <= not b(25) and not w48830;
w48832 <= not w48096 and w48394;
w48833 <= not w48390 and w48832;
w48834 <= not w48391 and not w48394;
w48835 <= not w48833 and not w48834;
w48836 <= not w48559 and not w48835;
w48837 <= not w48086 and not w48558;
w48838 <= not w48557 and w48837;
w48839 <= not w48836 and not w48838;
w48840 <= not b(24) and not w48839;
w48841 <= not w48105 and w48389;
w48842 <= not w48385 and w48841;
w48843 <= not w48386 and not w48389;
w48844 <= not w48842 and not w48843;
w48845 <= not w48559 and not w48844;
w48846 <= not w48095 and not w48558;
w48847 <= not w48557 and w48846;
w48848 <= not w48845 and not w48847;
w48849 <= not b(23) and not w48848;
w48850 <= not w48114 and w48384;
w48851 <= not w48380 and w48850;
w48852 <= not w48381 and not w48384;
w48853 <= not w48851 and not w48852;
w48854 <= not w48559 and not w48853;
w48855 <= not w48104 and not w48558;
w48856 <= not w48557 and w48855;
w48857 <= not w48854 and not w48856;
w48858 <= not b(22) and not w48857;
w48859 <= not w48123 and w48379;
w48860 <= not w48375 and w48859;
w48861 <= not w48376 and not w48379;
w48862 <= not w48860 and not w48861;
w48863 <= not w48559 and not w48862;
w48864 <= not w48113 and not w48558;
w48865 <= not w48557 and w48864;
w48866 <= not w48863 and not w48865;
w48867 <= not b(21) and not w48866;
w48868 <= not w48132 and w48374;
w48869 <= not w48370 and w48868;
w48870 <= not w48371 and not w48374;
w48871 <= not w48869 and not w48870;
w48872 <= not w48559 and not w48871;
w48873 <= not w48122 and not w48558;
w48874 <= not w48557 and w48873;
w48875 <= not w48872 and not w48874;
w48876 <= not b(20) and not w48875;
w48877 <= not w48141 and w48369;
w48878 <= not w48365 and w48877;
w48879 <= not w48366 and not w48369;
w48880 <= not w48878 and not w48879;
w48881 <= not w48559 and not w48880;
w48882 <= not w48131 and not w48558;
w48883 <= not w48557 and w48882;
w48884 <= not w48881 and not w48883;
w48885 <= not b(19) and not w48884;
w48886 <= not w48150 and w48364;
w48887 <= not w48360 and w48886;
w48888 <= not w48361 and not w48364;
w48889 <= not w48887 and not w48888;
w48890 <= not w48559 and not w48889;
w48891 <= not w48140 and not w48558;
w48892 <= not w48557 and w48891;
w48893 <= not w48890 and not w48892;
w48894 <= not b(18) and not w48893;
w48895 <= not w48159 and w48359;
w48896 <= not w48355 and w48895;
w48897 <= not w48356 and not w48359;
w48898 <= not w48896 and not w48897;
w48899 <= not w48559 and not w48898;
w48900 <= not w48149 and not w48558;
w48901 <= not w48557 and w48900;
w48902 <= not w48899 and not w48901;
w48903 <= not b(17) and not w48902;
w48904 <= not w48168 and w48354;
w48905 <= not w48350 and w48904;
w48906 <= not w48351 and not w48354;
w48907 <= not w48905 and not w48906;
w48908 <= not w48559 and not w48907;
w48909 <= not w48158 and not w48558;
w48910 <= not w48557 and w48909;
w48911 <= not w48908 and not w48910;
w48912 <= not b(16) and not w48911;
w48913 <= not w48177 and w48349;
w48914 <= not w48345 and w48913;
w48915 <= not w48346 and not w48349;
w48916 <= not w48914 and not w48915;
w48917 <= not w48559 and not w48916;
w48918 <= not w48167 and not w48558;
w48919 <= not w48557 and w48918;
w48920 <= not w48917 and not w48919;
w48921 <= not b(15) and not w48920;
w48922 <= not w48186 and w48344;
w48923 <= not w48340 and w48922;
w48924 <= not w48341 and not w48344;
w48925 <= not w48923 and not w48924;
w48926 <= not w48559 and not w48925;
w48927 <= not w48176 and not w48558;
w48928 <= not w48557 and w48927;
w48929 <= not w48926 and not w48928;
w48930 <= not b(14) and not w48929;
w48931 <= not w48195 and w48339;
w48932 <= not w48335 and w48931;
w48933 <= not w48336 and not w48339;
w48934 <= not w48932 and not w48933;
w48935 <= not w48559 and not w48934;
w48936 <= not w48185 and not w48558;
w48937 <= not w48557 and w48936;
w48938 <= not w48935 and not w48937;
w48939 <= not b(13) and not w48938;
w48940 <= not w48204 and w48334;
w48941 <= not w48330 and w48940;
w48942 <= not w48331 and not w48334;
w48943 <= not w48941 and not w48942;
w48944 <= not w48559 and not w48943;
w48945 <= not w48194 and not w48558;
w48946 <= not w48557 and w48945;
w48947 <= not w48944 and not w48946;
w48948 <= not b(12) and not w48947;
w48949 <= not w48213 and w48329;
w48950 <= not w48325 and w48949;
w48951 <= not w48326 and not w48329;
w48952 <= not w48950 and not w48951;
w48953 <= not w48559 and not w48952;
w48954 <= not w48203 and not w48558;
w48955 <= not w48557 and w48954;
w48956 <= not w48953 and not w48955;
w48957 <= not b(11) and not w48956;
w48958 <= not w48222 and w48324;
w48959 <= not w48320 and w48958;
w48960 <= not w48321 and not w48324;
w48961 <= not w48959 and not w48960;
w48962 <= not w48559 and not w48961;
w48963 <= not w48212 and not w48558;
w48964 <= not w48557 and w48963;
w48965 <= not w48962 and not w48964;
w48966 <= not b(10) and not w48965;
w48967 <= not w48231 and w48319;
w48968 <= not w48315 and w48967;
w48969 <= not w48316 and not w48319;
w48970 <= not w48968 and not w48969;
w48971 <= not w48559 and not w48970;
w48972 <= not w48221 and not w48558;
w48973 <= not w48557 and w48972;
w48974 <= not w48971 and not w48973;
w48975 <= not b(9) and not w48974;
w48976 <= not w48240 and w48314;
w48977 <= not w48310 and w48976;
w48978 <= not w48311 and not w48314;
w48979 <= not w48977 and not w48978;
w48980 <= not w48559 and not w48979;
w48981 <= not w48230 and not w48558;
w48982 <= not w48557 and w48981;
w48983 <= not w48980 and not w48982;
w48984 <= not b(8) and not w48983;
w48985 <= not w48249 and w48309;
w48986 <= not w48305 and w48985;
w48987 <= not w48306 and not w48309;
w48988 <= not w48986 and not w48987;
w48989 <= not w48559 and not w48988;
w48990 <= not w48239 and not w48558;
w48991 <= not w48557 and w48990;
w48992 <= not w48989 and not w48991;
w48993 <= not b(7) and not w48992;
w48994 <= not w48258 and w48304;
w48995 <= not w48300 and w48994;
w48996 <= not w48301 and not w48304;
w48997 <= not w48995 and not w48996;
w48998 <= not w48559 and not w48997;
w48999 <= not w48248 and not w48558;
w49000 <= not w48557 and w48999;
w49001 <= not w48998 and not w49000;
w49002 <= not b(6) and not w49001;
w49003 <= not w48267 and w48299;
w49004 <= not w48295 and w49003;
w49005 <= not w48296 and not w48299;
w49006 <= not w49004 and not w49005;
w49007 <= not w48559 and not w49006;
w49008 <= not w48257 and not w48558;
w49009 <= not w48557 and w49008;
w49010 <= not w49007 and not w49009;
w49011 <= not b(5) and not w49010;
w49012 <= not w48275 and w48294;
w49013 <= not w48290 and w49012;
w49014 <= not w48291 and not w48294;
w49015 <= not w49013 and not w49014;
w49016 <= not w48559 and not w49015;
w49017 <= not w48266 and not w48558;
w49018 <= not w48557 and w49017;
w49019 <= not w49016 and not w49018;
w49020 <= not b(4) and not w49019;
w49021 <= not w48285 and w48289;
w49022 <= not w48284 and w49021;
w49023 <= not w48286 and not w48289;
w49024 <= not w49022 and not w49023;
w49025 <= not w48559 and not w49024;
w49026 <= not w48274 and not w48558;
w49027 <= not w48557 and w49026;
w49028 <= not w49025 and not w49027;
w49029 <= not b(3) and not w49028;
w49030 <= w20245 and not w48282;
w49031 <= not w48280 and w49030;
w49032 <= not w48284 and not w49031;
w49033 <= not w48559 and w49032;
w49034 <= not w48279 and not w48558;
w49035 <= not w48557 and w49034;
w49036 <= not w49033 and not w49035;
w49037 <= not b(2) and not w49036;
w49038 <= b(0) and not w48559;
w49039 <= a(10) and not w49038;
w49040 <= w20245 and not w48559;
w49041 <= not w49039 and not w49040;
w49042 <= b(1) and not w49041;
w49043 <= not b(1) and not w49040;
w49044 <= not w49039 and w49043;
w49045 <= not w49042 and not w49044;
w49046 <= not w21010 and not w49045;
w49047 <= not b(1) and not w49041;
w49048 <= not w49046 and not w49047;
w49049 <= b(2) and not w49035;
w49050 <= not w49033 and w49049;
w49051 <= not w49037 and not w49050;
w49052 <= not w49048 and w49051;
w49053 <= not w49037 and not w49052;
w49054 <= b(3) and not w49027;
w49055 <= not w49025 and w49054;
w49056 <= not w49029 and not w49055;
w49057 <= not w49053 and w49056;
w49058 <= not w49029 and not w49057;
w49059 <= b(4) and not w49018;
w49060 <= not w49016 and w49059;
w49061 <= not w49020 and not w49060;
w49062 <= not w49058 and w49061;
w49063 <= not w49020 and not w49062;
w49064 <= b(5) and not w49009;
w49065 <= not w49007 and w49064;
w49066 <= not w49011 and not w49065;
w49067 <= not w49063 and w49066;
w49068 <= not w49011 and not w49067;
w49069 <= b(6) and not w49000;
w49070 <= not w48998 and w49069;
w49071 <= not w49002 and not w49070;
w49072 <= not w49068 and w49071;
w49073 <= not w49002 and not w49072;
w49074 <= b(7) and not w48991;
w49075 <= not w48989 and w49074;
w49076 <= not w48993 and not w49075;
w49077 <= not w49073 and w49076;
w49078 <= not w48993 and not w49077;
w49079 <= b(8) and not w48982;
w49080 <= not w48980 and w49079;
w49081 <= not w48984 and not w49080;
w49082 <= not w49078 and w49081;
w49083 <= not w48984 and not w49082;
w49084 <= b(9) and not w48973;
w49085 <= not w48971 and w49084;
w49086 <= not w48975 and not w49085;
w49087 <= not w49083 and w49086;
w49088 <= not w48975 and not w49087;
w49089 <= b(10) and not w48964;
w49090 <= not w48962 and w49089;
w49091 <= not w48966 and not w49090;
w49092 <= not w49088 and w49091;
w49093 <= not w48966 and not w49092;
w49094 <= b(11) and not w48955;
w49095 <= not w48953 and w49094;
w49096 <= not w48957 and not w49095;
w49097 <= not w49093 and w49096;
w49098 <= not w48957 and not w49097;
w49099 <= b(12) and not w48946;
w49100 <= not w48944 and w49099;
w49101 <= not w48948 and not w49100;
w49102 <= not w49098 and w49101;
w49103 <= not w48948 and not w49102;
w49104 <= b(13) and not w48937;
w49105 <= not w48935 and w49104;
w49106 <= not w48939 and not w49105;
w49107 <= not w49103 and w49106;
w49108 <= not w48939 and not w49107;
w49109 <= b(14) and not w48928;
w49110 <= not w48926 and w49109;
w49111 <= not w48930 and not w49110;
w49112 <= not w49108 and w49111;
w49113 <= not w48930 and not w49112;
w49114 <= b(15) and not w48919;
w49115 <= not w48917 and w49114;
w49116 <= not w48921 and not w49115;
w49117 <= not w49113 and w49116;
w49118 <= not w48921 and not w49117;
w49119 <= b(16) and not w48910;
w49120 <= not w48908 and w49119;
w49121 <= not w48912 and not w49120;
w49122 <= not w49118 and w49121;
w49123 <= not w48912 and not w49122;
w49124 <= b(17) and not w48901;
w49125 <= not w48899 and w49124;
w49126 <= not w48903 and not w49125;
w49127 <= not w49123 and w49126;
w49128 <= not w48903 and not w49127;
w49129 <= b(18) and not w48892;
w49130 <= not w48890 and w49129;
w49131 <= not w48894 and not w49130;
w49132 <= not w49128 and w49131;
w49133 <= not w48894 and not w49132;
w49134 <= b(19) and not w48883;
w49135 <= not w48881 and w49134;
w49136 <= not w48885 and not w49135;
w49137 <= not w49133 and w49136;
w49138 <= not w48885 and not w49137;
w49139 <= b(20) and not w48874;
w49140 <= not w48872 and w49139;
w49141 <= not w48876 and not w49140;
w49142 <= not w49138 and w49141;
w49143 <= not w48876 and not w49142;
w49144 <= b(21) and not w48865;
w49145 <= not w48863 and w49144;
w49146 <= not w48867 and not w49145;
w49147 <= not w49143 and w49146;
w49148 <= not w48867 and not w49147;
w49149 <= b(22) and not w48856;
w49150 <= not w48854 and w49149;
w49151 <= not w48858 and not w49150;
w49152 <= not w49148 and w49151;
w49153 <= not w48858 and not w49152;
w49154 <= b(23) and not w48847;
w49155 <= not w48845 and w49154;
w49156 <= not w48849 and not w49155;
w49157 <= not w49153 and w49156;
w49158 <= not w48849 and not w49157;
w49159 <= b(24) and not w48838;
w49160 <= not w48836 and w49159;
w49161 <= not w48840 and not w49160;
w49162 <= not w49158 and w49161;
w49163 <= not w48840 and not w49162;
w49164 <= b(25) and not w48829;
w49165 <= not w48827 and w49164;
w49166 <= not w48831 and not w49165;
w49167 <= not w49163 and w49166;
w49168 <= not w48831 and not w49167;
w49169 <= b(26) and not w48820;
w49170 <= not w48818 and w49169;
w49171 <= not w48822 and not w49170;
w49172 <= not w49168 and w49171;
w49173 <= not w48822 and not w49172;
w49174 <= b(27) and not w48811;
w49175 <= not w48809 and w49174;
w49176 <= not w48813 and not w49175;
w49177 <= not w49173 and w49176;
w49178 <= not w48813 and not w49177;
w49179 <= b(28) and not w48802;
w49180 <= not w48800 and w49179;
w49181 <= not w48804 and not w49180;
w49182 <= not w49178 and w49181;
w49183 <= not w48804 and not w49182;
w49184 <= b(29) and not w48793;
w49185 <= not w48791 and w49184;
w49186 <= not w48795 and not w49185;
w49187 <= not w49183 and w49186;
w49188 <= not w48795 and not w49187;
w49189 <= b(30) and not w48784;
w49190 <= not w48782 and w49189;
w49191 <= not w48786 and not w49190;
w49192 <= not w49188 and w49191;
w49193 <= not w48786 and not w49192;
w49194 <= b(31) and not w48775;
w49195 <= not w48773 and w49194;
w49196 <= not w48777 and not w49195;
w49197 <= not w49193 and w49196;
w49198 <= not w48777 and not w49197;
w49199 <= b(32) and not w48766;
w49200 <= not w48764 and w49199;
w49201 <= not w48768 and not w49200;
w49202 <= not w49198 and w49201;
w49203 <= not w48768 and not w49202;
w49204 <= b(33) and not w48757;
w49205 <= not w48755 and w49204;
w49206 <= not w48759 and not w49205;
w49207 <= not w49203 and w49206;
w49208 <= not w48759 and not w49207;
w49209 <= b(34) and not w48748;
w49210 <= not w48746 and w49209;
w49211 <= not w48750 and not w49210;
w49212 <= not w49208 and w49211;
w49213 <= not w48750 and not w49212;
w49214 <= b(35) and not w48739;
w49215 <= not w48737 and w49214;
w49216 <= not w48741 and not w49215;
w49217 <= not w49213 and w49216;
w49218 <= not w48741 and not w49217;
w49219 <= b(36) and not w48730;
w49220 <= not w48728 and w49219;
w49221 <= not w48732 and not w49220;
w49222 <= not w49218 and w49221;
w49223 <= not w48732 and not w49222;
w49224 <= b(37) and not w48721;
w49225 <= not w48719 and w49224;
w49226 <= not w48723 and not w49225;
w49227 <= not w49223 and w49226;
w49228 <= not w48723 and not w49227;
w49229 <= b(38) and not w48712;
w49230 <= not w48710 and w49229;
w49231 <= not w48714 and not w49230;
w49232 <= not w49228 and w49231;
w49233 <= not w48714 and not w49232;
w49234 <= b(39) and not w48703;
w49235 <= not w48701 and w49234;
w49236 <= not w48705 and not w49235;
w49237 <= not w49233 and w49236;
w49238 <= not w48705 and not w49237;
w49239 <= b(40) and not w48694;
w49240 <= not w48692 and w49239;
w49241 <= not w48696 and not w49240;
w49242 <= not w49238 and w49241;
w49243 <= not w48696 and not w49242;
w49244 <= b(41) and not w48685;
w49245 <= not w48683 and w49244;
w49246 <= not w48687 and not w49245;
w49247 <= not w49243 and w49246;
w49248 <= not w48687 and not w49247;
w49249 <= b(42) and not w48676;
w49250 <= not w48674 and w49249;
w49251 <= not w48678 and not w49250;
w49252 <= not w49248 and w49251;
w49253 <= not w48678 and not w49252;
w49254 <= b(43) and not w48667;
w49255 <= not w48665 and w49254;
w49256 <= not w48669 and not w49255;
w49257 <= not w49253 and w49256;
w49258 <= not w48669 and not w49257;
w49259 <= b(44) and not w48658;
w49260 <= not w48656 and w49259;
w49261 <= not w48660 and not w49260;
w49262 <= not w49258 and w49261;
w49263 <= not w48660 and not w49262;
w49264 <= b(45) and not w48649;
w49265 <= not w48647 and w49264;
w49266 <= not w48651 and not w49265;
w49267 <= not w49263 and w49266;
w49268 <= not w48651 and not w49267;
w49269 <= b(46) and not w48640;
w49270 <= not w48638 and w49269;
w49271 <= not w48642 and not w49270;
w49272 <= not w49268 and w49271;
w49273 <= not w48642 and not w49272;
w49274 <= b(47) and not w48631;
w49275 <= not w48629 and w49274;
w49276 <= not w48633 and not w49275;
w49277 <= not w49273 and w49276;
w49278 <= not w48633 and not w49277;
w49279 <= b(48) and not w48622;
w49280 <= not w48620 and w49279;
w49281 <= not w48624 and not w49280;
w49282 <= not w49278 and w49281;
w49283 <= not w48624 and not w49282;
w49284 <= b(49) and not w48613;
w49285 <= not w48611 and w49284;
w49286 <= not w48615 and not w49285;
w49287 <= not w49283 and w49286;
w49288 <= not w48615 and not w49287;
w49289 <= b(50) and not w48604;
w49290 <= not w48602 and w49289;
w49291 <= not w48606 and not w49290;
w49292 <= not w49288 and w49291;
w49293 <= not w48606 and not w49292;
w49294 <= b(51) and not w48595;
w49295 <= not w48593 and w49294;
w49296 <= not w48597 and not w49295;
w49297 <= not w49293 and w49296;
w49298 <= not w48597 and not w49297;
w49299 <= b(52) and not w48586;
w49300 <= not w48584 and w49299;
w49301 <= not w48588 and not w49300;
w49302 <= not w49298 and w49301;
w49303 <= not w48588 and not w49302;
w49304 <= b(53) and not w48566;
w49305 <= not w48564 and w49304;
w49306 <= not w48579 and not w49305;
w49307 <= not w49303 and w49306;
w49308 <= not w48579 and not w49307;
w49309 <= b(54) and not w48576;
w49310 <= not w48574 and w49309;
w49311 <= not w48578 and not w49310;
w49312 <= not w49308 and w49311;
w49313 <= not w48578 and not w49312;
w49314 <= w21280 and not w49313;
w49315 <= not w48567 and not w49314;
w49316 <= not w48588 and w49306;
w49317 <= not w49302 and w49316;
w49318 <= not w49303 and not w49306;
w49319 <= not w49317 and not w49318;
w49320 <= w21280 and not w49319;
w49321 <= not w49313 and w49320;
w49322 <= not w49315 and not w49321;
w49323 <= not b(54) and not w49322;
w49324 <= not w48587 and not w49314;
w49325 <= not w48597 and w49301;
w49326 <= not w49297 and w49325;
w49327 <= not w49298 and not w49301;
w49328 <= not w49326 and not w49327;
w49329 <= w21280 and not w49328;
w49330 <= not w49313 and w49329;
w49331 <= not w49324 and not w49330;
w49332 <= not b(53) and not w49331;
w49333 <= not w48596 and not w49314;
w49334 <= not w48606 and w49296;
w49335 <= not w49292 and w49334;
w49336 <= not w49293 and not w49296;
w49337 <= not w49335 and not w49336;
w49338 <= w21280 and not w49337;
w49339 <= not w49313 and w49338;
w49340 <= not w49333 and not w49339;
w49341 <= not b(52) and not w49340;
w49342 <= not w48605 and not w49314;
w49343 <= not w48615 and w49291;
w49344 <= not w49287 and w49343;
w49345 <= not w49288 and not w49291;
w49346 <= not w49344 and not w49345;
w49347 <= w21280 and not w49346;
w49348 <= not w49313 and w49347;
w49349 <= not w49342 and not w49348;
w49350 <= not b(51) and not w49349;
w49351 <= not w48614 and not w49314;
w49352 <= not w48624 and w49286;
w49353 <= not w49282 and w49352;
w49354 <= not w49283 and not w49286;
w49355 <= not w49353 and not w49354;
w49356 <= w21280 and not w49355;
w49357 <= not w49313 and w49356;
w49358 <= not w49351 and not w49357;
w49359 <= not b(50) and not w49358;
w49360 <= not w48623 and not w49314;
w49361 <= not w48633 and w49281;
w49362 <= not w49277 and w49361;
w49363 <= not w49278 and not w49281;
w49364 <= not w49362 and not w49363;
w49365 <= w21280 and not w49364;
w49366 <= not w49313 and w49365;
w49367 <= not w49360 and not w49366;
w49368 <= not b(49) and not w49367;
w49369 <= not w48632 and not w49314;
w49370 <= not w48642 and w49276;
w49371 <= not w49272 and w49370;
w49372 <= not w49273 and not w49276;
w49373 <= not w49371 and not w49372;
w49374 <= w21280 and not w49373;
w49375 <= not w49313 and w49374;
w49376 <= not w49369 and not w49375;
w49377 <= not b(48) and not w49376;
w49378 <= not w48641 and not w49314;
w49379 <= not w48651 and w49271;
w49380 <= not w49267 and w49379;
w49381 <= not w49268 and not w49271;
w49382 <= not w49380 and not w49381;
w49383 <= w21280 and not w49382;
w49384 <= not w49313 and w49383;
w49385 <= not w49378 and not w49384;
w49386 <= not b(47) and not w49385;
w49387 <= not w48650 and not w49314;
w49388 <= not w48660 and w49266;
w49389 <= not w49262 and w49388;
w49390 <= not w49263 and not w49266;
w49391 <= not w49389 and not w49390;
w49392 <= w21280 and not w49391;
w49393 <= not w49313 and w49392;
w49394 <= not w49387 and not w49393;
w49395 <= not b(46) and not w49394;
w49396 <= not w48659 and not w49314;
w49397 <= not w48669 and w49261;
w49398 <= not w49257 and w49397;
w49399 <= not w49258 and not w49261;
w49400 <= not w49398 and not w49399;
w49401 <= w21280 and not w49400;
w49402 <= not w49313 and w49401;
w49403 <= not w49396 and not w49402;
w49404 <= not b(45) and not w49403;
w49405 <= not w48668 and not w49314;
w49406 <= not w48678 and w49256;
w49407 <= not w49252 and w49406;
w49408 <= not w49253 and not w49256;
w49409 <= not w49407 and not w49408;
w49410 <= w21280 and not w49409;
w49411 <= not w49313 and w49410;
w49412 <= not w49405 and not w49411;
w49413 <= not b(44) and not w49412;
w49414 <= not w48677 and not w49314;
w49415 <= not w48687 and w49251;
w49416 <= not w49247 and w49415;
w49417 <= not w49248 and not w49251;
w49418 <= not w49416 and not w49417;
w49419 <= w21280 and not w49418;
w49420 <= not w49313 and w49419;
w49421 <= not w49414 and not w49420;
w49422 <= not b(43) and not w49421;
w49423 <= not w48686 and not w49314;
w49424 <= not w48696 and w49246;
w49425 <= not w49242 and w49424;
w49426 <= not w49243 and not w49246;
w49427 <= not w49425 and not w49426;
w49428 <= w21280 and not w49427;
w49429 <= not w49313 and w49428;
w49430 <= not w49423 and not w49429;
w49431 <= not b(42) and not w49430;
w49432 <= not w48695 and not w49314;
w49433 <= not w48705 and w49241;
w49434 <= not w49237 and w49433;
w49435 <= not w49238 and not w49241;
w49436 <= not w49434 and not w49435;
w49437 <= w21280 and not w49436;
w49438 <= not w49313 and w49437;
w49439 <= not w49432 and not w49438;
w49440 <= not b(41) and not w49439;
w49441 <= not w48704 and not w49314;
w49442 <= not w48714 and w49236;
w49443 <= not w49232 and w49442;
w49444 <= not w49233 and not w49236;
w49445 <= not w49443 and not w49444;
w49446 <= w21280 and not w49445;
w49447 <= not w49313 and w49446;
w49448 <= not w49441 and not w49447;
w49449 <= not b(40) and not w49448;
w49450 <= not w48713 and not w49314;
w49451 <= not w48723 and w49231;
w49452 <= not w49227 and w49451;
w49453 <= not w49228 and not w49231;
w49454 <= not w49452 and not w49453;
w49455 <= w21280 and not w49454;
w49456 <= not w49313 and w49455;
w49457 <= not w49450 and not w49456;
w49458 <= not b(39) and not w49457;
w49459 <= not w48722 and not w49314;
w49460 <= not w48732 and w49226;
w49461 <= not w49222 and w49460;
w49462 <= not w49223 and not w49226;
w49463 <= not w49461 and not w49462;
w49464 <= w21280 and not w49463;
w49465 <= not w49313 and w49464;
w49466 <= not w49459 and not w49465;
w49467 <= not b(38) and not w49466;
w49468 <= not w48731 and not w49314;
w49469 <= not w48741 and w49221;
w49470 <= not w49217 and w49469;
w49471 <= not w49218 and not w49221;
w49472 <= not w49470 and not w49471;
w49473 <= w21280 and not w49472;
w49474 <= not w49313 and w49473;
w49475 <= not w49468 and not w49474;
w49476 <= not b(37) and not w49475;
w49477 <= not w48740 and not w49314;
w49478 <= not w48750 and w49216;
w49479 <= not w49212 and w49478;
w49480 <= not w49213 and not w49216;
w49481 <= not w49479 and not w49480;
w49482 <= w21280 and not w49481;
w49483 <= not w49313 and w49482;
w49484 <= not w49477 and not w49483;
w49485 <= not b(36) and not w49484;
w49486 <= not w48749 and not w49314;
w49487 <= not w48759 and w49211;
w49488 <= not w49207 and w49487;
w49489 <= not w49208 and not w49211;
w49490 <= not w49488 and not w49489;
w49491 <= w21280 and not w49490;
w49492 <= not w49313 and w49491;
w49493 <= not w49486 and not w49492;
w49494 <= not b(35) and not w49493;
w49495 <= not w48758 and not w49314;
w49496 <= not w48768 and w49206;
w49497 <= not w49202 and w49496;
w49498 <= not w49203 and not w49206;
w49499 <= not w49497 and not w49498;
w49500 <= w21280 and not w49499;
w49501 <= not w49313 and w49500;
w49502 <= not w49495 and not w49501;
w49503 <= not b(34) and not w49502;
w49504 <= not w48767 and not w49314;
w49505 <= not w48777 and w49201;
w49506 <= not w49197 and w49505;
w49507 <= not w49198 and not w49201;
w49508 <= not w49506 and not w49507;
w49509 <= w21280 and not w49508;
w49510 <= not w49313 and w49509;
w49511 <= not w49504 and not w49510;
w49512 <= not b(33) and not w49511;
w49513 <= not w48776 and not w49314;
w49514 <= not w48786 and w49196;
w49515 <= not w49192 and w49514;
w49516 <= not w49193 and not w49196;
w49517 <= not w49515 and not w49516;
w49518 <= w21280 and not w49517;
w49519 <= not w49313 and w49518;
w49520 <= not w49513 and not w49519;
w49521 <= not b(32) and not w49520;
w49522 <= not w48785 and not w49314;
w49523 <= not w48795 and w49191;
w49524 <= not w49187 and w49523;
w49525 <= not w49188 and not w49191;
w49526 <= not w49524 and not w49525;
w49527 <= w21280 and not w49526;
w49528 <= not w49313 and w49527;
w49529 <= not w49522 and not w49528;
w49530 <= not b(31) and not w49529;
w49531 <= not w48794 and not w49314;
w49532 <= not w48804 and w49186;
w49533 <= not w49182 and w49532;
w49534 <= not w49183 and not w49186;
w49535 <= not w49533 and not w49534;
w49536 <= w21280 and not w49535;
w49537 <= not w49313 and w49536;
w49538 <= not w49531 and not w49537;
w49539 <= not b(30) and not w49538;
w49540 <= not w48803 and not w49314;
w49541 <= not w48813 and w49181;
w49542 <= not w49177 and w49541;
w49543 <= not w49178 and not w49181;
w49544 <= not w49542 and not w49543;
w49545 <= w21280 and not w49544;
w49546 <= not w49313 and w49545;
w49547 <= not w49540 and not w49546;
w49548 <= not b(29) and not w49547;
w49549 <= not w48812 and not w49314;
w49550 <= not w48822 and w49176;
w49551 <= not w49172 and w49550;
w49552 <= not w49173 and not w49176;
w49553 <= not w49551 and not w49552;
w49554 <= w21280 and not w49553;
w49555 <= not w49313 and w49554;
w49556 <= not w49549 and not w49555;
w49557 <= not b(28) and not w49556;
w49558 <= not w48821 and not w49314;
w49559 <= not w48831 and w49171;
w49560 <= not w49167 and w49559;
w49561 <= not w49168 and not w49171;
w49562 <= not w49560 and not w49561;
w49563 <= w21280 and not w49562;
w49564 <= not w49313 and w49563;
w49565 <= not w49558 and not w49564;
w49566 <= not b(27) and not w49565;
w49567 <= not w48830 and not w49314;
w49568 <= not w48840 and w49166;
w49569 <= not w49162 and w49568;
w49570 <= not w49163 and not w49166;
w49571 <= not w49569 and not w49570;
w49572 <= w21280 and not w49571;
w49573 <= not w49313 and w49572;
w49574 <= not w49567 and not w49573;
w49575 <= not b(26) and not w49574;
w49576 <= not w48839 and not w49314;
w49577 <= not w48849 and w49161;
w49578 <= not w49157 and w49577;
w49579 <= not w49158 and not w49161;
w49580 <= not w49578 and not w49579;
w49581 <= w21280 and not w49580;
w49582 <= not w49313 and w49581;
w49583 <= not w49576 and not w49582;
w49584 <= not b(25) and not w49583;
w49585 <= not w48848 and not w49314;
w49586 <= not w48858 and w49156;
w49587 <= not w49152 and w49586;
w49588 <= not w49153 and not w49156;
w49589 <= not w49587 and not w49588;
w49590 <= w21280 and not w49589;
w49591 <= not w49313 and w49590;
w49592 <= not w49585 and not w49591;
w49593 <= not b(24) and not w49592;
w49594 <= not w48857 and not w49314;
w49595 <= not w48867 and w49151;
w49596 <= not w49147 and w49595;
w49597 <= not w49148 and not w49151;
w49598 <= not w49596 and not w49597;
w49599 <= w21280 and not w49598;
w49600 <= not w49313 and w49599;
w49601 <= not w49594 and not w49600;
w49602 <= not b(23) and not w49601;
w49603 <= not w48866 and not w49314;
w49604 <= not w48876 and w49146;
w49605 <= not w49142 and w49604;
w49606 <= not w49143 and not w49146;
w49607 <= not w49605 and not w49606;
w49608 <= w21280 and not w49607;
w49609 <= not w49313 and w49608;
w49610 <= not w49603 and not w49609;
w49611 <= not b(22) and not w49610;
w49612 <= not w48875 and not w49314;
w49613 <= not w48885 and w49141;
w49614 <= not w49137 and w49613;
w49615 <= not w49138 and not w49141;
w49616 <= not w49614 and not w49615;
w49617 <= w21280 and not w49616;
w49618 <= not w49313 and w49617;
w49619 <= not w49612 and not w49618;
w49620 <= not b(21) and not w49619;
w49621 <= not w48884 and not w49314;
w49622 <= not w48894 and w49136;
w49623 <= not w49132 and w49622;
w49624 <= not w49133 and not w49136;
w49625 <= not w49623 and not w49624;
w49626 <= w21280 and not w49625;
w49627 <= not w49313 and w49626;
w49628 <= not w49621 and not w49627;
w49629 <= not b(20) and not w49628;
w49630 <= not w48893 and not w49314;
w49631 <= not w48903 and w49131;
w49632 <= not w49127 and w49631;
w49633 <= not w49128 and not w49131;
w49634 <= not w49632 and not w49633;
w49635 <= w21280 and not w49634;
w49636 <= not w49313 and w49635;
w49637 <= not w49630 and not w49636;
w49638 <= not b(19) and not w49637;
w49639 <= not w48902 and not w49314;
w49640 <= not w48912 and w49126;
w49641 <= not w49122 and w49640;
w49642 <= not w49123 and not w49126;
w49643 <= not w49641 and not w49642;
w49644 <= w21280 and not w49643;
w49645 <= not w49313 and w49644;
w49646 <= not w49639 and not w49645;
w49647 <= not b(18) and not w49646;
w49648 <= not w48911 and not w49314;
w49649 <= not w48921 and w49121;
w49650 <= not w49117 and w49649;
w49651 <= not w49118 and not w49121;
w49652 <= not w49650 and not w49651;
w49653 <= w21280 and not w49652;
w49654 <= not w49313 and w49653;
w49655 <= not w49648 and not w49654;
w49656 <= not b(17) and not w49655;
w49657 <= not w48920 and not w49314;
w49658 <= not w48930 and w49116;
w49659 <= not w49112 and w49658;
w49660 <= not w49113 and not w49116;
w49661 <= not w49659 and not w49660;
w49662 <= w21280 and not w49661;
w49663 <= not w49313 and w49662;
w49664 <= not w49657 and not w49663;
w49665 <= not b(16) and not w49664;
w49666 <= not w48929 and not w49314;
w49667 <= not w48939 and w49111;
w49668 <= not w49107 and w49667;
w49669 <= not w49108 and not w49111;
w49670 <= not w49668 and not w49669;
w49671 <= w21280 and not w49670;
w49672 <= not w49313 and w49671;
w49673 <= not w49666 and not w49672;
w49674 <= not b(15) and not w49673;
w49675 <= not w48938 and not w49314;
w49676 <= not w48948 and w49106;
w49677 <= not w49102 and w49676;
w49678 <= not w49103 and not w49106;
w49679 <= not w49677 and not w49678;
w49680 <= w21280 and not w49679;
w49681 <= not w49313 and w49680;
w49682 <= not w49675 and not w49681;
w49683 <= not b(14) and not w49682;
w49684 <= not w48947 and not w49314;
w49685 <= not w48957 and w49101;
w49686 <= not w49097 and w49685;
w49687 <= not w49098 and not w49101;
w49688 <= not w49686 and not w49687;
w49689 <= w21280 and not w49688;
w49690 <= not w49313 and w49689;
w49691 <= not w49684 and not w49690;
w49692 <= not b(13) and not w49691;
w49693 <= not w48956 and not w49314;
w49694 <= not w48966 and w49096;
w49695 <= not w49092 and w49694;
w49696 <= not w49093 and not w49096;
w49697 <= not w49695 and not w49696;
w49698 <= w21280 and not w49697;
w49699 <= not w49313 and w49698;
w49700 <= not w49693 and not w49699;
w49701 <= not b(12) and not w49700;
w49702 <= not w48965 and not w49314;
w49703 <= not w48975 and w49091;
w49704 <= not w49087 and w49703;
w49705 <= not w49088 and not w49091;
w49706 <= not w49704 and not w49705;
w49707 <= w21280 and not w49706;
w49708 <= not w49313 and w49707;
w49709 <= not w49702 and not w49708;
w49710 <= not b(11) and not w49709;
w49711 <= not w48974 and not w49314;
w49712 <= not w48984 and w49086;
w49713 <= not w49082 and w49712;
w49714 <= not w49083 and not w49086;
w49715 <= not w49713 and not w49714;
w49716 <= w21280 and not w49715;
w49717 <= not w49313 and w49716;
w49718 <= not w49711 and not w49717;
w49719 <= not b(10) and not w49718;
w49720 <= not w48983 and not w49314;
w49721 <= not w48993 and w49081;
w49722 <= not w49077 and w49721;
w49723 <= not w49078 and not w49081;
w49724 <= not w49722 and not w49723;
w49725 <= w21280 and not w49724;
w49726 <= not w49313 and w49725;
w49727 <= not w49720 and not w49726;
w49728 <= not b(9) and not w49727;
w49729 <= not w48992 and not w49314;
w49730 <= not w49002 and w49076;
w49731 <= not w49072 and w49730;
w49732 <= not w49073 and not w49076;
w49733 <= not w49731 and not w49732;
w49734 <= w21280 and not w49733;
w49735 <= not w49313 and w49734;
w49736 <= not w49729 and not w49735;
w49737 <= not b(8) and not w49736;
w49738 <= not w49001 and not w49314;
w49739 <= not w49011 and w49071;
w49740 <= not w49067 and w49739;
w49741 <= not w49068 and not w49071;
w49742 <= not w49740 and not w49741;
w49743 <= w21280 and not w49742;
w49744 <= not w49313 and w49743;
w49745 <= not w49738 and not w49744;
w49746 <= not b(7) and not w49745;
w49747 <= not w49010 and not w49314;
w49748 <= not w49020 and w49066;
w49749 <= not w49062 and w49748;
w49750 <= not w49063 and not w49066;
w49751 <= not w49749 and not w49750;
w49752 <= w21280 and not w49751;
w49753 <= not w49313 and w49752;
w49754 <= not w49747 and not w49753;
w49755 <= not b(6) and not w49754;
w49756 <= not w49019 and not w49314;
w49757 <= not w49029 and w49061;
w49758 <= not w49057 and w49757;
w49759 <= not w49058 and not w49061;
w49760 <= not w49758 and not w49759;
w49761 <= w21280 and not w49760;
w49762 <= not w49313 and w49761;
w49763 <= not w49756 and not w49762;
w49764 <= not b(5) and not w49763;
w49765 <= not w49028 and not w49314;
w49766 <= not w49037 and w49056;
w49767 <= not w49052 and w49766;
w49768 <= not w49053 and not w49056;
w49769 <= not w49767 and not w49768;
w49770 <= w21280 and not w49769;
w49771 <= not w49313 and w49770;
w49772 <= not w49765 and not w49771;
w49773 <= not b(4) and not w49772;
w49774 <= not w49036 and not w49314;
w49775 <= not w49047 and w49051;
w49776 <= not w49046 and w49775;
w49777 <= not w49048 and not w49051;
w49778 <= not w49776 and not w49777;
w49779 <= w21280 and not w49778;
w49780 <= not w49313 and w49779;
w49781 <= not w49774 and not w49780;
w49782 <= not b(3) and not w49781;
w49783 <= not w49041 and not w49314;
w49784 <= w21010 and not w49044;
w49785 <= not w49042 and w49784;
w49786 <= w21280 and not w49785;
w49787 <= not w49046 and w49786;
w49788 <= not w49313 and w49787;
w49789 <= not w49783 and not w49788;
w49790 <= not b(2) and not w49789;
w49791 <= w21760 and not w49313;
w49792 <= a(9) and not w49791;
w49793 <= w21765 and not w49313;
w49794 <= not w49792 and not w49793;
w49795 <= b(1) and not w49794;
w49796 <= not b(1) and not w49793;
w49797 <= not w49792 and w49796;
w49798 <= not w49795 and not w49797;
w49799 <= not w21772 and not w49798;
w49800 <= not b(1) and not w49794;
w49801 <= not w49799 and not w49800;
w49802 <= b(2) and not w49788;
w49803 <= not w49783 and w49802;
w49804 <= not w49790 and not w49803;
w49805 <= not w49801 and w49804;
w49806 <= not w49790 and not w49805;
w49807 <= b(3) and not w49780;
w49808 <= not w49774 and w49807;
w49809 <= not w49782 and not w49808;
w49810 <= not w49806 and w49809;
w49811 <= not w49782 and not w49810;
w49812 <= b(4) and not w49771;
w49813 <= not w49765 and w49812;
w49814 <= not w49773 and not w49813;
w49815 <= not w49811 and w49814;
w49816 <= not w49773 and not w49815;
w49817 <= b(5) and not w49762;
w49818 <= not w49756 and w49817;
w49819 <= not w49764 and not w49818;
w49820 <= not w49816 and w49819;
w49821 <= not w49764 and not w49820;
w49822 <= b(6) and not w49753;
w49823 <= not w49747 and w49822;
w49824 <= not w49755 and not w49823;
w49825 <= not w49821 and w49824;
w49826 <= not w49755 and not w49825;
w49827 <= b(7) and not w49744;
w49828 <= not w49738 and w49827;
w49829 <= not w49746 and not w49828;
w49830 <= not w49826 and w49829;
w49831 <= not w49746 and not w49830;
w49832 <= b(8) and not w49735;
w49833 <= not w49729 and w49832;
w49834 <= not w49737 and not w49833;
w49835 <= not w49831 and w49834;
w49836 <= not w49737 and not w49835;
w49837 <= b(9) and not w49726;
w49838 <= not w49720 and w49837;
w49839 <= not w49728 and not w49838;
w49840 <= not w49836 and w49839;
w49841 <= not w49728 and not w49840;
w49842 <= b(10) and not w49717;
w49843 <= not w49711 and w49842;
w49844 <= not w49719 and not w49843;
w49845 <= not w49841 and w49844;
w49846 <= not w49719 and not w49845;
w49847 <= b(11) and not w49708;
w49848 <= not w49702 and w49847;
w49849 <= not w49710 and not w49848;
w49850 <= not w49846 and w49849;
w49851 <= not w49710 and not w49850;
w49852 <= b(12) and not w49699;
w49853 <= not w49693 and w49852;
w49854 <= not w49701 and not w49853;
w49855 <= not w49851 and w49854;
w49856 <= not w49701 and not w49855;
w49857 <= b(13) and not w49690;
w49858 <= not w49684 and w49857;
w49859 <= not w49692 and not w49858;
w49860 <= not w49856 and w49859;
w49861 <= not w49692 and not w49860;
w49862 <= b(14) and not w49681;
w49863 <= not w49675 and w49862;
w49864 <= not w49683 and not w49863;
w49865 <= not w49861 and w49864;
w49866 <= not w49683 and not w49865;
w49867 <= b(15) and not w49672;
w49868 <= not w49666 and w49867;
w49869 <= not w49674 and not w49868;
w49870 <= not w49866 and w49869;
w49871 <= not w49674 and not w49870;
w49872 <= b(16) and not w49663;
w49873 <= not w49657 and w49872;
w49874 <= not w49665 and not w49873;
w49875 <= not w49871 and w49874;
w49876 <= not w49665 and not w49875;
w49877 <= b(17) and not w49654;
w49878 <= not w49648 and w49877;
w49879 <= not w49656 and not w49878;
w49880 <= not w49876 and w49879;
w49881 <= not w49656 and not w49880;
w49882 <= b(18) and not w49645;
w49883 <= not w49639 and w49882;
w49884 <= not w49647 and not w49883;
w49885 <= not w49881 and w49884;
w49886 <= not w49647 and not w49885;
w49887 <= b(19) and not w49636;
w49888 <= not w49630 and w49887;
w49889 <= not w49638 and not w49888;
w49890 <= not w49886 and w49889;
w49891 <= not w49638 and not w49890;
w49892 <= b(20) and not w49627;
w49893 <= not w49621 and w49892;
w49894 <= not w49629 and not w49893;
w49895 <= not w49891 and w49894;
w49896 <= not w49629 and not w49895;
w49897 <= b(21) and not w49618;
w49898 <= not w49612 and w49897;
w49899 <= not w49620 and not w49898;
w49900 <= not w49896 and w49899;
w49901 <= not w49620 and not w49900;
w49902 <= b(22) and not w49609;
w49903 <= not w49603 and w49902;
w49904 <= not w49611 and not w49903;
w49905 <= not w49901 and w49904;
w49906 <= not w49611 and not w49905;
w49907 <= b(23) and not w49600;
w49908 <= not w49594 and w49907;
w49909 <= not w49602 and not w49908;
w49910 <= not w49906 and w49909;
w49911 <= not w49602 and not w49910;
w49912 <= b(24) and not w49591;
w49913 <= not w49585 and w49912;
w49914 <= not w49593 and not w49913;
w49915 <= not w49911 and w49914;
w49916 <= not w49593 and not w49915;
w49917 <= b(25) and not w49582;
w49918 <= not w49576 and w49917;
w49919 <= not w49584 and not w49918;
w49920 <= not w49916 and w49919;
w49921 <= not w49584 and not w49920;
w49922 <= b(26) and not w49573;
w49923 <= not w49567 and w49922;
w49924 <= not w49575 and not w49923;
w49925 <= not w49921 and w49924;
w49926 <= not w49575 and not w49925;
w49927 <= b(27) and not w49564;
w49928 <= not w49558 and w49927;
w49929 <= not w49566 and not w49928;
w49930 <= not w49926 and w49929;
w49931 <= not w49566 and not w49930;
w49932 <= b(28) and not w49555;
w49933 <= not w49549 and w49932;
w49934 <= not w49557 and not w49933;
w49935 <= not w49931 and w49934;
w49936 <= not w49557 and not w49935;
w49937 <= b(29) and not w49546;
w49938 <= not w49540 and w49937;
w49939 <= not w49548 and not w49938;
w49940 <= not w49936 and w49939;
w49941 <= not w49548 and not w49940;
w49942 <= b(30) and not w49537;
w49943 <= not w49531 and w49942;
w49944 <= not w49539 and not w49943;
w49945 <= not w49941 and w49944;
w49946 <= not w49539 and not w49945;
w49947 <= b(31) and not w49528;
w49948 <= not w49522 and w49947;
w49949 <= not w49530 and not w49948;
w49950 <= not w49946 and w49949;
w49951 <= not w49530 and not w49950;
w49952 <= b(32) and not w49519;
w49953 <= not w49513 and w49952;
w49954 <= not w49521 and not w49953;
w49955 <= not w49951 and w49954;
w49956 <= not w49521 and not w49955;
w49957 <= b(33) and not w49510;
w49958 <= not w49504 and w49957;
w49959 <= not w49512 and not w49958;
w49960 <= not w49956 and w49959;
w49961 <= not w49512 and not w49960;
w49962 <= b(34) and not w49501;
w49963 <= not w49495 and w49962;
w49964 <= not w49503 and not w49963;
w49965 <= not w49961 and w49964;
w49966 <= not w49503 and not w49965;
w49967 <= b(35) and not w49492;
w49968 <= not w49486 and w49967;
w49969 <= not w49494 and not w49968;
w49970 <= not w49966 and w49969;
w49971 <= not w49494 and not w49970;
w49972 <= b(36) and not w49483;
w49973 <= not w49477 and w49972;
w49974 <= not w49485 and not w49973;
w49975 <= not w49971 and w49974;
w49976 <= not w49485 and not w49975;
w49977 <= b(37) and not w49474;
w49978 <= not w49468 and w49977;
w49979 <= not w49476 and not w49978;
w49980 <= not w49976 and w49979;
w49981 <= not w49476 and not w49980;
w49982 <= b(38) and not w49465;
w49983 <= not w49459 and w49982;
w49984 <= not w49467 and not w49983;
w49985 <= not w49981 and w49984;
w49986 <= not w49467 and not w49985;
w49987 <= b(39) and not w49456;
w49988 <= not w49450 and w49987;
w49989 <= not w49458 and not w49988;
w49990 <= not w49986 and w49989;
w49991 <= not w49458 and not w49990;
w49992 <= b(40) and not w49447;
w49993 <= not w49441 and w49992;
w49994 <= not w49449 and not w49993;
w49995 <= not w49991 and w49994;
w49996 <= not w49449 and not w49995;
w49997 <= b(41) and not w49438;
w49998 <= not w49432 and w49997;
w49999 <= not w49440 and not w49998;
w50000 <= not w49996 and w49999;
w50001 <= not w49440 and not w50000;
w50002 <= b(42) and not w49429;
w50003 <= not w49423 and w50002;
w50004 <= not w49431 and not w50003;
w50005 <= not w50001 and w50004;
w50006 <= not w49431 and not w50005;
w50007 <= b(43) and not w49420;
w50008 <= not w49414 and w50007;
w50009 <= not w49422 and not w50008;
w50010 <= not w50006 and w50009;
w50011 <= not w49422 and not w50010;
w50012 <= b(44) and not w49411;
w50013 <= not w49405 and w50012;
w50014 <= not w49413 and not w50013;
w50015 <= not w50011 and w50014;
w50016 <= not w49413 and not w50015;
w50017 <= b(45) and not w49402;
w50018 <= not w49396 and w50017;
w50019 <= not w49404 and not w50018;
w50020 <= not w50016 and w50019;
w50021 <= not w49404 and not w50020;
w50022 <= b(46) and not w49393;
w50023 <= not w49387 and w50022;
w50024 <= not w49395 and not w50023;
w50025 <= not w50021 and w50024;
w50026 <= not w49395 and not w50025;
w50027 <= b(47) and not w49384;
w50028 <= not w49378 and w50027;
w50029 <= not w49386 and not w50028;
w50030 <= not w50026 and w50029;
w50031 <= not w49386 and not w50030;
w50032 <= b(48) and not w49375;
w50033 <= not w49369 and w50032;
w50034 <= not w49377 and not w50033;
w50035 <= not w50031 and w50034;
w50036 <= not w49377 and not w50035;
w50037 <= b(49) and not w49366;
w50038 <= not w49360 and w50037;
w50039 <= not w49368 and not w50038;
w50040 <= not w50036 and w50039;
w50041 <= not w49368 and not w50040;
w50042 <= b(50) and not w49357;
w50043 <= not w49351 and w50042;
w50044 <= not w49359 and not w50043;
w50045 <= not w50041 and w50044;
w50046 <= not w49359 and not w50045;
w50047 <= b(51) and not w49348;
w50048 <= not w49342 and w50047;
w50049 <= not w49350 and not w50048;
w50050 <= not w50046 and w50049;
w50051 <= not w49350 and not w50050;
w50052 <= b(52) and not w49339;
w50053 <= not w49333 and w50052;
w50054 <= not w49341 and not w50053;
w50055 <= not w50051 and w50054;
w50056 <= not w49341 and not w50055;
w50057 <= b(53) and not w49330;
w50058 <= not w49324 and w50057;
w50059 <= not w49332 and not w50058;
w50060 <= not w50056 and w50059;
w50061 <= not w49332 and not w50060;
w50062 <= b(54) and not w49321;
w50063 <= not w49315 and w50062;
w50064 <= not w49323 and not w50063;
w50065 <= not w50061 and w50064;
w50066 <= not w49323 and not w50065;
w50067 <= not w48577 and not w49314;
w50068 <= not w48579 and w49311;
w50069 <= not w49307 and w50068;
w50070 <= not w49308 and not w49311;
w50071 <= not w50069 and not w50070;
w50072 <= w49314 and not w50071;
w50073 <= not w50067 and not w50072;
w50074 <= not b(55) and not w50073;
w50075 <= b(55) and not w50067;
w50076 <= not w50072 and w50075;
w50077 <= w80 and not w50076;
w50078 <= not w50074 and w50077;
w50079 <= not w50066 and w50078;
w50080 <= w21280 and not w50073;
w50081 <= not w50079 and not w50080;
w50082 <= not w49332 and w50064;
w50083 <= not w50060 and w50082;
w50084 <= not w50061 and not w50064;
w50085 <= not w50083 and not w50084;
w50086 <= not w50081 and not w50085;
w50087 <= not w49322 and not w50080;
w50088 <= not w50079 and w50087;
w50089 <= not w50086 and not w50088;
w50090 <= not b(55) and not w50089;
w50091 <= not w49341 and w50059;
w50092 <= not w50055 and w50091;
w50093 <= not w50056 and not w50059;
w50094 <= not w50092 and not w50093;
w50095 <= not w50081 and not w50094;
w50096 <= not w49331 and not w50080;
w50097 <= not w50079 and w50096;
w50098 <= not w50095 and not w50097;
w50099 <= not b(54) and not w50098;
w50100 <= not w49350 and w50054;
w50101 <= not w50050 and w50100;
w50102 <= not w50051 and not w50054;
w50103 <= not w50101 and not w50102;
w50104 <= not w50081 and not w50103;
w50105 <= not w49340 and not w50080;
w50106 <= not w50079 and w50105;
w50107 <= not w50104 and not w50106;
w50108 <= not b(53) and not w50107;
w50109 <= not w49359 and w50049;
w50110 <= not w50045 and w50109;
w50111 <= not w50046 and not w50049;
w50112 <= not w50110 and not w50111;
w50113 <= not w50081 and not w50112;
w50114 <= not w49349 and not w50080;
w50115 <= not w50079 and w50114;
w50116 <= not w50113 and not w50115;
w50117 <= not b(52) and not w50116;
w50118 <= not w49368 and w50044;
w50119 <= not w50040 and w50118;
w50120 <= not w50041 and not w50044;
w50121 <= not w50119 and not w50120;
w50122 <= not w50081 and not w50121;
w50123 <= not w49358 and not w50080;
w50124 <= not w50079 and w50123;
w50125 <= not w50122 and not w50124;
w50126 <= not b(51) and not w50125;
w50127 <= not w49377 and w50039;
w50128 <= not w50035 and w50127;
w50129 <= not w50036 and not w50039;
w50130 <= not w50128 and not w50129;
w50131 <= not w50081 and not w50130;
w50132 <= not w49367 and not w50080;
w50133 <= not w50079 and w50132;
w50134 <= not w50131 and not w50133;
w50135 <= not b(50) and not w50134;
w50136 <= not w49386 and w50034;
w50137 <= not w50030 and w50136;
w50138 <= not w50031 and not w50034;
w50139 <= not w50137 and not w50138;
w50140 <= not w50081 and not w50139;
w50141 <= not w49376 and not w50080;
w50142 <= not w50079 and w50141;
w50143 <= not w50140 and not w50142;
w50144 <= not b(49) and not w50143;
w50145 <= not w49395 and w50029;
w50146 <= not w50025 and w50145;
w50147 <= not w50026 and not w50029;
w50148 <= not w50146 and not w50147;
w50149 <= not w50081 and not w50148;
w50150 <= not w49385 and not w50080;
w50151 <= not w50079 and w50150;
w50152 <= not w50149 and not w50151;
w50153 <= not b(48) and not w50152;
w50154 <= not w49404 and w50024;
w50155 <= not w50020 and w50154;
w50156 <= not w50021 and not w50024;
w50157 <= not w50155 and not w50156;
w50158 <= not w50081 and not w50157;
w50159 <= not w49394 and not w50080;
w50160 <= not w50079 and w50159;
w50161 <= not w50158 and not w50160;
w50162 <= not b(47) and not w50161;
w50163 <= not w49413 and w50019;
w50164 <= not w50015 and w50163;
w50165 <= not w50016 and not w50019;
w50166 <= not w50164 and not w50165;
w50167 <= not w50081 and not w50166;
w50168 <= not w49403 and not w50080;
w50169 <= not w50079 and w50168;
w50170 <= not w50167 and not w50169;
w50171 <= not b(46) and not w50170;
w50172 <= not w49422 and w50014;
w50173 <= not w50010 and w50172;
w50174 <= not w50011 and not w50014;
w50175 <= not w50173 and not w50174;
w50176 <= not w50081 and not w50175;
w50177 <= not w49412 and not w50080;
w50178 <= not w50079 and w50177;
w50179 <= not w50176 and not w50178;
w50180 <= not b(45) and not w50179;
w50181 <= not w49431 and w50009;
w50182 <= not w50005 and w50181;
w50183 <= not w50006 and not w50009;
w50184 <= not w50182 and not w50183;
w50185 <= not w50081 and not w50184;
w50186 <= not w49421 and not w50080;
w50187 <= not w50079 and w50186;
w50188 <= not w50185 and not w50187;
w50189 <= not b(44) and not w50188;
w50190 <= not w49440 and w50004;
w50191 <= not w50000 and w50190;
w50192 <= not w50001 and not w50004;
w50193 <= not w50191 and not w50192;
w50194 <= not w50081 and not w50193;
w50195 <= not w49430 and not w50080;
w50196 <= not w50079 and w50195;
w50197 <= not w50194 and not w50196;
w50198 <= not b(43) and not w50197;
w50199 <= not w49449 and w49999;
w50200 <= not w49995 and w50199;
w50201 <= not w49996 and not w49999;
w50202 <= not w50200 and not w50201;
w50203 <= not w50081 and not w50202;
w50204 <= not w49439 and not w50080;
w50205 <= not w50079 and w50204;
w50206 <= not w50203 and not w50205;
w50207 <= not b(42) and not w50206;
w50208 <= not w49458 and w49994;
w50209 <= not w49990 and w50208;
w50210 <= not w49991 and not w49994;
w50211 <= not w50209 and not w50210;
w50212 <= not w50081 and not w50211;
w50213 <= not w49448 and not w50080;
w50214 <= not w50079 and w50213;
w50215 <= not w50212 and not w50214;
w50216 <= not b(41) and not w50215;
w50217 <= not w49467 and w49989;
w50218 <= not w49985 and w50217;
w50219 <= not w49986 and not w49989;
w50220 <= not w50218 and not w50219;
w50221 <= not w50081 and not w50220;
w50222 <= not w49457 and not w50080;
w50223 <= not w50079 and w50222;
w50224 <= not w50221 and not w50223;
w50225 <= not b(40) and not w50224;
w50226 <= not w49476 and w49984;
w50227 <= not w49980 and w50226;
w50228 <= not w49981 and not w49984;
w50229 <= not w50227 and not w50228;
w50230 <= not w50081 and not w50229;
w50231 <= not w49466 and not w50080;
w50232 <= not w50079 and w50231;
w50233 <= not w50230 and not w50232;
w50234 <= not b(39) and not w50233;
w50235 <= not w49485 and w49979;
w50236 <= not w49975 and w50235;
w50237 <= not w49976 and not w49979;
w50238 <= not w50236 and not w50237;
w50239 <= not w50081 and not w50238;
w50240 <= not w49475 and not w50080;
w50241 <= not w50079 and w50240;
w50242 <= not w50239 and not w50241;
w50243 <= not b(38) and not w50242;
w50244 <= not w49494 and w49974;
w50245 <= not w49970 and w50244;
w50246 <= not w49971 and not w49974;
w50247 <= not w50245 and not w50246;
w50248 <= not w50081 and not w50247;
w50249 <= not w49484 and not w50080;
w50250 <= not w50079 and w50249;
w50251 <= not w50248 and not w50250;
w50252 <= not b(37) and not w50251;
w50253 <= not w49503 and w49969;
w50254 <= not w49965 and w50253;
w50255 <= not w49966 and not w49969;
w50256 <= not w50254 and not w50255;
w50257 <= not w50081 and not w50256;
w50258 <= not w49493 and not w50080;
w50259 <= not w50079 and w50258;
w50260 <= not w50257 and not w50259;
w50261 <= not b(36) and not w50260;
w50262 <= not w49512 and w49964;
w50263 <= not w49960 and w50262;
w50264 <= not w49961 and not w49964;
w50265 <= not w50263 and not w50264;
w50266 <= not w50081 and not w50265;
w50267 <= not w49502 and not w50080;
w50268 <= not w50079 and w50267;
w50269 <= not w50266 and not w50268;
w50270 <= not b(35) and not w50269;
w50271 <= not w49521 and w49959;
w50272 <= not w49955 and w50271;
w50273 <= not w49956 and not w49959;
w50274 <= not w50272 and not w50273;
w50275 <= not w50081 and not w50274;
w50276 <= not w49511 and not w50080;
w50277 <= not w50079 and w50276;
w50278 <= not w50275 and not w50277;
w50279 <= not b(34) and not w50278;
w50280 <= not w49530 and w49954;
w50281 <= not w49950 and w50280;
w50282 <= not w49951 and not w49954;
w50283 <= not w50281 and not w50282;
w50284 <= not w50081 and not w50283;
w50285 <= not w49520 and not w50080;
w50286 <= not w50079 and w50285;
w50287 <= not w50284 and not w50286;
w50288 <= not b(33) and not w50287;
w50289 <= not w49539 and w49949;
w50290 <= not w49945 and w50289;
w50291 <= not w49946 and not w49949;
w50292 <= not w50290 and not w50291;
w50293 <= not w50081 and not w50292;
w50294 <= not w49529 and not w50080;
w50295 <= not w50079 and w50294;
w50296 <= not w50293 and not w50295;
w50297 <= not b(32) and not w50296;
w50298 <= not w49548 and w49944;
w50299 <= not w49940 and w50298;
w50300 <= not w49941 and not w49944;
w50301 <= not w50299 and not w50300;
w50302 <= not w50081 and not w50301;
w50303 <= not w49538 and not w50080;
w50304 <= not w50079 and w50303;
w50305 <= not w50302 and not w50304;
w50306 <= not b(31) and not w50305;
w50307 <= not w49557 and w49939;
w50308 <= not w49935 and w50307;
w50309 <= not w49936 and not w49939;
w50310 <= not w50308 and not w50309;
w50311 <= not w50081 and not w50310;
w50312 <= not w49547 and not w50080;
w50313 <= not w50079 and w50312;
w50314 <= not w50311 and not w50313;
w50315 <= not b(30) and not w50314;
w50316 <= not w49566 and w49934;
w50317 <= not w49930 and w50316;
w50318 <= not w49931 and not w49934;
w50319 <= not w50317 and not w50318;
w50320 <= not w50081 and not w50319;
w50321 <= not w49556 and not w50080;
w50322 <= not w50079 and w50321;
w50323 <= not w50320 and not w50322;
w50324 <= not b(29) and not w50323;
w50325 <= not w49575 and w49929;
w50326 <= not w49925 and w50325;
w50327 <= not w49926 and not w49929;
w50328 <= not w50326 and not w50327;
w50329 <= not w50081 and not w50328;
w50330 <= not w49565 and not w50080;
w50331 <= not w50079 and w50330;
w50332 <= not w50329 and not w50331;
w50333 <= not b(28) and not w50332;
w50334 <= not w49584 and w49924;
w50335 <= not w49920 and w50334;
w50336 <= not w49921 and not w49924;
w50337 <= not w50335 and not w50336;
w50338 <= not w50081 and not w50337;
w50339 <= not w49574 and not w50080;
w50340 <= not w50079 and w50339;
w50341 <= not w50338 and not w50340;
w50342 <= not b(27) and not w50341;
w50343 <= not w49593 and w49919;
w50344 <= not w49915 and w50343;
w50345 <= not w49916 and not w49919;
w50346 <= not w50344 and not w50345;
w50347 <= not w50081 and not w50346;
w50348 <= not w49583 and not w50080;
w50349 <= not w50079 and w50348;
w50350 <= not w50347 and not w50349;
w50351 <= not b(26) and not w50350;
w50352 <= not w49602 and w49914;
w50353 <= not w49910 and w50352;
w50354 <= not w49911 and not w49914;
w50355 <= not w50353 and not w50354;
w50356 <= not w50081 and not w50355;
w50357 <= not w49592 and not w50080;
w50358 <= not w50079 and w50357;
w50359 <= not w50356 and not w50358;
w50360 <= not b(25) and not w50359;
w50361 <= not w49611 and w49909;
w50362 <= not w49905 and w50361;
w50363 <= not w49906 and not w49909;
w50364 <= not w50362 and not w50363;
w50365 <= not w50081 and not w50364;
w50366 <= not w49601 and not w50080;
w50367 <= not w50079 and w50366;
w50368 <= not w50365 and not w50367;
w50369 <= not b(24) and not w50368;
w50370 <= not w49620 and w49904;
w50371 <= not w49900 and w50370;
w50372 <= not w49901 and not w49904;
w50373 <= not w50371 and not w50372;
w50374 <= not w50081 and not w50373;
w50375 <= not w49610 and not w50080;
w50376 <= not w50079 and w50375;
w50377 <= not w50374 and not w50376;
w50378 <= not b(23) and not w50377;
w50379 <= not w49629 and w49899;
w50380 <= not w49895 and w50379;
w50381 <= not w49896 and not w49899;
w50382 <= not w50380 and not w50381;
w50383 <= not w50081 and not w50382;
w50384 <= not w49619 and not w50080;
w50385 <= not w50079 and w50384;
w50386 <= not w50383 and not w50385;
w50387 <= not b(22) and not w50386;
w50388 <= not w49638 and w49894;
w50389 <= not w49890 and w50388;
w50390 <= not w49891 and not w49894;
w50391 <= not w50389 and not w50390;
w50392 <= not w50081 and not w50391;
w50393 <= not w49628 and not w50080;
w50394 <= not w50079 and w50393;
w50395 <= not w50392 and not w50394;
w50396 <= not b(21) and not w50395;
w50397 <= not w49647 and w49889;
w50398 <= not w49885 and w50397;
w50399 <= not w49886 and not w49889;
w50400 <= not w50398 and not w50399;
w50401 <= not w50081 and not w50400;
w50402 <= not w49637 and not w50080;
w50403 <= not w50079 and w50402;
w50404 <= not w50401 and not w50403;
w50405 <= not b(20) and not w50404;
w50406 <= not w49656 and w49884;
w50407 <= not w49880 and w50406;
w50408 <= not w49881 and not w49884;
w50409 <= not w50407 and not w50408;
w50410 <= not w50081 and not w50409;
w50411 <= not w49646 and not w50080;
w50412 <= not w50079 and w50411;
w50413 <= not w50410 and not w50412;
w50414 <= not b(19) and not w50413;
w50415 <= not w49665 and w49879;
w50416 <= not w49875 and w50415;
w50417 <= not w49876 and not w49879;
w50418 <= not w50416 and not w50417;
w50419 <= not w50081 and not w50418;
w50420 <= not w49655 and not w50080;
w50421 <= not w50079 and w50420;
w50422 <= not w50419 and not w50421;
w50423 <= not b(18) and not w50422;
w50424 <= not w49674 and w49874;
w50425 <= not w49870 and w50424;
w50426 <= not w49871 and not w49874;
w50427 <= not w50425 and not w50426;
w50428 <= not w50081 and not w50427;
w50429 <= not w49664 and not w50080;
w50430 <= not w50079 and w50429;
w50431 <= not w50428 and not w50430;
w50432 <= not b(17) and not w50431;
w50433 <= not w49683 and w49869;
w50434 <= not w49865 and w50433;
w50435 <= not w49866 and not w49869;
w50436 <= not w50434 and not w50435;
w50437 <= not w50081 and not w50436;
w50438 <= not w49673 and not w50080;
w50439 <= not w50079 and w50438;
w50440 <= not w50437 and not w50439;
w50441 <= not b(16) and not w50440;
w50442 <= not w49692 and w49864;
w50443 <= not w49860 and w50442;
w50444 <= not w49861 and not w49864;
w50445 <= not w50443 and not w50444;
w50446 <= not w50081 and not w50445;
w50447 <= not w49682 and not w50080;
w50448 <= not w50079 and w50447;
w50449 <= not w50446 and not w50448;
w50450 <= not b(15) and not w50449;
w50451 <= not w49701 and w49859;
w50452 <= not w49855 and w50451;
w50453 <= not w49856 and not w49859;
w50454 <= not w50452 and not w50453;
w50455 <= not w50081 and not w50454;
w50456 <= not w49691 and not w50080;
w50457 <= not w50079 and w50456;
w50458 <= not w50455 and not w50457;
w50459 <= not b(14) and not w50458;
w50460 <= not w49710 and w49854;
w50461 <= not w49850 and w50460;
w50462 <= not w49851 and not w49854;
w50463 <= not w50461 and not w50462;
w50464 <= not w50081 and not w50463;
w50465 <= not w49700 and not w50080;
w50466 <= not w50079 and w50465;
w50467 <= not w50464 and not w50466;
w50468 <= not b(13) and not w50467;
w50469 <= not w49719 and w49849;
w50470 <= not w49845 and w50469;
w50471 <= not w49846 and not w49849;
w50472 <= not w50470 and not w50471;
w50473 <= not w50081 and not w50472;
w50474 <= not w49709 and not w50080;
w50475 <= not w50079 and w50474;
w50476 <= not w50473 and not w50475;
w50477 <= not b(12) and not w50476;
w50478 <= not w49728 and w49844;
w50479 <= not w49840 and w50478;
w50480 <= not w49841 and not w49844;
w50481 <= not w50479 and not w50480;
w50482 <= not w50081 and not w50481;
w50483 <= not w49718 and not w50080;
w50484 <= not w50079 and w50483;
w50485 <= not w50482 and not w50484;
w50486 <= not b(11) and not w50485;
w50487 <= not w49737 and w49839;
w50488 <= not w49835 and w50487;
w50489 <= not w49836 and not w49839;
w50490 <= not w50488 and not w50489;
w50491 <= not w50081 and not w50490;
w50492 <= not w49727 and not w50080;
w50493 <= not w50079 and w50492;
w50494 <= not w50491 and not w50493;
w50495 <= not b(10) and not w50494;
w50496 <= not w49746 and w49834;
w50497 <= not w49830 and w50496;
w50498 <= not w49831 and not w49834;
w50499 <= not w50497 and not w50498;
w50500 <= not w50081 and not w50499;
w50501 <= not w49736 and not w50080;
w50502 <= not w50079 and w50501;
w50503 <= not w50500 and not w50502;
w50504 <= not b(9) and not w50503;
w50505 <= not w49755 and w49829;
w50506 <= not w49825 and w50505;
w50507 <= not w49826 and not w49829;
w50508 <= not w50506 and not w50507;
w50509 <= not w50081 and not w50508;
w50510 <= not w49745 and not w50080;
w50511 <= not w50079 and w50510;
w50512 <= not w50509 and not w50511;
w50513 <= not b(8) and not w50512;
w50514 <= not w49764 and w49824;
w50515 <= not w49820 and w50514;
w50516 <= not w49821 and not w49824;
w50517 <= not w50515 and not w50516;
w50518 <= not w50081 and not w50517;
w50519 <= not w49754 and not w50080;
w50520 <= not w50079 and w50519;
w50521 <= not w50518 and not w50520;
w50522 <= not b(7) and not w50521;
w50523 <= not w49773 and w49819;
w50524 <= not w49815 and w50523;
w50525 <= not w49816 and not w49819;
w50526 <= not w50524 and not w50525;
w50527 <= not w50081 and not w50526;
w50528 <= not w49763 and not w50080;
w50529 <= not w50079 and w50528;
w50530 <= not w50527 and not w50529;
w50531 <= not b(6) and not w50530;
w50532 <= not w49782 and w49814;
w50533 <= not w49810 and w50532;
w50534 <= not w49811 and not w49814;
w50535 <= not w50533 and not w50534;
w50536 <= not w50081 and not w50535;
w50537 <= not w49772 and not w50080;
w50538 <= not w50079 and w50537;
w50539 <= not w50536 and not w50538;
w50540 <= not b(5) and not w50539;
w50541 <= not w49790 and w49809;
w50542 <= not w49805 and w50541;
w50543 <= not w49806 and not w49809;
w50544 <= not w50542 and not w50543;
w50545 <= not w50081 and not w50544;
w50546 <= not w49781 and not w50080;
w50547 <= not w50079 and w50546;
w50548 <= not w50545 and not w50547;
w50549 <= not b(4) and not w50548;
w50550 <= not w49800 and w49804;
w50551 <= not w49799 and w50550;
w50552 <= not w49801 and not w49804;
w50553 <= not w50551 and not w50552;
w50554 <= not w50081 and not w50553;
w50555 <= not w49789 and not w50080;
w50556 <= not w50079 and w50555;
w50557 <= not w50554 and not w50556;
w50558 <= not b(3) and not w50557;
w50559 <= w21772 and not w49797;
w50560 <= not w49795 and w50559;
w50561 <= not w49799 and not w50560;
w50562 <= not w50081 and w50561;
w50563 <= not w49794 and not w50080;
w50564 <= not w50079 and w50563;
w50565 <= not w50562 and not w50564;
w50566 <= not b(2) and not w50565;
w50567 <= b(0) and not w50081;
w50568 <= a(8) and not w50567;
w50569 <= w21772 and not w50081;
w50570 <= not w50568 and not w50569;
w50571 <= b(1) and not w50570;
w50572 <= not b(1) and not w50569;
w50573 <= not w50568 and w50572;
w50574 <= not w50571 and not w50573;
w50575 <= not w22549 and not w50574;
w50576 <= not b(1) and not w50570;
w50577 <= not w50575 and not w50576;
w50578 <= b(2) and not w50564;
w50579 <= not w50562 and w50578;
w50580 <= not w50566 and not w50579;
w50581 <= not w50577 and w50580;
w50582 <= not w50566 and not w50581;
w50583 <= b(3) and not w50556;
w50584 <= not w50554 and w50583;
w50585 <= not w50558 and not w50584;
w50586 <= not w50582 and w50585;
w50587 <= not w50558 and not w50586;
w50588 <= b(4) and not w50547;
w50589 <= not w50545 and w50588;
w50590 <= not w50549 and not w50589;
w50591 <= not w50587 and w50590;
w50592 <= not w50549 and not w50591;
w50593 <= b(5) and not w50538;
w50594 <= not w50536 and w50593;
w50595 <= not w50540 and not w50594;
w50596 <= not w50592 and w50595;
w50597 <= not w50540 and not w50596;
w50598 <= b(6) and not w50529;
w50599 <= not w50527 and w50598;
w50600 <= not w50531 and not w50599;
w50601 <= not w50597 and w50600;
w50602 <= not w50531 and not w50601;
w50603 <= b(7) and not w50520;
w50604 <= not w50518 and w50603;
w50605 <= not w50522 and not w50604;
w50606 <= not w50602 and w50605;
w50607 <= not w50522 and not w50606;
w50608 <= b(8) and not w50511;
w50609 <= not w50509 and w50608;
w50610 <= not w50513 and not w50609;
w50611 <= not w50607 and w50610;
w50612 <= not w50513 and not w50611;
w50613 <= b(9) and not w50502;
w50614 <= not w50500 and w50613;
w50615 <= not w50504 and not w50614;
w50616 <= not w50612 and w50615;
w50617 <= not w50504 and not w50616;
w50618 <= b(10) and not w50493;
w50619 <= not w50491 and w50618;
w50620 <= not w50495 and not w50619;
w50621 <= not w50617 and w50620;
w50622 <= not w50495 and not w50621;
w50623 <= b(11) and not w50484;
w50624 <= not w50482 and w50623;
w50625 <= not w50486 and not w50624;
w50626 <= not w50622 and w50625;
w50627 <= not w50486 and not w50626;
w50628 <= b(12) and not w50475;
w50629 <= not w50473 and w50628;
w50630 <= not w50477 and not w50629;
w50631 <= not w50627 and w50630;
w50632 <= not w50477 and not w50631;
w50633 <= b(13) and not w50466;
w50634 <= not w50464 and w50633;
w50635 <= not w50468 and not w50634;
w50636 <= not w50632 and w50635;
w50637 <= not w50468 and not w50636;
w50638 <= b(14) and not w50457;
w50639 <= not w50455 and w50638;
w50640 <= not w50459 and not w50639;
w50641 <= not w50637 and w50640;
w50642 <= not w50459 and not w50641;
w50643 <= b(15) and not w50448;
w50644 <= not w50446 and w50643;
w50645 <= not w50450 and not w50644;
w50646 <= not w50642 and w50645;
w50647 <= not w50450 and not w50646;
w50648 <= b(16) and not w50439;
w50649 <= not w50437 and w50648;
w50650 <= not w50441 and not w50649;
w50651 <= not w50647 and w50650;
w50652 <= not w50441 and not w50651;
w50653 <= b(17) and not w50430;
w50654 <= not w50428 and w50653;
w50655 <= not w50432 and not w50654;
w50656 <= not w50652 and w50655;
w50657 <= not w50432 and not w50656;
w50658 <= b(18) and not w50421;
w50659 <= not w50419 and w50658;
w50660 <= not w50423 and not w50659;
w50661 <= not w50657 and w50660;
w50662 <= not w50423 and not w50661;
w50663 <= b(19) and not w50412;
w50664 <= not w50410 and w50663;
w50665 <= not w50414 and not w50664;
w50666 <= not w50662 and w50665;
w50667 <= not w50414 and not w50666;
w50668 <= b(20) and not w50403;
w50669 <= not w50401 and w50668;
w50670 <= not w50405 and not w50669;
w50671 <= not w50667 and w50670;
w50672 <= not w50405 and not w50671;
w50673 <= b(21) and not w50394;
w50674 <= not w50392 and w50673;
w50675 <= not w50396 and not w50674;
w50676 <= not w50672 and w50675;
w50677 <= not w50396 and not w50676;
w50678 <= b(22) and not w50385;
w50679 <= not w50383 and w50678;
w50680 <= not w50387 and not w50679;
w50681 <= not w50677 and w50680;
w50682 <= not w50387 and not w50681;
w50683 <= b(23) and not w50376;
w50684 <= not w50374 and w50683;
w50685 <= not w50378 and not w50684;
w50686 <= not w50682 and w50685;
w50687 <= not w50378 and not w50686;
w50688 <= b(24) and not w50367;
w50689 <= not w50365 and w50688;
w50690 <= not w50369 and not w50689;
w50691 <= not w50687 and w50690;
w50692 <= not w50369 and not w50691;
w50693 <= b(25) and not w50358;
w50694 <= not w50356 and w50693;
w50695 <= not w50360 and not w50694;
w50696 <= not w50692 and w50695;
w50697 <= not w50360 and not w50696;
w50698 <= b(26) and not w50349;
w50699 <= not w50347 and w50698;
w50700 <= not w50351 and not w50699;
w50701 <= not w50697 and w50700;
w50702 <= not w50351 and not w50701;
w50703 <= b(27) and not w50340;
w50704 <= not w50338 and w50703;
w50705 <= not w50342 and not w50704;
w50706 <= not w50702 and w50705;
w50707 <= not w50342 and not w50706;
w50708 <= b(28) and not w50331;
w50709 <= not w50329 and w50708;
w50710 <= not w50333 and not w50709;
w50711 <= not w50707 and w50710;
w50712 <= not w50333 and not w50711;
w50713 <= b(29) and not w50322;
w50714 <= not w50320 and w50713;
w50715 <= not w50324 and not w50714;
w50716 <= not w50712 and w50715;
w50717 <= not w50324 and not w50716;
w50718 <= b(30) and not w50313;
w50719 <= not w50311 and w50718;
w50720 <= not w50315 and not w50719;
w50721 <= not w50717 and w50720;
w50722 <= not w50315 and not w50721;
w50723 <= b(31) and not w50304;
w50724 <= not w50302 and w50723;
w50725 <= not w50306 and not w50724;
w50726 <= not w50722 and w50725;
w50727 <= not w50306 and not w50726;
w50728 <= b(32) and not w50295;
w50729 <= not w50293 and w50728;
w50730 <= not w50297 and not w50729;
w50731 <= not w50727 and w50730;
w50732 <= not w50297 and not w50731;
w50733 <= b(33) and not w50286;
w50734 <= not w50284 and w50733;
w50735 <= not w50288 and not w50734;
w50736 <= not w50732 and w50735;
w50737 <= not w50288 and not w50736;
w50738 <= b(34) and not w50277;
w50739 <= not w50275 and w50738;
w50740 <= not w50279 and not w50739;
w50741 <= not w50737 and w50740;
w50742 <= not w50279 and not w50741;
w50743 <= b(35) and not w50268;
w50744 <= not w50266 and w50743;
w50745 <= not w50270 and not w50744;
w50746 <= not w50742 and w50745;
w50747 <= not w50270 and not w50746;
w50748 <= b(36) and not w50259;
w50749 <= not w50257 and w50748;
w50750 <= not w50261 and not w50749;
w50751 <= not w50747 and w50750;
w50752 <= not w50261 and not w50751;
w50753 <= b(37) and not w50250;
w50754 <= not w50248 and w50753;
w50755 <= not w50252 and not w50754;
w50756 <= not w50752 and w50755;
w50757 <= not w50252 and not w50756;
w50758 <= b(38) and not w50241;
w50759 <= not w50239 and w50758;
w50760 <= not w50243 and not w50759;
w50761 <= not w50757 and w50760;
w50762 <= not w50243 and not w50761;
w50763 <= b(39) and not w50232;
w50764 <= not w50230 and w50763;
w50765 <= not w50234 and not w50764;
w50766 <= not w50762 and w50765;
w50767 <= not w50234 and not w50766;
w50768 <= b(40) and not w50223;
w50769 <= not w50221 and w50768;
w50770 <= not w50225 and not w50769;
w50771 <= not w50767 and w50770;
w50772 <= not w50225 and not w50771;
w50773 <= b(41) and not w50214;
w50774 <= not w50212 and w50773;
w50775 <= not w50216 and not w50774;
w50776 <= not w50772 and w50775;
w50777 <= not w50216 and not w50776;
w50778 <= b(42) and not w50205;
w50779 <= not w50203 and w50778;
w50780 <= not w50207 and not w50779;
w50781 <= not w50777 and w50780;
w50782 <= not w50207 and not w50781;
w50783 <= b(43) and not w50196;
w50784 <= not w50194 and w50783;
w50785 <= not w50198 and not w50784;
w50786 <= not w50782 and w50785;
w50787 <= not w50198 and not w50786;
w50788 <= b(44) and not w50187;
w50789 <= not w50185 and w50788;
w50790 <= not w50189 and not w50789;
w50791 <= not w50787 and w50790;
w50792 <= not w50189 and not w50791;
w50793 <= b(45) and not w50178;
w50794 <= not w50176 and w50793;
w50795 <= not w50180 and not w50794;
w50796 <= not w50792 and w50795;
w50797 <= not w50180 and not w50796;
w50798 <= b(46) and not w50169;
w50799 <= not w50167 and w50798;
w50800 <= not w50171 and not w50799;
w50801 <= not w50797 and w50800;
w50802 <= not w50171 and not w50801;
w50803 <= b(47) and not w50160;
w50804 <= not w50158 and w50803;
w50805 <= not w50162 and not w50804;
w50806 <= not w50802 and w50805;
w50807 <= not w50162 and not w50806;
w50808 <= b(48) and not w50151;
w50809 <= not w50149 and w50808;
w50810 <= not w50153 and not w50809;
w50811 <= not w50807 and w50810;
w50812 <= not w50153 and not w50811;
w50813 <= b(49) and not w50142;
w50814 <= not w50140 and w50813;
w50815 <= not w50144 and not w50814;
w50816 <= not w50812 and w50815;
w50817 <= not w50144 and not w50816;
w50818 <= b(50) and not w50133;
w50819 <= not w50131 and w50818;
w50820 <= not w50135 and not w50819;
w50821 <= not w50817 and w50820;
w50822 <= not w50135 and not w50821;
w50823 <= b(51) and not w50124;
w50824 <= not w50122 and w50823;
w50825 <= not w50126 and not w50824;
w50826 <= not w50822 and w50825;
w50827 <= not w50126 and not w50826;
w50828 <= b(52) and not w50115;
w50829 <= not w50113 and w50828;
w50830 <= not w50117 and not w50829;
w50831 <= not w50827 and w50830;
w50832 <= not w50117 and not w50831;
w50833 <= b(53) and not w50106;
w50834 <= not w50104 and w50833;
w50835 <= not w50108 and not w50834;
w50836 <= not w50832 and w50835;
w50837 <= not w50108 and not w50836;
w50838 <= b(54) and not w50097;
w50839 <= not w50095 and w50838;
w50840 <= not w50099 and not w50839;
w50841 <= not w50837 and w50840;
w50842 <= not w50099 and not w50841;
w50843 <= b(55) and not w50088;
w50844 <= not w50086 and w50843;
w50845 <= not w50090 and not w50844;
w50846 <= not w50842 and w50845;
w50847 <= not w50090 and not w50846;
w50848 <= not w49323 and not w50076;
w50849 <= not w50074 and w50848;
w50850 <= not w50065 and w50849;
w50851 <= not w50074 and not w50076;
w50852 <= not w50066 and not w50851;
w50853 <= not w50850 and not w50852;
w50854 <= not w50081 and not w50853;
w50855 <= not w50073 and not w50080;
w50856 <= not w50079 and w50855;
w50857 <= not w50854 and not w50856;
w50858 <= not b(56) and not w50857;
w50859 <= b(56) and not w50856;
w50860 <= not w50854 and w50859;
w50861 <= w150 and not w50860;
w50862 <= not w50858 and w50861;
w50863 <= not w50847 and w50862;
w50864 <= w80 and not w50857;
w50865 <= not w50863 and not w50864;
w50866 <= not w50099 and w50845;
w50867 <= not w50841 and w50866;
w50868 <= not w50842 and not w50845;
w50869 <= not w50867 and not w50868;
w50870 <= not w50865 and not w50869;
w50871 <= not w50089 and not w50864;
w50872 <= not w50863 and w50871;
w50873 <= not w50870 and not w50872;
w50874 <= not w50090 and not w50860;
w50875 <= not w50858 and w50874;
w50876 <= not w50846 and w50875;
w50877 <= not w50858 and not w50860;
w50878 <= not w50847 and not w50877;
w50879 <= not w50876 and not w50878;
w50880 <= not w50865 and not w50879;
w50881 <= not w50857 and not w50864;
w50882 <= not w50863 and w50881;
w50883 <= not w50880 and not w50882;
w50884 <= not b(57) and not w50883;
w50885 <= not b(56) and not w50873;
w50886 <= not w50108 and w50840;
w50887 <= not w50836 and w50886;
w50888 <= not w50837 and not w50840;
w50889 <= not w50887 and not w50888;
w50890 <= not w50865 and not w50889;
w50891 <= not w50098 and not w50864;
w50892 <= not w50863 and w50891;
w50893 <= not w50890 and not w50892;
w50894 <= not b(55) and not w50893;
w50895 <= not w50117 and w50835;
w50896 <= not w50831 and w50895;
w50897 <= not w50832 and not w50835;
w50898 <= not w50896 and not w50897;
w50899 <= not w50865 and not w50898;
w50900 <= not w50107 and not w50864;
w50901 <= not w50863 and w50900;
w50902 <= not w50899 and not w50901;
w50903 <= not b(54) and not w50902;
w50904 <= not w50126 and w50830;
w50905 <= not w50826 and w50904;
w50906 <= not w50827 and not w50830;
w50907 <= not w50905 and not w50906;
w50908 <= not w50865 and not w50907;
w50909 <= not w50116 and not w50864;
w50910 <= not w50863 and w50909;
w50911 <= not w50908 and not w50910;
w50912 <= not b(53) and not w50911;
w50913 <= not w50135 and w50825;
w50914 <= not w50821 and w50913;
w50915 <= not w50822 and not w50825;
w50916 <= not w50914 and not w50915;
w50917 <= not w50865 and not w50916;
w50918 <= not w50125 and not w50864;
w50919 <= not w50863 and w50918;
w50920 <= not w50917 and not w50919;
w50921 <= not b(52) and not w50920;
w50922 <= not w50144 and w50820;
w50923 <= not w50816 and w50922;
w50924 <= not w50817 and not w50820;
w50925 <= not w50923 and not w50924;
w50926 <= not w50865 and not w50925;
w50927 <= not w50134 and not w50864;
w50928 <= not w50863 and w50927;
w50929 <= not w50926 and not w50928;
w50930 <= not b(51) and not w50929;
w50931 <= not w50153 and w50815;
w50932 <= not w50811 and w50931;
w50933 <= not w50812 and not w50815;
w50934 <= not w50932 and not w50933;
w50935 <= not w50865 and not w50934;
w50936 <= not w50143 and not w50864;
w50937 <= not w50863 and w50936;
w50938 <= not w50935 and not w50937;
w50939 <= not b(50) and not w50938;
w50940 <= not w50162 and w50810;
w50941 <= not w50806 and w50940;
w50942 <= not w50807 and not w50810;
w50943 <= not w50941 and not w50942;
w50944 <= not w50865 and not w50943;
w50945 <= not w50152 and not w50864;
w50946 <= not w50863 and w50945;
w50947 <= not w50944 and not w50946;
w50948 <= not b(49) and not w50947;
w50949 <= not w50171 and w50805;
w50950 <= not w50801 and w50949;
w50951 <= not w50802 and not w50805;
w50952 <= not w50950 and not w50951;
w50953 <= not w50865 and not w50952;
w50954 <= not w50161 and not w50864;
w50955 <= not w50863 and w50954;
w50956 <= not w50953 and not w50955;
w50957 <= not b(48) and not w50956;
w50958 <= not w50180 and w50800;
w50959 <= not w50796 and w50958;
w50960 <= not w50797 and not w50800;
w50961 <= not w50959 and not w50960;
w50962 <= not w50865 and not w50961;
w50963 <= not w50170 and not w50864;
w50964 <= not w50863 and w50963;
w50965 <= not w50962 and not w50964;
w50966 <= not b(47) and not w50965;
w50967 <= not w50189 and w50795;
w50968 <= not w50791 and w50967;
w50969 <= not w50792 and not w50795;
w50970 <= not w50968 and not w50969;
w50971 <= not w50865 and not w50970;
w50972 <= not w50179 and not w50864;
w50973 <= not w50863 and w50972;
w50974 <= not w50971 and not w50973;
w50975 <= not b(46) and not w50974;
w50976 <= not w50198 and w50790;
w50977 <= not w50786 and w50976;
w50978 <= not w50787 and not w50790;
w50979 <= not w50977 and not w50978;
w50980 <= not w50865 and not w50979;
w50981 <= not w50188 and not w50864;
w50982 <= not w50863 and w50981;
w50983 <= not w50980 and not w50982;
w50984 <= not b(45) and not w50983;
w50985 <= not w50207 and w50785;
w50986 <= not w50781 and w50985;
w50987 <= not w50782 and not w50785;
w50988 <= not w50986 and not w50987;
w50989 <= not w50865 and not w50988;
w50990 <= not w50197 and not w50864;
w50991 <= not w50863 and w50990;
w50992 <= not w50989 and not w50991;
w50993 <= not b(44) and not w50992;
w50994 <= not w50216 and w50780;
w50995 <= not w50776 and w50994;
w50996 <= not w50777 and not w50780;
w50997 <= not w50995 and not w50996;
w50998 <= not w50865 and not w50997;
w50999 <= not w50206 and not w50864;
w51000 <= not w50863 and w50999;
w51001 <= not w50998 and not w51000;
w51002 <= not b(43) and not w51001;
w51003 <= not w50225 and w50775;
w51004 <= not w50771 and w51003;
w51005 <= not w50772 and not w50775;
w51006 <= not w51004 and not w51005;
w51007 <= not w50865 and not w51006;
w51008 <= not w50215 and not w50864;
w51009 <= not w50863 and w51008;
w51010 <= not w51007 and not w51009;
w51011 <= not b(42) and not w51010;
w51012 <= not w50234 and w50770;
w51013 <= not w50766 and w51012;
w51014 <= not w50767 and not w50770;
w51015 <= not w51013 and not w51014;
w51016 <= not w50865 and not w51015;
w51017 <= not w50224 and not w50864;
w51018 <= not w50863 and w51017;
w51019 <= not w51016 and not w51018;
w51020 <= not b(41) and not w51019;
w51021 <= not w50243 and w50765;
w51022 <= not w50761 and w51021;
w51023 <= not w50762 and not w50765;
w51024 <= not w51022 and not w51023;
w51025 <= not w50865 and not w51024;
w51026 <= not w50233 and not w50864;
w51027 <= not w50863 and w51026;
w51028 <= not w51025 and not w51027;
w51029 <= not b(40) and not w51028;
w51030 <= not w50252 and w50760;
w51031 <= not w50756 and w51030;
w51032 <= not w50757 and not w50760;
w51033 <= not w51031 and not w51032;
w51034 <= not w50865 and not w51033;
w51035 <= not w50242 and not w50864;
w51036 <= not w50863 and w51035;
w51037 <= not w51034 and not w51036;
w51038 <= not b(39) and not w51037;
w51039 <= not w50261 and w50755;
w51040 <= not w50751 and w51039;
w51041 <= not w50752 and not w50755;
w51042 <= not w51040 and not w51041;
w51043 <= not w50865 and not w51042;
w51044 <= not w50251 and not w50864;
w51045 <= not w50863 and w51044;
w51046 <= not w51043 and not w51045;
w51047 <= not b(38) and not w51046;
w51048 <= not w50270 and w50750;
w51049 <= not w50746 and w51048;
w51050 <= not w50747 and not w50750;
w51051 <= not w51049 and not w51050;
w51052 <= not w50865 and not w51051;
w51053 <= not w50260 and not w50864;
w51054 <= not w50863 and w51053;
w51055 <= not w51052 and not w51054;
w51056 <= not b(37) and not w51055;
w51057 <= not w50279 and w50745;
w51058 <= not w50741 and w51057;
w51059 <= not w50742 and not w50745;
w51060 <= not w51058 and not w51059;
w51061 <= not w50865 and not w51060;
w51062 <= not w50269 and not w50864;
w51063 <= not w50863 and w51062;
w51064 <= not w51061 and not w51063;
w51065 <= not b(36) and not w51064;
w51066 <= not w50288 and w50740;
w51067 <= not w50736 and w51066;
w51068 <= not w50737 and not w50740;
w51069 <= not w51067 and not w51068;
w51070 <= not w50865 and not w51069;
w51071 <= not w50278 and not w50864;
w51072 <= not w50863 and w51071;
w51073 <= not w51070 and not w51072;
w51074 <= not b(35) and not w51073;
w51075 <= not w50297 and w50735;
w51076 <= not w50731 and w51075;
w51077 <= not w50732 and not w50735;
w51078 <= not w51076 and not w51077;
w51079 <= not w50865 and not w51078;
w51080 <= not w50287 and not w50864;
w51081 <= not w50863 and w51080;
w51082 <= not w51079 and not w51081;
w51083 <= not b(34) and not w51082;
w51084 <= not w50306 and w50730;
w51085 <= not w50726 and w51084;
w51086 <= not w50727 and not w50730;
w51087 <= not w51085 and not w51086;
w51088 <= not w50865 and not w51087;
w51089 <= not w50296 and not w50864;
w51090 <= not w50863 and w51089;
w51091 <= not w51088 and not w51090;
w51092 <= not b(33) and not w51091;
w51093 <= not w50315 and w50725;
w51094 <= not w50721 and w51093;
w51095 <= not w50722 and not w50725;
w51096 <= not w51094 and not w51095;
w51097 <= not w50865 and not w51096;
w51098 <= not w50305 and not w50864;
w51099 <= not w50863 and w51098;
w51100 <= not w51097 and not w51099;
w51101 <= not b(32) and not w51100;
w51102 <= not w50324 and w50720;
w51103 <= not w50716 and w51102;
w51104 <= not w50717 and not w50720;
w51105 <= not w51103 and not w51104;
w51106 <= not w50865 and not w51105;
w51107 <= not w50314 and not w50864;
w51108 <= not w50863 and w51107;
w51109 <= not w51106 and not w51108;
w51110 <= not b(31) and not w51109;
w51111 <= not w50333 and w50715;
w51112 <= not w50711 and w51111;
w51113 <= not w50712 and not w50715;
w51114 <= not w51112 and not w51113;
w51115 <= not w50865 and not w51114;
w51116 <= not w50323 and not w50864;
w51117 <= not w50863 and w51116;
w51118 <= not w51115 and not w51117;
w51119 <= not b(30) and not w51118;
w51120 <= not w50342 and w50710;
w51121 <= not w50706 and w51120;
w51122 <= not w50707 and not w50710;
w51123 <= not w51121 and not w51122;
w51124 <= not w50865 and not w51123;
w51125 <= not w50332 and not w50864;
w51126 <= not w50863 and w51125;
w51127 <= not w51124 and not w51126;
w51128 <= not b(29) and not w51127;
w51129 <= not w50351 and w50705;
w51130 <= not w50701 and w51129;
w51131 <= not w50702 and not w50705;
w51132 <= not w51130 and not w51131;
w51133 <= not w50865 and not w51132;
w51134 <= not w50341 and not w50864;
w51135 <= not w50863 and w51134;
w51136 <= not w51133 and not w51135;
w51137 <= not b(28) and not w51136;
w51138 <= not w50360 and w50700;
w51139 <= not w50696 and w51138;
w51140 <= not w50697 and not w50700;
w51141 <= not w51139 and not w51140;
w51142 <= not w50865 and not w51141;
w51143 <= not w50350 and not w50864;
w51144 <= not w50863 and w51143;
w51145 <= not w51142 and not w51144;
w51146 <= not b(27) and not w51145;
w51147 <= not w50369 and w50695;
w51148 <= not w50691 and w51147;
w51149 <= not w50692 and not w50695;
w51150 <= not w51148 and not w51149;
w51151 <= not w50865 and not w51150;
w51152 <= not w50359 and not w50864;
w51153 <= not w50863 and w51152;
w51154 <= not w51151 and not w51153;
w51155 <= not b(26) and not w51154;
w51156 <= not w50378 and w50690;
w51157 <= not w50686 and w51156;
w51158 <= not w50687 and not w50690;
w51159 <= not w51157 and not w51158;
w51160 <= not w50865 and not w51159;
w51161 <= not w50368 and not w50864;
w51162 <= not w50863 and w51161;
w51163 <= not w51160 and not w51162;
w51164 <= not b(25) and not w51163;
w51165 <= not w50387 and w50685;
w51166 <= not w50681 and w51165;
w51167 <= not w50682 and not w50685;
w51168 <= not w51166 and not w51167;
w51169 <= not w50865 and not w51168;
w51170 <= not w50377 and not w50864;
w51171 <= not w50863 and w51170;
w51172 <= not w51169 and not w51171;
w51173 <= not b(24) and not w51172;
w51174 <= not w50396 and w50680;
w51175 <= not w50676 and w51174;
w51176 <= not w50677 and not w50680;
w51177 <= not w51175 and not w51176;
w51178 <= not w50865 and not w51177;
w51179 <= not w50386 and not w50864;
w51180 <= not w50863 and w51179;
w51181 <= not w51178 and not w51180;
w51182 <= not b(23) and not w51181;
w51183 <= not w50405 and w50675;
w51184 <= not w50671 and w51183;
w51185 <= not w50672 and not w50675;
w51186 <= not w51184 and not w51185;
w51187 <= not w50865 and not w51186;
w51188 <= not w50395 and not w50864;
w51189 <= not w50863 and w51188;
w51190 <= not w51187 and not w51189;
w51191 <= not b(22) and not w51190;
w51192 <= not w50414 and w50670;
w51193 <= not w50666 and w51192;
w51194 <= not w50667 and not w50670;
w51195 <= not w51193 and not w51194;
w51196 <= not w50865 and not w51195;
w51197 <= not w50404 and not w50864;
w51198 <= not w50863 and w51197;
w51199 <= not w51196 and not w51198;
w51200 <= not b(21) and not w51199;
w51201 <= not w50423 and w50665;
w51202 <= not w50661 and w51201;
w51203 <= not w50662 and not w50665;
w51204 <= not w51202 and not w51203;
w51205 <= not w50865 and not w51204;
w51206 <= not w50413 and not w50864;
w51207 <= not w50863 and w51206;
w51208 <= not w51205 and not w51207;
w51209 <= not b(20) and not w51208;
w51210 <= not w50432 and w50660;
w51211 <= not w50656 and w51210;
w51212 <= not w50657 and not w50660;
w51213 <= not w51211 and not w51212;
w51214 <= not w50865 and not w51213;
w51215 <= not w50422 and not w50864;
w51216 <= not w50863 and w51215;
w51217 <= not w51214 and not w51216;
w51218 <= not b(19) and not w51217;
w51219 <= not w50441 and w50655;
w51220 <= not w50651 and w51219;
w51221 <= not w50652 and not w50655;
w51222 <= not w51220 and not w51221;
w51223 <= not w50865 and not w51222;
w51224 <= not w50431 and not w50864;
w51225 <= not w50863 and w51224;
w51226 <= not w51223 and not w51225;
w51227 <= not b(18) and not w51226;
w51228 <= not w50450 and w50650;
w51229 <= not w50646 and w51228;
w51230 <= not w50647 and not w50650;
w51231 <= not w51229 and not w51230;
w51232 <= not w50865 and not w51231;
w51233 <= not w50440 and not w50864;
w51234 <= not w50863 and w51233;
w51235 <= not w51232 and not w51234;
w51236 <= not b(17) and not w51235;
w51237 <= not w50459 and w50645;
w51238 <= not w50641 and w51237;
w51239 <= not w50642 and not w50645;
w51240 <= not w51238 and not w51239;
w51241 <= not w50865 and not w51240;
w51242 <= not w50449 and not w50864;
w51243 <= not w50863 and w51242;
w51244 <= not w51241 and not w51243;
w51245 <= not b(16) and not w51244;
w51246 <= not w50468 and w50640;
w51247 <= not w50636 and w51246;
w51248 <= not w50637 and not w50640;
w51249 <= not w51247 and not w51248;
w51250 <= not w50865 and not w51249;
w51251 <= not w50458 and not w50864;
w51252 <= not w50863 and w51251;
w51253 <= not w51250 and not w51252;
w51254 <= not b(15) and not w51253;
w51255 <= not w50477 and w50635;
w51256 <= not w50631 and w51255;
w51257 <= not w50632 and not w50635;
w51258 <= not w51256 and not w51257;
w51259 <= not w50865 and not w51258;
w51260 <= not w50467 and not w50864;
w51261 <= not w50863 and w51260;
w51262 <= not w51259 and not w51261;
w51263 <= not b(14) and not w51262;
w51264 <= not w50486 and w50630;
w51265 <= not w50626 and w51264;
w51266 <= not w50627 and not w50630;
w51267 <= not w51265 and not w51266;
w51268 <= not w50865 and not w51267;
w51269 <= not w50476 and not w50864;
w51270 <= not w50863 and w51269;
w51271 <= not w51268 and not w51270;
w51272 <= not b(13) and not w51271;
w51273 <= not w50495 and w50625;
w51274 <= not w50621 and w51273;
w51275 <= not w50622 and not w50625;
w51276 <= not w51274 and not w51275;
w51277 <= not w50865 and not w51276;
w51278 <= not w50485 and not w50864;
w51279 <= not w50863 and w51278;
w51280 <= not w51277 and not w51279;
w51281 <= not b(12) and not w51280;
w51282 <= not w50504 and w50620;
w51283 <= not w50616 and w51282;
w51284 <= not w50617 and not w50620;
w51285 <= not w51283 and not w51284;
w51286 <= not w50865 and not w51285;
w51287 <= not w50494 and not w50864;
w51288 <= not w50863 and w51287;
w51289 <= not w51286 and not w51288;
w51290 <= not b(11) and not w51289;
w51291 <= not w50513 and w50615;
w51292 <= not w50611 and w51291;
w51293 <= not w50612 and not w50615;
w51294 <= not w51292 and not w51293;
w51295 <= not w50865 and not w51294;
w51296 <= not w50503 and not w50864;
w51297 <= not w50863 and w51296;
w51298 <= not w51295 and not w51297;
w51299 <= not b(10) and not w51298;
w51300 <= not w50522 and w50610;
w51301 <= not w50606 and w51300;
w51302 <= not w50607 and not w50610;
w51303 <= not w51301 and not w51302;
w51304 <= not w50865 and not w51303;
w51305 <= not w50512 and not w50864;
w51306 <= not w50863 and w51305;
w51307 <= not w51304 and not w51306;
w51308 <= not b(9) and not w51307;
w51309 <= not w50531 and w50605;
w51310 <= not w50601 and w51309;
w51311 <= not w50602 and not w50605;
w51312 <= not w51310 and not w51311;
w51313 <= not w50865 and not w51312;
w51314 <= not w50521 and not w50864;
w51315 <= not w50863 and w51314;
w51316 <= not w51313 and not w51315;
w51317 <= not b(8) and not w51316;
w51318 <= not w50540 and w50600;
w51319 <= not w50596 and w51318;
w51320 <= not w50597 and not w50600;
w51321 <= not w51319 and not w51320;
w51322 <= not w50865 and not w51321;
w51323 <= not w50530 and not w50864;
w51324 <= not w50863 and w51323;
w51325 <= not w51322 and not w51324;
w51326 <= not b(7) and not w51325;
w51327 <= not w50549 and w50595;
w51328 <= not w50591 and w51327;
w51329 <= not w50592 and not w50595;
w51330 <= not w51328 and not w51329;
w51331 <= not w50865 and not w51330;
w51332 <= not w50539 and not w50864;
w51333 <= not w50863 and w51332;
w51334 <= not w51331 and not w51333;
w51335 <= not b(6) and not w51334;
w51336 <= not w50558 and w50590;
w51337 <= not w50586 and w51336;
w51338 <= not w50587 and not w50590;
w51339 <= not w51337 and not w51338;
w51340 <= not w50865 and not w51339;
w51341 <= not w50548 and not w50864;
w51342 <= not w50863 and w51341;
w51343 <= not w51340 and not w51342;
w51344 <= not b(5) and not w51343;
w51345 <= not w50566 and w50585;
w51346 <= not w50581 and w51345;
w51347 <= not w50582 and not w50585;
w51348 <= not w51346 and not w51347;
w51349 <= not w50865 and not w51348;
w51350 <= not w50557 and not w50864;
w51351 <= not w50863 and w51350;
w51352 <= not w51349 and not w51351;
w51353 <= not b(4) and not w51352;
w51354 <= not w50576 and w50580;
w51355 <= not w50575 and w51354;
w51356 <= not w50577 and not w50580;
w51357 <= not w51355 and not w51356;
w51358 <= not w50865 and not w51357;
w51359 <= not w50565 and not w50864;
w51360 <= not w50863 and w51359;
w51361 <= not w51358 and not w51360;
w51362 <= not b(3) and not w51361;
w51363 <= w22549 and not w50573;
w51364 <= not w50571 and w51363;
w51365 <= not w50575 and not w51364;
w51366 <= not w50865 and w51365;
w51367 <= not w50570 and not w50864;
w51368 <= not w50863 and w51367;
w51369 <= not w51366 and not w51368;
w51370 <= not b(2) and not w51369;
w51371 <= b(0) and not w50865;
w51372 <= a(7) and not w51371;
w51373 <= w22549 and not w50865;
w51374 <= not w51372 and not w51373;
w51375 <= b(1) and not w51374;
w51376 <= not b(1) and not w51373;
w51377 <= not w51372 and w51376;
w51378 <= not w51375 and not w51377;
w51379 <= not w23354 and not w51378;
w51380 <= not b(1) and not w51374;
w51381 <= not w51379 and not w51380;
w51382 <= b(2) and not w51368;
w51383 <= not w51366 and w51382;
w51384 <= not w51370 and not w51383;
w51385 <= not w51381 and w51384;
w51386 <= not w51370 and not w51385;
w51387 <= b(3) and not w51360;
w51388 <= not w51358 and w51387;
w51389 <= not w51362 and not w51388;
w51390 <= not w51386 and w51389;
w51391 <= not w51362 and not w51390;
w51392 <= b(4) and not w51351;
w51393 <= not w51349 and w51392;
w51394 <= not w51353 and not w51393;
w51395 <= not w51391 and w51394;
w51396 <= not w51353 and not w51395;
w51397 <= b(5) and not w51342;
w51398 <= not w51340 and w51397;
w51399 <= not w51344 and not w51398;
w51400 <= not w51396 and w51399;
w51401 <= not w51344 and not w51400;
w51402 <= b(6) and not w51333;
w51403 <= not w51331 and w51402;
w51404 <= not w51335 and not w51403;
w51405 <= not w51401 and w51404;
w51406 <= not w51335 and not w51405;
w51407 <= b(7) and not w51324;
w51408 <= not w51322 and w51407;
w51409 <= not w51326 and not w51408;
w51410 <= not w51406 and w51409;
w51411 <= not w51326 and not w51410;
w51412 <= b(8) and not w51315;
w51413 <= not w51313 and w51412;
w51414 <= not w51317 and not w51413;
w51415 <= not w51411 and w51414;
w51416 <= not w51317 and not w51415;
w51417 <= b(9) and not w51306;
w51418 <= not w51304 and w51417;
w51419 <= not w51308 and not w51418;
w51420 <= not w51416 and w51419;
w51421 <= not w51308 and not w51420;
w51422 <= b(10) and not w51297;
w51423 <= not w51295 and w51422;
w51424 <= not w51299 and not w51423;
w51425 <= not w51421 and w51424;
w51426 <= not w51299 and not w51425;
w51427 <= b(11) and not w51288;
w51428 <= not w51286 and w51427;
w51429 <= not w51290 and not w51428;
w51430 <= not w51426 and w51429;
w51431 <= not w51290 and not w51430;
w51432 <= b(12) and not w51279;
w51433 <= not w51277 and w51432;
w51434 <= not w51281 and not w51433;
w51435 <= not w51431 and w51434;
w51436 <= not w51281 and not w51435;
w51437 <= b(13) and not w51270;
w51438 <= not w51268 and w51437;
w51439 <= not w51272 and not w51438;
w51440 <= not w51436 and w51439;
w51441 <= not w51272 and not w51440;
w51442 <= b(14) and not w51261;
w51443 <= not w51259 and w51442;
w51444 <= not w51263 and not w51443;
w51445 <= not w51441 and w51444;
w51446 <= not w51263 and not w51445;
w51447 <= b(15) and not w51252;
w51448 <= not w51250 and w51447;
w51449 <= not w51254 and not w51448;
w51450 <= not w51446 and w51449;
w51451 <= not w51254 and not w51450;
w51452 <= b(16) and not w51243;
w51453 <= not w51241 and w51452;
w51454 <= not w51245 and not w51453;
w51455 <= not w51451 and w51454;
w51456 <= not w51245 and not w51455;
w51457 <= b(17) and not w51234;
w51458 <= not w51232 and w51457;
w51459 <= not w51236 and not w51458;
w51460 <= not w51456 and w51459;
w51461 <= not w51236 and not w51460;
w51462 <= b(18) and not w51225;
w51463 <= not w51223 and w51462;
w51464 <= not w51227 and not w51463;
w51465 <= not w51461 and w51464;
w51466 <= not w51227 and not w51465;
w51467 <= b(19) and not w51216;
w51468 <= not w51214 and w51467;
w51469 <= not w51218 and not w51468;
w51470 <= not w51466 and w51469;
w51471 <= not w51218 and not w51470;
w51472 <= b(20) and not w51207;
w51473 <= not w51205 and w51472;
w51474 <= not w51209 and not w51473;
w51475 <= not w51471 and w51474;
w51476 <= not w51209 and not w51475;
w51477 <= b(21) and not w51198;
w51478 <= not w51196 and w51477;
w51479 <= not w51200 and not w51478;
w51480 <= not w51476 and w51479;
w51481 <= not w51200 and not w51480;
w51482 <= b(22) and not w51189;
w51483 <= not w51187 and w51482;
w51484 <= not w51191 and not w51483;
w51485 <= not w51481 and w51484;
w51486 <= not w51191 and not w51485;
w51487 <= b(23) and not w51180;
w51488 <= not w51178 and w51487;
w51489 <= not w51182 and not w51488;
w51490 <= not w51486 and w51489;
w51491 <= not w51182 and not w51490;
w51492 <= b(24) and not w51171;
w51493 <= not w51169 and w51492;
w51494 <= not w51173 and not w51493;
w51495 <= not w51491 and w51494;
w51496 <= not w51173 and not w51495;
w51497 <= b(25) and not w51162;
w51498 <= not w51160 and w51497;
w51499 <= not w51164 and not w51498;
w51500 <= not w51496 and w51499;
w51501 <= not w51164 and not w51500;
w51502 <= b(26) and not w51153;
w51503 <= not w51151 and w51502;
w51504 <= not w51155 and not w51503;
w51505 <= not w51501 and w51504;
w51506 <= not w51155 and not w51505;
w51507 <= b(27) and not w51144;
w51508 <= not w51142 and w51507;
w51509 <= not w51146 and not w51508;
w51510 <= not w51506 and w51509;
w51511 <= not w51146 and not w51510;
w51512 <= b(28) and not w51135;
w51513 <= not w51133 and w51512;
w51514 <= not w51137 and not w51513;
w51515 <= not w51511 and w51514;
w51516 <= not w51137 and not w51515;
w51517 <= b(29) and not w51126;
w51518 <= not w51124 and w51517;
w51519 <= not w51128 and not w51518;
w51520 <= not w51516 and w51519;
w51521 <= not w51128 and not w51520;
w51522 <= b(30) and not w51117;
w51523 <= not w51115 and w51522;
w51524 <= not w51119 and not w51523;
w51525 <= not w51521 and w51524;
w51526 <= not w51119 and not w51525;
w51527 <= b(31) and not w51108;
w51528 <= not w51106 and w51527;
w51529 <= not w51110 and not w51528;
w51530 <= not w51526 and w51529;
w51531 <= not w51110 and not w51530;
w51532 <= b(32) and not w51099;
w51533 <= not w51097 and w51532;
w51534 <= not w51101 and not w51533;
w51535 <= not w51531 and w51534;
w51536 <= not w51101 and not w51535;
w51537 <= b(33) and not w51090;
w51538 <= not w51088 and w51537;
w51539 <= not w51092 and not w51538;
w51540 <= not w51536 and w51539;
w51541 <= not w51092 and not w51540;
w51542 <= b(34) and not w51081;
w51543 <= not w51079 and w51542;
w51544 <= not w51083 and not w51543;
w51545 <= not w51541 and w51544;
w51546 <= not w51083 and not w51545;
w51547 <= b(35) and not w51072;
w51548 <= not w51070 and w51547;
w51549 <= not w51074 and not w51548;
w51550 <= not w51546 and w51549;
w51551 <= not w51074 and not w51550;
w51552 <= b(36) and not w51063;
w51553 <= not w51061 and w51552;
w51554 <= not w51065 and not w51553;
w51555 <= not w51551 and w51554;
w51556 <= not w51065 and not w51555;
w51557 <= b(37) and not w51054;
w51558 <= not w51052 and w51557;
w51559 <= not w51056 and not w51558;
w51560 <= not w51556 and w51559;
w51561 <= not w51056 and not w51560;
w51562 <= b(38) and not w51045;
w51563 <= not w51043 and w51562;
w51564 <= not w51047 and not w51563;
w51565 <= not w51561 and w51564;
w51566 <= not w51047 and not w51565;
w51567 <= b(39) and not w51036;
w51568 <= not w51034 and w51567;
w51569 <= not w51038 and not w51568;
w51570 <= not w51566 and w51569;
w51571 <= not w51038 and not w51570;
w51572 <= b(40) and not w51027;
w51573 <= not w51025 and w51572;
w51574 <= not w51029 and not w51573;
w51575 <= not w51571 and w51574;
w51576 <= not w51029 and not w51575;
w51577 <= b(41) and not w51018;
w51578 <= not w51016 and w51577;
w51579 <= not w51020 and not w51578;
w51580 <= not w51576 and w51579;
w51581 <= not w51020 and not w51580;
w51582 <= b(42) and not w51009;
w51583 <= not w51007 and w51582;
w51584 <= not w51011 and not w51583;
w51585 <= not w51581 and w51584;
w51586 <= not w51011 and not w51585;
w51587 <= b(43) and not w51000;
w51588 <= not w50998 and w51587;
w51589 <= not w51002 and not w51588;
w51590 <= not w51586 and w51589;
w51591 <= not w51002 and not w51590;
w51592 <= b(44) and not w50991;
w51593 <= not w50989 and w51592;
w51594 <= not w50993 and not w51593;
w51595 <= not w51591 and w51594;
w51596 <= not w50993 and not w51595;
w51597 <= b(45) and not w50982;
w51598 <= not w50980 and w51597;
w51599 <= not w50984 and not w51598;
w51600 <= not w51596 and w51599;
w51601 <= not w50984 and not w51600;
w51602 <= b(46) and not w50973;
w51603 <= not w50971 and w51602;
w51604 <= not w50975 and not w51603;
w51605 <= not w51601 and w51604;
w51606 <= not w50975 and not w51605;
w51607 <= b(47) and not w50964;
w51608 <= not w50962 and w51607;
w51609 <= not w50966 and not w51608;
w51610 <= not w51606 and w51609;
w51611 <= not w50966 and not w51610;
w51612 <= b(48) and not w50955;
w51613 <= not w50953 and w51612;
w51614 <= not w50957 and not w51613;
w51615 <= not w51611 and w51614;
w51616 <= not w50957 and not w51615;
w51617 <= b(49) and not w50946;
w51618 <= not w50944 and w51617;
w51619 <= not w50948 and not w51618;
w51620 <= not w51616 and w51619;
w51621 <= not w50948 and not w51620;
w51622 <= b(50) and not w50937;
w51623 <= not w50935 and w51622;
w51624 <= not w50939 and not w51623;
w51625 <= not w51621 and w51624;
w51626 <= not w50939 and not w51625;
w51627 <= b(51) and not w50928;
w51628 <= not w50926 and w51627;
w51629 <= not w50930 and not w51628;
w51630 <= not w51626 and w51629;
w51631 <= not w50930 and not w51630;
w51632 <= b(52) and not w50919;
w51633 <= not w50917 and w51632;
w51634 <= not w50921 and not w51633;
w51635 <= not w51631 and w51634;
w51636 <= not w50921 and not w51635;
w51637 <= b(53) and not w50910;
w51638 <= not w50908 and w51637;
w51639 <= not w50912 and not w51638;
w51640 <= not w51636 and w51639;
w51641 <= not w50912 and not w51640;
w51642 <= b(54) and not w50901;
w51643 <= not w50899 and w51642;
w51644 <= not w50903 and not w51643;
w51645 <= not w51641 and w51644;
w51646 <= not w50903 and not w51645;
w51647 <= b(55) and not w50892;
w51648 <= not w50890 and w51647;
w51649 <= not w50894 and not w51648;
w51650 <= not w51646 and w51649;
w51651 <= not w50894 and not w51650;
w51652 <= b(56) and not w50872;
w51653 <= not w50870 and w51652;
w51654 <= not w50885 and not w51653;
w51655 <= not w51651 and w51654;
w51656 <= not w50885 and not w51655;
w51657 <= b(57) and not w50882;
w51658 <= not w50880 and w51657;
w51659 <= not w50884 and not w51658;
w51660 <= not w51656 and w51659;
w51661 <= not w50884 and not w51660;
w51662 <= w23638 and not w51661;
w51663 <= not w50873 and not w51662;
w51664 <= not w50894 and w51654;
w51665 <= not w51650 and w51664;
w51666 <= not w51651 and not w51654;
w51667 <= not w51665 and not w51666;
w51668 <= w23638 and not w51667;
w51669 <= not w51661 and w51668;
w51670 <= not w51663 and not w51669;
w51671 <= not b(57) and not w51670;
w51672 <= not w50893 and not w51662;
w51673 <= not w50903 and w51649;
w51674 <= not w51645 and w51673;
w51675 <= not w51646 and not w51649;
w51676 <= not w51674 and not w51675;
w51677 <= w23638 and not w51676;
w51678 <= not w51661 and w51677;
w51679 <= not w51672 and not w51678;
w51680 <= not b(56) and not w51679;
w51681 <= not w50902 and not w51662;
w51682 <= not w50912 and w51644;
w51683 <= not w51640 and w51682;
w51684 <= not w51641 and not w51644;
w51685 <= not w51683 and not w51684;
w51686 <= w23638 and not w51685;
w51687 <= not w51661 and w51686;
w51688 <= not w51681 and not w51687;
w51689 <= not b(55) and not w51688;
w51690 <= not w50911 and not w51662;
w51691 <= not w50921 and w51639;
w51692 <= not w51635 and w51691;
w51693 <= not w51636 and not w51639;
w51694 <= not w51692 and not w51693;
w51695 <= w23638 and not w51694;
w51696 <= not w51661 and w51695;
w51697 <= not w51690 and not w51696;
w51698 <= not b(54) and not w51697;
w51699 <= not w50920 and not w51662;
w51700 <= not w50930 and w51634;
w51701 <= not w51630 and w51700;
w51702 <= not w51631 and not w51634;
w51703 <= not w51701 and not w51702;
w51704 <= w23638 and not w51703;
w51705 <= not w51661 and w51704;
w51706 <= not w51699 and not w51705;
w51707 <= not b(53) and not w51706;
w51708 <= not w50929 and not w51662;
w51709 <= not w50939 and w51629;
w51710 <= not w51625 and w51709;
w51711 <= not w51626 and not w51629;
w51712 <= not w51710 and not w51711;
w51713 <= w23638 and not w51712;
w51714 <= not w51661 and w51713;
w51715 <= not w51708 and not w51714;
w51716 <= not b(52) and not w51715;
w51717 <= not w50938 and not w51662;
w51718 <= not w50948 and w51624;
w51719 <= not w51620 and w51718;
w51720 <= not w51621 and not w51624;
w51721 <= not w51719 and not w51720;
w51722 <= w23638 and not w51721;
w51723 <= not w51661 and w51722;
w51724 <= not w51717 and not w51723;
w51725 <= not b(51) and not w51724;
w51726 <= not w50947 and not w51662;
w51727 <= not w50957 and w51619;
w51728 <= not w51615 and w51727;
w51729 <= not w51616 and not w51619;
w51730 <= not w51728 and not w51729;
w51731 <= w23638 and not w51730;
w51732 <= not w51661 and w51731;
w51733 <= not w51726 and not w51732;
w51734 <= not b(50) and not w51733;
w51735 <= not w50956 and not w51662;
w51736 <= not w50966 and w51614;
w51737 <= not w51610 and w51736;
w51738 <= not w51611 and not w51614;
w51739 <= not w51737 and not w51738;
w51740 <= w23638 and not w51739;
w51741 <= not w51661 and w51740;
w51742 <= not w51735 and not w51741;
w51743 <= not b(49) and not w51742;
w51744 <= not w50965 and not w51662;
w51745 <= not w50975 and w51609;
w51746 <= not w51605 and w51745;
w51747 <= not w51606 and not w51609;
w51748 <= not w51746 and not w51747;
w51749 <= w23638 and not w51748;
w51750 <= not w51661 and w51749;
w51751 <= not w51744 and not w51750;
w51752 <= not b(48) and not w51751;
w51753 <= not w50974 and not w51662;
w51754 <= not w50984 and w51604;
w51755 <= not w51600 and w51754;
w51756 <= not w51601 and not w51604;
w51757 <= not w51755 and not w51756;
w51758 <= w23638 and not w51757;
w51759 <= not w51661 and w51758;
w51760 <= not w51753 and not w51759;
w51761 <= not b(47) and not w51760;
w51762 <= not w50983 and not w51662;
w51763 <= not w50993 and w51599;
w51764 <= not w51595 and w51763;
w51765 <= not w51596 and not w51599;
w51766 <= not w51764 and not w51765;
w51767 <= w23638 and not w51766;
w51768 <= not w51661 and w51767;
w51769 <= not w51762 and not w51768;
w51770 <= not b(46) and not w51769;
w51771 <= not w50992 and not w51662;
w51772 <= not w51002 and w51594;
w51773 <= not w51590 and w51772;
w51774 <= not w51591 and not w51594;
w51775 <= not w51773 and not w51774;
w51776 <= w23638 and not w51775;
w51777 <= not w51661 and w51776;
w51778 <= not w51771 and not w51777;
w51779 <= not b(45) and not w51778;
w51780 <= not w51001 and not w51662;
w51781 <= not w51011 and w51589;
w51782 <= not w51585 and w51781;
w51783 <= not w51586 and not w51589;
w51784 <= not w51782 and not w51783;
w51785 <= w23638 and not w51784;
w51786 <= not w51661 and w51785;
w51787 <= not w51780 and not w51786;
w51788 <= not b(44) and not w51787;
w51789 <= not w51010 and not w51662;
w51790 <= not w51020 and w51584;
w51791 <= not w51580 and w51790;
w51792 <= not w51581 and not w51584;
w51793 <= not w51791 and not w51792;
w51794 <= w23638 and not w51793;
w51795 <= not w51661 and w51794;
w51796 <= not w51789 and not w51795;
w51797 <= not b(43) and not w51796;
w51798 <= not w51019 and not w51662;
w51799 <= not w51029 and w51579;
w51800 <= not w51575 and w51799;
w51801 <= not w51576 and not w51579;
w51802 <= not w51800 and not w51801;
w51803 <= w23638 and not w51802;
w51804 <= not w51661 and w51803;
w51805 <= not w51798 and not w51804;
w51806 <= not b(42) and not w51805;
w51807 <= not w51028 and not w51662;
w51808 <= not w51038 and w51574;
w51809 <= not w51570 and w51808;
w51810 <= not w51571 and not w51574;
w51811 <= not w51809 and not w51810;
w51812 <= w23638 and not w51811;
w51813 <= not w51661 and w51812;
w51814 <= not w51807 and not w51813;
w51815 <= not b(41) and not w51814;
w51816 <= not w51037 and not w51662;
w51817 <= not w51047 and w51569;
w51818 <= not w51565 and w51817;
w51819 <= not w51566 and not w51569;
w51820 <= not w51818 and not w51819;
w51821 <= w23638 and not w51820;
w51822 <= not w51661 and w51821;
w51823 <= not w51816 and not w51822;
w51824 <= not b(40) and not w51823;
w51825 <= not w51046 and not w51662;
w51826 <= not w51056 and w51564;
w51827 <= not w51560 and w51826;
w51828 <= not w51561 and not w51564;
w51829 <= not w51827 and not w51828;
w51830 <= w23638 and not w51829;
w51831 <= not w51661 and w51830;
w51832 <= not w51825 and not w51831;
w51833 <= not b(39) and not w51832;
w51834 <= not w51055 and not w51662;
w51835 <= not w51065 and w51559;
w51836 <= not w51555 and w51835;
w51837 <= not w51556 and not w51559;
w51838 <= not w51836 and not w51837;
w51839 <= w23638 and not w51838;
w51840 <= not w51661 and w51839;
w51841 <= not w51834 and not w51840;
w51842 <= not b(38) and not w51841;
w51843 <= not w51064 and not w51662;
w51844 <= not w51074 and w51554;
w51845 <= not w51550 and w51844;
w51846 <= not w51551 and not w51554;
w51847 <= not w51845 and not w51846;
w51848 <= w23638 and not w51847;
w51849 <= not w51661 and w51848;
w51850 <= not w51843 and not w51849;
w51851 <= not b(37) and not w51850;
w51852 <= not w51073 and not w51662;
w51853 <= not w51083 and w51549;
w51854 <= not w51545 and w51853;
w51855 <= not w51546 and not w51549;
w51856 <= not w51854 and not w51855;
w51857 <= w23638 and not w51856;
w51858 <= not w51661 and w51857;
w51859 <= not w51852 and not w51858;
w51860 <= not b(36) and not w51859;
w51861 <= not w51082 and not w51662;
w51862 <= not w51092 and w51544;
w51863 <= not w51540 and w51862;
w51864 <= not w51541 and not w51544;
w51865 <= not w51863 and not w51864;
w51866 <= w23638 and not w51865;
w51867 <= not w51661 and w51866;
w51868 <= not w51861 and not w51867;
w51869 <= not b(35) and not w51868;
w51870 <= not w51091 and not w51662;
w51871 <= not w51101 and w51539;
w51872 <= not w51535 and w51871;
w51873 <= not w51536 and not w51539;
w51874 <= not w51872 and not w51873;
w51875 <= w23638 and not w51874;
w51876 <= not w51661 and w51875;
w51877 <= not w51870 and not w51876;
w51878 <= not b(34) and not w51877;
w51879 <= not w51100 and not w51662;
w51880 <= not w51110 and w51534;
w51881 <= not w51530 and w51880;
w51882 <= not w51531 and not w51534;
w51883 <= not w51881 and not w51882;
w51884 <= w23638 and not w51883;
w51885 <= not w51661 and w51884;
w51886 <= not w51879 and not w51885;
w51887 <= not b(33) and not w51886;
w51888 <= not w51109 and not w51662;
w51889 <= not w51119 and w51529;
w51890 <= not w51525 and w51889;
w51891 <= not w51526 and not w51529;
w51892 <= not w51890 and not w51891;
w51893 <= w23638 and not w51892;
w51894 <= not w51661 and w51893;
w51895 <= not w51888 and not w51894;
w51896 <= not b(32) and not w51895;
w51897 <= not w51118 and not w51662;
w51898 <= not w51128 and w51524;
w51899 <= not w51520 and w51898;
w51900 <= not w51521 and not w51524;
w51901 <= not w51899 and not w51900;
w51902 <= w23638 and not w51901;
w51903 <= not w51661 and w51902;
w51904 <= not w51897 and not w51903;
w51905 <= not b(31) and not w51904;
w51906 <= not w51127 and not w51662;
w51907 <= not w51137 and w51519;
w51908 <= not w51515 and w51907;
w51909 <= not w51516 and not w51519;
w51910 <= not w51908 and not w51909;
w51911 <= w23638 and not w51910;
w51912 <= not w51661 and w51911;
w51913 <= not w51906 and not w51912;
w51914 <= not b(30) and not w51913;
w51915 <= not w51136 and not w51662;
w51916 <= not w51146 and w51514;
w51917 <= not w51510 and w51916;
w51918 <= not w51511 and not w51514;
w51919 <= not w51917 and not w51918;
w51920 <= w23638 and not w51919;
w51921 <= not w51661 and w51920;
w51922 <= not w51915 and not w51921;
w51923 <= not b(29) and not w51922;
w51924 <= not w51145 and not w51662;
w51925 <= not w51155 and w51509;
w51926 <= not w51505 and w51925;
w51927 <= not w51506 and not w51509;
w51928 <= not w51926 and not w51927;
w51929 <= w23638 and not w51928;
w51930 <= not w51661 and w51929;
w51931 <= not w51924 and not w51930;
w51932 <= not b(28) and not w51931;
w51933 <= not w51154 and not w51662;
w51934 <= not w51164 and w51504;
w51935 <= not w51500 and w51934;
w51936 <= not w51501 and not w51504;
w51937 <= not w51935 and not w51936;
w51938 <= w23638 and not w51937;
w51939 <= not w51661 and w51938;
w51940 <= not w51933 and not w51939;
w51941 <= not b(27) and not w51940;
w51942 <= not w51163 and not w51662;
w51943 <= not w51173 and w51499;
w51944 <= not w51495 and w51943;
w51945 <= not w51496 and not w51499;
w51946 <= not w51944 and not w51945;
w51947 <= w23638 and not w51946;
w51948 <= not w51661 and w51947;
w51949 <= not w51942 and not w51948;
w51950 <= not b(26) and not w51949;
w51951 <= not w51172 and not w51662;
w51952 <= not w51182 and w51494;
w51953 <= not w51490 and w51952;
w51954 <= not w51491 and not w51494;
w51955 <= not w51953 and not w51954;
w51956 <= w23638 and not w51955;
w51957 <= not w51661 and w51956;
w51958 <= not w51951 and not w51957;
w51959 <= not b(25) and not w51958;
w51960 <= not w51181 and not w51662;
w51961 <= not w51191 and w51489;
w51962 <= not w51485 and w51961;
w51963 <= not w51486 and not w51489;
w51964 <= not w51962 and not w51963;
w51965 <= w23638 and not w51964;
w51966 <= not w51661 and w51965;
w51967 <= not w51960 and not w51966;
w51968 <= not b(24) and not w51967;
w51969 <= not w51190 and not w51662;
w51970 <= not w51200 and w51484;
w51971 <= not w51480 and w51970;
w51972 <= not w51481 and not w51484;
w51973 <= not w51971 and not w51972;
w51974 <= w23638 and not w51973;
w51975 <= not w51661 and w51974;
w51976 <= not w51969 and not w51975;
w51977 <= not b(23) and not w51976;
w51978 <= not w51199 and not w51662;
w51979 <= not w51209 and w51479;
w51980 <= not w51475 and w51979;
w51981 <= not w51476 and not w51479;
w51982 <= not w51980 and not w51981;
w51983 <= w23638 and not w51982;
w51984 <= not w51661 and w51983;
w51985 <= not w51978 and not w51984;
w51986 <= not b(22) and not w51985;
w51987 <= not w51208 and not w51662;
w51988 <= not w51218 and w51474;
w51989 <= not w51470 and w51988;
w51990 <= not w51471 and not w51474;
w51991 <= not w51989 and not w51990;
w51992 <= w23638 and not w51991;
w51993 <= not w51661 and w51992;
w51994 <= not w51987 and not w51993;
w51995 <= not b(21) and not w51994;
w51996 <= not w51217 and not w51662;
w51997 <= not w51227 and w51469;
w51998 <= not w51465 and w51997;
w51999 <= not w51466 and not w51469;
w52000 <= not w51998 and not w51999;
w52001 <= w23638 and not w52000;
w52002 <= not w51661 and w52001;
w52003 <= not w51996 and not w52002;
w52004 <= not b(20) and not w52003;
w52005 <= not w51226 and not w51662;
w52006 <= not w51236 and w51464;
w52007 <= not w51460 and w52006;
w52008 <= not w51461 and not w51464;
w52009 <= not w52007 and not w52008;
w52010 <= w23638 and not w52009;
w52011 <= not w51661 and w52010;
w52012 <= not w52005 and not w52011;
w52013 <= not b(19) and not w52012;
w52014 <= not w51235 and not w51662;
w52015 <= not w51245 and w51459;
w52016 <= not w51455 and w52015;
w52017 <= not w51456 and not w51459;
w52018 <= not w52016 and not w52017;
w52019 <= w23638 and not w52018;
w52020 <= not w51661 and w52019;
w52021 <= not w52014 and not w52020;
w52022 <= not b(18) and not w52021;
w52023 <= not w51244 and not w51662;
w52024 <= not w51254 and w51454;
w52025 <= not w51450 and w52024;
w52026 <= not w51451 and not w51454;
w52027 <= not w52025 and not w52026;
w52028 <= w23638 and not w52027;
w52029 <= not w51661 and w52028;
w52030 <= not w52023 and not w52029;
w52031 <= not b(17) and not w52030;
w52032 <= not w51253 and not w51662;
w52033 <= not w51263 and w51449;
w52034 <= not w51445 and w52033;
w52035 <= not w51446 and not w51449;
w52036 <= not w52034 and not w52035;
w52037 <= w23638 and not w52036;
w52038 <= not w51661 and w52037;
w52039 <= not w52032 and not w52038;
w52040 <= not b(16) and not w52039;
w52041 <= not w51262 and not w51662;
w52042 <= not w51272 and w51444;
w52043 <= not w51440 and w52042;
w52044 <= not w51441 and not w51444;
w52045 <= not w52043 and not w52044;
w52046 <= w23638 and not w52045;
w52047 <= not w51661 and w52046;
w52048 <= not w52041 and not w52047;
w52049 <= not b(15) and not w52048;
w52050 <= not w51271 and not w51662;
w52051 <= not w51281 and w51439;
w52052 <= not w51435 and w52051;
w52053 <= not w51436 and not w51439;
w52054 <= not w52052 and not w52053;
w52055 <= w23638 and not w52054;
w52056 <= not w51661 and w52055;
w52057 <= not w52050 and not w52056;
w52058 <= not b(14) and not w52057;
w52059 <= not w51280 and not w51662;
w52060 <= not w51290 and w51434;
w52061 <= not w51430 and w52060;
w52062 <= not w51431 and not w51434;
w52063 <= not w52061 and not w52062;
w52064 <= w23638 and not w52063;
w52065 <= not w51661 and w52064;
w52066 <= not w52059 and not w52065;
w52067 <= not b(13) and not w52066;
w52068 <= not w51289 and not w51662;
w52069 <= not w51299 and w51429;
w52070 <= not w51425 and w52069;
w52071 <= not w51426 and not w51429;
w52072 <= not w52070 and not w52071;
w52073 <= w23638 and not w52072;
w52074 <= not w51661 and w52073;
w52075 <= not w52068 and not w52074;
w52076 <= not b(12) and not w52075;
w52077 <= not w51298 and not w51662;
w52078 <= not w51308 and w51424;
w52079 <= not w51420 and w52078;
w52080 <= not w51421 and not w51424;
w52081 <= not w52079 and not w52080;
w52082 <= w23638 and not w52081;
w52083 <= not w51661 and w52082;
w52084 <= not w52077 and not w52083;
w52085 <= not b(11) and not w52084;
w52086 <= not w51307 and not w51662;
w52087 <= not w51317 and w51419;
w52088 <= not w51415 and w52087;
w52089 <= not w51416 and not w51419;
w52090 <= not w52088 and not w52089;
w52091 <= w23638 and not w52090;
w52092 <= not w51661 and w52091;
w52093 <= not w52086 and not w52092;
w52094 <= not b(10) and not w52093;
w52095 <= not w51316 and not w51662;
w52096 <= not w51326 and w51414;
w52097 <= not w51410 and w52096;
w52098 <= not w51411 and not w51414;
w52099 <= not w52097 and not w52098;
w52100 <= w23638 and not w52099;
w52101 <= not w51661 and w52100;
w52102 <= not w52095 and not w52101;
w52103 <= not b(9) and not w52102;
w52104 <= not w51325 and not w51662;
w52105 <= not w51335 and w51409;
w52106 <= not w51405 and w52105;
w52107 <= not w51406 and not w51409;
w52108 <= not w52106 and not w52107;
w52109 <= w23638 and not w52108;
w52110 <= not w51661 and w52109;
w52111 <= not w52104 and not w52110;
w52112 <= not b(8) and not w52111;
w52113 <= not w51334 and not w51662;
w52114 <= not w51344 and w51404;
w52115 <= not w51400 and w52114;
w52116 <= not w51401 and not w51404;
w52117 <= not w52115 and not w52116;
w52118 <= w23638 and not w52117;
w52119 <= not w51661 and w52118;
w52120 <= not w52113 and not w52119;
w52121 <= not b(7) and not w52120;
w52122 <= not w51343 and not w51662;
w52123 <= not w51353 and w51399;
w52124 <= not w51395 and w52123;
w52125 <= not w51396 and not w51399;
w52126 <= not w52124 and not w52125;
w52127 <= w23638 and not w52126;
w52128 <= not w51661 and w52127;
w52129 <= not w52122 and not w52128;
w52130 <= not b(6) and not w52129;
w52131 <= not w51352 and not w51662;
w52132 <= not w51362 and w51394;
w52133 <= not w51390 and w52132;
w52134 <= not w51391 and not w51394;
w52135 <= not w52133 and not w52134;
w52136 <= w23638 and not w52135;
w52137 <= not w51661 and w52136;
w52138 <= not w52131 and not w52137;
w52139 <= not b(5) and not w52138;
w52140 <= not w51361 and not w51662;
w52141 <= not w51370 and w51389;
w52142 <= not w51385 and w52141;
w52143 <= not w51386 and not w51389;
w52144 <= not w52142 and not w52143;
w52145 <= w23638 and not w52144;
w52146 <= not w51661 and w52145;
w52147 <= not w52140 and not w52146;
w52148 <= not b(4) and not w52147;
w52149 <= not w51369 and not w51662;
w52150 <= not w51380 and w51384;
w52151 <= not w51379 and w52150;
w52152 <= not w51381 and not w51384;
w52153 <= not w52151 and not w52152;
w52154 <= w23638 and not w52153;
w52155 <= not w51661 and w52154;
w52156 <= not w52149 and not w52155;
w52157 <= not b(3) and not w52156;
w52158 <= not w51374 and not w51662;
w52159 <= w23354 and not w51377;
w52160 <= not w51375 and w52159;
w52161 <= w23638 and not w52160;
w52162 <= not w51379 and w52161;
w52163 <= not w51661 and w52162;
w52164 <= not w52158 and not w52163;
w52165 <= not b(2) and not w52164;
w52166 <= w24145 and not w51661;
w52167 <= a(6) and not w52166;
w52168 <= w24149 and not w51661;
w52169 <= not w52167 and not w52168;
w52170 <= b(1) and not w52169;
w52171 <= not b(1) and not w52168;
w52172 <= not w52167 and w52171;
w52173 <= not w52170 and not w52172;
w52174 <= not w24156 and not w52173;
w52175 <= not b(1) and not w52169;
w52176 <= not w52174 and not w52175;
w52177 <= b(2) and not w52163;
w52178 <= not w52158 and w52177;
w52179 <= not w52165 and not w52178;
w52180 <= not w52176 and w52179;
w52181 <= not w52165 and not w52180;
w52182 <= b(3) and not w52155;
w52183 <= not w52149 and w52182;
w52184 <= not w52157 and not w52183;
w52185 <= not w52181 and w52184;
w52186 <= not w52157 and not w52185;
w52187 <= b(4) and not w52146;
w52188 <= not w52140 and w52187;
w52189 <= not w52148 and not w52188;
w52190 <= not w52186 and w52189;
w52191 <= not w52148 and not w52190;
w52192 <= b(5) and not w52137;
w52193 <= not w52131 and w52192;
w52194 <= not w52139 and not w52193;
w52195 <= not w52191 and w52194;
w52196 <= not w52139 and not w52195;
w52197 <= b(6) and not w52128;
w52198 <= not w52122 and w52197;
w52199 <= not w52130 and not w52198;
w52200 <= not w52196 and w52199;
w52201 <= not w52130 and not w52200;
w52202 <= b(7) and not w52119;
w52203 <= not w52113 and w52202;
w52204 <= not w52121 and not w52203;
w52205 <= not w52201 and w52204;
w52206 <= not w52121 and not w52205;
w52207 <= b(8) and not w52110;
w52208 <= not w52104 and w52207;
w52209 <= not w52112 and not w52208;
w52210 <= not w52206 and w52209;
w52211 <= not w52112 and not w52210;
w52212 <= b(9) and not w52101;
w52213 <= not w52095 and w52212;
w52214 <= not w52103 and not w52213;
w52215 <= not w52211 and w52214;
w52216 <= not w52103 and not w52215;
w52217 <= b(10) and not w52092;
w52218 <= not w52086 and w52217;
w52219 <= not w52094 and not w52218;
w52220 <= not w52216 and w52219;
w52221 <= not w52094 and not w52220;
w52222 <= b(11) and not w52083;
w52223 <= not w52077 and w52222;
w52224 <= not w52085 and not w52223;
w52225 <= not w52221 and w52224;
w52226 <= not w52085 and not w52225;
w52227 <= b(12) and not w52074;
w52228 <= not w52068 and w52227;
w52229 <= not w52076 and not w52228;
w52230 <= not w52226 and w52229;
w52231 <= not w52076 and not w52230;
w52232 <= b(13) and not w52065;
w52233 <= not w52059 and w52232;
w52234 <= not w52067 and not w52233;
w52235 <= not w52231 and w52234;
w52236 <= not w52067 and not w52235;
w52237 <= b(14) and not w52056;
w52238 <= not w52050 and w52237;
w52239 <= not w52058 and not w52238;
w52240 <= not w52236 and w52239;
w52241 <= not w52058 and not w52240;
w52242 <= b(15) and not w52047;
w52243 <= not w52041 and w52242;
w52244 <= not w52049 and not w52243;
w52245 <= not w52241 and w52244;
w52246 <= not w52049 and not w52245;
w52247 <= b(16) and not w52038;
w52248 <= not w52032 and w52247;
w52249 <= not w52040 and not w52248;
w52250 <= not w52246 and w52249;
w52251 <= not w52040 and not w52250;
w52252 <= b(17) and not w52029;
w52253 <= not w52023 and w52252;
w52254 <= not w52031 and not w52253;
w52255 <= not w52251 and w52254;
w52256 <= not w52031 and not w52255;
w52257 <= b(18) and not w52020;
w52258 <= not w52014 and w52257;
w52259 <= not w52022 and not w52258;
w52260 <= not w52256 and w52259;
w52261 <= not w52022 and not w52260;
w52262 <= b(19) and not w52011;
w52263 <= not w52005 and w52262;
w52264 <= not w52013 and not w52263;
w52265 <= not w52261 and w52264;
w52266 <= not w52013 and not w52265;
w52267 <= b(20) and not w52002;
w52268 <= not w51996 and w52267;
w52269 <= not w52004 and not w52268;
w52270 <= not w52266 and w52269;
w52271 <= not w52004 and not w52270;
w52272 <= b(21) and not w51993;
w52273 <= not w51987 and w52272;
w52274 <= not w51995 and not w52273;
w52275 <= not w52271 and w52274;
w52276 <= not w51995 and not w52275;
w52277 <= b(22) and not w51984;
w52278 <= not w51978 and w52277;
w52279 <= not w51986 and not w52278;
w52280 <= not w52276 and w52279;
w52281 <= not w51986 and not w52280;
w52282 <= b(23) and not w51975;
w52283 <= not w51969 and w52282;
w52284 <= not w51977 and not w52283;
w52285 <= not w52281 and w52284;
w52286 <= not w51977 and not w52285;
w52287 <= b(24) and not w51966;
w52288 <= not w51960 and w52287;
w52289 <= not w51968 and not w52288;
w52290 <= not w52286 and w52289;
w52291 <= not w51968 and not w52290;
w52292 <= b(25) and not w51957;
w52293 <= not w51951 and w52292;
w52294 <= not w51959 and not w52293;
w52295 <= not w52291 and w52294;
w52296 <= not w51959 and not w52295;
w52297 <= b(26) and not w51948;
w52298 <= not w51942 and w52297;
w52299 <= not w51950 and not w52298;
w52300 <= not w52296 and w52299;
w52301 <= not w51950 and not w52300;
w52302 <= b(27) and not w51939;
w52303 <= not w51933 and w52302;
w52304 <= not w51941 and not w52303;
w52305 <= not w52301 and w52304;
w52306 <= not w51941 and not w52305;
w52307 <= b(28) and not w51930;
w52308 <= not w51924 and w52307;
w52309 <= not w51932 and not w52308;
w52310 <= not w52306 and w52309;
w52311 <= not w51932 and not w52310;
w52312 <= b(29) and not w51921;
w52313 <= not w51915 and w52312;
w52314 <= not w51923 and not w52313;
w52315 <= not w52311 and w52314;
w52316 <= not w51923 and not w52315;
w52317 <= b(30) and not w51912;
w52318 <= not w51906 and w52317;
w52319 <= not w51914 and not w52318;
w52320 <= not w52316 and w52319;
w52321 <= not w51914 and not w52320;
w52322 <= b(31) and not w51903;
w52323 <= not w51897 and w52322;
w52324 <= not w51905 and not w52323;
w52325 <= not w52321 and w52324;
w52326 <= not w51905 and not w52325;
w52327 <= b(32) and not w51894;
w52328 <= not w51888 and w52327;
w52329 <= not w51896 and not w52328;
w52330 <= not w52326 and w52329;
w52331 <= not w51896 and not w52330;
w52332 <= b(33) and not w51885;
w52333 <= not w51879 and w52332;
w52334 <= not w51887 and not w52333;
w52335 <= not w52331 and w52334;
w52336 <= not w51887 and not w52335;
w52337 <= b(34) and not w51876;
w52338 <= not w51870 and w52337;
w52339 <= not w51878 and not w52338;
w52340 <= not w52336 and w52339;
w52341 <= not w51878 and not w52340;
w52342 <= b(35) and not w51867;
w52343 <= not w51861 and w52342;
w52344 <= not w51869 and not w52343;
w52345 <= not w52341 and w52344;
w52346 <= not w51869 and not w52345;
w52347 <= b(36) and not w51858;
w52348 <= not w51852 and w52347;
w52349 <= not w51860 and not w52348;
w52350 <= not w52346 and w52349;
w52351 <= not w51860 and not w52350;
w52352 <= b(37) and not w51849;
w52353 <= not w51843 and w52352;
w52354 <= not w51851 and not w52353;
w52355 <= not w52351 and w52354;
w52356 <= not w51851 and not w52355;
w52357 <= b(38) and not w51840;
w52358 <= not w51834 and w52357;
w52359 <= not w51842 and not w52358;
w52360 <= not w52356 and w52359;
w52361 <= not w51842 and not w52360;
w52362 <= b(39) and not w51831;
w52363 <= not w51825 and w52362;
w52364 <= not w51833 and not w52363;
w52365 <= not w52361 and w52364;
w52366 <= not w51833 and not w52365;
w52367 <= b(40) and not w51822;
w52368 <= not w51816 and w52367;
w52369 <= not w51824 and not w52368;
w52370 <= not w52366 and w52369;
w52371 <= not w51824 and not w52370;
w52372 <= b(41) and not w51813;
w52373 <= not w51807 and w52372;
w52374 <= not w51815 and not w52373;
w52375 <= not w52371 and w52374;
w52376 <= not w51815 and not w52375;
w52377 <= b(42) and not w51804;
w52378 <= not w51798 and w52377;
w52379 <= not w51806 and not w52378;
w52380 <= not w52376 and w52379;
w52381 <= not w51806 and not w52380;
w52382 <= b(43) and not w51795;
w52383 <= not w51789 and w52382;
w52384 <= not w51797 and not w52383;
w52385 <= not w52381 and w52384;
w52386 <= not w51797 and not w52385;
w52387 <= b(44) and not w51786;
w52388 <= not w51780 and w52387;
w52389 <= not w51788 and not w52388;
w52390 <= not w52386 and w52389;
w52391 <= not w51788 and not w52390;
w52392 <= b(45) and not w51777;
w52393 <= not w51771 and w52392;
w52394 <= not w51779 and not w52393;
w52395 <= not w52391 and w52394;
w52396 <= not w51779 and not w52395;
w52397 <= b(46) and not w51768;
w52398 <= not w51762 and w52397;
w52399 <= not w51770 and not w52398;
w52400 <= not w52396 and w52399;
w52401 <= not w51770 and not w52400;
w52402 <= b(47) and not w51759;
w52403 <= not w51753 and w52402;
w52404 <= not w51761 and not w52403;
w52405 <= not w52401 and w52404;
w52406 <= not w51761 and not w52405;
w52407 <= b(48) and not w51750;
w52408 <= not w51744 and w52407;
w52409 <= not w51752 and not w52408;
w52410 <= not w52406 and w52409;
w52411 <= not w51752 and not w52410;
w52412 <= b(49) and not w51741;
w52413 <= not w51735 and w52412;
w52414 <= not w51743 and not w52413;
w52415 <= not w52411 and w52414;
w52416 <= not w51743 and not w52415;
w52417 <= b(50) and not w51732;
w52418 <= not w51726 and w52417;
w52419 <= not w51734 and not w52418;
w52420 <= not w52416 and w52419;
w52421 <= not w51734 and not w52420;
w52422 <= b(51) and not w51723;
w52423 <= not w51717 and w52422;
w52424 <= not w51725 and not w52423;
w52425 <= not w52421 and w52424;
w52426 <= not w51725 and not w52425;
w52427 <= b(52) and not w51714;
w52428 <= not w51708 and w52427;
w52429 <= not w51716 and not w52428;
w52430 <= not w52426 and w52429;
w52431 <= not w51716 and not w52430;
w52432 <= b(53) and not w51705;
w52433 <= not w51699 and w52432;
w52434 <= not w51707 and not w52433;
w52435 <= not w52431 and w52434;
w52436 <= not w51707 and not w52435;
w52437 <= b(54) and not w51696;
w52438 <= not w51690 and w52437;
w52439 <= not w51698 and not w52438;
w52440 <= not w52436 and w52439;
w52441 <= not w51698 and not w52440;
w52442 <= b(55) and not w51687;
w52443 <= not w51681 and w52442;
w52444 <= not w51689 and not w52443;
w52445 <= not w52441 and w52444;
w52446 <= not w51689 and not w52445;
w52447 <= b(56) and not w51678;
w52448 <= not w51672 and w52447;
w52449 <= not w51680 and not w52448;
w52450 <= not w52446 and w52449;
w52451 <= not w51680 and not w52450;
w52452 <= b(57) and not w51669;
w52453 <= not w51663 and w52452;
w52454 <= not w51671 and not w52453;
w52455 <= not w52451 and w52454;
w52456 <= not w51671 and not w52455;
w52457 <= not w50883 and not w51662;
w52458 <= not w50885 and w51659;
w52459 <= not w51655 and w52458;
w52460 <= not w51656 and not w51659;
w52461 <= not w52459 and not w52460;
w52462 <= w51662 and not w52461;
w52463 <= not w52457 and not w52462;
w52464 <= not b(58) and not w52463;
w52465 <= b(58) and not w52457;
w52466 <= not w52462 and w52465;
w52467 <= w24450 and not w52466;
w52468 <= not w52464 and w52467;
w52469 <= not w52456 and w52468;
w52470 <= w23638 and not w52463;
w52471 <= not w52469 and not w52470;
w52472 <= not w51680 and w52454;
w52473 <= not w52450 and w52472;
w52474 <= not w52451 and not w52454;
w52475 <= not w52473 and not w52474;
w52476 <= not w52471 and not w52475;
w52477 <= not w51670 and not w52470;
w52478 <= not w52469 and w52477;
w52479 <= not w52476 and not w52478;
w52480 <= not b(58) and not w52479;
w52481 <= not w51689 and w52449;
w52482 <= not w52445 and w52481;
w52483 <= not w52446 and not w52449;
w52484 <= not w52482 and not w52483;
w52485 <= not w52471 and not w52484;
w52486 <= not w51679 and not w52470;
w52487 <= not w52469 and w52486;
w52488 <= not w52485 and not w52487;
w52489 <= not b(57) and not w52488;
w52490 <= not w51698 and w52444;
w52491 <= not w52440 and w52490;
w52492 <= not w52441 and not w52444;
w52493 <= not w52491 and not w52492;
w52494 <= not w52471 and not w52493;
w52495 <= not w51688 and not w52470;
w52496 <= not w52469 and w52495;
w52497 <= not w52494 and not w52496;
w52498 <= not b(56) and not w52497;
w52499 <= not w51707 and w52439;
w52500 <= not w52435 and w52499;
w52501 <= not w52436 and not w52439;
w52502 <= not w52500 and not w52501;
w52503 <= not w52471 and not w52502;
w52504 <= not w51697 and not w52470;
w52505 <= not w52469 and w52504;
w52506 <= not w52503 and not w52505;
w52507 <= not b(55) and not w52506;
w52508 <= not w51716 and w52434;
w52509 <= not w52430 and w52508;
w52510 <= not w52431 and not w52434;
w52511 <= not w52509 and not w52510;
w52512 <= not w52471 and not w52511;
w52513 <= not w51706 and not w52470;
w52514 <= not w52469 and w52513;
w52515 <= not w52512 and not w52514;
w52516 <= not b(54) and not w52515;
w52517 <= not w51725 and w52429;
w52518 <= not w52425 and w52517;
w52519 <= not w52426 and not w52429;
w52520 <= not w52518 and not w52519;
w52521 <= not w52471 and not w52520;
w52522 <= not w51715 and not w52470;
w52523 <= not w52469 and w52522;
w52524 <= not w52521 and not w52523;
w52525 <= not b(53) and not w52524;
w52526 <= not w51734 and w52424;
w52527 <= not w52420 and w52526;
w52528 <= not w52421 and not w52424;
w52529 <= not w52527 and not w52528;
w52530 <= not w52471 and not w52529;
w52531 <= not w51724 and not w52470;
w52532 <= not w52469 and w52531;
w52533 <= not w52530 and not w52532;
w52534 <= not b(52) and not w52533;
w52535 <= not w51743 and w52419;
w52536 <= not w52415 and w52535;
w52537 <= not w52416 and not w52419;
w52538 <= not w52536 and not w52537;
w52539 <= not w52471 and not w52538;
w52540 <= not w51733 and not w52470;
w52541 <= not w52469 and w52540;
w52542 <= not w52539 and not w52541;
w52543 <= not b(51) and not w52542;
w52544 <= not w51752 and w52414;
w52545 <= not w52410 and w52544;
w52546 <= not w52411 and not w52414;
w52547 <= not w52545 and not w52546;
w52548 <= not w52471 and not w52547;
w52549 <= not w51742 and not w52470;
w52550 <= not w52469 and w52549;
w52551 <= not w52548 and not w52550;
w52552 <= not b(50) and not w52551;
w52553 <= not w51761 and w52409;
w52554 <= not w52405 and w52553;
w52555 <= not w52406 and not w52409;
w52556 <= not w52554 and not w52555;
w52557 <= not w52471 and not w52556;
w52558 <= not w51751 and not w52470;
w52559 <= not w52469 and w52558;
w52560 <= not w52557 and not w52559;
w52561 <= not b(49) and not w52560;
w52562 <= not w51770 and w52404;
w52563 <= not w52400 and w52562;
w52564 <= not w52401 and not w52404;
w52565 <= not w52563 and not w52564;
w52566 <= not w52471 and not w52565;
w52567 <= not w51760 and not w52470;
w52568 <= not w52469 and w52567;
w52569 <= not w52566 and not w52568;
w52570 <= not b(48) and not w52569;
w52571 <= not w51779 and w52399;
w52572 <= not w52395 and w52571;
w52573 <= not w52396 and not w52399;
w52574 <= not w52572 and not w52573;
w52575 <= not w52471 and not w52574;
w52576 <= not w51769 and not w52470;
w52577 <= not w52469 and w52576;
w52578 <= not w52575 and not w52577;
w52579 <= not b(47) and not w52578;
w52580 <= not w51788 and w52394;
w52581 <= not w52390 and w52580;
w52582 <= not w52391 and not w52394;
w52583 <= not w52581 and not w52582;
w52584 <= not w52471 and not w52583;
w52585 <= not w51778 and not w52470;
w52586 <= not w52469 and w52585;
w52587 <= not w52584 and not w52586;
w52588 <= not b(46) and not w52587;
w52589 <= not w51797 and w52389;
w52590 <= not w52385 and w52589;
w52591 <= not w52386 and not w52389;
w52592 <= not w52590 and not w52591;
w52593 <= not w52471 and not w52592;
w52594 <= not w51787 and not w52470;
w52595 <= not w52469 and w52594;
w52596 <= not w52593 and not w52595;
w52597 <= not b(45) and not w52596;
w52598 <= not w51806 and w52384;
w52599 <= not w52380 and w52598;
w52600 <= not w52381 and not w52384;
w52601 <= not w52599 and not w52600;
w52602 <= not w52471 and not w52601;
w52603 <= not w51796 and not w52470;
w52604 <= not w52469 and w52603;
w52605 <= not w52602 and not w52604;
w52606 <= not b(44) and not w52605;
w52607 <= not w51815 and w52379;
w52608 <= not w52375 and w52607;
w52609 <= not w52376 and not w52379;
w52610 <= not w52608 and not w52609;
w52611 <= not w52471 and not w52610;
w52612 <= not w51805 and not w52470;
w52613 <= not w52469 and w52612;
w52614 <= not w52611 and not w52613;
w52615 <= not b(43) and not w52614;
w52616 <= not w51824 and w52374;
w52617 <= not w52370 and w52616;
w52618 <= not w52371 and not w52374;
w52619 <= not w52617 and not w52618;
w52620 <= not w52471 and not w52619;
w52621 <= not w51814 and not w52470;
w52622 <= not w52469 and w52621;
w52623 <= not w52620 and not w52622;
w52624 <= not b(42) and not w52623;
w52625 <= not w51833 and w52369;
w52626 <= not w52365 and w52625;
w52627 <= not w52366 and not w52369;
w52628 <= not w52626 and not w52627;
w52629 <= not w52471 and not w52628;
w52630 <= not w51823 and not w52470;
w52631 <= not w52469 and w52630;
w52632 <= not w52629 and not w52631;
w52633 <= not b(41) and not w52632;
w52634 <= not w51842 and w52364;
w52635 <= not w52360 and w52634;
w52636 <= not w52361 and not w52364;
w52637 <= not w52635 and not w52636;
w52638 <= not w52471 and not w52637;
w52639 <= not w51832 and not w52470;
w52640 <= not w52469 and w52639;
w52641 <= not w52638 and not w52640;
w52642 <= not b(40) and not w52641;
w52643 <= not w51851 and w52359;
w52644 <= not w52355 and w52643;
w52645 <= not w52356 and not w52359;
w52646 <= not w52644 and not w52645;
w52647 <= not w52471 and not w52646;
w52648 <= not w51841 and not w52470;
w52649 <= not w52469 and w52648;
w52650 <= not w52647 and not w52649;
w52651 <= not b(39) and not w52650;
w52652 <= not w51860 and w52354;
w52653 <= not w52350 and w52652;
w52654 <= not w52351 and not w52354;
w52655 <= not w52653 and not w52654;
w52656 <= not w52471 and not w52655;
w52657 <= not w51850 and not w52470;
w52658 <= not w52469 and w52657;
w52659 <= not w52656 and not w52658;
w52660 <= not b(38) and not w52659;
w52661 <= not w51869 and w52349;
w52662 <= not w52345 and w52661;
w52663 <= not w52346 and not w52349;
w52664 <= not w52662 and not w52663;
w52665 <= not w52471 and not w52664;
w52666 <= not w51859 and not w52470;
w52667 <= not w52469 and w52666;
w52668 <= not w52665 and not w52667;
w52669 <= not b(37) and not w52668;
w52670 <= not w51878 and w52344;
w52671 <= not w52340 and w52670;
w52672 <= not w52341 and not w52344;
w52673 <= not w52671 and not w52672;
w52674 <= not w52471 and not w52673;
w52675 <= not w51868 and not w52470;
w52676 <= not w52469 and w52675;
w52677 <= not w52674 and not w52676;
w52678 <= not b(36) and not w52677;
w52679 <= not w51887 and w52339;
w52680 <= not w52335 and w52679;
w52681 <= not w52336 and not w52339;
w52682 <= not w52680 and not w52681;
w52683 <= not w52471 and not w52682;
w52684 <= not w51877 and not w52470;
w52685 <= not w52469 and w52684;
w52686 <= not w52683 and not w52685;
w52687 <= not b(35) and not w52686;
w52688 <= not w51896 and w52334;
w52689 <= not w52330 and w52688;
w52690 <= not w52331 and not w52334;
w52691 <= not w52689 and not w52690;
w52692 <= not w52471 and not w52691;
w52693 <= not w51886 and not w52470;
w52694 <= not w52469 and w52693;
w52695 <= not w52692 and not w52694;
w52696 <= not b(34) and not w52695;
w52697 <= not w51905 and w52329;
w52698 <= not w52325 and w52697;
w52699 <= not w52326 and not w52329;
w52700 <= not w52698 and not w52699;
w52701 <= not w52471 and not w52700;
w52702 <= not w51895 and not w52470;
w52703 <= not w52469 and w52702;
w52704 <= not w52701 and not w52703;
w52705 <= not b(33) and not w52704;
w52706 <= not w51914 and w52324;
w52707 <= not w52320 and w52706;
w52708 <= not w52321 and not w52324;
w52709 <= not w52707 and not w52708;
w52710 <= not w52471 and not w52709;
w52711 <= not w51904 and not w52470;
w52712 <= not w52469 and w52711;
w52713 <= not w52710 and not w52712;
w52714 <= not b(32) and not w52713;
w52715 <= not w51923 and w52319;
w52716 <= not w52315 and w52715;
w52717 <= not w52316 and not w52319;
w52718 <= not w52716 and not w52717;
w52719 <= not w52471 and not w52718;
w52720 <= not w51913 and not w52470;
w52721 <= not w52469 and w52720;
w52722 <= not w52719 and not w52721;
w52723 <= not b(31) and not w52722;
w52724 <= not w51932 and w52314;
w52725 <= not w52310 and w52724;
w52726 <= not w52311 and not w52314;
w52727 <= not w52725 and not w52726;
w52728 <= not w52471 and not w52727;
w52729 <= not w51922 and not w52470;
w52730 <= not w52469 and w52729;
w52731 <= not w52728 and not w52730;
w52732 <= not b(30) and not w52731;
w52733 <= not w51941 and w52309;
w52734 <= not w52305 and w52733;
w52735 <= not w52306 and not w52309;
w52736 <= not w52734 and not w52735;
w52737 <= not w52471 and not w52736;
w52738 <= not w51931 and not w52470;
w52739 <= not w52469 and w52738;
w52740 <= not w52737 and not w52739;
w52741 <= not b(29) and not w52740;
w52742 <= not w51950 and w52304;
w52743 <= not w52300 and w52742;
w52744 <= not w52301 and not w52304;
w52745 <= not w52743 and not w52744;
w52746 <= not w52471 and not w52745;
w52747 <= not w51940 and not w52470;
w52748 <= not w52469 and w52747;
w52749 <= not w52746 and not w52748;
w52750 <= not b(28) and not w52749;
w52751 <= not w51959 and w52299;
w52752 <= not w52295 and w52751;
w52753 <= not w52296 and not w52299;
w52754 <= not w52752 and not w52753;
w52755 <= not w52471 and not w52754;
w52756 <= not w51949 and not w52470;
w52757 <= not w52469 and w52756;
w52758 <= not w52755 and not w52757;
w52759 <= not b(27) and not w52758;
w52760 <= not w51968 and w52294;
w52761 <= not w52290 and w52760;
w52762 <= not w52291 and not w52294;
w52763 <= not w52761 and not w52762;
w52764 <= not w52471 and not w52763;
w52765 <= not w51958 and not w52470;
w52766 <= not w52469 and w52765;
w52767 <= not w52764 and not w52766;
w52768 <= not b(26) and not w52767;
w52769 <= not w51977 and w52289;
w52770 <= not w52285 and w52769;
w52771 <= not w52286 and not w52289;
w52772 <= not w52770 and not w52771;
w52773 <= not w52471 and not w52772;
w52774 <= not w51967 and not w52470;
w52775 <= not w52469 and w52774;
w52776 <= not w52773 and not w52775;
w52777 <= not b(25) and not w52776;
w52778 <= not w51986 and w52284;
w52779 <= not w52280 and w52778;
w52780 <= not w52281 and not w52284;
w52781 <= not w52779 and not w52780;
w52782 <= not w52471 and not w52781;
w52783 <= not w51976 and not w52470;
w52784 <= not w52469 and w52783;
w52785 <= not w52782 and not w52784;
w52786 <= not b(24) and not w52785;
w52787 <= not w51995 and w52279;
w52788 <= not w52275 and w52787;
w52789 <= not w52276 and not w52279;
w52790 <= not w52788 and not w52789;
w52791 <= not w52471 and not w52790;
w52792 <= not w51985 and not w52470;
w52793 <= not w52469 and w52792;
w52794 <= not w52791 and not w52793;
w52795 <= not b(23) and not w52794;
w52796 <= not w52004 and w52274;
w52797 <= not w52270 and w52796;
w52798 <= not w52271 and not w52274;
w52799 <= not w52797 and not w52798;
w52800 <= not w52471 and not w52799;
w52801 <= not w51994 and not w52470;
w52802 <= not w52469 and w52801;
w52803 <= not w52800 and not w52802;
w52804 <= not b(22) and not w52803;
w52805 <= not w52013 and w52269;
w52806 <= not w52265 and w52805;
w52807 <= not w52266 and not w52269;
w52808 <= not w52806 and not w52807;
w52809 <= not w52471 and not w52808;
w52810 <= not w52003 and not w52470;
w52811 <= not w52469 and w52810;
w52812 <= not w52809 and not w52811;
w52813 <= not b(21) and not w52812;
w52814 <= not w52022 and w52264;
w52815 <= not w52260 and w52814;
w52816 <= not w52261 and not w52264;
w52817 <= not w52815 and not w52816;
w52818 <= not w52471 and not w52817;
w52819 <= not w52012 and not w52470;
w52820 <= not w52469 and w52819;
w52821 <= not w52818 and not w52820;
w52822 <= not b(20) and not w52821;
w52823 <= not w52031 and w52259;
w52824 <= not w52255 and w52823;
w52825 <= not w52256 and not w52259;
w52826 <= not w52824 and not w52825;
w52827 <= not w52471 and not w52826;
w52828 <= not w52021 and not w52470;
w52829 <= not w52469 and w52828;
w52830 <= not w52827 and not w52829;
w52831 <= not b(19) and not w52830;
w52832 <= not w52040 and w52254;
w52833 <= not w52250 and w52832;
w52834 <= not w52251 and not w52254;
w52835 <= not w52833 and not w52834;
w52836 <= not w52471 and not w52835;
w52837 <= not w52030 and not w52470;
w52838 <= not w52469 and w52837;
w52839 <= not w52836 and not w52838;
w52840 <= not b(18) and not w52839;
w52841 <= not w52049 and w52249;
w52842 <= not w52245 and w52841;
w52843 <= not w52246 and not w52249;
w52844 <= not w52842 and not w52843;
w52845 <= not w52471 and not w52844;
w52846 <= not w52039 and not w52470;
w52847 <= not w52469 and w52846;
w52848 <= not w52845 and not w52847;
w52849 <= not b(17) and not w52848;
w52850 <= not w52058 and w52244;
w52851 <= not w52240 and w52850;
w52852 <= not w52241 and not w52244;
w52853 <= not w52851 and not w52852;
w52854 <= not w52471 and not w52853;
w52855 <= not w52048 and not w52470;
w52856 <= not w52469 and w52855;
w52857 <= not w52854 and not w52856;
w52858 <= not b(16) and not w52857;
w52859 <= not w52067 and w52239;
w52860 <= not w52235 and w52859;
w52861 <= not w52236 and not w52239;
w52862 <= not w52860 and not w52861;
w52863 <= not w52471 and not w52862;
w52864 <= not w52057 and not w52470;
w52865 <= not w52469 and w52864;
w52866 <= not w52863 and not w52865;
w52867 <= not b(15) and not w52866;
w52868 <= not w52076 and w52234;
w52869 <= not w52230 and w52868;
w52870 <= not w52231 and not w52234;
w52871 <= not w52869 and not w52870;
w52872 <= not w52471 and not w52871;
w52873 <= not w52066 and not w52470;
w52874 <= not w52469 and w52873;
w52875 <= not w52872 and not w52874;
w52876 <= not b(14) and not w52875;
w52877 <= not w52085 and w52229;
w52878 <= not w52225 and w52877;
w52879 <= not w52226 and not w52229;
w52880 <= not w52878 and not w52879;
w52881 <= not w52471 and not w52880;
w52882 <= not w52075 and not w52470;
w52883 <= not w52469 and w52882;
w52884 <= not w52881 and not w52883;
w52885 <= not b(13) and not w52884;
w52886 <= not w52094 and w52224;
w52887 <= not w52220 and w52886;
w52888 <= not w52221 and not w52224;
w52889 <= not w52887 and not w52888;
w52890 <= not w52471 and not w52889;
w52891 <= not w52084 and not w52470;
w52892 <= not w52469 and w52891;
w52893 <= not w52890 and not w52892;
w52894 <= not b(12) and not w52893;
w52895 <= not w52103 and w52219;
w52896 <= not w52215 and w52895;
w52897 <= not w52216 and not w52219;
w52898 <= not w52896 and not w52897;
w52899 <= not w52471 and not w52898;
w52900 <= not w52093 and not w52470;
w52901 <= not w52469 and w52900;
w52902 <= not w52899 and not w52901;
w52903 <= not b(11) and not w52902;
w52904 <= not w52112 and w52214;
w52905 <= not w52210 and w52904;
w52906 <= not w52211 and not w52214;
w52907 <= not w52905 and not w52906;
w52908 <= not w52471 and not w52907;
w52909 <= not w52102 and not w52470;
w52910 <= not w52469 and w52909;
w52911 <= not w52908 and not w52910;
w52912 <= not b(10) and not w52911;
w52913 <= not w52121 and w52209;
w52914 <= not w52205 and w52913;
w52915 <= not w52206 and not w52209;
w52916 <= not w52914 and not w52915;
w52917 <= not w52471 and not w52916;
w52918 <= not w52111 and not w52470;
w52919 <= not w52469 and w52918;
w52920 <= not w52917 and not w52919;
w52921 <= not b(9) and not w52920;
w52922 <= not w52130 and w52204;
w52923 <= not w52200 and w52922;
w52924 <= not w52201 and not w52204;
w52925 <= not w52923 and not w52924;
w52926 <= not w52471 and not w52925;
w52927 <= not w52120 and not w52470;
w52928 <= not w52469 and w52927;
w52929 <= not w52926 and not w52928;
w52930 <= not b(8) and not w52929;
w52931 <= not w52139 and w52199;
w52932 <= not w52195 and w52931;
w52933 <= not w52196 and not w52199;
w52934 <= not w52932 and not w52933;
w52935 <= not w52471 and not w52934;
w52936 <= not w52129 and not w52470;
w52937 <= not w52469 and w52936;
w52938 <= not w52935 and not w52937;
w52939 <= not b(7) and not w52938;
w52940 <= not w52148 and w52194;
w52941 <= not w52190 and w52940;
w52942 <= not w52191 and not w52194;
w52943 <= not w52941 and not w52942;
w52944 <= not w52471 and not w52943;
w52945 <= not w52138 and not w52470;
w52946 <= not w52469 and w52945;
w52947 <= not w52944 and not w52946;
w52948 <= not b(6) and not w52947;
w52949 <= not w52157 and w52189;
w52950 <= not w52185 and w52949;
w52951 <= not w52186 and not w52189;
w52952 <= not w52950 and not w52951;
w52953 <= not w52471 and not w52952;
w52954 <= not w52147 and not w52470;
w52955 <= not w52469 and w52954;
w52956 <= not w52953 and not w52955;
w52957 <= not b(5) and not w52956;
w52958 <= not w52165 and w52184;
w52959 <= not w52180 and w52958;
w52960 <= not w52181 and not w52184;
w52961 <= not w52959 and not w52960;
w52962 <= not w52471 and not w52961;
w52963 <= not w52156 and not w52470;
w52964 <= not w52469 and w52963;
w52965 <= not w52962 and not w52964;
w52966 <= not b(4) and not w52965;
w52967 <= not w52175 and w52179;
w52968 <= not w52174 and w52967;
w52969 <= not w52176 and not w52179;
w52970 <= not w52968 and not w52969;
w52971 <= not w52471 and not w52970;
w52972 <= not w52164 and not w52470;
w52973 <= not w52469 and w52972;
w52974 <= not w52971 and not w52973;
w52975 <= not b(3) and not w52974;
w52976 <= w24156 and not w52172;
w52977 <= not w52170 and w52976;
w52978 <= not w52174 and not w52977;
w52979 <= not w52471 and w52978;
w52980 <= not w52169 and not w52470;
w52981 <= not w52469 and w52980;
w52982 <= not w52979 and not w52981;
w52983 <= not b(2) and not w52982;
w52984 <= b(0) and not w52471;
w52985 <= a(5) and not w52984;
w52986 <= w24156 and not w52471;
w52987 <= not w52985 and not w52986;
w52988 <= b(1) and not w52987;
w52989 <= not b(1) and not w52986;
w52990 <= not w52985 and w52989;
w52991 <= not w52988 and not w52990;
w52992 <= not w24976 and not w52991;
w52993 <= not b(1) and not w52987;
w52994 <= not w52992 and not w52993;
w52995 <= b(2) and not w52981;
w52996 <= not w52979 and w52995;
w52997 <= not w52983 and not w52996;
w52998 <= not w52994 and w52997;
w52999 <= not w52983 and not w52998;
w53000 <= b(3) and not w52973;
w53001 <= not w52971 and w53000;
w53002 <= not w52975 and not w53001;
w53003 <= not w52999 and w53002;
w53004 <= not w52975 and not w53003;
w53005 <= b(4) and not w52964;
w53006 <= not w52962 and w53005;
w53007 <= not w52966 and not w53006;
w53008 <= not w53004 and w53007;
w53009 <= not w52966 and not w53008;
w53010 <= b(5) and not w52955;
w53011 <= not w52953 and w53010;
w53012 <= not w52957 and not w53011;
w53013 <= not w53009 and w53012;
w53014 <= not w52957 and not w53013;
w53015 <= b(6) and not w52946;
w53016 <= not w52944 and w53015;
w53017 <= not w52948 and not w53016;
w53018 <= not w53014 and w53017;
w53019 <= not w52948 and not w53018;
w53020 <= b(7) and not w52937;
w53021 <= not w52935 and w53020;
w53022 <= not w52939 and not w53021;
w53023 <= not w53019 and w53022;
w53024 <= not w52939 and not w53023;
w53025 <= b(8) and not w52928;
w53026 <= not w52926 and w53025;
w53027 <= not w52930 and not w53026;
w53028 <= not w53024 and w53027;
w53029 <= not w52930 and not w53028;
w53030 <= b(9) and not w52919;
w53031 <= not w52917 and w53030;
w53032 <= not w52921 and not w53031;
w53033 <= not w53029 and w53032;
w53034 <= not w52921 and not w53033;
w53035 <= b(10) and not w52910;
w53036 <= not w52908 and w53035;
w53037 <= not w52912 and not w53036;
w53038 <= not w53034 and w53037;
w53039 <= not w52912 and not w53038;
w53040 <= b(11) and not w52901;
w53041 <= not w52899 and w53040;
w53042 <= not w52903 and not w53041;
w53043 <= not w53039 and w53042;
w53044 <= not w52903 and not w53043;
w53045 <= b(12) and not w52892;
w53046 <= not w52890 and w53045;
w53047 <= not w52894 and not w53046;
w53048 <= not w53044 and w53047;
w53049 <= not w52894 and not w53048;
w53050 <= b(13) and not w52883;
w53051 <= not w52881 and w53050;
w53052 <= not w52885 and not w53051;
w53053 <= not w53049 and w53052;
w53054 <= not w52885 and not w53053;
w53055 <= b(14) and not w52874;
w53056 <= not w52872 and w53055;
w53057 <= not w52876 and not w53056;
w53058 <= not w53054 and w53057;
w53059 <= not w52876 and not w53058;
w53060 <= b(15) and not w52865;
w53061 <= not w52863 and w53060;
w53062 <= not w52867 and not w53061;
w53063 <= not w53059 and w53062;
w53064 <= not w52867 and not w53063;
w53065 <= b(16) and not w52856;
w53066 <= not w52854 and w53065;
w53067 <= not w52858 and not w53066;
w53068 <= not w53064 and w53067;
w53069 <= not w52858 and not w53068;
w53070 <= b(17) and not w52847;
w53071 <= not w52845 and w53070;
w53072 <= not w52849 and not w53071;
w53073 <= not w53069 and w53072;
w53074 <= not w52849 and not w53073;
w53075 <= b(18) and not w52838;
w53076 <= not w52836 and w53075;
w53077 <= not w52840 and not w53076;
w53078 <= not w53074 and w53077;
w53079 <= not w52840 and not w53078;
w53080 <= b(19) and not w52829;
w53081 <= not w52827 and w53080;
w53082 <= not w52831 and not w53081;
w53083 <= not w53079 and w53082;
w53084 <= not w52831 and not w53083;
w53085 <= b(20) and not w52820;
w53086 <= not w52818 and w53085;
w53087 <= not w52822 and not w53086;
w53088 <= not w53084 and w53087;
w53089 <= not w52822 and not w53088;
w53090 <= b(21) and not w52811;
w53091 <= not w52809 and w53090;
w53092 <= not w52813 and not w53091;
w53093 <= not w53089 and w53092;
w53094 <= not w52813 and not w53093;
w53095 <= b(22) and not w52802;
w53096 <= not w52800 and w53095;
w53097 <= not w52804 and not w53096;
w53098 <= not w53094 and w53097;
w53099 <= not w52804 and not w53098;
w53100 <= b(23) and not w52793;
w53101 <= not w52791 and w53100;
w53102 <= not w52795 and not w53101;
w53103 <= not w53099 and w53102;
w53104 <= not w52795 and not w53103;
w53105 <= b(24) and not w52784;
w53106 <= not w52782 and w53105;
w53107 <= not w52786 and not w53106;
w53108 <= not w53104 and w53107;
w53109 <= not w52786 and not w53108;
w53110 <= b(25) and not w52775;
w53111 <= not w52773 and w53110;
w53112 <= not w52777 and not w53111;
w53113 <= not w53109 and w53112;
w53114 <= not w52777 and not w53113;
w53115 <= b(26) and not w52766;
w53116 <= not w52764 and w53115;
w53117 <= not w52768 and not w53116;
w53118 <= not w53114 and w53117;
w53119 <= not w52768 and not w53118;
w53120 <= b(27) and not w52757;
w53121 <= not w52755 and w53120;
w53122 <= not w52759 and not w53121;
w53123 <= not w53119 and w53122;
w53124 <= not w52759 and not w53123;
w53125 <= b(28) and not w52748;
w53126 <= not w52746 and w53125;
w53127 <= not w52750 and not w53126;
w53128 <= not w53124 and w53127;
w53129 <= not w52750 and not w53128;
w53130 <= b(29) and not w52739;
w53131 <= not w52737 and w53130;
w53132 <= not w52741 and not w53131;
w53133 <= not w53129 and w53132;
w53134 <= not w52741 and not w53133;
w53135 <= b(30) and not w52730;
w53136 <= not w52728 and w53135;
w53137 <= not w52732 and not w53136;
w53138 <= not w53134 and w53137;
w53139 <= not w52732 and not w53138;
w53140 <= b(31) and not w52721;
w53141 <= not w52719 and w53140;
w53142 <= not w52723 and not w53141;
w53143 <= not w53139 and w53142;
w53144 <= not w52723 and not w53143;
w53145 <= b(32) and not w52712;
w53146 <= not w52710 and w53145;
w53147 <= not w52714 and not w53146;
w53148 <= not w53144 and w53147;
w53149 <= not w52714 and not w53148;
w53150 <= b(33) and not w52703;
w53151 <= not w52701 and w53150;
w53152 <= not w52705 and not w53151;
w53153 <= not w53149 and w53152;
w53154 <= not w52705 and not w53153;
w53155 <= b(34) and not w52694;
w53156 <= not w52692 and w53155;
w53157 <= not w52696 and not w53156;
w53158 <= not w53154 and w53157;
w53159 <= not w52696 and not w53158;
w53160 <= b(35) and not w52685;
w53161 <= not w52683 and w53160;
w53162 <= not w52687 and not w53161;
w53163 <= not w53159 and w53162;
w53164 <= not w52687 and not w53163;
w53165 <= b(36) and not w52676;
w53166 <= not w52674 and w53165;
w53167 <= not w52678 and not w53166;
w53168 <= not w53164 and w53167;
w53169 <= not w52678 and not w53168;
w53170 <= b(37) and not w52667;
w53171 <= not w52665 and w53170;
w53172 <= not w52669 and not w53171;
w53173 <= not w53169 and w53172;
w53174 <= not w52669 and not w53173;
w53175 <= b(38) and not w52658;
w53176 <= not w52656 and w53175;
w53177 <= not w52660 and not w53176;
w53178 <= not w53174 and w53177;
w53179 <= not w52660 and not w53178;
w53180 <= b(39) and not w52649;
w53181 <= not w52647 and w53180;
w53182 <= not w52651 and not w53181;
w53183 <= not w53179 and w53182;
w53184 <= not w52651 and not w53183;
w53185 <= b(40) and not w52640;
w53186 <= not w52638 and w53185;
w53187 <= not w52642 and not w53186;
w53188 <= not w53184 and w53187;
w53189 <= not w52642 and not w53188;
w53190 <= b(41) and not w52631;
w53191 <= not w52629 and w53190;
w53192 <= not w52633 and not w53191;
w53193 <= not w53189 and w53192;
w53194 <= not w52633 and not w53193;
w53195 <= b(42) and not w52622;
w53196 <= not w52620 and w53195;
w53197 <= not w52624 and not w53196;
w53198 <= not w53194 and w53197;
w53199 <= not w52624 and not w53198;
w53200 <= b(43) and not w52613;
w53201 <= not w52611 and w53200;
w53202 <= not w52615 and not w53201;
w53203 <= not w53199 and w53202;
w53204 <= not w52615 and not w53203;
w53205 <= b(44) and not w52604;
w53206 <= not w52602 and w53205;
w53207 <= not w52606 and not w53206;
w53208 <= not w53204 and w53207;
w53209 <= not w52606 and not w53208;
w53210 <= b(45) and not w52595;
w53211 <= not w52593 and w53210;
w53212 <= not w52597 and not w53211;
w53213 <= not w53209 and w53212;
w53214 <= not w52597 and not w53213;
w53215 <= b(46) and not w52586;
w53216 <= not w52584 and w53215;
w53217 <= not w52588 and not w53216;
w53218 <= not w53214 and w53217;
w53219 <= not w52588 and not w53218;
w53220 <= b(47) and not w52577;
w53221 <= not w52575 and w53220;
w53222 <= not w52579 and not w53221;
w53223 <= not w53219 and w53222;
w53224 <= not w52579 and not w53223;
w53225 <= b(48) and not w52568;
w53226 <= not w52566 and w53225;
w53227 <= not w52570 and not w53226;
w53228 <= not w53224 and w53227;
w53229 <= not w52570 and not w53228;
w53230 <= b(49) and not w52559;
w53231 <= not w52557 and w53230;
w53232 <= not w52561 and not w53231;
w53233 <= not w53229 and w53232;
w53234 <= not w52561 and not w53233;
w53235 <= b(50) and not w52550;
w53236 <= not w52548 and w53235;
w53237 <= not w52552 and not w53236;
w53238 <= not w53234 and w53237;
w53239 <= not w52552 and not w53238;
w53240 <= b(51) and not w52541;
w53241 <= not w52539 and w53240;
w53242 <= not w52543 and not w53241;
w53243 <= not w53239 and w53242;
w53244 <= not w52543 and not w53243;
w53245 <= b(52) and not w52532;
w53246 <= not w52530 and w53245;
w53247 <= not w52534 and not w53246;
w53248 <= not w53244 and w53247;
w53249 <= not w52534 and not w53248;
w53250 <= b(53) and not w52523;
w53251 <= not w52521 and w53250;
w53252 <= not w52525 and not w53251;
w53253 <= not w53249 and w53252;
w53254 <= not w52525 and not w53253;
w53255 <= b(54) and not w52514;
w53256 <= not w52512 and w53255;
w53257 <= not w52516 and not w53256;
w53258 <= not w53254 and w53257;
w53259 <= not w52516 and not w53258;
w53260 <= b(55) and not w52505;
w53261 <= not w52503 and w53260;
w53262 <= not w52507 and not w53261;
w53263 <= not w53259 and w53262;
w53264 <= not w52507 and not w53263;
w53265 <= b(56) and not w52496;
w53266 <= not w52494 and w53265;
w53267 <= not w52498 and not w53266;
w53268 <= not w53264 and w53267;
w53269 <= not w52498 and not w53268;
w53270 <= b(57) and not w52487;
w53271 <= not w52485 and w53270;
w53272 <= not w52489 and not w53271;
w53273 <= not w53269 and w53272;
w53274 <= not w52489 and not w53273;
w53275 <= b(58) and not w52478;
w53276 <= not w52476 and w53275;
w53277 <= not w52480 and not w53276;
w53278 <= not w53274 and w53277;
w53279 <= not w52480 and not w53278;
w53280 <= not w51671 and not w52466;
w53281 <= not w52464 and w53280;
w53282 <= not w52455 and w53281;
w53283 <= not w52464 and not w52466;
w53284 <= not w52456 and not w53283;
w53285 <= not w53282 and not w53284;
w53286 <= not w52471 and not w53285;
w53287 <= not w52463 and not w52470;
w53288 <= not w52469 and w53287;
w53289 <= not w53286 and not w53288;
w53290 <= not b(59) and not w53289;
w53291 <= b(59) and not w53288;
w53292 <= not w53286 and w53291;
w53293 <= w23 and not w53292;
w53294 <= not w53290 and w53293;
w53295 <= not w53279 and w53294;
w53296 <= w24450 and not w53289;
w53297 <= not w53295 and not w53296;
w53298 <= not w52489 and w53277;
w53299 <= not w53273 and w53298;
w53300 <= not w53274 and not w53277;
w53301 <= not w53299 and not w53300;
w53302 <= not w53297 and not w53301;
w53303 <= not w52479 and not w53296;
w53304 <= not w53295 and w53303;
w53305 <= not w53302 and not w53304;
w53306 <= not b(59) and not w53305;
w53307 <= not w52498 and w53272;
w53308 <= not w53268 and w53307;
w53309 <= not w53269 and not w53272;
w53310 <= not w53308 and not w53309;
w53311 <= not w53297 and not w53310;
w53312 <= not w52488 and not w53296;
w53313 <= not w53295 and w53312;
w53314 <= not w53311 and not w53313;
w53315 <= not b(58) and not w53314;
w53316 <= not w52507 and w53267;
w53317 <= not w53263 and w53316;
w53318 <= not w53264 and not w53267;
w53319 <= not w53317 and not w53318;
w53320 <= not w53297 and not w53319;
w53321 <= not w52497 and not w53296;
w53322 <= not w53295 and w53321;
w53323 <= not w53320 and not w53322;
w53324 <= not b(57) and not w53323;
w53325 <= not w52516 and w53262;
w53326 <= not w53258 and w53325;
w53327 <= not w53259 and not w53262;
w53328 <= not w53326 and not w53327;
w53329 <= not w53297 and not w53328;
w53330 <= not w52506 and not w53296;
w53331 <= not w53295 and w53330;
w53332 <= not w53329 and not w53331;
w53333 <= not b(56) and not w53332;
w53334 <= not w52525 and w53257;
w53335 <= not w53253 and w53334;
w53336 <= not w53254 and not w53257;
w53337 <= not w53335 and not w53336;
w53338 <= not w53297 and not w53337;
w53339 <= not w52515 and not w53296;
w53340 <= not w53295 and w53339;
w53341 <= not w53338 and not w53340;
w53342 <= not b(55) and not w53341;
w53343 <= not w52534 and w53252;
w53344 <= not w53248 and w53343;
w53345 <= not w53249 and not w53252;
w53346 <= not w53344 and not w53345;
w53347 <= not w53297 and not w53346;
w53348 <= not w52524 and not w53296;
w53349 <= not w53295 and w53348;
w53350 <= not w53347 and not w53349;
w53351 <= not b(54) and not w53350;
w53352 <= not w52543 and w53247;
w53353 <= not w53243 and w53352;
w53354 <= not w53244 and not w53247;
w53355 <= not w53353 and not w53354;
w53356 <= not w53297 and not w53355;
w53357 <= not w52533 and not w53296;
w53358 <= not w53295 and w53357;
w53359 <= not w53356 and not w53358;
w53360 <= not b(53) and not w53359;
w53361 <= not w52552 and w53242;
w53362 <= not w53238 and w53361;
w53363 <= not w53239 and not w53242;
w53364 <= not w53362 and not w53363;
w53365 <= not w53297 and not w53364;
w53366 <= not w52542 and not w53296;
w53367 <= not w53295 and w53366;
w53368 <= not w53365 and not w53367;
w53369 <= not b(52) and not w53368;
w53370 <= not w52561 and w53237;
w53371 <= not w53233 and w53370;
w53372 <= not w53234 and not w53237;
w53373 <= not w53371 and not w53372;
w53374 <= not w53297 and not w53373;
w53375 <= not w52551 and not w53296;
w53376 <= not w53295 and w53375;
w53377 <= not w53374 and not w53376;
w53378 <= not b(51) and not w53377;
w53379 <= not w52570 and w53232;
w53380 <= not w53228 and w53379;
w53381 <= not w53229 and not w53232;
w53382 <= not w53380 and not w53381;
w53383 <= not w53297 and not w53382;
w53384 <= not w52560 and not w53296;
w53385 <= not w53295 and w53384;
w53386 <= not w53383 and not w53385;
w53387 <= not b(50) and not w53386;
w53388 <= not w52579 and w53227;
w53389 <= not w53223 and w53388;
w53390 <= not w53224 and not w53227;
w53391 <= not w53389 and not w53390;
w53392 <= not w53297 and not w53391;
w53393 <= not w52569 and not w53296;
w53394 <= not w53295 and w53393;
w53395 <= not w53392 and not w53394;
w53396 <= not b(49) and not w53395;
w53397 <= not w52588 and w53222;
w53398 <= not w53218 and w53397;
w53399 <= not w53219 and not w53222;
w53400 <= not w53398 and not w53399;
w53401 <= not w53297 and not w53400;
w53402 <= not w52578 and not w53296;
w53403 <= not w53295 and w53402;
w53404 <= not w53401 and not w53403;
w53405 <= not b(48) and not w53404;
w53406 <= not w52597 and w53217;
w53407 <= not w53213 and w53406;
w53408 <= not w53214 and not w53217;
w53409 <= not w53407 and not w53408;
w53410 <= not w53297 and not w53409;
w53411 <= not w52587 and not w53296;
w53412 <= not w53295 and w53411;
w53413 <= not w53410 and not w53412;
w53414 <= not b(47) and not w53413;
w53415 <= not w52606 and w53212;
w53416 <= not w53208 and w53415;
w53417 <= not w53209 and not w53212;
w53418 <= not w53416 and not w53417;
w53419 <= not w53297 and not w53418;
w53420 <= not w52596 and not w53296;
w53421 <= not w53295 and w53420;
w53422 <= not w53419 and not w53421;
w53423 <= not b(46) and not w53422;
w53424 <= not w52615 and w53207;
w53425 <= not w53203 and w53424;
w53426 <= not w53204 and not w53207;
w53427 <= not w53425 and not w53426;
w53428 <= not w53297 and not w53427;
w53429 <= not w52605 and not w53296;
w53430 <= not w53295 and w53429;
w53431 <= not w53428 and not w53430;
w53432 <= not b(45) and not w53431;
w53433 <= not w52624 and w53202;
w53434 <= not w53198 and w53433;
w53435 <= not w53199 and not w53202;
w53436 <= not w53434 and not w53435;
w53437 <= not w53297 and not w53436;
w53438 <= not w52614 and not w53296;
w53439 <= not w53295 and w53438;
w53440 <= not w53437 and not w53439;
w53441 <= not b(44) and not w53440;
w53442 <= not w52633 and w53197;
w53443 <= not w53193 and w53442;
w53444 <= not w53194 and not w53197;
w53445 <= not w53443 and not w53444;
w53446 <= not w53297 and not w53445;
w53447 <= not w52623 and not w53296;
w53448 <= not w53295 and w53447;
w53449 <= not w53446 and not w53448;
w53450 <= not b(43) and not w53449;
w53451 <= not w52642 and w53192;
w53452 <= not w53188 and w53451;
w53453 <= not w53189 and not w53192;
w53454 <= not w53452 and not w53453;
w53455 <= not w53297 and not w53454;
w53456 <= not w52632 and not w53296;
w53457 <= not w53295 and w53456;
w53458 <= not w53455 and not w53457;
w53459 <= not b(42) and not w53458;
w53460 <= not w52651 and w53187;
w53461 <= not w53183 and w53460;
w53462 <= not w53184 and not w53187;
w53463 <= not w53461 and not w53462;
w53464 <= not w53297 and not w53463;
w53465 <= not w52641 and not w53296;
w53466 <= not w53295 and w53465;
w53467 <= not w53464 and not w53466;
w53468 <= not b(41) and not w53467;
w53469 <= not w52660 and w53182;
w53470 <= not w53178 and w53469;
w53471 <= not w53179 and not w53182;
w53472 <= not w53470 and not w53471;
w53473 <= not w53297 and not w53472;
w53474 <= not w52650 and not w53296;
w53475 <= not w53295 and w53474;
w53476 <= not w53473 and not w53475;
w53477 <= not b(40) and not w53476;
w53478 <= not w52669 and w53177;
w53479 <= not w53173 and w53478;
w53480 <= not w53174 and not w53177;
w53481 <= not w53479 and not w53480;
w53482 <= not w53297 and not w53481;
w53483 <= not w52659 and not w53296;
w53484 <= not w53295 and w53483;
w53485 <= not w53482 and not w53484;
w53486 <= not b(39) and not w53485;
w53487 <= not w52678 and w53172;
w53488 <= not w53168 and w53487;
w53489 <= not w53169 and not w53172;
w53490 <= not w53488 and not w53489;
w53491 <= not w53297 and not w53490;
w53492 <= not w52668 and not w53296;
w53493 <= not w53295 and w53492;
w53494 <= not w53491 and not w53493;
w53495 <= not b(38) and not w53494;
w53496 <= not w52687 and w53167;
w53497 <= not w53163 and w53496;
w53498 <= not w53164 and not w53167;
w53499 <= not w53497 and not w53498;
w53500 <= not w53297 and not w53499;
w53501 <= not w52677 and not w53296;
w53502 <= not w53295 and w53501;
w53503 <= not w53500 and not w53502;
w53504 <= not b(37) and not w53503;
w53505 <= not w52696 and w53162;
w53506 <= not w53158 and w53505;
w53507 <= not w53159 and not w53162;
w53508 <= not w53506 and not w53507;
w53509 <= not w53297 and not w53508;
w53510 <= not w52686 and not w53296;
w53511 <= not w53295 and w53510;
w53512 <= not w53509 and not w53511;
w53513 <= not b(36) and not w53512;
w53514 <= not w52705 and w53157;
w53515 <= not w53153 and w53514;
w53516 <= not w53154 and not w53157;
w53517 <= not w53515 and not w53516;
w53518 <= not w53297 and not w53517;
w53519 <= not w52695 and not w53296;
w53520 <= not w53295 and w53519;
w53521 <= not w53518 and not w53520;
w53522 <= not b(35) and not w53521;
w53523 <= not w52714 and w53152;
w53524 <= not w53148 and w53523;
w53525 <= not w53149 and not w53152;
w53526 <= not w53524 and not w53525;
w53527 <= not w53297 and not w53526;
w53528 <= not w52704 and not w53296;
w53529 <= not w53295 and w53528;
w53530 <= not w53527 and not w53529;
w53531 <= not b(34) and not w53530;
w53532 <= not w52723 and w53147;
w53533 <= not w53143 and w53532;
w53534 <= not w53144 and not w53147;
w53535 <= not w53533 and not w53534;
w53536 <= not w53297 and not w53535;
w53537 <= not w52713 and not w53296;
w53538 <= not w53295 and w53537;
w53539 <= not w53536 and not w53538;
w53540 <= not b(33) and not w53539;
w53541 <= not w52732 and w53142;
w53542 <= not w53138 and w53541;
w53543 <= not w53139 and not w53142;
w53544 <= not w53542 and not w53543;
w53545 <= not w53297 and not w53544;
w53546 <= not w52722 and not w53296;
w53547 <= not w53295 and w53546;
w53548 <= not w53545 and not w53547;
w53549 <= not b(32) and not w53548;
w53550 <= not w52741 and w53137;
w53551 <= not w53133 and w53550;
w53552 <= not w53134 and not w53137;
w53553 <= not w53551 and not w53552;
w53554 <= not w53297 and not w53553;
w53555 <= not w52731 and not w53296;
w53556 <= not w53295 and w53555;
w53557 <= not w53554 and not w53556;
w53558 <= not b(31) and not w53557;
w53559 <= not w52750 and w53132;
w53560 <= not w53128 and w53559;
w53561 <= not w53129 and not w53132;
w53562 <= not w53560 and not w53561;
w53563 <= not w53297 and not w53562;
w53564 <= not w52740 and not w53296;
w53565 <= not w53295 and w53564;
w53566 <= not w53563 and not w53565;
w53567 <= not b(30) and not w53566;
w53568 <= not w52759 and w53127;
w53569 <= not w53123 and w53568;
w53570 <= not w53124 and not w53127;
w53571 <= not w53569 and not w53570;
w53572 <= not w53297 and not w53571;
w53573 <= not w52749 and not w53296;
w53574 <= not w53295 and w53573;
w53575 <= not w53572 and not w53574;
w53576 <= not b(29) and not w53575;
w53577 <= not w52768 and w53122;
w53578 <= not w53118 and w53577;
w53579 <= not w53119 and not w53122;
w53580 <= not w53578 and not w53579;
w53581 <= not w53297 and not w53580;
w53582 <= not w52758 and not w53296;
w53583 <= not w53295 and w53582;
w53584 <= not w53581 and not w53583;
w53585 <= not b(28) and not w53584;
w53586 <= not w52777 and w53117;
w53587 <= not w53113 and w53586;
w53588 <= not w53114 and not w53117;
w53589 <= not w53587 and not w53588;
w53590 <= not w53297 and not w53589;
w53591 <= not w52767 and not w53296;
w53592 <= not w53295 and w53591;
w53593 <= not w53590 and not w53592;
w53594 <= not b(27) and not w53593;
w53595 <= not w52786 and w53112;
w53596 <= not w53108 and w53595;
w53597 <= not w53109 and not w53112;
w53598 <= not w53596 and not w53597;
w53599 <= not w53297 and not w53598;
w53600 <= not w52776 and not w53296;
w53601 <= not w53295 and w53600;
w53602 <= not w53599 and not w53601;
w53603 <= not b(26) and not w53602;
w53604 <= not w52795 and w53107;
w53605 <= not w53103 and w53604;
w53606 <= not w53104 and not w53107;
w53607 <= not w53605 and not w53606;
w53608 <= not w53297 and not w53607;
w53609 <= not w52785 and not w53296;
w53610 <= not w53295 and w53609;
w53611 <= not w53608 and not w53610;
w53612 <= not b(25) and not w53611;
w53613 <= not w52804 and w53102;
w53614 <= not w53098 and w53613;
w53615 <= not w53099 and not w53102;
w53616 <= not w53614 and not w53615;
w53617 <= not w53297 and not w53616;
w53618 <= not w52794 and not w53296;
w53619 <= not w53295 and w53618;
w53620 <= not w53617 and not w53619;
w53621 <= not b(24) and not w53620;
w53622 <= not w52813 and w53097;
w53623 <= not w53093 and w53622;
w53624 <= not w53094 and not w53097;
w53625 <= not w53623 and not w53624;
w53626 <= not w53297 and not w53625;
w53627 <= not w52803 and not w53296;
w53628 <= not w53295 and w53627;
w53629 <= not w53626 and not w53628;
w53630 <= not b(23) and not w53629;
w53631 <= not w52822 and w53092;
w53632 <= not w53088 and w53631;
w53633 <= not w53089 and not w53092;
w53634 <= not w53632 and not w53633;
w53635 <= not w53297 and not w53634;
w53636 <= not w52812 and not w53296;
w53637 <= not w53295 and w53636;
w53638 <= not w53635 and not w53637;
w53639 <= not b(22) and not w53638;
w53640 <= not w52831 and w53087;
w53641 <= not w53083 and w53640;
w53642 <= not w53084 and not w53087;
w53643 <= not w53641 and not w53642;
w53644 <= not w53297 and not w53643;
w53645 <= not w52821 and not w53296;
w53646 <= not w53295 and w53645;
w53647 <= not w53644 and not w53646;
w53648 <= not b(21) and not w53647;
w53649 <= not w52840 and w53082;
w53650 <= not w53078 and w53649;
w53651 <= not w53079 and not w53082;
w53652 <= not w53650 and not w53651;
w53653 <= not w53297 and not w53652;
w53654 <= not w52830 and not w53296;
w53655 <= not w53295 and w53654;
w53656 <= not w53653 and not w53655;
w53657 <= not b(20) and not w53656;
w53658 <= not w52849 and w53077;
w53659 <= not w53073 and w53658;
w53660 <= not w53074 and not w53077;
w53661 <= not w53659 and not w53660;
w53662 <= not w53297 and not w53661;
w53663 <= not w52839 and not w53296;
w53664 <= not w53295 and w53663;
w53665 <= not w53662 and not w53664;
w53666 <= not b(19) and not w53665;
w53667 <= not w52858 and w53072;
w53668 <= not w53068 and w53667;
w53669 <= not w53069 and not w53072;
w53670 <= not w53668 and not w53669;
w53671 <= not w53297 and not w53670;
w53672 <= not w52848 and not w53296;
w53673 <= not w53295 and w53672;
w53674 <= not w53671 and not w53673;
w53675 <= not b(18) and not w53674;
w53676 <= not w52867 and w53067;
w53677 <= not w53063 and w53676;
w53678 <= not w53064 and not w53067;
w53679 <= not w53677 and not w53678;
w53680 <= not w53297 and not w53679;
w53681 <= not w52857 and not w53296;
w53682 <= not w53295 and w53681;
w53683 <= not w53680 and not w53682;
w53684 <= not b(17) and not w53683;
w53685 <= not w52876 and w53062;
w53686 <= not w53058 and w53685;
w53687 <= not w53059 and not w53062;
w53688 <= not w53686 and not w53687;
w53689 <= not w53297 and not w53688;
w53690 <= not w52866 and not w53296;
w53691 <= not w53295 and w53690;
w53692 <= not w53689 and not w53691;
w53693 <= not b(16) and not w53692;
w53694 <= not w52885 and w53057;
w53695 <= not w53053 and w53694;
w53696 <= not w53054 and not w53057;
w53697 <= not w53695 and not w53696;
w53698 <= not w53297 and not w53697;
w53699 <= not w52875 and not w53296;
w53700 <= not w53295 and w53699;
w53701 <= not w53698 and not w53700;
w53702 <= not b(15) and not w53701;
w53703 <= not w52894 and w53052;
w53704 <= not w53048 and w53703;
w53705 <= not w53049 and not w53052;
w53706 <= not w53704 and not w53705;
w53707 <= not w53297 and not w53706;
w53708 <= not w52884 and not w53296;
w53709 <= not w53295 and w53708;
w53710 <= not w53707 and not w53709;
w53711 <= not b(14) and not w53710;
w53712 <= not w52903 and w53047;
w53713 <= not w53043 and w53712;
w53714 <= not w53044 and not w53047;
w53715 <= not w53713 and not w53714;
w53716 <= not w53297 and not w53715;
w53717 <= not w52893 and not w53296;
w53718 <= not w53295 and w53717;
w53719 <= not w53716 and not w53718;
w53720 <= not b(13) and not w53719;
w53721 <= not w52912 and w53042;
w53722 <= not w53038 and w53721;
w53723 <= not w53039 and not w53042;
w53724 <= not w53722 and not w53723;
w53725 <= not w53297 and not w53724;
w53726 <= not w52902 and not w53296;
w53727 <= not w53295 and w53726;
w53728 <= not w53725 and not w53727;
w53729 <= not b(12) and not w53728;
w53730 <= not w52921 and w53037;
w53731 <= not w53033 and w53730;
w53732 <= not w53034 and not w53037;
w53733 <= not w53731 and not w53732;
w53734 <= not w53297 and not w53733;
w53735 <= not w52911 and not w53296;
w53736 <= not w53295 and w53735;
w53737 <= not w53734 and not w53736;
w53738 <= not b(11) and not w53737;
w53739 <= not w52930 and w53032;
w53740 <= not w53028 and w53739;
w53741 <= not w53029 and not w53032;
w53742 <= not w53740 and not w53741;
w53743 <= not w53297 and not w53742;
w53744 <= not w52920 and not w53296;
w53745 <= not w53295 and w53744;
w53746 <= not w53743 and not w53745;
w53747 <= not b(10) and not w53746;
w53748 <= not w52939 and w53027;
w53749 <= not w53023 and w53748;
w53750 <= not w53024 and not w53027;
w53751 <= not w53749 and not w53750;
w53752 <= not w53297 and not w53751;
w53753 <= not w52929 and not w53296;
w53754 <= not w53295 and w53753;
w53755 <= not w53752 and not w53754;
w53756 <= not b(9) and not w53755;
w53757 <= not w52948 and w53022;
w53758 <= not w53018 and w53757;
w53759 <= not w53019 and not w53022;
w53760 <= not w53758 and not w53759;
w53761 <= not w53297 and not w53760;
w53762 <= not w52938 and not w53296;
w53763 <= not w53295 and w53762;
w53764 <= not w53761 and not w53763;
w53765 <= not b(8) and not w53764;
w53766 <= not w52957 and w53017;
w53767 <= not w53013 and w53766;
w53768 <= not w53014 and not w53017;
w53769 <= not w53767 and not w53768;
w53770 <= not w53297 and not w53769;
w53771 <= not w52947 and not w53296;
w53772 <= not w53295 and w53771;
w53773 <= not w53770 and not w53772;
w53774 <= not b(7) and not w53773;
w53775 <= not w52966 and w53012;
w53776 <= not w53008 and w53775;
w53777 <= not w53009 and not w53012;
w53778 <= not w53776 and not w53777;
w53779 <= not w53297 and not w53778;
w53780 <= not w52956 and not w53296;
w53781 <= not w53295 and w53780;
w53782 <= not w53779 and not w53781;
w53783 <= not b(6) and not w53782;
w53784 <= not w52975 and w53007;
w53785 <= not w53003 and w53784;
w53786 <= not w53004 and not w53007;
w53787 <= not w53785 and not w53786;
w53788 <= not w53297 and not w53787;
w53789 <= not w52965 and not w53296;
w53790 <= not w53295 and w53789;
w53791 <= not w53788 and not w53790;
w53792 <= not b(5) and not w53791;
w53793 <= not w52983 and w53002;
w53794 <= not w52998 and w53793;
w53795 <= not w52999 and not w53002;
w53796 <= not w53794 and not w53795;
w53797 <= not w53297 and not w53796;
w53798 <= not w52974 and not w53296;
w53799 <= not w53295 and w53798;
w53800 <= not w53797 and not w53799;
w53801 <= not b(4) and not w53800;
w53802 <= not w52993 and w52997;
w53803 <= not w52992 and w53802;
w53804 <= not w52994 and not w52997;
w53805 <= not w53803 and not w53804;
w53806 <= not w53297 and not w53805;
w53807 <= not w52982 and not w53296;
w53808 <= not w53295 and w53807;
w53809 <= not w53806 and not w53808;
w53810 <= not b(3) and not w53809;
w53811 <= w24976 and not w52990;
w53812 <= not w52988 and w53811;
w53813 <= not w52992 and not w53812;
w53814 <= not w53297 and w53813;
w53815 <= not w52987 and not w53296;
w53816 <= not w53295 and w53815;
w53817 <= not w53814 and not w53816;
w53818 <= not b(2) and not w53817;
w53819 <= b(0) and not w53297;
w53820 <= a(4) and not w53819;
w53821 <= w24976 and not w53297;
w53822 <= not w53820 and not w53821;
w53823 <= b(1) and not w53822;
w53824 <= not b(1) and not w53821;
w53825 <= not w53820 and w53824;
w53826 <= not w53823 and not w53825;
w53827 <= not w25812 and not w53826;
w53828 <= not b(1) and not w53822;
w53829 <= not w53827 and not w53828;
w53830 <= b(2) and not w53816;
w53831 <= not w53814 and w53830;
w53832 <= not w53818 and not w53831;
w53833 <= not w53829 and w53832;
w53834 <= not w53818 and not w53833;
w53835 <= b(3) and not w53808;
w53836 <= not w53806 and w53835;
w53837 <= not w53810 and not w53836;
w53838 <= not w53834 and w53837;
w53839 <= not w53810 and not w53838;
w53840 <= b(4) and not w53799;
w53841 <= not w53797 and w53840;
w53842 <= not w53801 and not w53841;
w53843 <= not w53839 and w53842;
w53844 <= not w53801 and not w53843;
w53845 <= b(5) and not w53790;
w53846 <= not w53788 and w53845;
w53847 <= not w53792 and not w53846;
w53848 <= not w53844 and w53847;
w53849 <= not w53792 and not w53848;
w53850 <= b(6) and not w53781;
w53851 <= not w53779 and w53850;
w53852 <= not w53783 and not w53851;
w53853 <= not w53849 and w53852;
w53854 <= not w53783 and not w53853;
w53855 <= b(7) and not w53772;
w53856 <= not w53770 and w53855;
w53857 <= not w53774 and not w53856;
w53858 <= not w53854 and w53857;
w53859 <= not w53774 and not w53858;
w53860 <= b(8) and not w53763;
w53861 <= not w53761 and w53860;
w53862 <= not w53765 and not w53861;
w53863 <= not w53859 and w53862;
w53864 <= not w53765 and not w53863;
w53865 <= b(9) and not w53754;
w53866 <= not w53752 and w53865;
w53867 <= not w53756 and not w53866;
w53868 <= not w53864 and w53867;
w53869 <= not w53756 and not w53868;
w53870 <= b(10) and not w53745;
w53871 <= not w53743 and w53870;
w53872 <= not w53747 and not w53871;
w53873 <= not w53869 and w53872;
w53874 <= not w53747 and not w53873;
w53875 <= b(11) and not w53736;
w53876 <= not w53734 and w53875;
w53877 <= not w53738 and not w53876;
w53878 <= not w53874 and w53877;
w53879 <= not w53738 and not w53878;
w53880 <= b(12) and not w53727;
w53881 <= not w53725 and w53880;
w53882 <= not w53729 and not w53881;
w53883 <= not w53879 and w53882;
w53884 <= not w53729 and not w53883;
w53885 <= b(13) and not w53718;
w53886 <= not w53716 and w53885;
w53887 <= not w53720 and not w53886;
w53888 <= not w53884 and w53887;
w53889 <= not w53720 and not w53888;
w53890 <= b(14) and not w53709;
w53891 <= not w53707 and w53890;
w53892 <= not w53711 and not w53891;
w53893 <= not w53889 and w53892;
w53894 <= not w53711 and not w53893;
w53895 <= b(15) and not w53700;
w53896 <= not w53698 and w53895;
w53897 <= not w53702 and not w53896;
w53898 <= not w53894 and w53897;
w53899 <= not w53702 and not w53898;
w53900 <= b(16) and not w53691;
w53901 <= not w53689 and w53900;
w53902 <= not w53693 and not w53901;
w53903 <= not w53899 and w53902;
w53904 <= not w53693 and not w53903;
w53905 <= b(17) and not w53682;
w53906 <= not w53680 and w53905;
w53907 <= not w53684 and not w53906;
w53908 <= not w53904 and w53907;
w53909 <= not w53684 and not w53908;
w53910 <= b(18) and not w53673;
w53911 <= not w53671 and w53910;
w53912 <= not w53675 and not w53911;
w53913 <= not w53909 and w53912;
w53914 <= not w53675 and not w53913;
w53915 <= b(19) and not w53664;
w53916 <= not w53662 and w53915;
w53917 <= not w53666 and not w53916;
w53918 <= not w53914 and w53917;
w53919 <= not w53666 and not w53918;
w53920 <= b(20) and not w53655;
w53921 <= not w53653 and w53920;
w53922 <= not w53657 and not w53921;
w53923 <= not w53919 and w53922;
w53924 <= not w53657 and not w53923;
w53925 <= b(21) and not w53646;
w53926 <= not w53644 and w53925;
w53927 <= not w53648 and not w53926;
w53928 <= not w53924 and w53927;
w53929 <= not w53648 and not w53928;
w53930 <= b(22) and not w53637;
w53931 <= not w53635 and w53930;
w53932 <= not w53639 and not w53931;
w53933 <= not w53929 and w53932;
w53934 <= not w53639 and not w53933;
w53935 <= b(23) and not w53628;
w53936 <= not w53626 and w53935;
w53937 <= not w53630 and not w53936;
w53938 <= not w53934 and w53937;
w53939 <= not w53630 and not w53938;
w53940 <= b(24) and not w53619;
w53941 <= not w53617 and w53940;
w53942 <= not w53621 and not w53941;
w53943 <= not w53939 and w53942;
w53944 <= not w53621 and not w53943;
w53945 <= b(25) and not w53610;
w53946 <= not w53608 and w53945;
w53947 <= not w53612 and not w53946;
w53948 <= not w53944 and w53947;
w53949 <= not w53612 and not w53948;
w53950 <= b(26) and not w53601;
w53951 <= not w53599 and w53950;
w53952 <= not w53603 and not w53951;
w53953 <= not w53949 and w53952;
w53954 <= not w53603 and not w53953;
w53955 <= b(27) and not w53592;
w53956 <= not w53590 and w53955;
w53957 <= not w53594 and not w53956;
w53958 <= not w53954 and w53957;
w53959 <= not w53594 and not w53958;
w53960 <= b(28) and not w53583;
w53961 <= not w53581 and w53960;
w53962 <= not w53585 and not w53961;
w53963 <= not w53959 and w53962;
w53964 <= not w53585 and not w53963;
w53965 <= b(29) and not w53574;
w53966 <= not w53572 and w53965;
w53967 <= not w53576 and not w53966;
w53968 <= not w53964 and w53967;
w53969 <= not w53576 and not w53968;
w53970 <= b(30) and not w53565;
w53971 <= not w53563 and w53970;
w53972 <= not w53567 and not w53971;
w53973 <= not w53969 and w53972;
w53974 <= not w53567 and not w53973;
w53975 <= b(31) and not w53556;
w53976 <= not w53554 and w53975;
w53977 <= not w53558 and not w53976;
w53978 <= not w53974 and w53977;
w53979 <= not w53558 and not w53978;
w53980 <= b(32) and not w53547;
w53981 <= not w53545 and w53980;
w53982 <= not w53549 and not w53981;
w53983 <= not w53979 and w53982;
w53984 <= not w53549 and not w53983;
w53985 <= b(33) and not w53538;
w53986 <= not w53536 and w53985;
w53987 <= not w53540 and not w53986;
w53988 <= not w53984 and w53987;
w53989 <= not w53540 and not w53988;
w53990 <= b(34) and not w53529;
w53991 <= not w53527 and w53990;
w53992 <= not w53531 and not w53991;
w53993 <= not w53989 and w53992;
w53994 <= not w53531 and not w53993;
w53995 <= b(35) and not w53520;
w53996 <= not w53518 and w53995;
w53997 <= not w53522 and not w53996;
w53998 <= not w53994 and w53997;
w53999 <= not w53522 and not w53998;
w54000 <= b(36) and not w53511;
w54001 <= not w53509 and w54000;
w54002 <= not w53513 and not w54001;
w54003 <= not w53999 and w54002;
w54004 <= not w53513 and not w54003;
w54005 <= b(37) and not w53502;
w54006 <= not w53500 and w54005;
w54007 <= not w53504 and not w54006;
w54008 <= not w54004 and w54007;
w54009 <= not w53504 and not w54008;
w54010 <= b(38) and not w53493;
w54011 <= not w53491 and w54010;
w54012 <= not w53495 and not w54011;
w54013 <= not w54009 and w54012;
w54014 <= not w53495 and not w54013;
w54015 <= b(39) and not w53484;
w54016 <= not w53482 and w54015;
w54017 <= not w53486 and not w54016;
w54018 <= not w54014 and w54017;
w54019 <= not w53486 and not w54018;
w54020 <= b(40) and not w53475;
w54021 <= not w53473 and w54020;
w54022 <= not w53477 and not w54021;
w54023 <= not w54019 and w54022;
w54024 <= not w53477 and not w54023;
w54025 <= b(41) and not w53466;
w54026 <= not w53464 and w54025;
w54027 <= not w53468 and not w54026;
w54028 <= not w54024 and w54027;
w54029 <= not w53468 and not w54028;
w54030 <= b(42) and not w53457;
w54031 <= not w53455 and w54030;
w54032 <= not w53459 and not w54031;
w54033 <= not w54029 and w54032;
w54034 <= not w53459 and not w54033;
w54035 <= b(43) and not w53448;
w54036 <= not w53446 and w54035;
w54037 <= not w53450 and not w54036;
w54038 <= not w54034 and w54037;
w54039 <= not w53450 and not w54038;
w54040 <= b(44) and not w53439;
w54041 <= not w53437 and w54040;
w54042 <= not w53441 and not w54041;
w54043 <= not w54039 and w54042;
w54044 <= not w53441 and not w54043;
w54045 <= b(45) and not w53430;
w54046 <= not w53428 and w54045;
w54047 <= not w53432 and not w54046;
w54048 <= not w54044 and w54047;
w54049 <= not w53432 and not w54048;
w54050 <= b(46) and not w53421;
w54051 <= not w53419 and w54050;
w54052 <= not w53423 and not w54051;
w54053 <= not w54049 and w54052;
w54054 <= not w53423 and not w54053;
w54055 <= b(47) and not w53412;
w54056 <= not w53410 and w54055;
w54057 <= not w53414 and not w54056;
w54058 <= not w54054 and w54057;
w54059 <= not w53414 and not w54058;
w54060 <= b(48) and not w53403;
w54061 <= not w53401 and w54060;
w54062 <= not w53405 and not w54061;
w54063 <= not w54059 and w54062;
w54064 <= not w53405 and not w54063;
w54065 <= b(49) and not w53394;
w54066 <= not w53392 and w54065;
w54067 <= not w53396 and not w54066;
w54068 <= not w54064 and w54067;
w54069 <= not w53396 and not w54068;
w54070 <= b(50) and not w53385;
w54071 <= not w53383 and w54070;
w54072 <= not w53387 and not w54071;
w54073 <= not w54069 and w54072;
w54074 <= not w53387 and not w54073;
w54075 <= b(51) and not w53376;
w54076 <= not w53374 and w54075;
w54077 <= not w53378 and not w54076;
w54078 <= not w54074 and w54077;
w54079 <= not w53378 and not w54078;
w54080 <= b(52) and not w53367;
w54081 <= not w53365 and w54080;
w54082 <= not w53369 and not w54081;
w54083 <= not w54079 and w54082;
w54084 <= not w53369 and not w54083;
w54085 <= b(53) and not w53358;
w54086 <= not w53356 and w54085;
w54087 <= not w53360 and not w54086;
w54088 <= not w54084 and w54087;
w54089 <= not w53360 and not w54088;
w54090 <= b(54) and not w53349;
w54091 <= not w53347 and w54090;
w54092 <= not w53351 and not w54091;
w54093 <= not w54089 and w54092;
w54094 <= not w53351 and not w54093;
w54095 <= b(55) and not w53340;
w54096 <= not w53338 and w54095;
w54097 <= not w53342 and not w54096;
w54098 <= not w54094 and w54097;
w54099 <= not w53342 and not w54098;
w54100 <= b(56) and not w53331;
w54101 <= not w53329 and w54100;
w54102 <= not w53333 and not w54101;
w54103 <= not w54099 and w54102;
w54104 <= not w53333 and not w54103;
w54105 <= b(57) and not w53322;
w54106 <= not w53320 and w54105;
w54107 <= not w53324 and not w54106;
w54108 <= not w54104 and w54107;
w54109 <= not w53324 and not w54108;
w54110 <= b(58) and not w53313;
w54111 <= not w53311 and w54110;
w54112 <= not w53315 and not w54111;
w54113 <= not w54109 and w54112;
w54114 <= not w53315 and not w54113;
w54115 <= b(59) and not w53304;
w54116 <= not w53302 and w54115;
w54117 <= not w53306 and not w54116;
w54118 <= not w54114 and w54117;
w54119 <= not w53306 and not w54118;
w54120 <= not w52480 and not w53292;
w54121 <= not w53290 and w54120;
w54122 <= not w53278 and w54121;
w54123 <= not w53290 and not w53292;
w54124 <= not w53279 and not w54123;
w54125 <= not w54122 and not w54124;
w54126 <= not w53297 and not w54125;
w54127 <= not w53289 and not w53296;
w54128 <= not w53295 and w54127;
w54129 <= not w54126 and not w54128;
w54130 <= not b(60) and not w54129;
w54131 <= b(60) and not w54128;
w54132 <= not w54126 and w54131;
w54133 <= w146 and not w54132;
w54134 <= not w54130 and w54133;
w54135 <= not w54119 and w54134;
w54136 <= w23 and not w54129;
w54137 <= not w54135 and not w54136;
w54138 <= not w53315 and w54117;
w54139 <= not w54113 and w54138;
w54140 <= not w54114 and not w54117;
w54141 <= not w54139 and not w54140;
w54142 <= not w54137 and not w54141;
w54143 <= not w53305 and not w54136;
w54144 <= not w54135 and w54143;
w54145 <= not w54142 and not w54144;
w54146 <= not b(60) and not w54145;
w54147 <= not w53324 and w54112;
w54148 <= not w54108 and w54147;
w54149 <= not w54109 and not w54112;
w54150 <= not w54148 and not w54149;
w54151 <= not w54137 and not w54150;
w54152 <= not w53314 and not w54136;
w54153 <= not w54135 and w54152;
w54154 <= not w54151 and not w54153;
w54155 <= not b(59) and not w54154;
w54156 <= not w53333 and w54107;
w54157 <= not w54103 and w54156;
w54158 <= not w54104 and not w54107;
w54159 <= not w54157 and not w54158;
w54160 <= not w54137 and not w54159;
w54161 <= not w53323 and not w54136;
w54162 <= not w54135 and w54161;
w54163 <= not w54160 and not w54162;
w54164 <= not b(58) and not w54163;
w54165 <= not w53342 and w54102;
w54166 <= not w54098 and w54165;
w54167 <= not w54099 and not w54102;
w54168 <= not w54166 and not w54167;
w54169 <= not w54137 and not w54168;
w54170 <= not w53332 and not w54136;
w54171 <= not w54135 and w54170;
w54172 <= not w54169 and not w54171;
w54173 <= not b(57) and not w54172;
w54174 <= not w53351 and w54097;
w54175 <= not w54093 and w54174;
w54176 <= not w54094 and not w54097;
w54177 <= not w54175 and not w54176;
w54178 <= not w54137 and not w54177;
w54179 <= not w53341 and not w54136;
w54180 <= not w54135 and w54179;
w54181 <= not w54178 and not w54180;
w54182 <= not b(56) and not w54181;
w54183 <= not w53360 and w54092;
w54184 <= not w54088 and w54183;
w54185 <= not w54089 and not w54092;
w54186 <= not w54184 and not w54185;
w54187 <= not w54137 and not w54186;
w54188 <= not w53350 and not w54136;
w54189 <= not w54135 and w54188;
w54190 <= not w54187 and not w54189;
w54191 <= not b(55) and not w54190;
w54192 <= not w53369 and w54087;
w54193 <= not w54083 and w54192;
w54194 <= not w54084 and not w54087;
w54195 <= not w54193 and not w54194;
w54196 <= not w54137 and not w54195;
w54197 <= not w53359 and not w54136;
w54198 <= not w54135 and w54197;
w54199 <= not w54196 and not w54198;
w54200 <= not b(54) and not w54199;
w54201 <= not w53378 and w54082;
w54202 <= not w54078 and w54201;
w54203 <= not w54079 and not w54082;
w54204 <= not w54202 and not w54203;
w54205 <= not w54137 and not w54204;
w54206 <= not w53368 and not w54136;
w54207 <= not w54135 and w54206;
w54208 <= not w54205 and not w54207;
w54209 <= not b(53) and not w54208;
w54210 <= not w53387 and w54077;
w54211 <= not w54073 and w54210;
w54212 <= not w54074 and not w54077;
w54213 <= not w54211 and not w54212;
w54214 <= not w54137 and not w54213;
w54215 <= not w53377 and not w54136;
w54216 <= not w54135 and w54215;
w54217 <= not w54214 and not w54216;
w54218 <= not b(52) and not w54217;
w54219 <= not w53396 and w54072;
w54220 <= not w54068 and w54219;
w54221 <= not w54069 and not w54072;
w54222 <= not w54220 and not w54221;
w54223 <= not w54137 and not w54222;
w54224 <= not w53386 and not w54136;
w54225 <= not w54135 and w54224;
w54226 <= not w54223 and not w54225;
w54227 <= not b(51) and not w54226;
w54228 <= not w53405 and w54067;
w54229 <= not w54063 and w54228;
w54230 <= not w54064 and not w54067;
w54231 <= not w54229 and not w54230;
w54232 <= not w54137 and not w54231;
w54233 <= not w53395 and not w54136;
w54234 <= not w54135 and w54233;
w54235 <= not w54232 and not w54234;
w54236 <= not b(50) and not w54235;
w54237 <= not w53414 and w54062;
w54238 <= not w54058 and w54237;
w54239 <= not w54059 and not w54062;
w54240 <= not w54238 and not w54239;
w54241 <= not w54137 and not w54240;
w54242 <= not w53404 and not w54136;
w54243 <= not w54135 and w54242;
w54244 <= not w54241 and not w54243;
w54245 <= not b(49) and not w54244;
w54246 <= not w53423 and w54057;
w54247 <= not w54053 and w54246;
w54248 <= not w54054 and not w54057;
w54249 <= not w54247 and not w54248;
w54250 <= not w54137 and not w54249;
w54251 <= not w53413 and not w54136;
w54252 <= not w54135 and w54251;
w54253 <= not w54250 and not w54252;
w54254 <= not b(48) and not w54253;
w54255 <= not w53432 and w54052;
w54256 <= not w54048 and w54255;
w54257 <= not w54049 and not w54052;
w54258 <= not w54256 and not w54257;
w54259 <= not w54137 and not w54258;
w54260 <= not w53422 and not w54136;
w54261 <= not w54135 and w54260;
w54262 <= not w54259 and not w54261;
w54263 <= not b(47) and not w54262;
w54264 <= not w53441 and w54047;
w54265 <= not w54043 and w54264;
w54266 <= not w54044 and not w54047;
w54267 <= not w54265 and not w54266;
w54268 <= not w54137 and not w54267;
w54269 <= not w53431 and not w54136;
w54270 <= not w54135 and w54269;
w54271 <= not w54268 and not w54270;
w54272 <= not b(46) and not w54271;
w54273 <= not w53450 and w54042;
w54274 <= not w54038 and w54273;
w54275 <= not w54039 and not w54042;
w54276 <= not w54274 and not w54275;
w54277 <= not w54137 and not w54276;
w54278 <= not w53440 and not w54136;
w54279 <= not w54135 and w54278;
w54280 <= not w54277 and not w54279;
w54281 <= not b(45) and not w54280;
w54282 <= not w53459 and w54037;
w54283 <= not w54033 and w54282;
w54284 <= not w54034 and not w54037;
w54285 <= not w54283 and not w54284;
w54286 <= not w54137 and not w54285;
w54287 <= not w53449 and not w54136;
w54288 <= not w54135 and w54287;
w54289 <= not w54286 and not w54288;
w54290 <= not b(44) and not w54289;
w54291 <= not w53468 and w54032;
w54292 <= not w54028 and w54291;
w54293 <= not w54029 and not w54032;
w54294 <= not w54292 and not w54293;
w54295 <= not w54137 and not w54294;
w54296 <= not w53458 and not w54136;
w54297 <= not w54135 and w54296;
w54298 <= not w54295 and not w54297;
w54299 <= not b(43) and not w54298;
w54300 <= not w53477 and w54027;
w54301 <= not w54023 and w54300;
w54302 <= not w54024 and not w54027;
w54303 <= not w54301 and not w54302;
w54304 <= not w54137 and not w54303;
w54305 <= not w53467 and not w54136;
w54306 <= not w54135 and w54305;
w54307 <= not w54304 and not w54306;
w54308 <= not b(42) and not w54307;
w54309 <= not w53486 and w54022;
w54310 <= not w54018 and w54309;
w54311 <= not w54019 and not w54022;
w54312 <= not w54310 and not w54311;
w54313 <= not w54137 and not w54312;
w54314 <= not w53476 and not w54136;
w54315 <= not w54135 and w54314;
w54316 <= not w54313 and not w54315;
w54317 <= not b(41) and not w54316;
w54318 <= not w53495 and w54017;
w54319 <= not w54013 and w54318;
w54320 <= not w54014 and not w54017;
w54321 <= not w54319 and not w54320;
w54322 <= not w54137 and not w54321;
w54323 <= not w53485 and not w54136;
w54324 <= not w54135 and w54323;
w54325 <= not w54322 and not w54324;
w54326 <= not b(40) and not w54325;
w54327 <= not w53504 and w54012;
w54328 <= not w54008 and w54327;
w54329 <= not w54009 and not w54012;
w54330 <= not w54328 and not w54329;
w54331 <= not w54137 and not w54330;
w54332 <= not w53494 and not w54136;
w54333 <= not w54135 and w54332;
w54334 <= not w54331 and not w54333;
w54335 <= not b(39) and not w54334;
w54336 <= not w53513 and w54007;
w54337 <= not w54003 and w54336;
w54338 <= not w54004 and not w54007;
w54339 <= not w54337 and not w54338;
w54340 <= not w54137 and not w54339;
w54341 <= not w53503 and not w54136;
w54342 <= not w54135 and w54341;
w54343 <= not w54340 and not w54342;
w54344 <= not b(38) and not w54343;
w54345 <= not w53522 and w54002;
w54346 <= not w53998 and w54345;
w54347 <= not w53999 and not w54002;
w54348 <= not w54346 and not w54347;
w54349 <= not w54137 and not w54348;
w54350 <= not w53512 and not w54136;
w54351 <= not w54135 and w54350;
w54352 <= not w54349 and not w54351;
w54353 <= not b(37) and not w54352;
w54354 <= not w53531 and w53997;
w54355 <= not w53993 and w54354;
w54356 <= not w53994 and not w53997;
w54357 <= not w54355 and not w54356;
w54358 <= not w54137 and not w54357;
w54359 <= not w53521 and not w54136;
w54360 <= not w54135 and w54359;
w54361 <= not w54358 and not w54360;
w54362 <= not b(36) and not w54361;
w54363 <= not w53540 and w53992;
w54364 <= not w53988 and w54363;
w54365 <= not w53989 and not w53992;
w54366 <= not w54364 and not w54365;
w54367 <= not w54137 and not w54366;
w54368 <= not w53530 and not w54136;
w54369 <= not w54135 and w54368;
w54370 <= not w54367 and not w54369;
w54371 <= not b(35) and not w54370;
w54372 <= not w53549 and w53987;
w54373 <= not w53983 and w54372;
w54374 <= not w53984 and not w53987;
w54375 <= not w54373 and not w54374;
w54376 <= not w54137 and not w54375;
w54377 <= not w53539 and not w54136;
w54378 <= not w54135 and w54377;
w54379 <= not w54376 and not w54378;
w54380 <= not b(34) and not w54379;
w54381 <= not w53558 and w53982;
w54382 <= not w53978 and w54381;
w54383 <= not w53979 and not w53982;
w54384 <= not w54382 and not w54383;
w54385 <= not w54137 and not w54384;
w54386 <= not w53548 and not w54136;
w54387 <= not w54135 and w54386;
w54388 <= not w54385 and not w54387;
w54389 <= not b(33) and not w54388;
w54390 <= not w53567 and w53977;
w54391 <= not w53973 and w54390;
w54392 <= not w53974 and not w53977;
w54393 <= not w54391 and not w54392;
w54394 <= not w54137 and not w54393;
w54395 <= not w53557 and not w54136;
w54396 <= not w54135 and w54395;
w54397 <= not w54394 and not w54396;
w54398 <= not b(32) and not w54397;
w54399 <= not w53576 and w53972;
w54400 <= not w53968 and w54399;
w54401 <= not w53969 and not w53972;
w54402 <= not w54400 and not w54401;
w54403 <= not w54137 and not w54402;
w54404 <= not w53566 and not w54136;
w54405 <= not w54135 and w54404;
w54406 <= not w54403 and not w54405;
w54407 <= not b(31) and not w54406;
w54408 <= not w53585 and w53967;
w54409 <= not w53963 and w54408;
w54410 <= not w53964 and not w53967;
w54411 <= not w54409 and not w54410;
w54412 <= not w54137 and not w54411;
w54413 <= not w53575 and not w54136;
w54414 <= not w54135 and w54413;
w54415 <= not w54412 and not w54414;
w54416 <= not b(30) and not w54415;
w54417 <= not w53594 and w53962;
w54418 <= not w53958 and w54417;
w54419 <= not w53959 and not w53962;
w54420 <= not w54418 and not w54419;
w54421 <= not w54137 and not w54420;
w54422 <= not w53584 and not w54136;
w54423 <= not w54135 and w54422;
w54424 <= not w54421 and not w54423;
w54425 <= not b(29) and not w54424;
w54426 <= not w53603 and w53957;
w54427 <= not w53953 and w54426;
w54428 <= not w53954 and not w53957;
w54429 <= not w54427 and not w54428;
w54430 <= not w54137 and not w54429;
w54431 <= not w53593 and not w54136;
w54432 <= not w54135 and w54431;
w54433 <= not w54430 and not w54432;
w54434 <= not b(28) and not w54433;
w54435 <= not w53612 and w53952;
w54436 <= not w53948 and w54435;
w54437 <= not w53949 and not w53952;
w54438 <= not w54436 and not w54437;
w54439 <= not w54137 and not w54438;
w54440 <= not w53602 and not w54136;
w54441 <= not w54135 and w54440;
w54442 <= not w54439 and not w54441;
w54443 <= not b(27) and not w54442;
w54444 <= not w53621 and w53947;
w54445 <= not w53943 and w54444;
w54446 <= not w53944 and not w53947;
w54447 <= not w54445 and not w54446;
w54448 <= not w54137 and not w54447;
w54449 <= not w53611 and not w54136;
w54450 <= not w54135 and w54449;
w54451 <= not w54448 and not w54450;
w54452 <= not b(26) and not w54451;
w54453 <= not w53630 and w53942;
w54454 <= not w53938 and w54453;
w54455 <= not w53939 and not w53942;
w54456 <= not w54454 and not w54455;
w54457 <= not w54137 and not w54456;
w54458 <= not w53620 and not w54136;
w54459 <= not w54135 and w54458;
w54460 <= not w54457 and not w54459;
w54461 <= not b(25) and not w54460;
w54462 <= not w53639 and w53937;
w54463 <= not w53933 and w54462;
w54464 <= not w53934 and not w53937;
w54465 <= not w54463 and not w54464;
w54466 <= not w54137 and not w54465;
w54467 <= not w53629 and not w54136;
w54468 <= not w54135 and w54467;
w54469 <= not w54466 and not w54468;
w54470 <= not b(24) and not w54469;
w54471 <= not w53648 and w53932;
w54472 <= not w53928 and w54471;
w54473 <= not w53929 and not w53932;
w54474 <= not w54472 and not w54473;
w54475 <= not w54137 and not w54474;
w54476 <= not w53638 and not w54136;
w54477 <= not w54135 and w54476;
w54478 <= not w54475 and not w54477;
w54479 <= not b(23) and not w54478;
w54480 <= not w53657 and w53927;
w54481 <= not w53923 and w54480;
w54482 <= not w53924 and not w53927;
w54483 <= not w54481 and not w54482;
w54484 <= not w54137 and not w54483;
w54485 <= not w53647 and not w54136;
w54486 <= not w54135 and w54485;
w54487 <= not w54484 and not w54486;
w54488 <= not b(22) and not w54487;
w54489 <= not w53666 and w53922;
w54490 <= not w53918 and w54489;
w54491 <= not w53919 and not w53922;
w54492 <= not w54490 and not w54491;
w54493 <= not w54137 and not w54492;
w54494 <= not w53656 and not w54136;
w54495 <= not w54135 and w54494;
w54496 <= not w54493 and not w54495;
w54497 <= not b(21) and not w54496;
w54498 <= not w53675 and w53917;
w54499 <= not w53913 and w54498;
w54500 <= not w53914 and not w53917;
w54501 <= not w54499 and not w54500;
w54502 <= not w54137 and not w54501;
w54503 <= not w53665 and not w54136;
w54504 <= not w54135 and w54503;
w54505 <= not w54502 and not w54504;
w54506 <= not b(20) and not w54505;
w54507 <= not w53684 and w53912;
w54508 <= not w53908 and w54507;
w54509 <= not w53909 and not w53912;
w54510 <= not w54508 and not w54509;
w54511 <= not w54137 and not w54510;
w54512 <= not w53674 and not w54136;
w54513 <= not w54135 and w54512;
w54514 <= not w54511 and not w54513;
w54515 <= not b(19) and not w54514;
w54516 <= not w53693 and w53907;
w54517 <= not w53903 and w54516;
w54518 <= not w53904 and not w53907;
w54519 <= not w54517 and not w54518;
w54520 <= not w54137 and not w54519;
w54521 <= not w53683 and not w54136;
w54522 <= not w54135 and w54521;
w54523 <= not w54520 and not w54522;
w54524 <= not b(18) and not w54523;
w54525 <= not w53702 and w53902;
w54526 <= not w53898 and w54525;
w54527 <= not w53899 and not w53902;
w54528 <= not w54526 and not w54527;
w54529 <= not w54137 and not w54528;
w54530 <= not w53692 and not w54136;
w54531 <= not w54135 and w54530;
w54532 <= not w54529 and not w54531;
w54533 <= not b(17) and not w54532;
w54534 <= not w53711 and w53897;
w54535 <= not w53893 and w54534;
w54536 <= not w53894 and not w53897;
w54537 <= not w54535 and not w54536;
w54538 <= not w54137 and not w54537;
w54539 <= not w53701 and not w54136;
w54540 <= not w54135 and w54539;
w54541 <= not w54538 and not w54540;
w54542 <= not b(16) and not w54541;
w54543 <= not w53720 and w53892;
w54544 <= not w53888 and w54543;
w54545 <= not w53889 and not w53892;
w54546 <= not w54544 and not w54545;
w54547 <= not w54137 and not w54546;
w54548 <= not w53710 and not w54136;
w54549 <= not w54135 and w54548;
w54550 <= not w54547 and not w54549;
w54551 <= not b(15) and not w54550;
w54552 <= not w53729 and w53887;
w54553 <= not w53883 and w54552;
w54554 <= not w53884 and not w53887;
w54555 <= not w54553 and not w54554;
w54556 <= not w54137 and not w54555;
w54557 <= not w53719 and not w54136;
w54558 <= not w54135 and w54557;
w54559 <= not w54556 and not w54558;
w54560 <= not b(14) and not w54559;
w54561 <= not w53738 and w53882;
w54562 <= not w53878 and w54561;
w54563 <= not w53879 and not w53882;
w54564 <= not w54562 and not w54563;
w54565 <= not w54137 and not w54564;
w54566 <= not w53728 and not w54136;
w54567 <= not w54135 and w54566;
w54568 <= not w54565 and not w54567;
w54569 <= not b(13) and not w54568;
w54570 <= not w53747 and w53877;
w54571 <= not w53873 and w54570;
w54572 <= not w53874 and not w53877;
w54573 <= not w54571 and not w54572;
w54574 <= not w54137 and not w54573;
w54575 <= not w53737 and not w54136;
w54576 <= not w54135 and w54575;
w54577 <= not w54574 and not w54576;
w54578 <= not b(12) and not w54577;
w54579 <= not w53756 and w53872;
w54580 <= not w53868 and w54579;
w54581 <= not w53869 and not w53872;
w54582 <= not w54580 and not w54581;
w54583 <= not w54137 and not w54582;
w54584 <= not w53746 and not w54136;
w54585 <= not w54135 and w54584;
w54586 <= not w54583 and not w54585;
w54587 <= not b(11) and not w54586;
w54588 <= not w53765 and w53867;
w54589 <= not w53863 and w54588;
w54590 <= not w53864 and not w53867;
w54591 <= not w54589 and not w54590;
w54592 <= not w54137 and not w54591;
w54593 <= not w53755 and not w54136;
w54594 <= not w54135 and w54593;
w54595 <= not w54592 and not w54594;
w54596 <= not b(10) and not w54595;
w54597 <= not w53774 and w53862;
w54598 <= not w53858 and w54597;
w54599 <= not w53859 and not w53862;
w54600 <= not w54598 and not w54599;
w54601 <= not w54137 and not w54600;
w54602 <= not w53764 and not w54136;
w54603 <= not w54135 and w54602;
w54604 <= not w54601 and not w54603;
w54605 <= not b(9) and not w54604;
w54606 <= not w53783 and w53857;
w54607 <= not w53853 and w54606;
w54608 <= not w53854 and not w53857;
w54609 <= not w54607 and not w54608;
w54610 <= not w54137 and not w54609;
w54611 <= not w53773 and not w54136;
w54612 <= not w54135 and w54611;
w54613 <= not w54610 and not w54612;
w54614 <= not b(8) and not w54613;
w54615 <= not w53792 and w53852;
w54616 <= not w53848 and w54615;
w54617 <= not w53849 and not w53852;
w54618 <= not w54616 and not w54617;
w54619 <= not w54137 and not w54618;
w54620 <= not w53782 and not w54136;
w54621 <= not w54135 and w54620;
w54622 <= not w54619 and not w54621;
w54623 <= not b(7) and not w54622;
w54624 <= not w53801 and w53847;
w54625 <= not w53843 and w54624;
w54626 <= not w53844 and not w53847;
w54627 <= not w54625 and not w54626;
w54628 <= not w54137 and not w54627;
w54629 <= not w53791 and not w54136;
w54630 <= not w54135 and w54629;
w54631 <= not w54628 and not w54630;
w54632 <= not b(6) and not w54631;
w54633 <= not w53810 and w53842;
w54634 <= not w53838 and w54633;
w54635 <= not w53839 and not w53842;
w54636 <= not w54634 and not w54635;
w54637 <= not w54137 and not w54636;
w54638 <= not w53800 and not w54136;
w54639 <= not w54135 and w54638;
w54640 <= not w54637 and not w54639;
w54641 <= not b(5) and not w54640;
w54642 <= not w53818 and w53837;
w54643 <= not w53833 and w54642;
w54644 <= not w53834 and not w53837;
w54645 <= not w54643 and not w54644;
w54646 <= not w54137 and not w54645;
w54647 <= not w53809 and not w54136;
w54648 <= not w54135 and w54647;
w54649 <= not w54646 and not w54648;
w54650 <= not b(4) and not w54649;
w54651 <= not w53828 and w53832;
w54652 <= not w53827 and w54651;
w54653 <= not w53829 and not w53832;
w54654 <= not w54652 and not w54653;
w54655 <= not w54137 and not w54654;
w54656 <= not w53817 and not w54136;
w54657 <= not w54135 and w54656;
w54658 <= not w54655 and not w54657;
w54659 <= not b(3) and not w54658;
w54660 <= w25812 and not w53825;
w54661 <= not w53823 and w54660;
w54662 <= not w53827 and not w54661;
w54663 <= not w54137 and w54662;
w54664 <= not w53822 and not w54136;
w54665 <= not w54135 and w54664;
w54666 <= not w54663 and not w54665;
w54667 <= not b(2) and not w54666;
w54668 <= b(0) and not w54137;
w54669 <= a(3) and not w54668;
w54670 <= w25812 and not w54137;
w54671 <= not w54669 and not w54670;
w54672 <= b(1) and not w54671;
w54673 <= not b(1) and not w54670;
w54674 <= not w54669 and w54673;
w54675 <= not w54672 and not w54674;
w54676 <= not w26662 and not w54675;
w54677 <= not b(1) and not w54671;
w54678 <= not w54676 and not w54677;
w54679 <= b(2) and not w54665;
w54680 <= not w54663 and w54679;
w54681 <= not w54667 and not w54680;
w54682 <= not w54678 and w54681;
w54683 <= not w54667 and not w54682;
w54684 <= b(3) and not w54657;
w54685 <= not w54655 and w54684;
w54686 <= not w54659 and not w54685;
w54687 <= not w54683 and w54686;
w54688 <= not w54659 and not w54687;
w54689 <= b(4) and not w54648;
w54690 <= not w54646 and w54689;
w54691 <= not w54650 and not w54690;
w54692 <= not w54688 and w54691;
w54693 <= not w54650 and not w54692;
w54694 <= b(5) and not w54639;
w54695 <= not w54637 and w54694;
w54696 <= not w54641 and not w54695;
w54697 <= not w54693 and w54696;
w54698 <= not w54641 and not w54697;
w54699 <= b(6) and not w54630;
w54700 <= not w54628 and w54699;
w54701 <= not w54632 and not w54700;
w54702 <= not w54698 and w54701;
w54703 <= not w54632 and not w54702;
w54704 <= b(7) and not w54621;
w54705 <= not w54619 and w54704;
w54706 <= not w54623 and not w54705;
w54707 <= not w54703 and w54706;
w54708 <= not w54623 and not w54707;
w54709 <= b(8) and not w54612;
w54710 <= not w54610 and w54709;
w54711 <= not w54614 and not w54710;
w54712 <= not w54708 and w54711;
w54713 <= not w54614 and not w54712;
w54714 <= b(9) and not w54603;
w54715 <= not w54601 and w54714;
w54716 <= not w54605 and not w54715;
w54717 <= not w54713 and w54716;
w54718 <= not w54605 and not w54717;
w54719 <= b(10) and not w54594;
w54720 <= not w54592 and w54719;
w54721 <= not w54596 and not w54720;
w54722 <= not w54718 and w54721;
w54723 <= not w54596 and not w54722;
w54724 <= b(11) and not w54585;
w54725 <= not w54583 and w54724;
w54726 <= not w54587 and not w54725;
w54727 <= not w54723 and w54726;
w54728 <= not w54587 and not w54727;
w54729 <= b(12) and not w54576;
w54730 <= not w54574 and w54729;
w54731 <= not w54578 and not w54730;
w54732 <= not w54728 and w54731;
w54733 <= not w54578 and not w54732;
w54734 <= b(13) and not w54567;
w54735 <= not w54565 and w54734;
w54736 <= not w54569 and not w54735;
w54737 <= not w54733 and w54736;
w54738 <= not w54569 and not w54737;
w54739 <= b(14) and not w54558;
w54740 <= not w54556 and w54739;
w54741 <= not w54560 and not w54740;
w54742 <= not w54738 and w54741;
w54743 <= not w54560 and not w54742;
w54744 <= b(15) and not w54549;
w54745 <= not w54547 and w54744;
w54746 <= not w54551 and not w54745;
w54747 <= not w54743 and w54746;
w54748 <= not w54551 and not w54747;
w54749 <= b(16) and not w54540;
w54750 <= not w54538 and w54749;
w54751 <= not w54542 and not w54750;
w54752 <= not w54748 and w54751;
w54753 <= not w54542 and not w54752;
w54754 <= b(17) and not w54531;
w54755 <= not w54529 and w54754;
w54756 <= not w54533 and not w54755;
w54757 <= not w54753 and w54756;
w54758 <= not w54533 and not w54757;
w54759 <= b(18) and not w54522;
w54760 <= not w54520 and w54759;
w54761 <= not w54524 and not w54760;
w54762 <= not w54758 and w54761;
w54763 <= not w54524 and not w54762;
w54764 <= b(19) and not w54513;
w54765 <= not w54511 and w54764;
w54766 <= not w54515 and not w54765;
w54767 <= not w54763 and w54766;
w54768 <= not w54515 and not w54767;
w54769 <= b(20) and not w54504;
w54770 <= not w54502 and w54769;
w54771 <= not w54506 and not w54770;
w54772 <= not w54768 and w54771;
w54773 <= not w54506 and not w54772;
w54774 <= b(21) and not w54495;
w54775 <= not w54493 and w54774;
w54776 <= not w54497 and not w54775;
w54777 <= not w54773 and w54776;
w54778 <= not w54497 and not w54777;
w54779 <= b(22) and not w54486;
w54780 <= not w54484 and w54779;
w54781 <= not w54488 and not w54780;
w54782 <= not w54778 and w54781;
w54783 <= not w54488 and not w54782;
w54784 <= b(23) and not w54477;
w54785 <= not w54475 and w54784;
w54786 <= not w54479 and not w54785;
w54787 <= not w54783 and w54786;
w54788 <= not w54479 and not w54787;
w54789 <= b(24) and not w54468;
w54790 <= not w54466 and w54789;
w54791 <= not w54470 and not w54790;
w54792 <= not w54788 and w54791;
w54793 <= not w54470 and not w54792;
w54794 <= b(25) and not w54459;
w54795 <= not w54457 and w54794;
w54796 <= not w54461 and not w54795;
w54797 <= not w54793 and w54796;
w54798 <= not w54461 and not w54797;
w54799 <= b(26) and not w54450;
w54800 <= not w54448 and w54799;
w54801 <= not w54452 and not w54800;
w54802 <= not w54798 and w54801;
w54803 <= not w54452 and not w54802;
w54804 <= b(27) and not w54441;
w54805 <= not w54439 and w54804;
w54806 <= not w54443 and not w54805;
w54807 <= not w54803 and w54806;
w54808 <= not w54443 and not w54807;
w54809 <= b(28) and not w54432;
w54810 <= not w54430 and w54809;
w54811 <= not w54434 and not w54810;
w54812 <= not w54808 and w54811;
w54813 <= not w54434 and not w54812;
w54814 <= b(29) and not w54423;
w54815 <= not w54421 and w54814;
w54816 <= not w54425 and not w54815;
w54817 <= not w54813 and w54816;
w54818 <= not w54425 and not w54817;
w54819 <= b(30) and not w54414;
w54820 <= not w54412 and w54819;
w54821 <= not w54416 and not w54820;
w54822 <= not w54818 and w54821;
w54823 <= not w54416 and not w54822;
w54824 <= b(31) and not w54405;
w54825 <= not w54403 and w54824;
w54826 <= not w54407 and not w54825;
w54827 <= not w54823 and w54826;
w54828 <= not w54407 and not w54827;
w54829 <= b(32) and not w54396;
w54830 <= not w54394 and w54829;
w54831 <= not w54398 and not w54830;
w54832 <= not w54828 and w54831;
w54833 <= not w54398 and not w54832;
w54834 <= b(33) and not w54387;
w54835 <= not w54385 and w54834;
w54836 <= not w54389 and not w54835;
w54837 <= not w54833 and w54836;
w54838 <= not w54389 and not w54837;
w54839 <= b(34) and not w54378;
w54840 <= not w54376 and w54839;
w54841 <= not w54380 and not w54840;
w54842 <= not w54838 and w54841;
w54843 <= not w54380 and not w54842;
w54844 <= b(35) and not w54369;
w54845 <= not w54367 and w54844;
w54846 <= not w54371 and not w54845;
w54847 <= not w54843 and w54846;
w54848 <= not w54371 and not w54847;
w54849 <= b(36) and not w54360;
w54850 <= not w54358 and w54849;
w54851 <= not w54362 and not w54850;
w54852 <= not w54848 and w54851;
w54853 <= not w54362 and not w54852;
w54854 <= b(37) and not w54351;
w54855 <= not w54349 and w54854;
w54856 <= not w54353 and not w54855;
w54857 <= not w54853 and w54856;
w54858 <= not w54353 and not w54857;
w54859 <= b(38) and not w54342;
w54860 <= not w54340 and w54859;
w54861 <= not w54344 and not w54860;
w54862 <= not w54858 and w54861;
w54863 <= not w54344 and not w54862;
w54864 <= b(39) and not w54333;
w54865 <= not w54331 and w54864;
w54866 <= not w54335 and not w54865;
w54867 <= not w54863 and w54866;
w54868 <= not w54335 and not w54867;
w54869 <= b(40) and not w54324;
w54870 <= not w54322 and w54869;
w54871 <= not w54326 and not w54870;
w54872 <= not w54868 and w54871;
w54873 <= not w54326 and not w54872;
w54874 <= b(41) and not w54315;
w54875 <= not w54313 and w54874;
w54876 <= not w54317 and not w54875;
w54877 <= not w54873 and w54876;
w54878 <= not w54317 and not w54877;
w54879 <= b(42) and not w54306;
w54880 <= not w54304 and w54879;
w54881 <= not w54308 and not w54880;
w54882 <= not w54878 and w54881;
w54883 <= not w54308 and not w54882;
w54884 <= b(43) and not w54297;
w54885 <= not w54295 and w54884;
w54886 <= not w54299 and not w54885;
w54887 <= not w54883 and w54886;
w54888 <= not w54299 and not w54887;
w54889 <= b(44) and not w54288;
w54890 <= not w54286 and w54889;
w54891 <= not w54290 and not w54890;
w54892 <= not w54888 and w54891;
w54893 <= not w54290 and not w54892;
w54894 <= b(45) and not w54279;
w54895 <= not w54277 and w54894;
w54896 <= not w54281 and not w54895;
w54897 <= not w54893 and w54896;
w54898 <= not w54281 and not w54897;
w54899 <= b(46) and not w54270;
w54900 <= not w54268 and w54899;
w54901 <= not w54272 and not w54900;
w54902 <= not w54898 and w54901;
w54903 <= not w54272 and not w54902;
w54904 <= b(47) and not w54261;
w54905 <= not w54259 and w54904;
w54906 <= not w54263 and not w54905;
w54907 <= not w54903 and w54906;
w54908 <= not w54263 and not w54907;
w54909 <= b(48) and not w54252;
w54910 <= not w54250 and w54909;
w54911 <= not w54254 and not w54910;
w54912 <= not w54908 and w54911;
w54913 <= not w54254 and not w54912;
w54914 <= b(49) and not w54243;
w54915 <= not w54241 and w54914;
w54916 <= not w54245 and not w54915;
w54917 <= not w54913 and w54916;
w54918 <= not w54245 and not w54917;
w54919 <= b(50) and not w54234;
w54920 <= not w54232 and w54919;
w54921 <= not w54236 and not w54920;
w54922 <= not w54918 and w54921;
w54923 <= not w54236 and not w54922;
w54924 <= b(51) and not w54225;
w54925 <= not w54223 and w54924;
w54926 <= not w54227 and not w54925;
w54927 <= not w54923 and w54926;
w54928 <= not w54227 and not w54927;
w54929 <= b(52) and not w54216;
w54930 <= not w54214 and w54929;
w54931 <= not w54218 and not w54930;
w54932 <= not w54928 and w54931;
w54933 <= not w54218 and not w54932;
w54934 <= b(53) and not w54207;
w54935 <= not w54205 and w54934;
w54936 <= not w54209 and not w54935;
w54937 <= not w54933 and w54936;
w54938 <= not w54209 and not w54937;
w54939 <= b(54) and not w54198;
w54940 <= not w54196 and w54939;
w54941 <= not w54200 and not w54940;
w54942 <= not w54938 and w54941;
w54943 <= not w54200 and not w54942;
w54944 <= b(55) and not w54189;
w54945 <= not w54187 and w54944;
w54946 <= not w54191 and not w54945;
w54947 <= not w54943 and w54946;
w54948 <= not w54191 and not w54947;
w54949 <= b(56) and not w54180;
w54950 <= not w54178 and w54949;
w54951 <= not w54182 and not w54950;
w54952 <= not w54948 and w54951;
w54953 <= not w54182 and not w54952;
w54954 <= b(57) and not w54171;
w54955 <= not w54169 and w54954;
w54956 <= not w54173 and not w54955;
w54957 <= not w54953 and w54956;
w54958 <= not w54173 and not w54957;
w54959 <= b(58) and not w54162;
w54960 <= not w54160 and w54959;
w54961 <= not w54164 and not w54960;
w54962 <= not w54958 and w54961;
w54963 <= not w54164 and not w54962;
w54964 <= b(59) and not w54153;
w54965 <= not w54151 and w54964;
w54966 <= not w54155 and not w54965;
w54967 <= not w54963 and w54966;
w54968 <= not w54155 and not w54967;
w54969 <= b(60) and not w54144;
w54970 <= not w54142 and w54969;
w54971 <= not w54146 and not w54970;
w54972 <= not w54968 and w54971;
w54973 <= not w54146 and not w54972;
w54974 <= not w53306 and not w54132;
w54975 <= not w54130 and w54974;
w54976 <= not w54118 and w54975;
w54977 <= not w54130 and not w54132;
w54978 <= not w54119 and not w54977;
w54979 <= not w54976 and not w54978;
w54980 <= not w54137 and not w54979;
w54981 <= not w54129 and not w54136;
w54982 <= not w54135 and w54981;
w54983 <= not w54980 and not w54982;
w54984 <= not b(61) and not w54983;
w54985 <= b(61) and not w54982;
w54986 <= not w54980 and w54985;
w54987 <= w22 and not w54986;
w54988 <= not w54984 and w54987;
w54989 <= not w54973 and w54988;
w54990 <= w146 and not w54983;
w54991 <= not w54989 and not w54990;
w54992 <= not w54155 and w54971;
w54993 <= not w54967 and w54992;
w54994 <= not w54968 and not w54971;
w54995 <= not w54993 and not w54994;
w54996 <= not w54991 and not w54995;
w54997 <= not w54145 and not w54990;
w54998 <= not w54989 and w54997;
w54999 <= not w54996 and not w54998;
w55000 <= not b(61) and not w54999;
w55001 <= not w54164 and w54966;
w55002 <= not w54962 and w55001;
w55003 <= not w54963 and not w54966;
w55004 <= not w55002 and not w55003;
w55005 <= not w54991 and not w55004;
w55006 <= not w54154 and not w54990;
w55007 <= not w54989 and w55006;
w55008 <= not w55005 and not w55007;
w55009 <= not b(60) and not w55008;
w55010 <= not w54173 and w54961;
w55011 <= not w54957 and w55010;
w55012 <= not w54958 and not w54961;
w55013 <= not w55011 and not w55012;
w55014 <= not w54991 and not w55013;
w55015 <= not w54163 and not w54990;
w55016 <= not w54989 and w55015;
w55017 <= not w55014 and not w55016;
w55018 <= not b(59) and not w55017;
w55019 <= not w54182 and w54956;
w55020 <= not w54952 and w55019;
w55021 <= not w54953 and not w54956;
w55022 <= not w55020 and not w55021;
w55023 <= not w54991 and not w55022;
w55024 <= not w54172 and not w54990;
w55025 <= not w54989 and w55024;
w55026 <= not w55023 and not w55025;
w55027 <= not b(58) and not w55026;
w55028 <= not w54191 and w54951;
w55029 <= not w54947 and w55028;
w55030 <= not w54948 and not w54951;
w55031 <= not w55029 and not w55030;
w55032 <= not w54991 and not w55031;
w55033 <= not w54181 and not w54990;
w55034 <= not w54989 and w55033;
w55035 <= not w55032 and not w55034;
w55036 <= not b(57) and not w55035;
w55037 <= not w54200 and w54946;
w55038 <= not w54942 and w55037;
w55039 <= not w54943 and not w54946;
w55040 <= not w55038 and not w55039;
w55041 <= not w54991 and not w55040;
w55042 <= not w54190 and not w54990;
w55043 <= not w54989 and w55042;
w55044 <= not w55041 and not w55043;
w55045 <= not b(56) and not w55044;
w55046 <= not w54209 and w54941;
w55047 <= not w54937 and w55046;
w55048 <= not w54938 and not w54941;
w55049 <= not w55047 and not w55048;
w55050 <= not w54991 and not w55049;
w55051 <= not w54199 and not w54990;
w55052 <= not w54989 and w55051;
w55053 <= not w55050 and not w55052;
w55054 <= not b(55) and not w55053;
w55055 <= not w54218 and w54936;
w55056 <= not w54932 and w55055;
w55057 <= not w54933 and not w54936;
w55058 <= not w55056 and not w55057;
w55059 <= not w54991 and not w55058;
w55060 <= not w54208 and not w54990;
w55061 <= not w54989 and w55060;
w55062 <= not w55059 and not w55061;
w55063 <= not b(54) and not w55062;
w55064 <= not w54227 and w54931;
w55065 <= not w54927 and w55064;
w55066 <= not w54928 and not w54931;
w55067 <= not w55065 and not w55066;
w55068 <= not w54991 and not w55067;
w55069 <= not w54217 and not w54990;
w55070 <= not w54989 and w55069;
w55071 <= not w55068 and not w55070;
w55072 <= not b(53) and not w55071;
w55073 <= not w54236 and w54926;
w55074 <= not w54922 and w55073;
w55075 <= not w54923 and not w54926;
w55076 <= not w55074 and not w55075;
w55077 <= not w54991 and not w55076;
w55078 <= not w54226 and not w54990;
w55079 <= not w54989 and w55078;
w55080 <= not w55077 and not w55079;
w55081 <= not b(52) and not w55080;
w55082 <= not w54245 and w54921;
w55083 <= not w54917 and w55082;
w55084 <= not w54918 and not w54921;
w55085 <= not w55083 and not w55084;
w55086 <= not w54991 and not w55085;
w55087 <= not w54235 and not w54990;
w55088 <= not w54989 and w55087;
w55089 <= not w55086 and not w55088;
w55090 <= not b(51) and not w55089;
w55091 <= not w54254 and w54916;
w55092 <= not w54912 and w55091;
w55093 <= not w54913 and not w54916;
w55094 <= not w55092 and not w55093;
w55095 <= not w54991 and not w55094;
w55096 <= not w54244 and not w54990;
w55097 <= not w54989 and w55096;
w55098 <= not w55095 and not w55097;
w55099 <= not b(50) and not w55098;
w55100 <= not w54263 and w54911;
w55101 <= not w54907 and w55100;
w55102 <= not w54908 and not w54911;
w55103 <= not w55101 and not w55102;
w55104 <= not w54991 and not w55103;
w55105 <= not w54253 and not w54990;
w55106 <= not w54989 and w55105;
w55107 <= not w55104 and not w55106;
w55108 <= not b(49) and not w55107;
w55109 <= not w54272 and w54906;
w55110 <= not w54902 and w55109;
w55111 <= not w54903 and not w54906;
w55112 <= not w55110 and not w55111;
w55113 <= not w54991 and not w55112;
w55114 <= not w54262 and not w54990;
w55115 <= not w54989 and w55114;
w55116 <= not w55113 and not w55115;
w55117 <= not b(48) and not w55116;
w55118 <= not w54281 and w54901;
w55119 <= not w54897 and w55118;
w55120 <= not w54898 and not w54901;
w55121 <= not w55119 and not w55120;
w55122 <= not w54991 and not w55121;
w55123 <= not w54271 and not w54990;
w55124 <= not w54989 and w55123;
w55125 <= not w55122 and not w55124;
w55126 <= not b(47) and not w55125;
w55127 <= not w54290 and w54896;
w55128 <= not w54892 and w55127;
w55129 <= not w54893 and not w54896;
w55130 <= not w55128 and not w55129;
w55131 <= not w54991 and not w55130;
w55132 <= not w54280 and not w54990;
w55133 <= not w54989 and w55132;
w55134 <= not w55131 and not w55133;
w55135 <= not b(46) and not w55134;
w55136 <= not w54299 and w54891;
w55137 <= not w54887 and w55136;
w55138 <= not w54888 and not w54891;
w55139 <= not w55137 and not w55138;
w55140 <= not w54991 and not w55139;
w55141 <= not w54289 and not w54990;
w55142 <= not w54989 and w55141;
w55143 <= not w55140 and not w55142;
w55144 <= not b(45) and not w55143;
w55145 <= not w54308 and w54886;
w55146 <= not w54882 and w55145;
w55147 <= not w54883 and not w54886;
w55148 <= not w55146 and not w55147;
w55149 <= not w54991 and not w55148;
w55150 <= not w54298 and not w54990;
w55151 <= not w54989 and w55150;
w55152 <= not w55149 and not w55151;
w55153 <= not b(44) and not w55152;
w55154 <= not w54317 and w54881;
w55155 <= not w54877 and w55154;
w55156 <= not w54878 and not w54881;
w55157 <= not w55155 and not w55156;
w55158 <= not w54991 and not w55157;
w55159 <= not w54307 and not w54990;
w55160 <= not w54989 and w55159;
w55161 <= not w55158 and not w55160;
w55162 <= not b(43) and not w55161;
w55163 <= not w54326 and w54876;
w55164 <= not w54872 and w55163;
w55165 <= not w54873 and not w54876;
w55166 <= not w55164 and not w55165;
w55167 <= not w54991 and not w55166;
w55168 <= not w54316 and not w54990;
w55169 <= not w54989 and w55168;
w55170 <= not w55167 and not w55169;
w55171 <= not b(42) and not w55170;
w55172 <= not w54335 and w54871;
w55173 <= not w54867 and w55172;
w55174 <= not w54868 and not w54871;
w55175 <= not w55173 and not w55174;
w55176 <= not w54991 and not w55175;
w55177 <= not w54325 and not w54990;
w55178 <= not w54989 and w55177;
w55179 <= not w55176 and not w55178;
w55180 <= not b(41) and not w55179;
w55181 <= not w54344 and w54866;
w55182 <= not w54862 and w55181;
w55183 <= not w54863 and not w54866;
w55184 <= not w55182 and not w55183;
w55185 <= not w54991 and not w55184;
w55186 <= not w54334 and not w54990;
w55187 <= not w54989 and w55186;
w55188 <= not w55185 and not w55187;
w55189 <= not b(40) and not w55188;
w55190 <= not w54353 and w54861;
w55191 <= not w54857 and w55190;
w55192 <= not w54858 and not w54861;
w55193 <= not w55191 and not w55192;
w55194 <= not w54991 and not w55193;
w55195 <= not w54343 and not w54990;
w55196 <= not w54989 and w55195;
w55197 <= not w55194 and not w55196;
w55198 <= not b(39) and not w55197;
w55199 <= not w54362 and w54856;
w55200 <= not w54852 and w55199;
w55201 <= not w54853 and not w54856;
w55202 <= not w55200 and not w55201;
w55203 <= not w54991 and not w55202;
w55204 <= not w54352 and not w54990;
w55205 <= not w54989 and w55204;
w55206 <= not w55203 and not w55205;
w55207 <= not b(38) and not w55206;
w55208 <= not w54371 and w54851;
w55209 <= not w54847 and w55208;
w55210 <= not w54848 and not w54851;
w55211 <= not w55209 and not w55210;
w55212 <= not w54991 and not w55211;
w55213 <= not w54361 and not w54990;
w55214 <= not w54989 and w55213;
w55215 <= not w55212 and not w55214;
w55216 <= not b(37) and not w55215;
w55217 <= not w54380 and w54846;
w55218 <= not w54842 and w55217;
w55219 <= not w54843 and not w54846;
w55220 <= not w55218 and not w55219;
w55221 <= not w54991 and not w55220;
w55222 <= not w54370 and not w54990;
w55223 <= not w54989 and w55222;
w55224 <= not w55221 and not w55223;
w55225 <= not b(36) and not w55224;
w55226 <= not w54389 and w54841;
w55227 <= not w54837 and w55226;
w55228 <= not w54838 and not w54841;
w55229 <= not w55227 and not w55228;
w55230 <= not w54991 and not w55229;
w55231 <= not w54379 and not w54990;
w55232 <= not w54989 and w55231;
w55233 <= not w55230 and not w55232;
w55234 <= not b(35) and not w55233;
w55235 <= not w54398 and w54836;
w55236 <= not w54832 and w55235;
w55237 <= not w54833 and not w54836;
w55238 <= not w55236 and not w55237;
w55239 <= not w54991 and not w55238;
w55240 <= not w54388 and not w54990;
w55241 <= not w54989 and w55240;
w55242 <= not w55239 and not w55241;
w55243 <= not b(34) and not w55242;
w55244 <= not w54407 and w54831;
w55245 <= not w54827 and w55244;
w55246 <= not w54828 and not w54831;
w55247 <= not w55245 and not w55246;
w55248 <= not w54991 and not w55247;
w55249 <= not w54397 and not w54990;
w55250 <= not w54989 and w55249;
w55251 <= not w55248 and not w55250;
w55252 <= not b(33) and not w55251;
w55253 <= not w54416 and w54826;
w55254 <= not w54822 and w55253;
w55255 <= not w54823 and not w54826;
w55256 <= not w55254 and not w55255;
w55257 <= not w54991 and not w55256;
w55258 <= not w54406 and not w54990;
w55259 <= not w54989 and w55258;
w55260 <= not w55257 and not w55259;
w55261 <= not b(32) and not w55260;
w55262 <= not w54425 and w54821;
w55263 <= not w54817 and w55262;
w55264 <= not w54818 and not w54821;
w55265 <= not w55263 and not w55264;
w55266 <= not w54991 and not w55265;
w55267 <= not w54415 and not w54990;
w55268 <= not w54989 and w55267;
w55269 <= not w55266 and not w55268;
w55270 <= not b(31) and not w55269;
w55271 <= not w54434 and w54816;
w55272 <= not w54812 and w55271;
w55273 <= not w54813 and not w54816;
w55274 <= not w55272 and not w55273;
w55275 <= not w54991 and not w55274;
w55276 <= not w54424 and not w54990;
w55277 <= not w54989 and w55276;
w55278 <= not w55275 and not w55277;
w55279 <= not b(30) and not w55278;
w55280 <= not w54443 and w54811;
w55281 <= not w54807 and w55280;
w55282 <= not w54808 and not w54811;
w55283 <= not w55281 and not w55282;
w55284 <= not w54991 and not w55283;
w55285 <= not w54433 and not w54990;
w55286 <= not w54989 and w55285;
w55287 <= not w55284 and not w55286;
w55288 <= not b(29) and not w55287;
w55289 <= not w54452 and w54806;
w55290 <= not w54802 and w55289;
w55291 <= not w54803 and not w54806;
w55292 <= not w55290 and not w55291;
w55293 <= not w54991 and not w55292;
w55294 <= not w54442 and not w54990;
w55295 <= not w54989 and w55294;
w55296 <= not w55293 and not w55295;
w55297 <= not b(28) and not w55296;
w55298 <= not w54461 and w54801;
w55299 <= not w54797 and w55298;
w55300 <= not w54798 and not w54801;
w55301 <= not w55299 and not w55300;
w55302 <= not w54991 and not w55301;
w55303 <= not w54451 and not w54990;
w55304 <= not w54989 and w55303;
w55305 <= not w55302 and not w55304;
w55306 <= not b(27) and not w55305;
w55307 <= not w54470 and w54796;
w55308 <= not w54792 and w55307;
w55309 <= not w54793 and not w54796;
w55310 <= not w55308 and not w55309;
w55311 <= not w54991 and not w55310;
w55312 <= not w54460 and not w54990;
w55313 <= not w54989 and w55312;
w55314 <= not w55311 and not w55313;
w55315 <= not b(26) and not w55314;
w55316 <= not w54479 and w54791;
w55317 <= not w54787 and w55316;
w55318 <= not w54788 and not w54791;
w55319 <= not w55317 and not w55318;
w55320 <= not w54991 and not w55319;
w55321 <= not w54469 and not w54990;
w55322 <= not w54989 and w55321;
w55323 <= not w55320 and not w55322;
w55324 <= not b(25) and not w55323;
w55325 <= not w54488 and w54786;
w55326 <= not w54782 and w55325;
w55327 <= not w54783 and not w54786;
w55328 <= not w55326 and not w55327;
w55329 <= not w54991 and not w55328;
w55330 <= not w54478 and not w54990;
w55331 <= not w54989 and w55330;
w55332 <= not w55329 and not w55331;
w55333 <= not b(24) and not w55332;
w55334 <= not w54497 and w54781;
w55335 <= not w54777 and w55334;
w55336 <= not w54778 and not w54781;
w55337 <= not w55335 and not w55336;
w55338 <= not w54991 and not w55337;
w55339 <= not w54487 and not w54990;
w55340 <= not w54989 and w55339;
w55341 <= not w55338 and not w55340;
w55342 <= not b(23) and not w55341;
w55343 <= not w54506 and w54776;
w55344 <= not w54772 and w55343;
w55345 <= not w54773 and not w54776;
w55346 <= not w55344 and not w55345;
w55347 <= not w54991 and not w55346;
w55348 <= not w54496 and not w54990;
w55349 <= not w54989 and w55348;
w55350 <= not w55347 and not w55349;
w55351 <= not b(22) and not w55350;
w55352 <= not w54515 and w54771;
w55353 <= not w54767 and w55352;
w55354 <= not w54768 and not w54771;
w55355 <= not w55353 and not w55354;
w55356 <= not w54991 and not w55355;
w55357 <= not w54505 and not w54990;
w55358 <= not w54989 and w55357;
w55359 <= not w55356 and not w55358;
w55360 <= not b(21) and not w55359;
w55361 <= not w54524 and w54766;
w55362 <= not w54762 and w55361;
w55363 <= not w54763 and not w54766;
w55364 <= not w55362 and not w55363;
w55365 <= not w54991 and not w55364;
w55366 <= not w54514 and not w54990;
w55367 <= not w54989 and w55366;
w55368 <= not w55365 and not w55367;
w55369 <= not b(20) and not w55368;
w55370 <= not w54533 and w54761;
w55371 <= not w54757 and w55370;
w55372 <= not w54758 and not w54761;
w55373 <= not w55371 and not w55372;
w55374 <= not w54991 and not w55373;
w55375 <= not w54523 and not w54990;
w55376 <= not w54989 and w55375;
w55377 <= not w55374 and not w55376;
w55378 <= not b(19) and not w55377;
w55379 <= not w54542 and w54756;
w55380 <= not w54752 and w55379;
w55381 <= not w54753 and not w54756;
w55382 <= not w55380 and not w55381;
w55383 <= not w54991 and not w55382;
w55384 <= not w54532 and not w54990;
w55385 <= not w54989 and w55384;
w55386 <= not w55383 and not w55385;
w55387 <= not b(18) and not w55386;
w55388 <= not w54551 and w54751;
w55389 <= not w54747 and w55388;
w55390 <= not w54748 and not w54751;
w55391 <= not w55389 and not w55390;
w55392 <= not w54991 and not w55391;
w55393 <= not w54541 and not w54990;
w55394 <= not w54989 and w55393;
w55395 <= not w55392 and not w55394;
w55396 <= not b(17) and not w55395;
w55397 <= not w54560 and w54746;
w55398 <= not w54742 and w55397;
w55399 <= not w54743 and not w54746;
w55400 <= not w55398 and not w55399;
w55401 <= not w54991 and not w55400;
w55402 <= not w54550 and not w54990;
w55403 <= not w54989 and w55402;
w55404 <= not w55401 and not w55403;
w55405 <= not b(16) and not w55404;
w55406 <= not w54569 and w54741;
w55407 <= not w54737 and w55406;
w55408 <= not w54738 and not w54741;
w55409 <= not w55407 and not w55408;
w55410 <= not w54991 and not w55409;
w55411 <= not w54559 and not w54990;
w55412 <= not w54989 and w55411;
w55413 <= not w55410 and not w55412;
w55414 <= not b(15) and not w55413;
w55415 <= not w54578 and w54736;
w55416 <= not w54732 and w55415;
w55417 <= not w54733 and not w54736;
w55418 <= not w55416 and not w55417;
w55419 <= not w54991 and not w55418;
w55420 <= not w54568 and not w54990;
w55421 <= not w54989 and w55420;
w55422 <= not w55419 and not w55421;
w55423 <= not b(14) and not w55422;
w55424 <= not w54587 and w54731;
w55425 <= not w54727 and w55424;
w55426 <= not w54728 and not w54731;
w55427 <= not w55425 and not w55426;
w55428 <= not w54991 and not w55427;
w55429 <= not w54577 and not w54990;
w55430 <= not w54989 and w55429;
w55431 <= not w55428 and not w55430;
w55432 <= not b(13) and not w55431;
w55433 <= not w54596 and w54726;
w55434 <= not w54722 and w55433;
w55435 <= not w54723 and not w54726;
w55436 <= not w55434 and not w55435;
w55437 <= not w54991 and not w55436;
w55438 <= not w54586 and not w54990;
w55439 <= not w54989 and w55438;
w55440 <= not w55437 and not w55439;
w55441 <= not b(12) and not w55440;
w55442 <= not w54605 and w54721;
w55443 <= not w54717 and w55442;
w55444 <= not w54718 and not w54721;
w55445 <= not w55443 and not w55444;
w55446 <= not w54991 and not w55445;
w55447 <= not w54595 and not w54990;
w55448 <= not w54989 and w55447;
w55449 <= not w55446 and not w55448;
w55450 <= not b(11) and not w55449;
w55451 <= not w54614 and w54716;
w55452 <= not w54712 and w55451;
w55453 <= not w54713 and not w54716;
w55454 <= not w55452 and not w55453;
w55455 <= not w54991 and not w55454;
w55456 <= not w54604 and not w54990;
w55457 <= not w54989 and w55456;
w55458 <= not w55455 and not w55457;
w55459 <= not b(10) and not w55458;
w55460 <= not w54623 and w54711;
w55461 <= not w54707 and w55460;
w55462 <= not w54708 and not w54711;
w55463 <= not w55461 and not w55462;
w55464 <= not w54991 and not w55463;
w55465 <= not w54613 and not w54990;
w55466 <= not w54989 and w55465;
w55467 <= not w55464 and not w55466;
w55468 <= not b(9) and not w55467;
w55469 <= not w54632 and w54706;
w55470 <= not w54702 and w55469;
w55471 <= not w54703 and not w54706;
w55472 <= not w55470 and not w55471;
w55473 <= not w54991 and not w55472;
w55474 <= not w54622 and not w54990;
w55475 <= not w54989 and w55474;
w55476 <= not w55473 and not w55475;
w55477 <= not b(8) and not w55476;
w55478 <= not w54641 and w54701;
w55479 <= not w54697 and w55478;
w55480 <= not w54698 and not w54701;
w55481 <= not w55479 and not w55480;
w55482 <= not w54991 and not w55481;
w55483 <= not w54631 and not w54990;
w55484 <= not w54989 and w55483;
w55485 <= not w55482 and not w55484;
w55486 <= not b(7) and not w55485;
w55487 <= not w54650 and w54696;
w55488 <= not w54692 and w55487;
w55489 <= not w54693 and not w54696;
w55490 <= not w55488 and not w55489;
w55491 <= not w54991 and not w55490;
w55492 <= not w54640 and not w54990;
w55493 <= not w54989 and w55492;
w55494 <= not w55491 and not w55493;
w55495 <= not b(6) and not w55494;
w55496 <= not w54659 and w54691;
w55497 <= not w54687 and w55496;
w55498 <= not w54688 and not w54691;
w55499 <= not w55497 and not w55498;
w55500 <= not w54991 and not w55499;
w55501 <= not w54649 and not w54990;
w55502 <= not w54989 and w55501;
w55503 <= not w55500 and not w55502;
w55504 <= not b(5) and not w55503;
w55505 <= not w54667 and w54686;
w55506 <= not w54682 and w55505;
w55507 <= not w54683 and not w54686;
w55508 <= not w55506 and not w55507;
w55509 <= not w54991 and not w55508;
w55510 <= not w54658 and not w54990;
w55511 <= not w54989 and w55510;
w55512 <= not w55509 and not w55511;
w55513 <= not b(4) and not w55512;
w55514 <= not w54677 and w54681;
w55515 <= not w54676 and w55514;
w55516 <= not w54678 and not w54681;
w55517 <= not w55515 and not w55516;
w55518 <= not w54991 and not w55517;
w55519 <= not w54666 and not w54990;
w55520 <= not w54989 and w55519;
w55521 <= not w55518 and not w55520;
w55522 <= not b(3) and not w55521;
w55523 <= w26662 and not w54674;
w55524 <= not w54672 and w55523;
w55525 <= not w54676 and not w55524;
w55526 <= not w54991 and w55525;
w55527 <= not w54671 and not w54990;
w55528 <= not w54989 and w55527;
w55529 <= not w55526 and not w55528;
w55530 <= not b(2) and not w55529;
w55531 <= b(0) and not w54991;
w55532 <= a(2) and not w55531;
w55533 <= w26662 and not w54991;
w55534 <= not w55532 and not w55533;
w55535 <= b(1) and not w55534;
w55536 <= not b(1) and not w55533;
w55537 <= not w55532 and w55536;
w55538 <= not w55535 and not w55537;
w55539 <= not w27526 and not w55538;
w55540 <= not b(1) and not w55534;
w55541 <= not w55539 and not w55540;
w55542 <= b(2) and not w55528;
w55543 <= not w55526 and w55542;
w55544 <= not w55530 and not w55543;
w55545 <= not w55541 and w55544;
w55546 <= not w55530 and not w55545;
w55547 <= b(3) and not w55520;
w55548 <= not w55518 and w55547;
w55549 <= not w55522 and not w55548;
w55550 <= not w55546 and w55549;
w55551 <= not w55522 and not w55550;
w55552 <= b(4) and not w55511;
w55553 <= not w55509 and w55552;
w55554 <= not w55513 and not w55553;
w55555 <= not w55551 and w55554;
w55556 <= not w55513 and not w55555;
w55557 <= b(5) and not w55502;
w55558 <= not w55500 and w55557;
w55559 <= not w55504 and not w55558;
w55560 <= not w55556 and w55559;
w55561 <= not w55504 and not w55560;
w55562 <= b(6) and not w55493;
w55563 <= not w55491 and w55562;
w55564 <= not w55495 and not w55563;
w55565 <= not w55561 and w55564;
w55566 <= not w55495 and not w55565;
w55567 <= b(7) and not w55484;
w55568 <= not w55482 and w55567;
w55569 <= not w55486 and not w55568;
w55570 <= not w55566 and w55569;
w55571 <= not w55486 and not w55570;
w55572 <= b(8) and not w55475;
w55573 <= not w55473 and w55572;
w55574 <= not w55477 and not w55573;
w55575 <= not w55571 and w55574;
w55576 <= not w55477 and not w55575;
w55577 <= b(9) and not w55466;
w55578 <= not w55464 and w55577;
w55579 <= not w55468 and not w55578;
w55580 <= not w55576 and w55579;
w55581 <= not w55468 and not w55580;
w55582 <= b(10) and not w55457;
w55583 <= not w55455 and w55582;
w55584 <= not w55459 and not w55583;
w55585 <= not w55581 and w55584;
w55586 <= not w55459 and not w55585;
w55587 <= b(11) and not w55448;
w55588 <= not w55446 and w55587;
w55589 <= not w55450 and not w55588;
w55590 <= not w55586 and w55589;
w55591 <= not w55450 and not w55590;
w55592 <= b(12) and not w55439;
w55593 <= not w55437 and w55592;
w55594 <= not w55441 and not w55593;
w55595 <= not w55591 and w55594;
w55596 <= not w55441 and not w55595;
w55597 <= b(13) and not w55430;
w55598 <= not w55428 and w55597;
w55599 <= not w55432 and not w55598;
w55600 <= not w55596 and w55599;
w55601 <= not w55432 and not w55600;
w55602 <= b(14) and not w55421;
w55603 <= not w55419 and w55602;
w55604 <= not w55423 and not w55603;
w55605 <= not w55601 and w55604;
w55606 <= not w55423 and not w55605;
w55607 <= b(15) and not w55412;
w55608 <= not w55410 and w55607;
w55609 <= not w55414 and not w55608;
w55610 <= not w55606 and w55609;
w55611 <= not w55414 and not w55610;
w55612 <= b(16) and not w55403;
w55613 <= not w55401 and w55612;
w55614 <= not w55405 and not w55613;
w55615 <= not w55611 and w55614;
w55616 <= not w55405 and not w55615;
w55617 <= b(17) and not w55394;
w55618 <= not w55392 and w55617;
w55619 <= not w55396 and not w55618;
w55620 <= not w55616 and w55619;
w55621 <= not w55396 and not w55620;
w55622 <= b(18) and not w55385;
w55623 <= not w55383 and w55622;
w55624 <= not w55387 and not w55623;
w55625 <= not w55621 and w55624;
w55626 <= not w55387 and not w55625;
w55627 <= b(19) and not w55376;
w55628 <= not w55374 and w55627;
w55629 <= not w55378 and not w55628;
w55630 <= not w55626 and w55629;
w55631 <= not w55378 and not w55630;
w55632 <= b(20) and not w55367;
w55633 <= not w55365 and w55632;
w55634 <= not w55369 and not w55633;
w55635 <= not w55631 and w55634;
w55636 <= not w55369 and not w55635;
w55637 <= b(21) and not w55358;
w55638 <= not w55356 and w55637;
w55639 <= not w55360 and not w55638;
w55640 <= not w55636 and w55639;
w55641 <= not w55360 and not w55640;
w55642 <= b(22) and not w55349;
w55643 <= not w55347 and w55642;
w55644 <= not w55351 and not w55643;
w55645 <= not w55641 and w55644;
w55646 <= not w55351 and not w55645;
w55647 <= b(23) and not w55340;
w55648 <= not w55338 and w55647;
w55649 <= not w55342 and not w55648;
w55650 <= not w55646 and w55649;
w55651 <= not w55342 and not w55650;
w55652 <= b(24) and not w55331;
w55653 <= not w55329 and w55652;
w55654 <= not w55333 and not w55653;
w55655 <= not w55651 and w55654;
w55656 <= not w55333 and not w55655;
w55657 <= b(25) and not w55322;
w55658 <= not w55320 and w55657;
w55659 <= not w55324 and not w55658;
w55660 <= not w55656 and w55659;
w55661 <= not w55324 and not w55660;
w55662 <= b(26) and not w55313;
w55663 <= not w55311 and w55662;
w55664 <= not w55315 and not w55663;
w55665 <= not w55661 and w55664;
w55666 <= not w55315 and not w55665;
w55667 <= b(27) and not w55304;
w55668 <= not w55302 and w55667;
w55669 <= not w55306 and not w55668;
w55670 <= not w55666 and w55669;
w55671 <= not w55306 and not w55670;
w55672 <= b(28) and not w55295;
w55673 <= not w55293 and w55672;
w55674 <= not w55297 and not w55673;
w55675 <= not w55671 and w55674;
w55676 <= not w55297 and not w55675;
w55677 <= b(29) and not w55286;
w55678 <= not w55284 and w55677;
w55679 <= not w55288 and not w55678;
w55680 <= not w55676 and w55679;
w55681 <= not w55288 and not w55680;
w55682 <= b(30) and not w55277;
w55683 <= not w55275 and w55682;
w55684 <= not w55279 and not w55683;
w55685 <= not w55681 and w55684;
w55686 <= not w55279 and not w55685;
w55687 <= b(31) and not w55268;
w55688 <= not w55266 and w55687;
w55689 <= not w55270 and not w55688;
w55690 <= not w55686 and w55689;
w55691 <= not w55270 and not w55690;
w55692 <= b(32) and not w55259;
w55693 <= not w55257 and w55692;
w55694 <= not w55261 and not w55693;
w55695 <= not w55691 and w55694;
w55696 <= not w55261 and not w55695;
w55697 <= b(33) and not w55250;
w55698 <= not w55248 and w55697;
w55699 <= not w55252 and not w55698;
w55700 <= not w55696 and w55699;
w55701 <= not w55252 and not w55700;
w55702 <= b(34) and not w55241;
w55703 <= not w55239 and w55702;
w55704 <= not w55243 and not w55703;
w55705 <= not w55701 and w55704;
w55706 <= not w55243 and not w55705;
w55707 <= b(35) and not w55232;
w55708 <= not w55230 and w55707;
w55709 <= not w55234 and not w55708;
w55710 <= not w55706 and w55709;
w55711 <= not w55234 and not w55710;
w55712 <= b(36) and not w55223;
w55713 <= not w55221 and w55712;
w55714 <= not w55225 and not w55713;
w55715 <= not w55711 and w55714;
w55716 <= not w55225 and not w55715;
w55717 <= b(37) and not w55214;
w55718 <= not w55212 and w55717;
w55719 <= not w55216 and not w55718;
w55720 <= not w55716 and w55719;
w55721 <= not w55216 and not w55720;
w55722 <= b(38) and not w55205;
w55723 <= not w55203 and w55722;
w55724 <= not w55207 and not w55723;
w55725 <= not w55721 and w55724;
w55726 <= not w55207 and not w55725;
w55727 <= b(39) and not w55196;
w55728 <= not w55194 and w55727;
w55729 <= not w55198 and not w55728;
w55730 <= not w55726 and w55729;
w55731 <= not w55198 and not w55730;
w55732 <= b(40) and not w55187;
w55733 <= not w55185 and w55732;
w55734 <= not w55189 and not w55733;
w55735 <= not w55731 and w55734;
w55736 <= not w55189 and not w55735;
w55737 <= b(41) and not w55178;
w55738 <= not w55176 and w55737;
w55739 <= not w55180 and not w55738;
w55740 <= not w55736 and w55739;
w55741 <= not w55180 and not w55740;
w55742 <= b(42) and not w55169;
w55743 <= not w55167 and w55742;
w55744 <= not w55171 and not w55743;
w55745 <= not w55741 and w55744;
w55746 <= not w55171 and not w55745;
w55747 <= b(43) and not w55160;
w55748 <= not w55158 and w55747;
w55749 <= not w55162 and not w55748;
w55750 <= not w55746 and w55749;
w55751 <= not w55162 and not w55750;
w55752 <= b(44) and not w55151;
w55753 <= not w55149 and w55752;
w55754 <= not w55153 and not w55753;
w55755 <= not w55751 and w55754;
w55756 <= not w55153 and not w55755;
w55757 <= b(45) and not w55142;
w55758 <= not w55140 and w55757;
w55759 <= not w55144 and not w55758;
w55760 <= not w55756 and w55759;
w55761 <= not w55144 and not w55760;
w55762 <= b(46) and not w55133;
w55763 <= not w55131 and w55762;
w55764 <= not w55135 and not w55763;
w55765 <= not w55761 and w55764;
w55766 <= not w55135 and not w55765;
w55767 <= b(47) and not w55124;
w55768 <= not w55122 and w55767;
w55769 <= not w55126 and not w55768;
w55770 <= not w55766 and w55769;
w55771 <= not w55126 and not w55770;
w55772 <= b(48) and not w55115;
w55773 <= not w55113 and w55772;
w55774 <= not w55117 and not w55773;
w55775 <= not w55771 and w55774;
w55776 <= not w55117 and not w55775;
w55777 <= b(49) and not w55106;
w55778 <= not w55104 and w55777;
w55779 <= not w55108 and not w55778;
w55780 <= not w55776 and w55779;
w55781 <= not w55108 and not w55780;
w55782 <= b(50) and not w55097;
w55783 <= not w55095 and w55782;
w55784 <= not w55099 and not w55783;
w55785 <= not w55781 and w55784;
w55786 <= not w55099 and not w55785;
w55787 <= b(51) and not w55088;
w55788 <= not w55086 and w55787;
w55789 <= not w55090 and not w55788;
w55790 <= not w55786 and w55789;
w55791 <= not w55090 and not w55790;
w55792 <= b(52) and not w55079;
w55793 <= not w55077 and w55792;
w55794 <= not w55081 and not w55793;
w55795 <= not w55791 and w55794;
w55796 <= not w55081 and not w55795;
w55797 <= b(53) and not w55070;
w55798 <= not w55068 and w55797;
w55799 <= not w55072 and not w55798;
w55800 <= not w55796 and w55799;
w55801 <= not w55072 and not w55800;
w55802 <= b(54) and not w55061;
w55803 <= not w55059 and w55802;
w55804 <= not w55063 and not w55803;
w55805 <= not w55801 and w55804;
w55806 <= not w55063 and not w55805;
w55807 <= b(55) and not w55052;
w55808 <= not w55050 and w55807;
w55809 <= not w55054 and not w55808;
w55810 <= not w55806 and w55809;
w55811 <= not w55054 and not w55810;
w55812 <= b(56) and not w55043;
w55813 <= not w55041 and w55812;
w55814 <= not w55045 and not w55813;
w55815 <= not w55811 and w55814;
w55816 <= not w55045 and not w55815;
w55817 <= b(57) and not w55034;
w55818 <= not w55032 and w55817;
w55819 <= not w55036 and not w55818;
w55820 <= not w55816 and w55819;
w55821 <= not w55036 and not w55820;
w55822 <= b(58) and not w55025;
w55823 <= not w55023 and w55822;
w55824 <= not w55027 and not w55823;
w55825 <= not w55821 and w55824;
w55826 <= not w55027 and not w55825;
w55827 <= b(59) and not w55016;
w55828 <= not w55014 and w55827;
w55829 <= not w55018 and not w55828;
w55830 <= not w55826 and w55829;
w55831 <= not w55018 and not w55830;
w55832 <= b(60) and not w55007;
w55833 <= not w55005 and w55832;
w55834 <= not w55009 and not w55833;
w55835 <= not w55831 and w55834;
w55836 <= not w55009 and not w55835;
w55837 <= b(61) and not w54998;
w55838 <= not w54996 and w55837;
w55839 <= not w55000 and not w55838;
w55840 <= not w55836 and w55839;
w55841 <= not w55000 and not w55840;
w55842 <= not w54146 and not w54986;
w55843 <= not w54984 and w55842;
w55844 <= not w54972 and w55843;
w55845 <= not w54984 and not w54986;
w55846 <= not w54973 and not w55845;
w55847 <= not w55844 and not w55846;
w55848 <= not w54991 and not w55847;
w55849 <= not w54983 and not w54990;
w55850 <= not w54989 and w55849;
w55851 <= not w55848 and not w55850;
w55852 <= not b(62) and not w55851;
w55853 <= b(62) and not w55850;
w55854 <= not w55848 and w55853;
w55855 <= not b(63) and not w55854;
w55856 <= not w55852 and w55855;
w55857 <= not w55841 and w55856;
w55858 <= w22 and not w55851;
w55859 <= not w55857 and not w55858;
w55860 <= not w55000 and not w55854;
w55861 <= not w55852 and w55860;
w55862 <= not w55840 and w55861;
w55863 <= not w55852 and not w55854;
w55864 <= not w55841 and not w55863;
w55865 <= not w55862 and not w55864;
w55866 <= not w55859 and not w55865;
w55867 <= not w55851 and not w55858;
w55868 <= not w55857 and w55867;
w55869 <= not w55866 and not w55868;
w55870 <= not b(63) and not w55869;
w55871 <= not w55009 and w55839;
w55872 <= not w55835 and w55871;
w55873 <= not w55836 and not w55839;
w55874 <= not w55872 and not w55873;
w55875 <= not w55859 and not w55874;
w55876 <= not w54999 and not w55858;
w55877 <= not w55857 and w55876;
w55878 <= not w55875 and not w55877;
w55879 <= not b(62) and not w55878;
w55880 <= not w55018 and w55834;
w55881 <= not w55830 and w55880;
w55882 <= not w55831 and not w55834;
w55883 <= not w55881 and not w55882;
w55884 <= not w55859 and not w55883;
w55885 <= not w55008 and not w55858;
w55886 <= not w55857 and w55885;
w55887 <= not w55884 and not w55886;
w55888 <= not b(61) and not w55887;
w55889 <= not w55027 and w55829;
w55890 <= not w55825 and w55889;
w55891 <= not w55826 and not w55829;
w55892 <= not w55890 and not w55891;
w55893 <= not w55859 and not w55892;
w55894 <= not w55017 and not w55858;
w55895 <= not w55857 and w55894;
w55896 <= not w55893 and not w55895;
w55897 <= not b(60) and not w55896;
w55898 <= not w55036 and w55824;
w55899 <= not w55820 and w55898;
w55900 <= not w55821 and not w55824;
w55901 <= not w55899 and not w55900;
w55902 <= not w55859 and not w55901;
w55903 <= not w55026 and not w55858;
w55904 <= not w55857 and w55903;
w55905 <= not w55902 and not w55904;
w55906 <= not b(59) and not w55905;
w55907 <= not w55045 and w55819;
w55908 <= not w55815 and w55907;
w55909 <= not w55816 and not w55819;
w55910 <= not w55908 and not w55909;
w55911 <= not w55859 and not w55910;
w55912 <= not w55035 and not w55858;
w55913 <= not w55857 and w55912;
w55914 <= not w55911 and not w55913;
w55915 <= not b(58) and not w55914;
w55916 <= not w55054 and w55814;
w55917 <= not w55810 and w55916;
w55918 <= not w55811 and not w55814;
w55919 <= not w55917 and not w55918;
w55920 <= not w55859 and not w55919;
w55921 <= not w55044 and not w55858;
w55922 <= not w55857 and w55921;
w55923 <= not w55920 and not w55922;
w55924 <= not b(57) and not w55923;
w55925 <= not w55063 and w55809;
w55926 <= not w55805 and w55925;
w55927 <= not w55806 and not w55809;
w55928 <= not w55926 and not w55927;
w55929 <= not w55859 and not w55928;
w55930 <= not w55053 and not w55858;
w55931 <= not w55857 and w55930;
w55932 <= not w55929 and not w55931;
w55933 <= not b(56) and not w55932;
w55934 <= not w55072 and w55804;
w55935 <= not w55800 and w55934;
w55936 <= not w55801 and not w55804;
w55937 <= not w55935 and not w55936;
w55938 <= not w55859 and not w55937;
w55939 <= not w55062 and not w55858;
w55940 <= not w55857 and w55939;
w55941 <= not w55938 and not w55940;
w55942 <= not b(55) and not w55941;
w55943 <= not w55081 and w55799;
w55944 <= not w55795 and w55943;
w55945 <= not w55796 and not w55799;
w55946 <= not w55944 and not w55945;
w55947 <= not w55859 and not w55946;
w55948 <= not w55071 and not w55858;
w55949 <= not w55857 and w55948;
w55950 <= not w55947 and not w55949;
w55951 <= not b(54) and not w55950;
w55952 <= not w55090 and w55794;
w55953 <= not w55790 and w55952;
w55954 <= not w55791 and not w55794;
w55955 <= not w55953 and not w55954;
w55956 <= not w55859 and not w55955;
w55957 <= not w55080 and not w55858;
w55958 <= not w55857 and w55957;
w55959 <= not w55956 and not w55958;
w55960 <= not b(53) and not w55959;
w55961 <= not w55099 and w55789;
w55962 <= not w55785 and w55961;
w55963 <= not w55786 and not w55789;
w55964 <= not w55962 and not w55963;
w55965 <= not w55859 and not w55964;
w55966 <= not w55089 and not w55858;
w55967 <= not w55857 and w55966;
w55968 <= not w55965 and not w55967;
w55969 <= not b(52) and not w55968;
w55970 <= not w55108 and w55784;
w55971 <= not w55780 and w55970;
w55972 <= not w55781 and not w55784;
w55973 <= not w55971 and not w55972;
w55974 <= not w55859 and not w55973;
w55975 <= not w55098 and not w55858;
w55976 <= not w55857 and w55975;
w55977 <= not w55974 and not w55976;
w55978 <= not b(51) and not w55977;
w55979 <= not w55117 and w55779;
w55980 <= not w55775 and w55979;
w55981 <= not w55776 and not w55779;
w55982 <= not w55980 and not w55981;
w55983 <= not w55859 and not w55982;
w55984 <= not w55107 and not w55858;
w55985 <= not w55857 and w55984;
w55986 <= not w55983 and not w55985;
w55987 <= not b(50) and not w55986;
w55988 <= not w55126 and w55774;
w55989 <= not w55770 and w55988;
w55990 <= not w55771 and not w55774;
w55991 <= not w55989 and not w55990;
w55992 <= not w55859 and not w55991;
w55993 <= not w55116 and not w55858;
w55994 <= not w55857 and w55993;
w55995 <= not w55992 and not w55994;
w55996 <= not b(49) and not w55995;
w55997 <= not w55135 and w55769;
w55998 <= not w55765 and w55997;
w55999 <= not w55766 and not w55769;
w56000 <= not w55998 and not w55999;
w56001 <= not w55859 and not w56000;
w56002 <= not w55125 and not w55858;
w56003 <= not w55857 and w56002;
w56004 <= not w56001 and not w56003;
w56005 <= not b(48) and not w56004;
w56006 <= not w55144 and w55764;
w56007 <= not w55760 and w56006;
w56008 <= not w55761 and not w55764;
w56009 <= not w56007 and not w56008;
w56010 <= not w55859 and not w56009;
w56011 <= not w55134 and not w55858;
w56012 <= not w55857 and w56011;
w56013 <= not w56010 and not w56012;
w56014 <= not b(47) and not w56013;
w56015 <= not w55153 and w55759;
w56016 <= not w55755 and w56015;
w56017 <= not w55756 and not w55759;
w56018 <= not w56016 and not w56017;
w56019 <= not w55859 and not w56018;
w56020 <= not w55143 and not w55858;
w56021 <= not w55857 and w56020;
w56022 <= not w56019 and not w56021;
w56023 <= not b(46) and not w56022;
w56024 <= not w55162 and w55754;
w56025 <= not w55750 and w56024;
w56026 <= not w55751 and not w55754;
w56027 <= not w56025 and not w56026;
w56028 <= not w55859 and not w56027;
w56029 <= not w55152 and not w55858;
w56030 <= not w55857 and w56029;
w56031 <= not w56028 and not w56030;
w56032 <= not b(45) and not w56031;
w56033 <= not w55171 and w55749;
w56034 <= not w55745 and w56033;
w56035 <= not w55746 and not w55749;
w56036 <= not w56034 and not w56035;
w56037 <= not w55859 and not w56036;
w56038 <= not w55161 and not w55858;
w56039 <= not w55857 and w56038;
w56040 <= not w56037 and not w56039;
w56041 <= not b(44) and not w56040;
w56042 <= not w55180 and w55744;
w56043 <= not w55740 and w56042;
w56044 <= not w55741 and not w55744;
w56045 <= not w56043 and not w56044;
w56046 <= not w55859 and not w56045;
w56047 <= not w55170 and not w55858;
w56048 <= not w55857 and w56047;
w56049 <= not w56046 and not w56048;
w56050 <= not b(43) and not w56049;
w56051 <= not w55189 and w55739;
w56052 <= not w55735 and w56051;
w56053 <= not w55736 and not w55739;
w56054 <= not w56052 and not w56053;
w56055 <= not w55859 and not w56054;
w56056 <= not w55179 and not w55858;
w56057 <= not w55857 and w56056;
w56058 <= not w56055 and not w56057;
w56059 <= not b(42) and not w56058;
w56060 <= not w55198 and w55734;
w56061 <= not w55730 and w56060;
w56062 <= not w55731 and not w55734;
w56063 <= not w56061 and not w56062;
w56064 <= not w55859 and not w56063;
w56065 <= not w55188 and not w55858;
w56066 <= not w55857 and w56065;
w56067 <= not w56064 and not w56066;
w56068 <= not b(41) and not w56067;
w56069 <= not w55207 and w55729;
w56070 <= not w55725 and w56069;
w56071 <= not w55726 and not w55729;
w56072 <= not w56070 and not w56071;
w56073 <= not w55859 and not w56072;
w56074 <= not w55197 and not w55858;
w56075 <= not w55857 and w56074;
w56076 <= not w56073 and not w56075;
w56077 <= not b(40) and not w56076;
w56078 <= not w55216 and w55724;
w56079 <= not w55720 and w56078;
w56080 <= not w55721 and not w55724;
w56081 <= not w56079 and not w56080;
w56082 <= not w55859 and not w56081;
w56083 <= not w55206 and not w55858;
w56084 <= not w55857 and w56083;
w56085 <= not w56082 and not w56084;
w56086 <= not b(39) and not w56085;
w56087 <= not w55225 and w55719;
w56088 <= not w55715 and w56087;
w56089 <= not w55716 and not w55719;
w56090 <= not w56088 and not w56089;
w56091 <= not w55859 and not w56090;
w56092 <= not w55215 and not w55858;
w56093 <= not w55857 and w56092;
w56094 <= not w56091 and not w56093;
w56095 <= not b(38) and not w56094;
w56096 <= not w55234 and w55714;
w56097 <= not w55710 and w56096;
w56098 <= not w55711 and not w55714;
w56099 <= not w56097 and not w56098;
w56100 <= not w55859 and not w56099;
w56101 <= not w55224 and not w55858;
w56102 <= not w55857 and w56101;
w56103 <= not w56100 and not w56102;
w56104 <= not b(37) and not w56103;
w56105 <= not w55243 and w55709;
w56106 <= not w55705 and w56105;
w56107 <= not w55706 and not w55709;
w56108 <= not w56106 and not w56107;
w56109 <= not w55859 and not w56108;
w56110 <= not w55233 and not w55858;
w56111 <= not w55857 and w56110;
w56112 <= not w56109 and not w56111;
w56113 <= not b(36) and not w56112;
w56114 <= not w55252 and w55704;
w56115 <= not w55700 and w56114;
w56116 <= not w55701 and not w55704;
w56117 <= not w56115 and not w56116;
w56118 <= not w55859 and not w56117;
w56119 <= not w55242 and not w55858;
w56120 <= not w55857 and w56119;
w56121 <= not w56118 and not w56120;
w56122 <= not b(35) and not w56121;
w56123 <= not w55261 and w55699;
w56124 <= not w55695 and w56123;
w56125 <= not w55696 and not w55699;
w56126 <= not w56124 and not w56125;
w56127 <= not w55859 and not w56126;
w56128 <= not w55251 and not w55858;
w56129 <= not w55857 and w56128;
w56130 <= not w56127 and not w56129;
w56131 <= not b(34) and not w56130;
w56132 <= not w55270 and w55694;
w56133 <= not w55690 and w56132;
w56134 <= not w55691 and not w55694;
w56135 <= not w56133 and not w56134;
w56136 <= not w55859 and not w56135;
w56137 <= not w55260 and not w55858;
w56138 <= not w55857 and w56137;
w56139 <= not w56136 and not w56138;
w56140 <= not b(33) and not w56139;
w56141 <= not w55279 and w55689;
w56142 <= not w55685 and w56141;
w56143 <= not w55686 and not w55689;
w56144 <= not w56142 and not w56143;
w56145 <= not w55859 and not w56144;
w56146 <= not w55269 and not w55858;
w56147 <= not w55857 and w56146;
w56148 <= not w56145 and not w56147;
w56149 <= not b(32) and not w56148;
w56150 <= not w55288 and w55684;
w56151 <= not w55680 and w56150;
w56152 <= not w55681 and not w55684;
w56153 <= not w56151 and not w56152;
w56154 <= not w55859 and not w56153;
w56155 <= not w55278 and not w55858;
w56156 <= not w55857 and w56155;
w56157 <= not w56154 and not w56156;
w56158 <= not b(31) and not w56157;
w56159 <= not w55297 and w55679;
w56160 <= not w55675 and w56159;
w56161 <= not w55676 and not w55679;
w56162 <= not w56160 and not w56161;
w56163 <= not w55859 and not w56162;
w56164 <= not w55287 and not w55858;
w56165 <= not w55857 and w56164;
w56166 <= not w56163 and not w56165;
w56167 <= not b(30) and not w56166;
w56168 <= not w55306 and w55674;
w56169 <= not w55670 and w56168;
w56170 <= not w55671 and not w55674;
w56171 <= not w56169 and not w56170;
w56172 <= not w55859 and not w56171;
w56173 <= not w55296 and not w55858;
w56174 <= not w55857 and w56173;
w56175 <= not w56172 and not w56174;
w56176 <= not b(29) and not w56175;
w56177 <= not w55315 and w55669;
w56178 <= not w55665 and w56177;
w56179 <= not w55666 and not w55669;
w56180 <= not w56178 and not w56179;
w56181 <= not w55859 and not w56180;
w56182 <= not w55305 and not w55858;
w56183 <= not w55857 and w56182;
w56184 <= not w56181 and not w56183;
w56185 <= not b(28) and not w56184;
w56186 <= not w55324 and w55664;
w56187 <= not w55660 and w56186;
w56188 <= not w55661 and not w55664;
w56189 <= not w56187 and not w56188;
w56190 <= not w55859 and not w56189;
w56191 <= not w55314 and not w55858;
w56192 <= not w55857 and w56191;
w56193 <= not w56190 and not w56192;
w56194 <= not b(27) and not w56193;
w56195 <= not w55333 and w55659;
w56196 <= not w55655 and w56195;
w56197 <= not w55656 and not w55659;
w56198 <= not w56196 and not w56197;
w56199 <= not w55859 and not w56198;
w56200 <= not w55323 and not w55858;
w56201 <= not w55857 and w56200;
w56202 <= not w56199 and not w56201;
w56203 <= not b(26) and not w56202;
w56204 <= not w55342 and w55654;
w56205 <= not w55650 and w56204;
w56206 <= not w55651 and not w55654;
w56207 <= not w56205 and not w56206;
w56208 <= not w55859 and not w56207;
w56209 <= not w55332 and not w55858;
w56210 <= not w55857 and w56209;
w56211 <= not w56208 and not w56210;
w56212 <= not b(25) and not w56211;
w56213 <= not w55351 and w55649;
w56214 <= not w55645 and w56213;
w56215 <= not w55646 and not w55649;
w56216 <= not w56214 and not w56215;
w56217 <= not w55859 and not w56216;
w56218 <= not w55341 and not w55858;
w56219 <= not w55857 and w56218;
w56220 <= not w56217 and not w56219;
w56221 <= not b(24) and not w56220;
w56222 <= not w55360 and w55644;
w56223 <= not w55640 and w56222;
w56224 <= not w55641 and not w55644;
w56225 <= not w56223 and not w56224;
w56226 <= not w55859 and not w56225;
w56227 <= not w55350 and not w55858;
w56228 <= not w55857 and w56227;
w56229 <= not w56226 and not w56228;
w56230 <= not b(23) and not w56229;
w56231 <= not w55369 and w55639;
w56232 <= not w55635 and w56231;
w56233 <= not w55636 and not w55639;
w56234 <= not w56232 and not w56233;
w56235 <= not w55859 and not w56234;
w56236 <= not w55359 and not w55858;
w56237 <= not w55857 and w56236;
w56238 <= not w56235 and not w56237;
w56239 <= not b(22) and not w56238;
w56240 <= not w55378 and w55634;
w56241 <= not w55630 and w56240;
w56242 <= not w55631 and not w55634;
w56243 <= not w56241 and not w56242;
w56244 <= not w55859 and not w56243;
w56245 <= not w55368 and not w55858;
w56246 <= not w55857 and w56245;
w56247 <= not w56244 and not w56246;
w56248 <= not b(21) and not w56247;
w56249 <= not w55387 and w55629;
w56250 <= not w55625 and w56249;
w56251 <= not w55626 and not w55629;
w56252 <= not w56250 and not w56251;
w56253 <= not w55859 and not w56252;
w56254 <= not w55377 and not w55858;
w56255 <= not w55857 and w56254;
w56256 <= not w56253 and not w56255;
w56257 <= not b(20) and not w56256;
w56258 <= not w55396 and w55624;
w56259 <= not w55620 and w56258;
w56260 <= not w55621 and not w55624;
w56261 <= not w56259 and not w56260;
w56262 <= not w55859 and not w56261;
w56263 <= not w55386 and not w55858;
w56264 <= not w55857 and w56263;
w56265 <= not w56262 and not w56264;
w56266 <= not b(19) and not w56265;
w56267 <= not w55405 and w55619;
w56268 <= not w55615 and w56267;
w56269 <= not w55616 and not w55619;
w56270 <= not w56268 and not w56269;
w56271 <= not w55859 and not w56270;
w56272 <= not w55395 and not w55858;
w56273 <= not w55857 and w56272;
w56274 <= not w56271 and not w56273;
w56275 <= not b(18) and not w56274;
w56276 <= not w55414 and w55614;
w56277 <= not w55610 and w56276;
w56278 <= not w55611 and not w55614;
w56279 <= not w56277 and not w56278;
w56280 <= not w55859 and not w56279;
w56281 <= not w55404 and not w55858;
w56282 <= not w55857 and w56281;
w56283 <= not w56280 and not w56282;
w56284 <= not b(17) and not w56283;
w56285 <= not w55423 and w55609;
w56286 <= not w55605 and w56285;
w56287 <= not w55606 and not w55609;
w56288 <= not w56286 and not w56287;
w56289 <= not w55859 and not w56288;
w56290 <= not w55413 and not w55858;
w56291 <= not w55857 and w56290;
w56292 <= not w56289 and not w56291;
w56293 <= not b(16) and not w56292;
w56294 <= not w55432 and w55604;
w56295 <= not w55600 and w56294;
w56296 <= not w55601 and not w55604;
w56297 <= not w56295 and not w56296;
w56298 <= not w55859 and not w56297;
w56299 <= not w55422 and not w55858;
w56300 <= not w55857 and w56299;
w56301 <= not w56298 and not w56300;
w56302 <= not b(15) and not w56301;
w56303 <= not w55441 and w55599;
w56304 <= not w55595 and w56303;
w56305 <= not w55596 and not w55599;
w56306 <= not w56304 and not w56305;
w56307 <= not w55859 and not w56306;
w56308 <= not w55431 and not w55858;
w56309 <= not w55857 and w56308;
w56310 <= not w56307 and not w56309;
w56311 <= not b(14) and not w56310;
w56312 <= not w55450 and w55594;
w56313 <= not w55590 and w56312;
w56314 <= not w55591 and not w55594;
w56315 <= not w56313 and not w56314;
w56316 <= not w55859 and not w56315;
w56317 <= not w55440 and not w55858;
w56318 <= not w55857 and w56317;
w56319 <= not w56316 and not w56318;
w56320 <= not b(13) and not w56319;
w56321 <= not w55459 and w55589;
w56322 <= not w55585 and w56321;
w56323 <= not w55586 and not w55589;
w56324 <= not w56322 and not w56323;
w56325 <= not w55859 and not w56324;
w56326 <= not w55449 and not w55858;
w56327 <= not w55857 and w56326;
w56328 <= not w56325 and not w56327;
w56329 <= not b(12) and not w56328;
w56330 <= not w55468 and w55584;
w56331 <= not w55580 and w56330;
w56332 <= not w55581 and not w55584;
w56333 <= not w56331 and not w56332;
w56334 <= not w55859 and not w56333;
w56335 <= not w55458 and not w55858;
w56336 <= not w55857 and w56335;
w56337 <= not w56334 and not w56336;
w56338 <= not b(11) and not w56337;
w56339 <= not w55477 and w55579;
w56340 <= not w55575 and w56339;
w56341 <= not w55576 and not w55579;
w56342 <= not w56340 and not w56341;
w56343 <= not w55859 and not w56342;
w56344 <= not w55467 and not w55858;
w56345 <= not w55857 and w56344;
w56346 <= not w56343 and not w56345;
w56347 <= not b(10) and not w56346;
w56348 <= not w55486 and w55574;
w56349 <= not w55570 and w56348;
w56350 <= not w55571 and not w55574;
w56351 <= not w56349 and not w56350;
w56352 <= not w55859 and not w56351;
w56353 <= not w55476 and not w55858;
w56354 <= not w55857 and w56353;
w56355 <= not w56352 and not w56354;
w56356 <= not b(9) and not w56355;
w56357 <= not w55495 and w55569;
w56358 <= not w55565 and w56357;
w56359 <= not w55566 and not w55569;
w56360 <= not w56358 and not w56359;
w56361 <= not w55859 and not w56360;
w56362 <= not w55485 and not w55858;
w56363 <= not w55857 and w56362;
w56364 <= not w56361 and not w56363;
w56365 <= not b(8) and not w56364;
w56366 <= not w55504 and w55564;
w56367 <= not w55560 and w56366;
w56368 <= not w55561 and not w55564;
w56369 <= not w56367 and not w56368;
w56370 <= not w55859 and not w56369;
w56371 <= not w55494 and not w55858;
w56372 <= not w55857 and w56371;
w56373 <= not w56370 and not w56372;
w56374 <= not b(7) and not w56373;
w56375 <= not w55513 and w55559;
w56376 <= not w55555 and w56375;
w56377 <= not w55556 and not w55559;
w56378 <= not w56376 and not w56377;
w56379 <= not w55859 and not w56378;
w56380 <= not w55503 and not w55858;
w56381 <= not w55857 and w56380;
w56382 <= not w56379 and not w56381;
w56383 <= not b(6) and not w56382;
w56384 <= not w55522 and w55554;
w56385 <= not w55550 and w56384;
w56386 <= not w55551 and not w55554;
w56387 <= not w56385 and not w56386;
w56388 <= not w55859 and not w56387;
w56389 <= not w55512 and not w55858;
w56390 <= not w55857 and w56389;
w56391 <= not w56388 and not w56390;
w56392 <= not b(5) and not w56391;
w56393 <= not w55530 and w55549;
w56394 <= not w55545 and w56393;
w56395 <= not w55546 and not w55549;
w56396 <= not w56394 and not w56395;
w56397 <= not w55859 and not w56396;
w56398 <= not w55521 and not w55858;
w56399 <= not w55857 and w56398;
w56400 <= not w56397 and not w56399;
w56401 <= not b(4) and not w56400;
w56402 <= not w55540 and w55544;
w56403 <= not w55539 and w56402;
w56404 <= not w55541 and not w55544;
w56405 <= not w56403 and not w56404;
w56406 <= not w55859 and not w56405;
w56407 <= not w55529 and not w55858;
w56408 <= not w55857 and w56407;
w56409 <= not w56406 and not w56408;
w56410 <= not b(3) and not w56409;
w56411 <= w27526 and not w55537;
w56412 <= not w55535 and w56411;
w56413 <= not w55539 and not w56412;
w56414 <= not w55859 and w56413;
w56415 <= not w55534 and not w55858;
w56416 <= not w55857 and w56415;
w56417 <= not w56414 and not w56416;
w56418 <= not b(2) and not w56417;
w56419 <= b(0) and not w55859;
w56420 <= a(1) and not w56419;
w56421 <= w27526 and not w55859;
w56422 <= not w56420 and not w56421;
w56423 <= b(1) and not w56422;
w56424 <= not b(1) and not w56421;
w56425 <= not w56420 and w56424;
w56426 <= not w56423 and not w56425;
w56427 <= not w28088 and not w56426;
w56428 <= not b(1) and not w56422;
w56429 <= not w56427 and not w56428;
w56430 <= b(2) and not w56416;
w56431 <= not w56414 and w56430;
w56432 <= not w56418 and not w56431;
w56433 <= not w56429 and w56432;
w56434 <= not w56418 and not w56433;
w56435 <= b(3) and not w56408;
w56436 <= not w56406 and w56435;
w56437 <= not w56410 and not w56436;
w56438 <= not w56434 and w56437;
w56439 <= not w56410 and not w56438;
w56440 <= b(4) and not w56399;
w56441 <= not w56397 and w56440;
w56442 <= not w56401 and not w56441;
w56443 <= not w56439 and w56442;
w56444 <= not w56401 and not w56443;
w56445 <= b(5) and not w56390;
w56446 <= not w56388 and w56445;
w56447 <= not w56392 and not w56446;
w56448 <= not w56444 and w56447;
w56449 <= not w56392 and not w56448;
w56450 <= b(6) and not w56381;
w56451 <= not w56379 and w56450;
w56452 <= not w56383 and not w56451;
w56453 <= not w56449 and w56452;
w56454 <= not w56383 and not w56453;
w56455 <= b(7) and not w56372;
w56456 <= not w56370 and w56455;
w56457 <= not w56374 and not w56456;
w56458 <= not w56454 and w56457;
w56459 <= not w56374 and not w56458;
w56460 <= b(8) and not w56363;
w56461 <= not w56361 and w56460;
w56462 <= not w56365 and not w56461;
w56463 <= not w56459 and w56462;
w56464 <= not w56365 and not w56463;
w56465 <= b(9) and not w56354;
w56466 <= not w56352 and w56465;
w56467 <= not w56356 and not w56466;
w56468 <= not w56464 and w56467;
w56469 <= not w56356 and not w56468;
w56470 <= b(10) and not w56345;
w56471 <= not w56343 and w56470;
w56472 <= not w56347 and not w56471;
w56473 <= not w56469 and w56472;
w56474 <= not w56347 and not w56473;
w56475 <= b(11) and not w56336;
w56476 <= not w56334 and w56475;
w56477 <= not w56338 and not w56476;
w56478 <= not w56474 and w56477;
w56479 <= not w56338 and not w56478;
w56480 <= b(12) and not w56327;
w56481 <= not w56325 and w56480;
w56482 <= not w56329 and not w56481;
w56483 <= not w56479 and w56482;
w56484 <= not w56329 and not w56483;
w56485 <= b(13) and not w56318;
w56486 <= not w56316 and w56485;
w56487 <= not w56320 and not w56486;
w56488 <= not w56484 and w56487;
w56489 <= not w56320 and not w56488;
w56490 <= b(14) and not w56309;
w56491 <= not w56307 and w56490;
w56492 <= not w56311 and not w56491;
w56493 <= not w56489 and w56492;
w56494 <= not w56311 and not w56493;
w56495 <= b(15) and not w56300;
w56496 <= not w56298 and w56495;
w56497 <= not w56302 and not w56496;
w56498 <= not w56494 and w56497;
w56499 <= not w56302 and not w56498;
w56500 <= b(16) and not w56291;
w56501 <= not w56289 and w56500;
w56502 <= not w56293 and not w56501;
w56503 <= not w56499 and w56502;
w56504 <= not w56293 and not w56503;
w56505 <= b(17) and not w56282;
w56506 <= not w56280 and w56505;
w56507 <= not w56284 and not w56506;
w56508 <= not w56504 and w56507;
w56509 <= not w56284 and not w56508;
w56510 <= b(18) and not w56273;
w56511 <= not w56271 and w56510;
w56512 <= not w56275 and not w56511;
w56513 <= not w56509 and w56512;
w56514 <= not w56275 and not w56513;
w56515 <= b(19) and not w56264;
w56516 <= not w56262 and w56515;
w56517 <= not w56266 and not w56516;
w56518 <= not w56514 and w56517;
w56519 <= not w56266 and not w56518;
w56520 <= b(20) and not w56255;
w56521 <= not w56253 and w56520;
w56522 <= not w56257 and not w56521;
w56523 <= not w56519 and w56522;
w56524 <= not w56257 and not w56523;
w56525 <= b(21) and not w56246;
w56526 <= not w56244 and w56525;
w56527 <= not w56248 and not w56526;
w56528 <= not w56524 and w56527;
w56529 <= not w56248 and not w56528;
w56530 <= b(22) and not w56237;
w56531 <= not w56235 and w56530;
w56532 <= not w56239 and not w56531;
w56533 <= not w56529 and w56532;
w56534 <= not w56239 and not w56533;
w56535 <= b(23) and not w56228;
w56536 <= not w56226 and w56535;
w56537 <= not w56230 and not w56536;
w56538 <= not w56534 and w56537;
w56539 <= not w56230 and not w56538;
w56540 <= b(24) and not w56219;
w56541 <= not w56217 and w56540;
w56542 <= not w56221 and not w56541;
w56543 <= not w56539 and w56542;
w56544 <= not w56221 and not w56543;
w56545 <= b(25) and not w56210;
w56546 <= not w56208 and w56545;
w56547 <= not w56212 and not w56546;
w56548 <= not w56544 and w56547;
w56549 <= not w56212 and not w56548;
w56550 <= b(26) and not w56201;
w56551 <= not w56199 and w56550;
w56552 <= not w56203 and not w56551;
w56553 <= not w56549 and w56552;
w56554 <= not w56203 and not w56553;
w56555 <= b(27) and not w56192;
w56556 <= not w56190 and w56555;
w56557 <= not w56194 and not w56556;
w56558 <= not w56554 and w56557;
w56559 <= not w56194 and not w56558;
w56560 <= b(28) and not w56183;
w56561 <= not w56181 and w56560;
w56562 <= not w56185 and not w56561;
w56563 <= not w56559 and w56562;
w56564 <= not w56185 and not w56563;
w56565 <= b(29) and not w56174;
w56566 <= not w56172 and w56565;
w56567 <= not w56176 and not w56566;
w56568 <= not w56564 and w56567;
w56569 <= not w56176 and not w56568;
w56570 <= b(30) and not w56165;
w56571 <= not w56163 and w56570;
w56572 <= not w56167 and not w56571;
w56573 <= not w56569 and w56572;
w56574 <= not w56167 and not w56573;
w56575 <= b(31) and not w56156;
w56576 <= not w56154 and w56575;
w56577 <= not w56158 and not w56576;
w56578 <= not w56574 and w56577;
w56579 <= not w56158 and not w56578;
w56580 <= b(32) and not w56147;
w56581 <= not w56145 and w56580;
w56582 <= not w56149 and not w56581;
w56583 <= not w56579 and w56582;
w56584 <= not w56149 and not w56583;
w56585 <= b(33) and not w56138;
w56586 <= not w56136 and w56585;
w56587 <= not w56140 and not w56586;
w56588 <= not w56584 and w56587;
w56589 <= not w56140 and not w56588;
w56590 <= b(34) and not w56129;
w56591 <= not w56127 and w56590;
w56592 <= not w56131 and not w56591;
w56593 <= not w56589 and w56592;
w56594 <= not w56131 and not w56593;
w56595 <= b(35) and not w56120;
w56596 <= not w56118 and w56595;
w56597 <= not w56122 and not w56596;
w56598 <= not w56594 and w56597;
w56599 <= not w56122 and not w56598;
w56600 <= b(36) and not w56111;
w56601 <= not w56109 and w56600;
w56602 <= not w56113 and not w56601;
w56603 <= not w56599 and w56602;
w56604 <= not w56113 and not w56603;
w56605 <= b(37) and not w56102;
w56606 <= not w56100 and w56605;
w56607 <= not w56104 and not w56606;
w56608 <= not w56604 and w56607;
w56609 <= not w56104 and not w56608;
w56610 <= b(38) and not w56093;
w56611 <= not w56091 and w56610;
w56612 <= not w56095 and not w56611;
w56613 <= not w56609 and w56612;
w56614 <= not w56095 and not w56613;
w56615 <= b(39) and not w56084;
w56616 <= not w56082 and w56615;
w56617 <= not w56086 and not w56616;
w56618 <= not w56614 and w56617;
w56619 <= not w56086 and not w56618;
w56620 <= b(40) and not w56075;
w56621 <= not w56073 and w56620;
w56622 <= not w56077 and not w56621;
w56623 <= not w56619 and w56622;
w56624 <= not w56077 and not w56623;
w56625 <= b(41) and not w56066;
w56626 <= not w56064 and w56625;
w56627 <= not w56068 and not w56626;
w56628 <= not w56624 and w56627;
w56629 <= not w56068 and not w56628;
w56630 <= b(42) and not w56057;
w56631 <= not w56055 and w56630;
w56632 <= not w56059 and not w56631;
w56633 <= not w56629 and w56632;
w56634 <= not w56059 and not w56633;
w56635 <= b(43) and not w56048;
w56636 <= not w56046 and w56635;
w56637 <= not w56050 and not w56636;
w56638 <= not w56634 and w56637;
w56639 <= not w56050 and not w56638;
w56640 <= b(44) and not w56039;
w56641 <= not w56037 and w56640;
w56642 <= not w56041 and not w56641;
w56643 <= not w56639 and w56642;
w56644 <= not w56041 and not w56643;
w56645 <= b(45) and not w56030;
w56646 <= not w56028 and w56645;
w56647 <= not w56032 and not w56646;
w56648 <= not w56644 and w56647;
w56649 <= not w56032 and not w56648;
w56650 <= b(46) and not w56021;
w56651 <= not w56019 and w56650;
w56652 <= not w56023 and not w56651;
w56653 <= not w56649 and w56652;
w56654 <= not w56023 and not w56653;
w56655 <= b(47) and not w56012;
w56656 <= not w56010 and w56655;
w56657 <= not w56014 and not w56656;
w56658 <= not w56654 and w56657;
w56659 <= not w56014 and not w56658;
w56660 <= b(48) and not w56003;
w56661 <= not w56001 and w56660;
w56662 <= not w56005 and not w56661;
w56663 <= not w56659 and w56662;
w56664 <= not w56005 and not w56663;
w56665 <= b(49) and not w55994;
w56666 <= not w55992 and w56665;
w56667 <= not w55996 and not w56666;
w56668 <= not w56664 and w56667;
w56669 <= not w55996 and not w56668;
w56670 <= b(50) and not w55985;
w56671 <= not w55983 and w56670;
w56672 <= not w55987 and not w56671;
w56673 <= not w56669 and w56672;
w56674 <= not w55987 and not w56673;
w56675 <= b(51) and not w55976;
w56676 <= not w55974 and w56675;
w56677 <= not w55978 and not w56676;
w56678 <= not w56674 and w56677;
w56679 <= not w55978 and not w56678;
w56680 <= b(52) and not w55967;
w56681 <= not w55965 and w56680;
w56682 <= not w55969 and not w56681;
w56683 <= not w56679 and w56682;
w56684 <= not w55969 and not w56683;
w56685 <= b(53) and not w55958;
w56686 <= not w55956 and w56685;
w56687 <= not w55960 and not w56686;
w56688 <= not w56684 and w56687;
w56689 <= not w55960 and not w56688;
w56690 <= b(54) and not w55949;
w56691 <= not w55947 and w56690;
w56692 <= not w55951 and not w56691;
w56693 <= not w56689 and w56692;
w56694 <= not w55951 and not w56693;
w56695 <= b(55) and not w55940;
w56696 <= not w55938 and w56695;
w56697 <= not w55942 and not w56696;
w56698 <= not w56694 and w56697;
w56699 <= not w55942 and not w56698;
w56700 <= b(56) and not w55931;
w56701 <= not w55929 and w56700;
w56702 <= not w55933 and not w56701;
w56703 <= not w56699 and w56702;
w56704 <= not w55933 and not w56703;
w56705 <= b(57) and not w55922;
w56706 <= not w55920 and w56705;
w56707 <= not w55924 and not w56706;
w56708 <= not w56704 and w56707;
w56709 <= not w55924 and not w56708;
w56710 <= b(58) and not w55913;
w56711 <= not w55911 and w56710;
w56712 <= not w55915 and not w56711;
w56713 <= not w56709 and w56712;
w56714 <= not w55915 and not w56713;
w56715 <= b(59) and not w55904;
w56716 <= not w55902 and w56715;
w56717 <= not w55906 and not w56716;
w56718 <= not w56714 and w56717;
w56719 <= not w55906 and not w56718;
w56720 <= b(60) and not w55895;
w56721 <= not w55893 and w56720;
w56722 <= not w55897 and not w56721;
w56723 <= not w56719 and w56722;
w56724 <= not w55897 and not w56723;
w56725 <= b(61) and not w55886;
w56726 <= not w55884 and w56725;
w56727 <= not w55888 and not w56726;
w56728 <= not w56724 and w56727;
w56729 <= not w55888 and not w56728;
w56730 <= b(62) and not w55877;
w56731 <= not w55875 and w56730;
w56732 <= not w55879 and not w56731;
w56733 <= not w56729 and w56732;
w56734 <= not w55879 and not w56733;
w56735 <= b(63) and not w55868;
w56736 <= not w55866 and w56735;
w56737 <= not w55870 and not w56736;
w56738 <= not w56734 and w56737;
w56739 <= not w55870 and not w56738;
w56740 <= b(0) and not w56739;
w56741 <= a(0) and not w56740;
w56742 <= w28088 and not w56739;
w56743 <= not w56741 and not w56742;
w56744 <= w28088 and not w56425;
w56745 <= not w56423 and w56744;
w56746 <= not w56427 and not w56745;
w56747 <= not w56739 and w56746;
w56748 <= not w55870 and not w56422;
w56749 <= not w56738 and w56748;
w56750 <= not w56747 and not w56749;
w56751 <= not w56428 and w56432;
w56752 <= not w56427 and w56751;
w56753 <= not w56429 and not w56432;
w56754 <= not w56752 and not w56753;
w56755 <= not w56739 and not w56754;
w56756 <= not w55870 and not w56417;
w56757 <= not w56738 and w56756;
w56758 <= not w56755 and not w56757;
w56759 <= not w56418 and w56437;
w56760 <= not w56433 and w56759;
w56761 <= not w56434 and not w56437;
w56762 <= not w56760 and not w56761;
w56763 <= not w56739 and not w56762;
w56764 <= not w55870 and not w56409;
w56765 <= not w56738 and w56764;
w56766 <= not w56763 and not w56765;
w56767 <= not w56410 and w56442;
w56768 <= not w56438 and w56767;
w56769 <= not w56439 and not w56442;
w56770 <= not w56768 and not w56769;
w56771 <= not w56739 and not w56770;
w56772 <= not w55870 and not w56400;
w56773 <= not w56738 and w56772;
w56774 <= not w56771 and not w56773;
w56775 <= not w56401 and w56447;
w56776 <= not w56443 and w56775;
w56777 <= not w56444 and not w56447;
w56778 <= not w56776 and not w56777;
w56779 <= not w56739 and not w56778;
w56780 <= not w55870 and not w56391;
w56781 <= not w56738 and w56780;
w56782 <= not w56779 and not w56781;
w56783 <= not w56392 and w56452;
w56784 <= not w56448 and w56783;
w56785 <= not w56449 and not w56452;
w56786 <= not w56784 and not w56785;
w56787 <= not w56739 and not w56786;
w56788 <= not w55870 and not w56382;
w56789 <= not w56738 and w56788;
w56790 <= not w56787 and not w56789;
w56791 <= not w56383 and w56457;
w56792 <= not w56453 and w56791;
w56793 <= not w56454 and not w56457;
w56794 <= not w56792 and not w56793;
w56795 <= not w56739 and not w56794;
w56796 <= not w55870 and not w56373;
w56797 <= not w56738 and w56796;
w56798 <= not w56795 and not w56797;
w56799 <= not w56374 and w56462;
w56800 <= not w56458 and w56799;
w56801 <= not w56459 and not w56462;
w56802 <= not w56800 and not w56801;
w56803 <= not w56739 and not w56802;
w56804 <= not w55870 and not w56364;
w56805 <= not w56738 and w56804;
w56806 <= not w56803 and not w56805;
w56807 <= not w56365 and w56467;
w56808 <= not w56463 and w56807;
w56809 <= not w56464 and not w56467;
w56810 <= not w56808 and not w56809;
w56811 <= not w56739 and not w56810;
w56812 <= not w55870 and not w56355;
w56813 <= not w56738 and w56812;
w56814 <= not w56811 and not w56813;
w56815 <= not w56356 and w56472;
w56816 <= not w56468 and w56815;
w56817 <= not w56469 and not w56472;
w56818 <= not w56816 and not w56817;
w56819 <= not w56739 and not w56818;
w56820 <= not w55870 and not w56346;
w56821 <= not w56738 and w56820;
w56822 <= not w56819 and not w56821;
w56823 <= not w56347 and w56477;
w56824 <= not w56473 and w56823;
w56825 <= not w56474 and not w56477;
w56826 <= not w56824 and not w56825;
w56827 <= not w56739 and not w56826;
w56828 <= not w55870 and not w56337;
w56829 <= not w56738 and w56828;
w56830 <= not w56827 and not w56829;
w56831 <= not w56338 and w56482;
w56832 <= not w56478 and w56831;
w56833 <= not w56479 and not w56482;
w56834 <= not w56832 and not w56833;
w56835 <= not w56739 and not w56834;
w56836 <= not w55870 and not w56328;
w56837 <= not w56738 and w56836;
w56838 <= not w56835 and not w56837;
w56839 <= not w56329 and w56487;
w56840 <= not w56483 and w56839;
w56841 <= not w56484 and not w56487;
w56842 <= not w56840 and not w56841;
w56843 <= not w56739 and not w56842;
w56844 <= not w55870 and not w56319;
w56845 <= not w56738 and w56844;
w56846 <= not w56843 and not w56845;
w56847 <= not w56320 and w56492;
w56848 <= not w56488 and w56847;
w56849 <= not w56489 and not w56492;
w56850 <= not w56848 and not w56849;
w56851 <= not w56739 and not w56850;
w56852 <= not w55870 and not w56310;
w56853 <= not w56738 and w56852;
w56854 <= not w56851 and not w56853;
w56855 <= not w56311 and w56497;
w56856 <= not w56493 and w56855;
w56857 <= not w56494 and not w56497;
w56858 <= not w56856 and not w56857;
w56859 <= not w56739 and not w56858;
w56860 <= not w55870 and not w56301;
w56861 <= not w56738 and w56860;
w56862 <= not w56859 and not w56861;
w56863 <= not w56302 and w56502;
w56864 <= not w56498 and w56863;
w56865 <= not w56499 and not w56502;
w56866 <= not w56864 and not w56865;
w56867 <= not w56739 and not w56866;
w56868 <= not w55870 and not w56292;
w56869 <= not w56738 and w56868;
w56870 <= not w56867 and not w56869;
w56871 <= not w56293 and w56507;
w56872 <= not w56503 and w56871;
w56873 <= not w56504 and not w56507;
w56874 <= not w56872 and not w56873;
w56875 <= not w56739 and not w56874;
w56876 <= not w55870 and not w56283;
w56877 <= not w56738 and w56876;
w56878 <= not w56875 and not w56877;
w56879 <= not w56284 and w56512;
w56880 <= not w56508 and w56879;
w56881 <= not w56509 and not w56512;
w56882 <= not w56880 and not w56881;
w56883 <= not w56739 and not w56882;
w56884 <= not w55870 and not w56274;
w56885 <= not w56738 and w56884;
w56886 <= not w56883 and not w56885;
w56887 <= not w56275 and w56517;
w56888 <= not w56513 and w56887;
w56889 <= not w56514 and not w56517;
w56890 <= not w56888 and not w56889;
w56891 <= not w56739 and not w56890;
w56892 <= not w55870 and not w56265;
w56893 <= not w56738 and w56892;
w56894 <= not w56891 and not w56893;
w56895 <= not w56266 and w56522;
w56896 <= not w56518 and w56895;
w56897 <= not w56519 and not w56522;
w56898 <= not w56896 and not w56897;
w56899 <= not w56739 and not w56898;
w56900 <= not w55870 and not w56256;
w56901 <= not w56738 and w56900;
w56902 <= not w56899 and not w56901;
w56903 <= not w56257 and w56527;
w56904 <= not w56523 and w56903;
w56905 <= not w56524 and not w56527;
w56906 <= not w56904 and not w56905;
w56907 <= not w56739 and not w56906;
w56908 <= not w55870 and not w56247;
w56909 <= not w56738 and w56908;
w56910 <= not w56907 and not w56909;
w56911 <= not w56248 and w56532;
w56912 <= not w56528 and w56911;
w56913 <= not w56529 and not w56532;
w56914 <= not w56912 and not w56913;
w56915 <= not w56739 and not w56914;
w56916 <= not w55870 and not w56238;
w56917 <= not w56738 and w56916;
w56918 <= not w56915 and not w56917;
w56919 <= not w56239 and w56537;
w56920 <= not w56533 and w56919;
w56921 <= not w56534 and not w56537;
w56922 <= not w56920 and not w56921;
w56923 <= not w56739 and not w56922;
w56924 <= not w55870 and not w56229;
w56925 <= not w56738 and w56924;
w56926 <= not w56923 and not w56925;
w56927 <= not w56230 and w56542;
w56928 <= not w56538 and w56927;
w56929 <= not w56539 and not w56542;
w56930 <= not w56928 and not w56929;
w56931 <= not w56739 and not w56930;
w56932 <= not w55870 and not w56220;
w56933 <= not w56738 and w56932;
w56934 <= not w56931 and not w56933;
w56935 <= not w56221 and w56547;
w56936 <= not w56543 and w56935;
w56937 <= not w56544 and not w56547;
w56938 <= not w56936 and not w56937;
w56939 <= not w56739 and not w56938;
w56940 <= not w55870 and not w56211;
w56941 <= not w56738 and w56940;
w56942 <= not w56939 and not w56941;
w56943 <= not w56212 and w56552;
w56944 <= not w56548 and w56943;
w56945 <= not w56549 and not w56552;
w56946 <= not w56944 and not w56945;
w56947 <= not w56739 and not w56946;
w56948 <= not w55870 and not w56202;
w56949 <= not w56738 and w56948;
w56950 <= not w56947 and not w56949;
w56951 <= not w56203 and w56557;
w56952 <= not w56553 and w56951;
w56953 <= not w56554 and not w56557;
w56954 <= not w56952 and not w56953;
w56955 <= not w56739 and not w56954;
w56956 <= not w55870 and not w56193;
w56957 <= not w56738 and w56956;
w56958 <= not w56955 and not w56957;
w56959 <= not w56194 and w56562;
w56960 <= not w56558 and w56959;
w56961 <= not w56559 and not w56562;
w56962 <= not w56960 and not w56961;
w56963 <= not w56739 and not w56962;
w56964 <= not w55870 and not w56184;
w56965 <= not w56738 and w56964;
w56966 <= not w56963 and not w56965;
w56967 <= not w56185 and w56567;
w56968 <= not w56563 and w56967;
w56969 <= not w56564 and not w56567;
w56970 <= not w56968 and not w56969;
w56971 <= not w56739 and not w56970;
w56972 <= not w55870 and not w56175;
w56973 <= not w56738 and w56972;
w56974 <= not w56971 and not w56973;
w56975 <= not w56176 and w56572;
w56976 <= not w56568 and w56975;
w56977 <= not w56569 and not w56572;
w56978 <= not w56976 and not w56977;
w56979 <= not w56739 and not w56978;
w56980 <= not w55870 and not w56166;
w56981 <= not w56738 and w56980;
w56982 <= not w56979 and not w56981;
w56983 <= not w56167 and w56577;
w56984 <= not w56573 and w56983;
w56985 <= not w56574 and not w56577;
w56986 <= not w56984 and not w56985;
w56987 <= not w56739 and not w56986;
w56988 <= not w55870 and not w56157;
w56989 <= not w56738 and w56988;
w56990 <= not w56987 and not w56989;
w56991 <= not w56158 and w56582;
w56992 <= not w56578 and w56991;
w56993 <= not w56579 and not w56582;
w56994 <= not w56992 and not w56993;
w56995 <= not w56739 and not w56994;
w56996 <= not w55870 and not w56148;
w56997 <= not w56738 and w56996;
w56998 <= not w56995 and not w56997;
w56999 <= not w56149 and w56587;
w57000 <= not w56583 and w56999;
w57001 <= not w56584 and not w56587;
w57002 <= not w57000 and not w57001;
w57003 <= not w56739 and not w57002;
w57004 <= not w55870 and not w56139;
w57005 <= not w56738 and w57004;
w57006 <= not w57003 and not w57005;
w57007 <= not w56140 and w56592;
w57008 <= not w56588 and w57007;
w57009 <= not w56589 and not w56592;
w57010 <= not w57008 and not w57009;
w57011 <= not w56739 and not w57010;
w57012 <= not w55870 and not w56130;
w57013 <= not w56738 and w57012;
w57014 <= not w57011 and not w57013;
w57015 <= not w56131 and w56597;
w57016 <= not w56593 and w57015;
w57017 <= not w56594 and not w56597;
w57018 <= not w57016 and not w57017;
w57019 <= not w56739 and not w57018;
w57020 <= not w55870 and not w56121;
w57021 <= not w56738 and w57020;
w57022 <= not w57019 and not w57021;
w57023 <= not w56122 and w56602;
w57024 <= not w56598 and w57023;
w57025 <= not w56599 and not w56602;
w57026 <= not w57024 and not w57025;
w57027 <= not w56739 and not w57026;
w57028 <= not w55870 and not w56112;
w57029 <= not w56738 and w57028;
w57030 <= not w57027 and not w57029;
w57031 <= not w56113 and w56607;
w57032 <= not w56603 and w57031;
w57033 <= not w56604 and not w56607;
w57034 <= not w57032 and not w57033;
w57035 <= not w56739 and not w57034;
w57036 <= not w55870 and not w56103;
w57037 <= not w56738 and w57036;
w57038 <= not w57035 and not w57037;
w57039 <= not w56104 and w56612;
w57040 <= not w56608 and w57039;
w57041 <= not w56609 and not w56612;
w57042 <= not w57040 and not w57041;
w57043 <= not w56739 and not w57042;
w57044 <= not w55870 and not w56094;
w57045 <= not w56738 and w57044;
w57046 <= not w57043 and not w57045;
w57047 <= not w56095 and w56617;
w57048 <= not w56613 and w57047;
w57049 <= not w56614 and not w56617;
w57050 <= not w57048 and not w57049;
w57051 <= not w56739 and not w57050;
w57052 <= not w55870 and not w56085;
w57053 <= not w56738 and w57052;
w57054 <= not w57051 and not w57053;
w57055 <= not w56086 and w56622;
w57056 <= not w56618 and w57055;
w57057 <= not w56619 and not w56622;
w57058 <= not w57056 and not w57057;
w57059 <= not w56739 and not w57058;
w57060 <= not w55870 and not w56076;
w57061 <= not w56738 and w57060;
w57062 <= not w57059 and not w57061;
w57063 <= not w56077 and w56627;
w57064 <= not w56623 and w57063;
w57065 <= not w56624 and not w56627;
w57066 <= not w57064 and not w57065;
w57067 <= not w56739 and not w57066;
w57068 <= not w55870 and not w56067;
w57069 <= not w56738 and w57068;
w57070 <= not w57067 and not w57069;
w57071 <= not w56068 and w56632;
w57072 <= not w56628 and w57071;
w57073 <= not w56629 and not w56632;
w57074 <= not w57072 and not w57073;
w57075 <= not w56739 and not w57074;
w57076 <= not w55870 and not w56058;
w57077 <= not w56738 and w57076;
w57078 <= not w57075 and not w57077;
w57079 <= not w56059 and w56637;
w57080 <= not w56633 and w57079;
w57081 <= not w56634 and not w56637;
w57082 <= not w57080 and not w57081;
w57083 <= not w56739 and not w57082;
w57084 <= not w55870 and not w56049;
w57085 <= not w56738 and w57084;
w57086 <= not w57083 and not w57085;
w57087 <= not w56050 and w56642;
w57088 <= not w56638 and w57087;
w57089 <= not w56639 and not w56642;
w57090 <= not w57088 and not w57089;
w57091 <= not w56739 and not w57090;
w57092 <= not w55870 and not w56040;
w57093 <= not w56738 and w57092;
w57094 <= not w57091 and not w57093;
w57095 <= not w56041 and w56647;
w57096 <= not w56643 and w57095;
w57097 <= not w56644 and not w56647;
w57098 <= not w57096 and not w57097;
w57099 <= not w56739 and not w57098;
w57100 <= not w55870 and not w56031;
w57101 <= not w56738 and w57100;
w57102 <= not w57099 and not w57101;
w57103 <= not w56032 and w56652;
w57104 <= not w56648 and w57103;
w57105 <= not w56649 and not w56652;
w57106 <= not w57104 and not w57105;
w57107 <= not w56739 and not w57106;
w57108 <= not w55870 and not w56022;
w57109 <= not w56738 and w57108;
w57110 <= not w57107 and not w57109;
w57111 <= not w56023 and w56657;
w57112 <= not w56653 and w57111;
w57113 <= not w56654 and not w56657;
w57114 <= not w57112 and not w57113;
w57115 <= not w56739 and not w57114;
w57116 <= not w55870 and not w56013;
w57117 <= not w56738 and w57116;
w57118 <= not w57115 and not w57117;
w57119 <= not w56014 and w56662;
w57120 <= not w56658 and w57119;
w57121 <= not w56659 and not w56662;
w57122 <= not w57120 and not w57121;
w57123 <= not w56739 and not w57122;
w57124 <= not w55870 and not w56004;
w57125 <= not w56738 and w57124;
w57126 <= not w57123 and not w57125;
w57127 <= not w56005 and w56667;
w57128 <= not w56663 and w57127;
w57129 <= not w56664 and not w56667;
w57130 <= not w57128 and not w57129;
w57131 <= not w56739 and not w57130;
w57132 <= not w55870 and not w55995;
w57133 <= not w56738 and w57132;
w57134 <= not w57131 and not w57133;
w57135 <= not w55996 and w56672;
w57136 <= not w56668 and w57135;
w57137 <= not w56669 and not w56672;
w57138 <= not w57136 and not w57137;
w57139 <= not w56739 and not w57138;
w57140 <= not w55870 and not w55986;
w57141 <= not w56738 and w57140;
w57142 <= not w57139 and not w57141;
w57143 <= not w55987 and w56677;
w57144 <= not w56673 and w57143;
w57145 <= not w56674 and not w56677;
w57146 <= not w57144 and not w57145;
w57147 <= not w56739 and not w57146;
w57148 <= not w55870 and not w55977;
w57149 <= not w56738 and w57148;
w57150 <= not w57147 and not w57149;
w57151 <= not w55978 and w56682;
w57152 <= not w56678 and w57151;
w57153 <= not w56679 and not w56682;
w57154 <= not w57152 and not w57153;
w57155 <= not w56739 and not w57154;
w57156 <= not w55870 and not w55968;
w57157 <= not w56738 and w57156;
w57158 <= not w57155 and not w57157;
w57159 <= not w55969 and w56687;
w57160 <= not w56683 and w57159;
w57161 <= not w56684 and not w56687;
w57162 <= not w57160 and not w57161;
w57163 <= not w56739 and not w57162;
w57164 <= not w55870 and not w55959;
w57165 <= not w56738 and w57164;
w57166 <= not w57163 and not w57165;
w57167 <= not w55960 and w56692;
w57168 <= not w56688 and w57167;
w57169 <= not w56689 and not w56692;
w57170 <= not w57168 and not w57169;
w57171 <= not w56739 and not w57170;
w57172 <= not w55870 and not w55950;
w57173 <= not w56738 and w57172;
w57174 <= not w57171 and not w57173;
w57175 <= not w55951 and w56697;
w57176 <= not w56693 and w57175;
w57177 <= not w56694 and not w56697;
w57178 <= not w57176 and not w57177;
w57179 <= not w56739 and not w57178;
w57180 <= not w55870 and not w55941;
w57181 <= not w56738 and w57180;
w57182 <= not w57179 and not w57181;
w57183 <= not w55942 and w56702;
w57184 <= not w56698 and w57183;
w57185 <= not w56699 and not w56702;
w57186 <= not w57184 and not w57185;
w57187 <= not w56739 and not w57186;
w57188 <= not w55870 and not w55932;
w57189 <= not w56738 and w57188;
w57190 <= not w57187 and not w57189;
w57191 <= not w55933 and w56707;
w57192 <= not w56703 and w57191;
w57193 <= not w56704 and not w56707;
w57194 <= not w57192 and not w57193;
w57195 <= not w56739 and not w57194;
w57196 <= not w55870 and not w55923;
w57197 <= not w56738 and w57196;
w57198 <= not w57195 and not w57197;
w57199 <= not w55924 and w56712;
w57200 <= not w56708 and w57199;
w57201 <= not w56709 and not w56712;
w57202 <= not w57200 and not w57201;
w57203 <= not w56739 and not w57202;
w57204 <= not w55870 and not w55914;
w57205 <= not w56738 and w57204;
w57206 <= not w57203 and not w57205;
w57207 <= not w55915 and w56717;
w57208 <= not w56713 and w57207;
w57209 <= not w56714 and not w56717;
w57210 <= not w57208 and not w57209;
w57211 <= not w56739 and not w57210;
w57212 <= not w55870 and not w55905;
w57213 <= not w56738 and w57212;
w57214 <= not w57211 and not w57213;
w57215 <= not w55906 and w56722;
w57216 <= not w56718 and w57215;
w57217 <= not w56719 and not w56722;
w57218 <= not w57216 and not w57217;
w57219 <= not w56739 and not w57218;
w57220 <= not w55870 and not w55896;
w57221 <= not w56738 and w57220;
w57222 <= not w57219 and not w57221;
w57223 <= not w55897 and w56727;
w57224 <= not w56723 and w57223;
w57225 <= not w56724 and not w56727;
w57226 <= not w57224 and not w57225;
w57227 <= not w56739 and not w57226;
w57228 <= not w55870 and not w55887;
w57229 <= not w56738 and w57228;
w57230 <= not w57227 and not w57229;
w57231 <= not w55888 and w56732;
w57232 <= not w56728 and w57231;
w57233 <= not w56729 and not w56732;
w57234 <= not w57232 and not w57233;
w57235 <= not w56739 and not w57234;
w57236 <= not w55870 and not w55878;
w57237 <= not w56738 and w57236;
w57238 <= not w57235 and not w57237;
w57239 <= not w55879 and w56737;
w57240 <= not w56733 and w57239;
w57241 <= not w56734 and not w56737;
w57242 <= not w57240 and not w57241;
w57243 <= not w56739 and not w57242;
w57244 <= not w55869 and not w55870;
w57245 <= not w56738 and w57244;
w57246 <= not w57243 and not w57245;
one <= '1';
quotient(0) <= not w28664;-- level 4372
quotient(1) <= not w27847;-- level 4212
quotient(2) <= not w26978;-- level 4083
quotient(3) <= not w26123;-- level 3956
quotient(4) <= not w25282;-- level 3831
quotient(5) <= not w24455;-- level 3708
quotient(6) <= w23639;-- level 3588
quotient(7) <= not w22840;-- level 3468
quotient(8) <= not w22055;-- level 3351
quotient(9) <= w21281;-- level 3237
quotient(10) <= not w20523;-- level 3123
quotient(11) <= not w19778;-- level 3012
quotient(12) <= w19047;-- level 2904
quotient(13) <= not w18333;-- level 2796
quotient(14) <= not w17630;-- level 2691
quotient(15) <= w16938;-- level 2589
quotient(16) <= not w16266;-- level 2487
quotient(17) <= not w15607;-- level 2388
quotient(18) <= w14956;-- level 2292
quotient(19) <= not w14324;-- level 2196
quotient(20) <= not w13706;-- level 2103
quotient(21) <= w13099;-- level 2013
quotient(22) <= not w12509;-- level 1923
quotient(23) <= w11928;-- level 1837
quotient(24) <= w11363;-- level 1752
quotient(25) <= not w10816;-- level 1668
quotient(26) <= w10274;-- level 1588
quotient(27) <= w9748;-- level 1509
quotient(28) <= not w9244;-- level 1431
quotient(29) <= w8748;-- level 1357
quotient(30) <= w8263;-- level 1284
quotient(31) <= not w7798;-- level 1212
quotient(32) <= w7345;-- level 1144
quotient(33) <= w6906;-- level 1077
quotient(34) <= not w6483;-- level 1011
quotient(35) <= w6068;-- level 949
quotient(36) <= w5670;-- level 888
quotient(37) <= not w5290;-- level 828
quotient(38) <= w4916;-- level 772
quotient(39) <= w4557;-- level 717
quotient(40) <= not w4219;-- level 663
quotient(41) <= w3887;-- level 613
quotient(42) <= w3567;-- level 564
quotient(43) <= not w3269;-- level 516
quotient(44) <= w2982;-- level 472
quotient(45) <= w2709;-- level 429
quotient(46) <= not w2453;-- level 387
quotient(47) <= w2204;-- level 349
quotient(48) <= w1976;-- level 312
quotient(49) <= not w1766;-- level 276
quotient(50) <= w1560;-- level 244
quotient(51) <= w1370;-- level 213
quotient(52) <= not w1200;-- level 183
quotient(53) <= w1038;-- level 157
quotient(54) <= w889;-- level 132
quotient(55) <= not w760;-- level 108
quotient(56) <= w639;-- level 88
quotient(57) <= w532;-- level 69
quotient(58) <= not w448;-- level 51
quotient(59) <= w28665;-- level 37
quotient(60) <= w261;-- level 26
quotient(61) <= w194;-- level 17
quotient(62) <= w28668;-- level 10
quotient(63) <= w28673;-- level 7
remainder(0) <= not w56743;-- level 4345
remainder(1) <= not w56750;-- level 4344
remainder(2) <= not w56758;-- level 4344
remainder(3) <= not w56766;-- level 4344
remainder(4) <= not w56774;-- level 4344
remainder(5) <= not w56782;-- level 4344
remainder(6) <= not w56790;-- level 4344
remainder(7) <= not w56798;-- level 4344
remainder(8) <= not w56806;-- level 4344
remainder(9) <= not w56814;-- level 4344
remainder(10) <= not w56822;-- level 4344
remainder(11) <= not w56830;-- level 4344
remainder(12) <= not w56838;-- level 4344
remainder(13) <= not w56846;-- level 4344
remainder(14) <= not w56854;-- level 4344
remainder(15) <= not w56862;-- level 4344
remainder(16) <= not w56870;-- level 4344
remainder(17) <= not w56878;-- level 4344
remainder(18) <= not w56886;-- level 4344
remainder(19) <= not w56894;-- level 4344
remainder(20) <= not w56902;-- level 4344
remainder(21) <= not w56910;-- level 4344
remainder(22) <= not w56918;-- level 4344
remainder(23) <= not w56926;-- level 4344
remainder(24) <= not w56934;-- level 4344
remainder(25) <= not w56942;-- level 4344
remainder(26) <= not w56950;-- level 4344
remainder(27) <= not w56958;-- level 4344
remainder(28) <= not w56966;-- level 4344
remainder(29) <= not w56974;-- level 4344
remainder(30) <= not w56982;-- level 4344
remainder(31) <= not w56990;-- level 4344
remainder(32) <= not w56998;-- level 4344
remainder(33) <= not w57006;-- level 4344
remainder(34) <= not w57014;-- level 4344
remainder(35) <= not w57022;-- level 4344
remainder(36) <= not w57030;-- level 4344
remainder(37) <= not w57038;-- level 4344
remainder(38) <= not w57046;-- level 4344
remainder(39) <= not w57054;-- level 4344
remainder(40) <= not w57062;-- level 4344
remainder(41) <= not w57070;-- level 4344
remainder(42) <= not w57078;-- level 4344
remainder(43) <= not w57086;-- level 4344
remainder(44) <= not w57094;-- level 4344
remainder(45) <= not w57102;-- level 4344
remainder(46) <= not w57110;-- level 4344
remainder(47) <= not w57118;-- level 4344
remainder(48) <= not w57126;-- level 4344
remainder(49) <= not w57134;-- level 4344
remainder(50) <= not w57142;-- level 4344
remainder(51) <= not w57150;-- level 4344
remainder(52) <= not w57158;-- level 4344
remainder(53) <= not w57166;-- level 4344
remainder(54) <= not w57174;-- level 4344
remainder(55) <= not w57182;-- level 4344
remainder(56) <= not w57190;-- level 4344
remainder(57) <= not w57198;-- level 4344
remainder(58) <= not w57206;-- level 4344
remainder(59) <= not w57214;-- level 4344
remainder(60) <= not w57222;-- level 4344
remainder(61) <= not w57230;-- level 4344
remainder(62) <= not w57238;-- level 4344
remainder(63) <= not w57246;-- level 4344
end Behavioral;
