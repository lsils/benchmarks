library ieee;
use ieee.std_logic_1164.all;

entity top is
	port (
totalcoeffs : in std_logic_vector(4 downto 0);
ctable : in std_logic_vector(2 downto 0);
trailingones : in std_logic_vector(1 downto 0);
coeff_token : out std_logic_vector(5 downto 0);
ctoken_len : out std_logic_vector(4 downto 0)
);
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692: std_logic;

begin

w0 <= not totalcoeffs(3) and not ctable(0);
w1 <= not totalcoeffs(1) and trailingones(1);
w2 <= not totalcoeffs(0) and trailingones(1);
w3 <= totalcoeffs(1) and not w2;
w4 <= not w1 and not w3;
w5 <= w0 and w4;
w6 <= totalcoeffs(0) and not trailingones(1);
w7 <= not totalcoeffs(1) and not w6;
w8 <= totalcoeffs(1) and not trailingones(1);
w9 <= not ctable(2) and not w8;
w10 <= not w7 and w9;
w11 <= not w5 and not w10;
w12 <= not totalcoeffs(2) and not w11;
w13 <= not totalcoeffs(2) and not ctable(0);
w14 <= not totalcoeffs(0) and not w13;
w15 <= totalcoeffs(1) and totalcoeffs(2);
w16 <= not w14 and not w15;
w17 <= not trailingones(1) and not w16;
w18 <= not totalcoeffs(2) and not totalcoeffs(3);
w19 <= trailingones(1) and not w18;
w20 <= totalcoeffs(0) and totalcoeffs(3);
w21 <= not w19 and not w20;
w22 <= not totalcoeffs(1) and not w21;
w23 <= totalcoeffs(1) and not totalcoeffs(3);
w24 <= not w22 and not w23;
w25 <= not w17 and w24;
w26 <= not ctable(2) and not w25;
w27 <= not w12 and not w26;
w28 <= not trailingones(0) and not w27;
w29 <= ctable(2) and trailingones(0);
w30 <= not ctable(0) and w29;
w31 <= not ctable(2) and trailingones(1);
w32 <= not w30 and not w31;
w33 <= totalcoeffs(1) and not w32;
w34 <= totalcoeffs(1) and not ctable(2);
w35 <= not ctable(0) and not trailingones(1);
w36 <= not w34 and w35;
w37 <= not w33 and not w36;
w38 <= totalcoeffs(0) and not totalcoeffs(2);
w39 <= not w37 and w38;
w40 <= totalcoeffs(2) and not trailingones(1);
w41 <= not totalcoeffs(0) and not totalcoeffs(1);
w42 <= w40 and w41;
w43 <= w30 and w42;
w44 <= not w39 and not w43;
w45 <= not totalcoeffs(3) and not w44;
w46 <= not w28 and not w45;
w47 <= not ctable(1) and not w46;
w48 <= not totalcoeffs(0) and not totalcoeffs(2);
w49 <= w1 and w48;
w50 <= not ctable(0) and not w49;
w51 <= ctable(1) and not w50;
w52 <= not totalcoeffs(0) and not trailingones(1);
w53 <= totalcoeffs(0) and trailingones(1);
w54 <= not w52 and not w53;
w55 <= totalcoeffs(1) and not w54;
w56 <= totalcoeffs(2) and w55;
w57 <= ctable(0) and w56;
w58 <= not w51 and not w57;
w59 <= trailingones(0) and not w58;
w60 <= not totalcoeffs(1) and not w2;
w61 <= not trailingones(0) and not w60;
w62 <= not totalcoeffs(1) and totalcoeffs(2);
w63 <= w6 and w62;
w64 <= not w61 and not w63;
w65 <= not ctable(0) and not w64;
w66 <= not w59 and not w65;
w67 <= totalcoeffs(3) and not w66;
w68 <= not totalcoeffs(2) and not w6;
w69 <= ctable(1) and not w68;
w70 <= w18 and w55;
w71 <= not w69 and not w70;
w72 <= ctable(0) and not w71;
w73 <= totalcoeffs(2) and trailingones(1);
w74 <= not totalcoeffs(2) and w8;
w75 <= not w73 and not w74;
w76 <= not totalcoeffs(0) and not totalcoeffs(3);
w77 <= not w75 and w76;
w78 <= ctable(1) and w77;
w79 <= not w72 and not w78;
w80 <= trailingones(0) and not w79;
w81 <= totalcoeffs(2) and not totalcoeffs(3);
w82 <= w1 and w81;
w83 <= totalcoeffs(1) and not trailingones(0);
w84 <= not w82 and not w83;
w85 <= not totalcoeffs(0) and not w84;
w86 <= not totalcoeffs(1) and not trailingones(1);
w87 <= not totalcoeffs(2) and ctable(1);
w88 <= totalcoeffs(3) and not w87;
w89 <= w86 and not w88;
w90 <= not w73 and not w89;
w91 <= not trailingones(0) and not w90;
w92 <= not w85 and not w91;
w93 <= not ctable(0) and not w92;
w94 <= not totalcoeffs(0) and w18;
w95 <= not trailingones(0) and w86;
w96 <= w94 and w95;
w97 <= not w93 and not w96;
w98 <= not w80 and w97;
w99 <= not w67 and w98;
w100 <= not ctable(2) and not w99;
w101 <= not w47 and not w100;
w102 <= not totalcoeffs(4) and not w101;
w103 <= not trailingones(0) and not trailingones(1);
w104 <= not ctable(1) and w103;
w105 <= totalcoeffs(4) and trailingones(0);
w106 <= ctable(1) and w105;
w107 <= not w104 and not w106;
w108 <= ctable(0) and not w107;
w109 <= ctable(1) and not trailingones(1);
w110 <= totalcoeffs(4) and trailingones(1);
w111 <= not w109 and not w110;
w112 <= ctable(0) and ctable(1);
w113 <= not w111 and not w112;
w114 <= not trailingones(0) and w113;
w115 <= not w108 and not w114;
w116 <= not ctable(2) and not w115;
w117 <= not totalcoeffs(1) and not totalcoeffs(3);
w118 <= not totalcoeffs(2) and w117;
w119 <= w116 and w118;
w120 <= not totalcoeffs(0) and w119;
w121 <= not w102 and not w120;
w122 <= totalcoeffs(0) and trailingones(0);
w123 <= w73 and w122;
w124 <= not totalcoeffs(2) and not trailingones(0);
w125 <= w52 and w124;
w126 <= not w123 and not w125;
w127 <= ctable(0) and not w126;
w128 <= not ctable(0) and trailingones(0);
w129 <= ctable(1) and trailingones(1);
w130 <= not w128 and not w129;
w131 <= not totalcoeffs(0) and not w130;
w132 <= trailingones(0) and w129;
w133 <= not trailingones(0) and w35;
w134 <= not w132 and not w133;
w135 <= not w131 and w134;
w136 <= totalcoeffs(2) and not w135;
w137 <= not w127 and not w136;
w138 <= not totalcoeffs(4) and not w137;
w139 <= not ctable(1) and trailingones(1);
w140 <= ctable(0) and not trailingones(0);
w141 <= not w105 and not w140;
w142 <= not ctable(1) and not w141;
w143 <= not w110 and not w142;
w144 <= not w139 and not w143;
w145 <= w48 and w144;
w146 <= not w138 and not w145;
w147 <= not totalcoeffs(1) and not w146;
w148 <= ctable(1) and trailingones(0);
w149 <= not w130 and not w148;
w150 <= totalcoeffs(0) and w149;
w151 <= not totalcoeffs(0) and ctable(0);
w152 <= not trailingones(0) and trailingones(1);
w153 <= w151 and w152;
w154 <= not w150 and not w153;
w155 <= not totalcoeffs(2) and not w154;
w156 <= not ctable(1) and not trailingones(0);
w157 <= not totalcoeffs(0) and ctable(1);
w158 <= not totalcoeffs(2) and not w157;
w159 <= w128 and not w158;
w160 <= not w156 and not w159;
w161 <= not trailingones(1) and not w160;
w162 <= not w155 and not w161;
w163 <= totalcoeffs(1) and not w162;
w164 <= not ctable(1) and trailingones(0);
w165 <= w40 and w164;
w166 <= not w163 and not w165;
w167 <= not totalcoeffs(4) and not w166;
w168 <= not w147 and not w167;
w169 <= not totalcoeffs(3) and not w168;
w170 <= ctable(0) and w124;
w171 <= not totalcoeffs(3) and not trailingones(0);
w172 <= not w128 and not w171;
w173 <= totalcoeffs(0) and w172;
w174 <= not w170 and not w173;
w175 <= not totalcoeffs(1) and not w174;
w176 <= totalcoeffs(3) and trailingones(0);
w177 <= not totalcoeffs(2) and not w176;
w178 <= not totalcoeffs(0) and not w177;
w179 <= not totalcoeffs(2) and trailingones(0);
w180 <= totalcoeffs(0) and w179;
w181 <= totalcoeffs(0) and not ctable(0);
w182 <= not w151 and not w181;
w183 <= not w180 and w182;
w184 <= totalcoeffs(1) and not w183;
w185 <= not w178 and not w184;
w186 <= not w175 and w185;
w187 <= not ctable(1) and not w186;
w188 <= not totalcoeffs(1) and ctable(1);
w189 <= totalcoeffs(2) and not w188;
w190 <= not totalcoeffs(1) and not trailingones(0);
w191 <= not w189 and not w190;
w192 <= totalcoeffs(3) and w191;
w193 <= not totalcoeffs(0) and trailingones(0);
w194 <= not totalcoeffs(1) and not ctable(1);
w195 <= totalcoeffs(0) and totalcoeffs(1);
w196 <= not w194 and not w195;
w197 <= not w193 and w196;
w198 <= not totalcoeffs(2) and w197;
w199 <= not w192 and not w198;
w200 <= not ctable(0) and not w199;
w201 <= not w187 and not w200;
w202 <= not trailingones(1) and not w201;
w203 <= totalcoeffs(1) and ctable(0);
w204 <= totalcoeffs(3) and not trailingones(0);
w205 <= not totalcoeffs(1) and not totalcoeffs(2);
w206 <= w204 and w205;
w207 <= not w203 and not w206;
w208 <= totalcoeffs(0) and not w207;
w209 <= ctable(0) and not w18;
w210 <= totalcoeffs(3) and w15;
w211 <= not w209 and not w210;
w212 <= not w208 and w211;
w213 <= ctable(1) and not w212;
w214 <= w140 and w210;
w215 <= not w213 and not w214;
w216 <= trailingones(1) and not w215;
w217 <= not w202 and not w216;
w218 <= not totalcoeffs(4) and not w217;
w219 <= not w169 and not w218;
w220 <= not ctable(2) and not w219;
w221 <= totalcoeffs(2) and not w41;
w222 <= w68 and not w195;
w223 <= not w221 and not w222;
w224 <= not trailingones(0) and w223;
w225 <= w8 and w179;
w226 <= not w224 and not w225;
w227 <= ctable(2) and not w226;
w228 <= not w42 and not w227;
w229 <= not totalcoeffs(4) and not w228;
w230 <= not ctable(1) and w229;
w231 <= w0 and w230;
w232 <= not w220 and not w231;
w233 <= not totalcoeffs(3) and trailingones(1);
w234 <= not w23 and not w152;
w235 <= not w233 and not w234;
w236 <= not ctable(1) and w235;
w237 <= totalcoeffs(3) and not w179;
w238 <= ctable(0) and not w237;
w239 <= totalcoeffs(2) and not ctable(0);
w240 <= totalcoeffs(3) and not w239;
w241 <= trailingones(0) and not w240;
w242 <= not w238 and not w241;
w243 <= totalcoeffs(1) and not w242;
w244 <= not ctable(0) and ctable(1);
w245 <= not trailingones(0) and w244;
w246 <= w117 and w245;
w247 <= not w243 and not w246;
w248 <= not trailingones(1) and not w247;
w249 <= not totalcoeffs(1) and not w177;
w250 <= totalcoeffs(2) and not w164;
w251 <= not w249 and not w250;
w252 <= ctable(0) and not w251;
w253 <= totalcoeffs(1) and trailingones(0);
w254 <= ctable(1) and not w253;
w255 <= not trailingones(1) and not w254;
w256 <= not totalcoeffs(2) and not w255;
w257 <= not totalcoeffs(1) and w152;
w258 <= not w256 and not w257;
w259 <= totalcoeffs(3) and not w258;
w260 <= ctable(1) and not trailingones(0);
w261 <= totalcoeffs(1) and w233;
w262 <= w260 and w261;
w263 <= not w259 and not w262;
w264 <= not w252 and w263;
w265 <= not w248 and w264;
w266 <= not w236 and w265;
w267 <= not totalcoeffs(4) and not w266;
w268 <= trailingones(0) and not trailingones(1);
w269 <= not w156 and not w268;
w270 <= not ctable(0) and w269;
w271 <= not totalcoeffs(3) and totalcoeffs(4);
w272 <= not totalcoeffs(1) and w271;
w273 <= not w270 and w272;
w274 <= not totalcoeffs(2) and w273;
w275 <= not w267 and not w274;
w276 <= not totalcoeffs(0) and not w275;
w277 <= trailingones(0) and w53;
w278 <= not w103 and not w277;
w279 <= ctable(0) and not w278;
w280 <= not ctable(0) and w73;
w281 <= not w279 and not w280;
w282 <= totalcoeffs(1) and not w281;
w283 <= not w152 and not w268;
w284 <= not w86 and w283;
w285 <= totalcoeffs(2) and not w284;
w286 <= not w282 and not w285;
w287 <= not totalcoeffs(3) and not w286;
w288 <= not totalcoeffs(1) and totalcoeffs(3);
w289 <= ctable(0) and not w288;
w290 <= not totalcoeffs(2) and w103;
w291 <= not w289 and w290;
w292 <= not totalcoeffs(1) and trailingones(0);
w293 <= w19 and w292;
w294 <= not w291 and not w293;
w295 <= totalcoeffs(0) and not w294;
w296 <= not w287 and not w295;
w297 <= not ctable(1) and not w296;
w298 <= totalcoeffs(1) and trailingones(1);
w299 <= totalcoeffs(2) and w298;
w300 <= not w292 and not w299;
w301 <= ctable(1) and not w300;
w302 <= trailingones(0) and not w40;
w303 <= totalcoeffs(2) and w103;
w304 <= not w302 and not w303;
w305 <= not w301 and w304;
w306 <= totalcoeffs(3) and not w305;
w307 <= ctable(1) and not w1;
w308 <= not w8 and not w307;
w309 <= trailingones(0) and not w308;
w310 <= not w86 and not w298;
w311 <= w171 and not w310;
w312 <= not w309 and not w311;
w313 <= not totalcoeffs(2) and not w312;
w314 <= not w306 and not w313;
w315 <= w181 and not w314;
w316 <= not w297 and not w315;
w317 <= not totalcoeffs(4) and not w316;
w318 <= not w276 and not w317;
w319 <= not ctable(2) and not w318;
w320 <= not ctable(0) and not ctable(1);
w321 <= w29 and w53;
w322 <= not w52 and not w321;
w323 <= totalcoeffs(1) and not w322;
w324 <= w6 and w190;
w325 <= not w323 and not w324;
w326 <= not totalcoeffs(4) and not w325;
w327 <= w18 and w326;
w328 <= w320 and w327;
w329 <= not w319 and not w328;
w330 <= totalcoeffs(3) and not w139;
w331 <= totalcoeffs(2) and ctable(1);
w332 <= not w330 and not w331;
w333 <= not totalcoeffs(4) and not w332;
w334 <= trailingones(0) and trailingones(1);
w335 <= w320 and w334;
w336 <= not w112 and not w335;
w337 <= not totalcoeffs(2) and w271;
w338 <= not w336 and w337;
w339 <= not w333 and not w338;
w340 <= not totalcoeffs(1) and not w339;
w341 <= ctable(0) and trailingones(0);
w342 <= w139 and w341;
w343 <= not w133 and not w342;
w344 <= totalcoeffs(2) and not w343;
w345 <= ctable(0) and not w164;
w346 <= totalcoeffs(3) and not w345;
w347 <= not w245 and not w346;
w348 <= not w344 and w347;
w349 <= totalcoeffs(1) and not w348;
w350 <= totalcoeffs(2) and w244;
w351 <= not w349 and not w350;
w352 <= not totalcoeffs(4) and not w351;
w353 <= not w340 and not w352;
w354 <= not totalcoeffs(0) and not w353;
w355 <= totalcoeffs(2) and not w172;
w356 <= not totalcoeffs(2) and w341;
w357 <= not w355 and not w356;
w358 <= not trailingones(1) and not w357;
w359 <= ctable(0) and trailingones(1);
w360 <= not trailingones(0) and w359;
w361 <= not totalcoeffs(3) and not w360;
w362 <= not totalcoeffs(2) and not w361;
w363 <= not ctable(1) and not w204;
w364 <= totalcoeffs(3) and not ctable(0);
w365 <= not w363 and not w364;
w366 <= not w362 and not w365;
w367 <= not w358 and w366;
w368 <= totalcoeffs(1) and not w367;
w369 <= not totalcoeffs(3) and w244;
w370 <= w170 and w194;
w371 <= not w369 and not w370;
w372 <= not trailingones(1) and not w371;
w373 <= not w368 and not w372;
w374 <= totalcoeffs(0) and not w373;
w375 <= not w18 and w244;
w376 <= totalcoeffs(3) and not ctable(1);
w377 <= totalcoeffs(2) and w376;
w378 <= not w375 and not w377;
w379 <= trailingones(1) and not w378;
w380 <= not trailingones(1) and w244;
w381 <= not w376 and not w380;
w382 <= not trailingones(0) and not w381;
w383 <= not w379 and not w382;
w384 <= not totalcoeffs(1) and not w383;
w385 <= not w35 and not w156;
w386 <= not totalcoeffs(2) and not w385;
w387 <= not ctable(1) and not w359;
w388 <= not w298 and not w341;
w389 <= w387 and not w388;
w390 <= not w386 and not w389;
w391 <= totalcoeffs(3) and not w390;
w392 <= totalcoeffs(1) and w268;
w393 <= w244 and w392;
w394 <= not w391 and not w393;
w395 <= not w384 and w394;
w396 <= not w374 and w395;
w397 <= not totalcoeffs(4) and not w396;
w398 <= not w354 and not w397;
w399 <= not ctable(2) and not w398;
w400 <= not totalcoeffs(4) and w221;
w401 <= totalcoeffs(3) and not totalcoeffs(4);
w402 <= not w271 and not w401;
w403 <= not totalcoeffs(0) and w205;
w404 <= not w402 and w403;
w405 <= not w400 and not w404;
w406 <= not ctable(2) and not w405;
w407 <= w112 and w406;
w408 <= w41 and w337;
w409 <= w401 and not w403;
w410 <= not w408 and not w409;
w411 <= not ctable(2) and not w410;
w412 <= w112 and w411;
w413 <= not totalcoeffs(1) and not ctable(0);
w414 <= totalcoeffs(2) and not w413;
w415 <= not trailingones(1) and not w414;
w416 <= not ctable(1) and w415;
w417 <= ctable(0) and w298;
w418 <= not w416 and not w417;
w419 <= totalcoeffs(0) and not w418;
w420 <= not totalcoeffs(0) and not w35;
w421 <= totalcoeffs(2) and w420;
w422 <= not w419 and not w421;
w423 <= trailingones(0) and not w422;
w424 <= totalcoeffs(2) and w2;
w425 <= not w95 and not w424;
w426 <= ctable(0) and not w425;
w427 <= not w423 and not w426;
w428 <= not w103 and not w334;
w429 <= ctable(1) and not w428;
w430 <= not totalcoeffs(2) and trailingones(1);
w431 <= not w40 and not w430;
w432 <= w429 and w431;
w433 <= w427 and not w432;
w434 <= not ctable(2) and not w433;
w435 <= ctable(2) and not trailingones(1);
w436 <= trailingones(0) and not w435;
w437 <= w62 and not w436;
w438 <= not w74 and not w437;
w439 <= not totalcoeffs(0) and not w438;
w440 <= w122 and w298;
w441 <= not w103 and not w440;
w442 <= ctable(2) and not w441;
w443 <= not totalcoeffs(2) and w442;
w444 <= not w439 and not w443;
w445 <= w320 and not w444;
w446 <= not w434 and not w445;
w447 <= not totalcoeffs(3) and not w446;
w448 <= not w95 and not w298;
w449 <= totalcoeffs(0) and not w448;
w450 <= totalcoeffs(2) and w8;
w451 <= not w449 and not w450;
w452 <= not totalcoeffs(0) and not ctable(1);
w453 <= not w190 and w310;
w454 <= w452 and w453;
w455 <= w451 and not w454;
w456 <= not ctable(0) and not w455;
w457 <= not trailingones(0) and w195;
w458 <= totalcoeffs(0) and w148;
w459 <= not w83 and not w458;
w460 <= not totalcoeffs(2) and not w459;
w461 <= not w457 and not w460;
w462 <= trailingones(1) and not w461;
w463 <= not totalcoeffs(0) and not trailingones(0);
w464 <= not w181 and not w463;
w465 <= w8 and w464;
w466 <= not w462 and not w465;
w467 <= not w456 and w466;
w468 <= totalcoeffs(3) and not w467;
w469 <= not totalcoeffs(2) and ctable(0);
w470 <= not w54 and w469;
w471 <= not ctable(1) and not w239;
w472 <= w2 and not w471;
w473 <= not w470 and not w472;
w474 <= not trailingones(0) and not w473;
w475 <= totalcoeffs(2) and not w103;
w476 <= not w277 and not w475;
w477 <= ctable(1) and not w476;
w478 <= not w474 and not w477;
w479 <= totalcoeffs(1) and not w478;
w480 <= not trailingones(0) and not w452;
w481 <= not w181 and not w480;
w482 <= not trailingones(1) and not w481;
w483 <= not totalcoeffs(2) and w482;
w484 <= totalcoeffs(2) and trailingones(0);
w485 <= w2 and w484;
w486 <= not w483 and not w485;
w487 <= not totalcoeffs(1) and not w486;
w488 <= not w479 and not w487;
w489 <= not w468 and w488;
w490 <= not ctable(2) and not w489;
w491 <= not w447 and not w490;
w492 <= not totalcoeffs(4) and not w491;
w493 <= not totalcoeffs(1) and totalcoeffs(4);
w494 <= w94 and w493;
w495 <= not w112 and not w494;
w496 <= not ctable(2) and not w495;
w497 <= not w492 and not w496;
w498 <= not totalcoeffs(3) and trailingones(0);
w499 <= not w129 and not w498;
w500 <= totalcoeffs(0) and not w499;
w501 <= w193 and w376;
w502 <= not w260 and not w501;
w503 <= trailingones(1) and not w502;
w504 <= not trailingones(1) and w148;
w505 <= not w503 and not w504;
w506 <= not w500 and w505;
w507 <= not totalcoeffs(2) and not w506;
w508 <= not totalcoeffs(3) and w334;
w509 <= totalcoeffs(3) and not w334;
w510 <= not w122 and not w509;
w511 <= not ctable(1) and not w510;
w512 <= not w508 and not w511;
w513 <= totalcoeffs(2) and not w512;
w514 <= not totalcoeffs(3) and w104;
w515 <= not w513 and not w514;
w516 <= not w507 and w515;
w517 <= totalcoeffs(1) and not w516;
w518 <= not w52 and not w152;
w519 <= not ctable(1) and not w518;
w520 <= not totalcoeffs(2) and w519;
w521 <= not totalcoeffs(0) and w429;
w522 <= not w520 and not w521;
w523 <= totalcoeffs(3) and not w522;
w524 <= not totalcoeffs(0) and w124;
w525 <= not w458 and not w524;
w526 <= not trailingones(1) and not w525;
w527 <= not ctable(1) and not w171;
w528 <= w475 and not w527;
w529 <= not w526 and not w528;
w530 <= not w523 and w529;
w531 <= not totalcoeffs(1) and not w530;
w532 <= not totalcoeffs(2) and totalcoeffs(3);
w533 <= not trailingones(1) and w260;
w534 <= w532 and w533;
w535 <= not w531 and not w534;
w536 <= not w517 and w535;
w537 <= not ctable(0) and not w536;
w538 <= totalcoeffs(0) and not w431;
w539 <= ctable(0) and not trailingones(1);
w540 <= not totalcoeffs(0) and w539;
w541 <= not w538 and not w540;
w542 <= trailingones(0) and not w541;
w543 <= w73 and w140;
w544 <= not w542 and not w543;
w545 <= not totalcoeffs(3) and not w544;
w546 <= totalcoeffs(3) and ctable(0);
w547 <= not w40 and not w546;
w548 <= not totalcoeffs(0) and not w547;
w549 <= totalcoeffs(3) and w469;
w550 <= not w548 and not w549;
w551 <= not trailingones(0) and not w550;
w552 <= w532 and w539;
w553 <= not w551 and not w552;
w554 <= not w545 and w553;
w555 <= totalcoeffs(1) and not w554;
w556 <= totalcoeffs(2) and totalcoeffs(3);
w557 <= not totalcoeffs(2) and not w20;
w558 <= not w428 and not w557;
w559 <= not w556 and not w558;
w560 <= ctable(0) and not w559;
w561 <= w20 and w303;
w562 <= not w560 and not w561;
w563 <= not totalcoeffs(1) and not w562;
w564 <= trailingones(0) and w359;
w565 <= w556 and w564;
w566 <= not w563 and not w565;
w567 <= not w555 and w566;
w568 <= not ctable(1) and not w567;
w569 <= not w537 and not w568;
w570 <= not ctable(2) and not w569;
w571 <= totalcoeffs(2) and not w283;
w572 <= not totalcoeffs(0) and w571;
w573 <= not trailingones(1) and w29;
w574 <= w38 and w573;
w575 <= not w572 and not w574;
w576 <= w194 and not w575;
w577 <= w0 and w576;
w578 <= not w570 and not w577;
w579 <= not totalcoeffs(4) and not w578;
w580 <= w13 and w76;
w581 <= totalcoeffs(4) and not ctable(2);
w582 <= w194 and w581;
w583 <= w580 and w582;
w584 <= not w579 and not w583;
w585 <= w205 and w539;
w586 <= not w261 and not w585;
w587 <= not totalcoeffs(0) and not w586;
w588 <= not totalcoeffs(1) and ctable(0);
w589 <= not w0 and not w588;
w590 <= not w86 and not w233;
w591 <= not w589 and w590;
w592 <= not totalcoeffs(2) and w591;
w593 <= w310 and not w413;
w594 <= w81 and not w593;
w595 <= not w592 and not w594;
w596 <= not w587 and w595;
w597 <= not trailingones(0) and not w596;
w598 <= not w76 and not w589;
w599 <= not totalcoeffs(2) and w598;
w600 <= w117 and w181;
w601 <= not w599 and not w600;
w602 <= trailingones(0) and not w601;
w603 <= not ctable(0) and not w193;
w604 <= not w546 and not w603;
w605 <= w15 and w604;
w606 <= not w602 and not w605;
w607 <= not trailingones(1) and not w606;
w608 <= not w239 and not w546;
w609 <= not w237 and not w608;
w610 <= totalcoeffs(1) and w609;
w611 <= not w151 and w288;
w612 <= w179 and w611;
w613 <= not w610 and not w612;
w614 <= trailingones(1) and not w613;
w615 <= not w607 and not w614;
w616 <= not w597 and w615;
w617 <= not ctable(1) and not w616;
w618 <= not totalcoeffs(1) and not w103;
w619 <= totalcoeffs(2) and not w618;
w620 <= not w307 and not w619;
w621 <= totalcoeffs(0) and not w620;
w622 <= not ctable(1) and not w83;
w623 <= totalcoeffs(2) and not w622;
w624 <= trailingones(0) and not w8;
w625 <= w307 and not w624;
w626 <= not w623 and not w625;
w627 <= not w621 and w626;
w628 <= w364 and not w627;
w629 <= not w617 and not w628;
w630 <= not ctable(2) and not w629;
w631 <= not w124 and not w484;
w632 <= not totalcoeffs(0) and not w631;
w633 <= not w180 and not w632;
w634 <= not trailingones(1) and not w633;
w635 <= w73 and w463;
w636 <= not w634 and not w635;
w637 <= not totalcoeffs(1) and not w636;
w638 <= w298 and w524;
w639 <= not w637 and not w638;
w640 <= w0 and not w639;
w641 <= not ctable(1) and w640;
w642 <= not w630 and not w641;
w643 <= not totalcoeffs(4) and not w642;
w644 <= w0 and w581;
w645 <= w403 and w644;
w646 <= not w643 and not w645;
w647 <= totalcoeffs(4) and not w118;
w648 <= w181 and w377;
w649 <= not ctable(2) and not w648;
w650 <= not w618 and not w649;
w651 <= not ctable(2) and not w118;
w652 <= totalcoeffs(0) and not w651;
w653 <= ctable(2) and not w81;
w654 <= not totalcoeffs(3) and not w35;
w655 <= totalcoeffs(3) and not w129;
w656 <= w193 and not w655;
w657 <= not w654 and not w656;
w658 <= not totalcoeffs(2) and not w657;
w659 <= not w334 and w377;
w660 <= not ctable(0) and w659;
w661 <= not ctable(1) and not w564;
w662 <= not totalcoeffs(3) and not w661;
w663 <= not w660 and not w662;
w664 <= not w658 and w663;
w665 <= totalcoeffs(1) and not w664;
w666 <= w193 and not w387;
w667 <= not w129 and not w666;
w668 <= totalcoeffs(3) and not w667;
w669 <= totalcoeffs(4) and not w320;
w670 <= not totalcoeffs(3) and not w669;
w671 <= not w668 and not w670;
w672 <= not totalcoeffs(2) and not w671;
w673 <= not trailingones(0) and not w359;
w674 <= w654 and not w673;
w675 <= totalcoeffs(2) and w674;
w676 <= not w672 and not w675;
w677 <= not totalcoeffs(1) and not w676;
w678 <= not ctable(0) and not w81;
w679 <= ctable(1) and not w678;
w680 <= not w677 and not w679;
w681 <= not w665 and w680;
w682 <= not w653 and w681;
w683 <= not w652 and w682;
w684 <= not w650 and w683;
w685 <= not w647 and w684;
w686 <= not trailingones(0) and not w7;
w687 <= not w3 and not w686;
w688 <= w401 and not w687;
w689 <= totalcoeffs(2) and w688;
w690 <= not w408 and not w689;
w691 <= not ctable(2) and not w690;
w692 <= w320 and w691;
one <= '1';
coeff_token(0) <= not w121;-- level 14
coeff_token(1) <= not w232;-- level 15
coeff_token(2) <= not w329;-- level 16
coeff_token(3) <= w399;-- level 13
coeff_token(4) <= w407;-- level 6
coeff_token(5) <= w412;-- level 6
ctoken_len(0) <= w497;-- level 16
ctoken_len(1) <= w584;-- level 16
ctoken_len(2) <= w646;-- level 16
ctoken_len(3) <= w685;-- level 15
ctoken_len(4) <= w692;-- level 9
end Behavioral;
